
module loss ( clk, reset, model, .yHat({\yHat[15][19] , \yHat[15][18] , 
        \yHat[15][17] , \yHat[15][16] , \yHat[15][15] , \yHat[15][14] , 
        \yHat[15][13] , \yHat[15][12] , \yHat[15][11] , \yHat[15][10] , 
        \yHat[15][9] , \yHat[15][8] , \yHat[15][7] , \yHat[15][6] , 
        \yHat[15][5] , \yHat[15][4] , \yHat[15][3] , \yHat[15][2] , 
        \yHat[15][1] , \yHat[15][0] , \yHat[14][19] , \yHat[14][18] , 
        \yHat[14][17] , \yHat[14][16] , \yHat[14][15] , \yHat[14][14] , 
        \yHat[14][13] , \yHat[14][12] , \yHat[14][11] , \yHat[14][10] , 
        \yHat[14][9] , \yHat[14][8] , \yHat[14][7] , \yHat[14][6] , 
        \yHat[14][5] , \yHat[14][4] , \yHat[14][3] , \yHat[14][2] , 
        \yHat[14][1] , \yHat[14][0] , \yHat[13][19] , \yHat[13][18] , 
        \yHat[13][17] , \yHat[13][16] , \yHat[13][15] , \yHat[13][14] , 
        \yHat[13][13] , \yHat[13][12] , \yHat[13][11] , \yHat[13][10] , 
        \yHat[13][9] , \yHat[13][8] , \yHat[13][7] , \yHat[13][6] , 
        \yHat[13][5] , \yHat[13][4] , \yHat[13][3] , \yHat[13][2] , 
        \yHat[13][1] , \yHat[13][0] , \yHat[12][19] , \yHat[12][18] , 
        \yHat[12][17] , \yHat[12][16] , \yHat[12][15] , \yHat[12][14] , 
        \yHat[12][13] , \yHat[12][12] , \yHat[12][11] , \yHat[12][10] , 
        \yHat[12][9] , \yHat[12][8] , \yHat[12][7] , \yHat[12][6] , 
        \yHat[12][5] , \yHat[12][4] , \yHat[12][3] , \yHat[12][2] , 
        \yHat[12][1] , \yHat[12][0] , \yHat[11][19] , \yHat[11][18] , 
        \yHat[11][17] , \yHat[11][16] , \yHat[11][15] , \yHat[11][14] , 
        \yHat[11][13] , \yHat[11][12] , \yHat[11][11] , \yHat[11][10] , 
        \yHat[11][9] , \yHat[11][8] , \yHat[11][7] , \yHat[11][6] , 
        \yHat[11][5] , \yHat[11][4] , \yHat[11][3] , \yHat[11][2] , 
        \yHat[11][1] , \yHat[11][0] , \yHat[10][19] , \yHat[10][18] , 
        \yHat[10][17] , \yHat[10][16] , \yHat[10][15] , \yHat[10][14] , 
        \yHat[10][13] , \yHat[10][12] , \yHat[10][11] , \yHat[10][10] , 
        \yHat[10][9] , \yHat[10][8] , \yHat[10][7] , \yHat[10][6] , 
        \yHat[10][5] , \yHat[10][4] , \yHat[10][3] , \yHat[10][2] , 
        \yHat[10][1] , \yHat[10][0] , \yHat[9][19] , \yHat[9][18] , 
        \yHat[9][17] , \yHat[9][16] , \yHat[9][15] , \yHat[9][14] , 
        \yHat[9][13] , \yHat[9][12] , \yHat[9][11] , \yHat[9][10] , 
        \yHat[9][9] , \yHat[9][8] , \yHat[9][7] , \yHat[9][6] , \yHat[9][5] , 
        \yHat[9][4] , \yHat[9][3] , \yHat[9][2] , \yHat[9][1] , \yHat[9][0] , 
        \yHat[8][19] , \yHat[8][18] , \yHat[8][17] , \yHat[8][16] , 
        \yHat[8][15] , \yHat[8][14] , \yHat[8][13] , \yHat[8][12] , 
        \yHat[8][11] , \yHat[8][10] , \yHat[8][9] , \yHat[8][8] , \yHat[8][7] , 
        \yHat[8][6] , \yHat[8][5] , \yHat[8][4] , \yHat[8][3] , \yHat[8][2] , 
        \yHat[8][1] , \yHat[8][0] , \yHat[7][19] , \yHat[7][18] , 
        \yHat[7][17] , \yHat[7][16] , \yHat[7][15] , \yHat[7][14] , 
        \yHat[7][13] , \yHat[7][12] , \yHat[7][11] , \yHat[7][10] , 
        \yHat[7][9] , \yHat[7][8] , \yHat[7][7] , \yHat[7][6] , \yHat[7][5] , 
        \yHat[7][4] , \yHat[7][3] , \yHat[7][2] , \yHat[7][1] , \yHat[7][0] , 
        \yHat[6][19] , \yHat[6][18] , \yHat[6][17] , \yHat[6][16] , 
        \yHat[6][15] , \yHat[6][14] , \yHat[6][13] , \yHat[6][12] , 
        \yHat[6][11] , \yHat[6][10] , \yHat[6][9] , \yHat[6][8] , \yHat[6][7] , 
        \yHat[6][6] , \yHat[6][5] , \yHat[6][4] , \yHat[6][3] , \yHat[6][2] , 
        \yHat[6][1] , \yHat[6][0] , \yHat[5][19] , \yHat[5][18] , 
        \yHat[5][17] , \yHat[5][16] , \yHat[5][15] , \yHat[5][14] , 
        \yHat[5][13] , \yHat[5][12] , \yHat[5][11] , \yHat[5][10] , 
        \yHat[5][9] , \yHat[5][8] , \yHat[5][7] , \yHat[5][6] , \yHat[5][5] , 
        \yHat[5][4] , \yHat[5][3] , \yHat[5][2] , \yHat[5][1] , \yHat[5][0] , 
        \yHat[4][19] , \yHat[4][18] , \yHat[4][17] , \yHat[4][16] , 
        \yHat[4][15] , \yHat[4][14] , \yHat[4][13] , \yHat[4][12] , 
        \yHat[4][11] , \yHat[4][10] , \yHat[4][9] , \yHat[4][8] , \yHat[4][7] , 
        \yHat[4][6] , \yHat[4][5] , \yHat[4][4] , \yHat[4][3] , \yHat[4][2] , 
        \yHat[4][1] , \yHat[4][0] , \yHat[3][19] , \yHat[3][18] , 
        \yHat[3][17] , \yHat[3][16] , \yHat[3][15] , \yHat[3][14] , 
        \yHat[3][13] , \yHat[3][12] , \yHat[3][11] , \yHat[3][10] , 
        \yHat[3][9] , \yHat[3][8] , \yHat[3][7] , \yHat[3][6] , \yHat[3][5] , 
        \yHat[3][4] , \yHat[3][3] , \yHat[3][2] , \yHat[3][1] , \yHat[3][0] , 
        \yHat[2][19] , \yHat[2][18] , \yHat[2][17] , \yHat[2][16] , 
        \yHat[2][15] , \yHat[2][14] , \yHat[2][13] , \yHat[2][12] , 
        \yHat[2][11] , \yHat[2][10] , \yHat[2][9] , \yHat[2][8] , \yHat[2][7] , 
        \yHat[2][6] , \yHat[2][5] , \yHat[2][4] , \yHat[2][3] , \yHat[2][2] , 
        \yHat[2][1] , \yHat[2][0] , \yHat[1][19] , \yHat[1][18] , 
        \yHat[1][17] , \yHat[1][16] , \yHat[1][15] , \yHat[1][14] , 
        \yHat[1][13] , \yHat[1][12] , \yHat[1][11] , \yHat[1][10] , 
        \yHat[1][9] , \yHat[1][8] , \yHat[1][7] , \yHat[1][6] , \yHat[1][5] , 
        \yHat[1][4] , \yHat[1][3] , \yHat[1][2] , \yHat[1][1] , \yHat[1][0] , 
        \yHat[0][19] , \yHat[0][18] , \yHat[0][17] , \yHat[0][16] , 
        \yHat[0][15] , \yHat[0][14] , \yHat[0][13] , \yHat[0][12] , 
        \yHat[0][11] , \yHat[0][10] , \yHat[0][9] , \yHat[0][8] , \yHat[0][7] , 
        \yHat[0][6] , \yHat[0][5] , \yHat[0][4] , \yHat[0][3] , \yHat[0][2] , 
        \yHat[0][1] , \yHat[0][0] }), .y({\y[15][19] , \y[15][18] , 
        \y[15][17] , \y[15][16] , \y[15][15] , \y[15][14] , \y[15][13] , 
        \y[15][12] , \y[15][11] , \y[15][10] , \y[15][9] , \y[15][8] , 
        \y[15][7] , \y[15][6] , \y[15][5] , \y[15][4] , \y[15][3] , \y[15][2] , 
        \y[15][1] , \y[15][0] , \y[14][19] , \y[14][18] , \y[14][17] , 
        \y[14][16] , \y[14][15] , \y[14][14] , \y[14][13] , \y[14][12] , 
        \y[14][11] , \y[14][10] , \y[14][9] , \y[14][8] , \y[14][7] , 
        \y[14][6] , \y[14][5] , \y[14][4] , \y[14][3] , \y[14][2] , \y[14][1] , 
        \y[14][0] , \y[13][19] , \y[13][18] , \y[13][17] , \y[13][16] , 
        \y[13][15] , \y[13][14] , \y[13][13] , \y[13][12] , \y[13][11] , 
        \y[13][10] , \y[13][9] , \y[13][8] , \y[13][7] , \y[13][6] , 
        \y[13][5] , \y[13][4] , \y[13][3] , \y[13][2] , \y[13][1] , \y[13][0] , 
        \y[12][19] , \y[12][18] , \y[12][17] , \y[12][16] , \y[12][15] , 
        \y[12][14] , \y[12][13] , \y[12][12] , \y[12][11] , \y[12][10] , 
        \y[12][9] , \y[12][8] , \y[12][7] , \y[12][6] , \y[12][5] , \y[12][4] , 
        \y[12][3] , \y[12][2] , \y[12][1] , \y[12][0] , \y[11][19] , 
        \y[11][18] , \y[11][17] , \y[11][16] , \y[11][15] , \y[11][14] , 
        \y[11][13] , \y[11][12] , \y[11][11] , \y[11][10] , \y[11][9] , 
        \y[11][8] , \y[11][7] , \y[11][6] , \y[11][5] , \y[11][4] , \y[11][3] , 
        \y[11][2] , \y[11][1] , \y[11][0] , \y[10][19] , \y[10][18] , 
        \y[10][17] , \y[10][16] , \y[10][15] , \y[10][14] , \y[10][13] , 
        \y[10][12] , \y[10][11] , \y[10][10] , \y[10][9] , \y[10][8] , 
        \y[10][7] , \y[10][6] , \y[10][5] , \y[10][4] , \y[10][3] , \y[10][2] , 
        \y[10][1] , \y[10][0] , \y[9][19] , \y[9][18] , \y[9][17] , \y[9][16] , 
        \y[9][15] , \y[9][14] , \y[9][13] , \y[9][12] , \y[9][11] , \y[9][10] , 
        \y[9][9] , \y[9][8] , \y[9][7] , \y[9][6] , \y[9][5] , \y[9][4] , 
        \y[9][3] , \y[9][2] , \y[9][1] , \y[9][0] , \y[8][19] , \y[8][18] , 
        \y[8][17] , \y[8][16] , \y[8][15] , \y[8][14] , \y[8][13] , \y[8][12] , 
        \y[8][11] , \y[8][10] , \y[8][9] , \y[8][8] , \y[8][7] , \y[8][6] , 
        \y[8][5] , \y[8][4] , \y[8][3] , \y[8][2] , \y[8][1] , \y[8][0] , 
        \y[7][19] , \y[7][18] , \y[7][17] , \y[7][16] , \y[7][15] , \y[7][14] , 
        \y[7][13] , \y[7][12] , \y[7][11] , \y[7][10] , \y[7][9] , \y[7][8] , 
        \y[7][7] , \y[7][6] , \y[7][5] , \y[7][4] , \y[7][3] , \y[7][2] , 
        \y[7][1] , \y[7][0] , \y[6][19] , \y[6][18] , \y[6][17] , \y[6][16] , 
        \y[6][15] , \y[6][14] , \y[6][13] , \y[6][12] , \y[6][11] , \y[6][10] , 
        \y[6][9] , \y[6][8] , \y[6][7] , \y[6][6] , \y[6][5] , \y[6][4] , 
        \y[6][3] , \y[6][2] , \y[6][1] , \y[6][0] , \y[5][19] , \y[5][18] , 
        \y[5][17] , \y[5][16] , \y[5][15] , \y[5][14] , \y[5][13] , \y[5][12] , 
        \y[5][11] , \y[5][10] , \y[5][9] , \y[5][8] , \y[5][7] , \y[5][6] , 
        \y[5][5] , \y[5][4] , \y[5][3] , \y[5][2] , \y[5][1] , \y[5][0] , 
        \y[4][19] , \y[4][18] , \y[4][17] , \y[4][16] , \y[4][15] , \y[4][14] , 
        \y[4][13] , \y[4][12] , \y[4][11] , \y[4][10] , \y[4][9] , \y[4][8] , 
        \y[4][7] , \y[4][6] , \y[4][5] , \y[4][4] , \y[4][3] , \y[4][2] , 
        \y[4][1] , \y[4][0] , \y[3][19] , \y[3][18] , \y[3][17] , \y[3][16] , 
        \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] , \y[3][10] , 
        \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] , \y[3][4] , 
        \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] , \y[2][19] , \y[2][18] , 
        \y[2][17] , \y[2][16] , \y[2][15] , \y[2][14] , \y[2][13] , \y[2][12] , 
        \y[2][11] , \y[2][10] , \y[2][9] , \y[2][8] , \y[2][7] , \y[2][6] , 
        \y[2][5] , \y[2][4] , \y[2][3] , \y[2][2] , \y[2][1] , \y[2][0] , 
        \y[1][19] , \y[1][18] , \y[1][17] , \y[1][16] , \y[1][15] , \y[1][14] , 
        \y[1][13] , \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] , \y[1][8] , 
        \y[1][7] , \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] , \y[1][2] , 
        \y[1][1] , \y[1][0] , \y[0][19] , \y[0][18] , \y[0][17] , \y[0][16] , 
        \y[0][15] , \y[0][14] , \y[0][13] , \y[0][12] , \y[0][11] , \y[0][10] , 
        \y[0][9] , \y[0][8] , \y[0][7] , \y[0][6] , \y[0][5] , \y[0][4] , 
        \y[0][3] , \y[0][2] , \y[0][1] , \y[0][0] }), num, input_ready, 
        output_taken, state, out );
  input [3:0] num;
  output [1:0] state;
  output [19:0] out;
  input clk, reset, model, \yHat[15][19] , \yHat[15][18] , \yHat[15][17] ,
         \yHat[15][16] , \yHat[15][15] , \yHat[15][14] , \yHat[15][13] ,
         \yHat[15][12] , \yHat[15][11] , \yHat[15][10] , \yHat[15][9] ,
         \yHat[15][8] , \yHat[15][7] , \yHat[15][6] , \yHat[15][5] ,
         \yHat[15][4] , \yHat[15][3] , \yHat[15][2] , \yHat[15][1] ,
         \yHat[15][0] , \yHat[14][19] , \yHat[14][18] , \yHat[14][17] ,
         \yHat[14][16] , \yHat[14][15] , \yHat[14][14] , \yHat[14][13] ,
         \yHat[14][12] , \yHat[14][11] , \yHat[14][10] , \yHat[14][9] ,
         \yHat[14][8] , \yHat[14][7] , \yHat[14][6] , \yHat[14][5] ,
         \yHat[14][4] , \yHat[14][3] , \yHat[14][2] , \yHat[14][1] ,
         \yHat[14][0] , \yHat[13][19] , \yHat[13][18] , \yHat[13][17] ,
         \yHat[13][16] , \yHat[13][15] , \yHat[13][14] , \yHat[13][13] ,
         \yHat[13][12] , \yHat[13][11] , \yHat[13][10] , \yHat[13][9] ,
         \yHat[13][8] , \yHat[13][7] , \yHat[13][6] , \yHat[13][5] ,
         \yHat[13][4] , \yHat[13][3] , \yHat[13][2] , \yHat[13][1] ,
         \yHat[13][0] , \yHat[12][19] , \yHat[12][18] , \yHat[12][17] ,
         \yHat[12][16] , \yHat[12][15] , \yHat[12][14] , \yHat[12][13] ,
         \yHat[12][12] , \yHat[12][11] , \yHat[12][10] , \yHat[12][9] ,
         \yHat[12][8] , \yHat[12][7] , \yHat[12][6] , \yHat[12][5] ,
         \yHat[12][4] , \yHat[12][3] , \yHat[12][2] , \yHat[12][1] ,
         \yHat[12][0] , \yHat[11][19] , \yHat[11][18] , \yHat[11][17] ,
         \yHat[11][16] , \yHat[11][15] , \yHat[11][14] , \yHat[11][13] ,
         \yHat[11][12] , \yHat[11][11] , \yHat[11][10] , \yHat[11][9] ,
         \yHat[11][8] , \yHat[11][7] , \yHat[11][6] , \yHat[11][5] ,
         \yHat[11][4] , \yHat[11][3] , \yHat[11][2] , \yHat[11][1] ,
         \yHat[11][0] , \yHat[10][19] , \yHat[10][18] , \yHat[10][17] ,
         \yHat[10][16] , \yHat[10][15] , \yHat[10][14] , \yHat[10][13] ,
         \yHat[10][12] , \yHat[10][11] , \yHat[10][10] , \yHat[10][9] ,
         \yHat[10][8] , \yHat[10][7] , \yHat[10][6] , \yHat[10][5] ,
         \yHat[10][4] , \yHat[10][3] , \yHat[10][2] , \yHat[10][1] ,
         \yHat[10][0] , \yHat[9][19] , \yHat[9][18] , \yHat[9][17] ,
         \yHat[9][16] , \yHat[9][15] , \yHat[9][14] , \yHat[9][13] ,
         \yHat[9][12] , \yHat[9][11] , \yHat[9][10] , \yHat[9][9] ,
         \yHat[9][8] , \yHat[9][7] , \yHat[9][6] , \yHat[9][5] , \yHat[9][4] ,
         \yHat[9][3] , \yHat[9][2] , \yHat[9][1] , \yHat[9][0] , \yHat[8][19] ,
         \yHat[8][18] , \yHat[8][17] , \yHat[8][16] , \yHat[8][15] ,
         \yHat[8][14] , \yHat[8][13] , \yHat[8][12] , \yHat[8][11] ,
         \yHat[8][10] , \yHat[8][9] , \yHat[8][8] , \yHat[8][7] , \yHat[8][6] ,
         \yHat[8][5] , \yHat[8][4] , \yHat[8][3] , \yHat[8][2] , \yHat[8][1] ,
         \yHat[8][0] , \yHat[7][19] , \yHat[7][18] , \yHat[7][17] ,
         \yHat[7][16] , \yHat[7][15] , \yHat[7][14] , \yHat[7][13] ,
         \yHat[7][12] , \yHat[7][11] , \yHat[7][10] , \yHat[7][9] ,
         \yHat[7][8] , \yHat[7][7] , \yHat[7][6] , \yHat[7][5] , \yHat[7][4] ,
         \yHat[7][3] , \yHat[7][2] , \yHat[7][1] , \yHat[7][0] , \yHat[6][19] ,
         \yHat[6][18] , \yHat[6][17] , \yHat[6][16] , \yHat[6][15] ,
         \yHat[6][14] , \yHat[6][13] , \yHat[6][12] , \yHat[6][11] ,
         \yHat[6][10] , \yHat[6][9] , \yHat[6][8] , \yHat[6][7] , \yHat[6][6] ,
         \yHat[6][5] , \yHat[6][4] , \yHat[6][3] , \yHat[6][2] , \yHat[6][1] ,
         \yHat[6][0] , \yHat[5][19] , \yHat[5][18] , \yHat[5][17] ,
         \yHat[5][16] , \yHat[5][15] , \yHat[5][14] , \yHat[5][13] ,
         \yHat[5][12] , \yHat[5][11] , \yHat[5][10] , \yHat[5][9] ,
         \yHat[5][8] , \yHat[5][7] , \yHat[5][6] , \yHat[5][5] , \yHat[5][4] ,
         \yHat[5][3] , \yHat[5][2] , \yHat[5][1] , \yHat[5][0] , \yHat[4][19] ,
         \yHat[4][18] , \yHat[4][17] , \yHat[4][16] , \yHat[4][15] ,
         \yHat[4][14] , \yHat[4][13] , \yHat[4][12] , \yHat[4][11] ,
         \yHat[4][10] , \yHat[4][9] , \yHat[4][8] , \yHat[4][7] , \yHat[4][6] ,
         \yHat[4][5] , \yHat[4][4] , \yHat[4][3] , \yHat[4][2] , \yHat[4][1] ,
         \yHat[4][0] , \yHat[3][19] , \yHat[3][18] , \yHat[3][17] ,
         \yHat[3][16] , \yHat[3][15] , \yHat[3][14] , \yHat[3][13] ,
         \yHat[3][12] , \yHat[3][11] , \yHat[3][10] , \yHat[3][9] ,
         \yHat[3][8] , \yHat[3][7] , \yHat[3][6] , \yHat[3][5] , \yHat[3][4] ,
         \yHat[3][3] , \yHat[3][2] , \yHat[3][1] , \yHat[3][0] , \yHat[2][19] ,
         \yHat[2][18] , \yHat[2][17] , \yHat[2][16] , \yHat[2][15] ,
         \yHat[2][14] , \yHat[2][13] , \yHat[2][12] , \yHat[2][11] ,
         \yHat[2][10] , \yHat[2][9] , \yHat[2][8] , \yHat[2][7] , \yHat[2][6] ,
         \yHat[2][5] , \yHat[2][4] , \yHat[2][3] , \yHat[2][2] , \yHat[2][1] ,
         \yHat[2][0] , \yHat[1][19] , \yHat[1][18] , \yHat[1][17] ,
         \yHat[1][16] , \yHat[1][15] , \yHat[1][14] , \yHat[1][13] ,
         \yHat[1][12] , \yHat[1][11] , \yHat[1][10] , \yHat[1][9] ,
         \yHat[1][8] , \yHat[1][7] , \yHat[1][6] , \yHat[1][5] , \yHat[1][4] ,
         \yHat[1][3] , \yHat[1][2] , \yHat[1][1] , \yHat[1][0] , \yHat[0][19] ,
         \yHat[0][18] , \yHat[0][17] , \yHat[0][16] , \yHat[0][15] ,
         \yHat[0][14] , \yHat[0][13] , \yHat[0][12] , \yHat[0][11] ,
         \yHat[0][10] , \yHat[0][9] , \yHat[0][8] , \yHat[0][7] , \yHat[0][6] ,
         \yHat[0][5] , \yHat[0][4] , \yHat[0][3] , \yHat[0][2] , \yHat[0][1] ,
         \yHat[0][0] , \y[15][19] , \y[15][18] , \y[15][17] , \y[15][16] ,
         \y[15][15] , \y[15][14] , \y[15][13] , \y[15][12] , \y[15][11] ,
         \y[15][10] , \y[15][9] , \y[15][8] , \y[15][7] , \y[15][6] ,
         \y[15][5] , \y[15][4] , \y[15][3] , \y[15][2] , \y[15][1] ,
         \y[15][0] , \y[14][19] , \y[14][18] , \y[14][17] , \y[14][16] ,
         \y[14][15] , \y[14][14] , \y[14][13] , \y[14][12] , \y[14][11] ,
         \y[14][10] , \y[14][9] , \y[14][8] , \y[14][7] , \y[14][6] ,
         \y[14][5] , \y[14][4] , \y[14][3] , \y[14][2] , \y[14][1] ,
         \y[14][0] , \y[13][19] , \y[13][18] , \y[13][17] , \y[13][16] ,
         \y[13][15] , \y[13][14] , \y[13][13] , \y[13][12] , \y[13][11] ,
         \y[13][10] , \y[13][9] , \y[13][8] , \y[13][7] , \y[13][6] ,
         \y[13][5] , \y[13][4] , \y[13][3] , \y[13][2] , \y[13][1] ,
         \y[13][0] , \y[12][19] , \y[12][18] , \y[12][17] , \y[12][16] ,
         \y[12][15] , \y[12][14] , \y[12][13] , \y[12][12] , \y[12][11] ,
         \y[12][10] , \y[12][9] , \y[12][8] , \y[12][7] , \y[12][6] ,
         \y[12][5] , \y[12][4] , \y[12][3] , \y[12][2] , \y[12][1] ,
         \y[12][0] , \y[11][19] , \y[11][18] , \y[11][17] , \y[11][16] ,
         \y[11][15] , \y[11][14] , \y[11][13] , \y[11][12] , \y[11][11] ,
         \y[11][10] , \y[11][9] , \y[11][8] , \y[11][7] , \y[11][6] ,
         \y[11][5] , \y[11][4] , \y[11][3] , \y[11][2] , \y[11][1] ,
         \y[11][0] , \y[10][19] , \y[10][18] , \y[10][17] , \y[10][16] ,
         \y[10][15] , \y[10][14] , \y[10][13] , \y[10][12] , \y[10][11] ,
         \y[10][10] , \y[10][9] , \y[10][8] , \y[10][7] , \y[10][6] ,
         \y[10][5] , \y[10][4] , \y[10][3] , \y[10][2] , \y[10][1] ,
         \y[10][0] , \y[9][19] , \y[9][18] , \y[9][17] , \y[9][16] ,
         \y[9][15] , \y[9][14] , \y[9][13] , \y[9][12] , \y[9][11] ,
         \y[9][10] , \y[9][9] , \y[9][8] , \y[9][7] , \y[9][6] , \y[9][5] ,
         \y[9][4] , \y[9][3] , \y[9][2] , \y[9][1] , \y[9][0] , \y[8][19] ,
         \y[8][18] , \y[8][17] , \y[8][16] , \y[8][15] , \y[8][14] ,
         \y[8][13] , \y[8][12] , \y[8][11] , \y[8][10] , \y[8][9] , \y[8][8] ,
         \y[8][7] , \y[8][6] , \y[8][5] , \y[8][4] , \y[8][3] , \y[8][2] ,
         \y[8][1] , \y[8][0] , \y[7][19] , \y[7][18] , \y[7][17] , \y[7][16] ,
         \y[7][15] , \y[7][14] , \y[7][13] , \y[7][12] , \y[7][11] ,
         \y[7][10] , \y[7][9] , \y[7][8] , \y[7][7] , \y[7][6] , \y[7][5] ,
         \y[7][4] , \y[7][3] , \y[7][2] , \y[7][1] , \y[7][0] , \y[6][19] ,
         \y[6][18] , \y[6][17] , \y[6][16] , \y[6][15] , \y[6][14] ,
         \y[6][13] , \y[6][12] , \y[6][11] , \y[6][10] , \y[6][9] , \y[6][8] ,
         \y[6][7] , \y[6][6] , \y[6][5] , \y[6][4] , \y[6][3] , \y[6][2] ,
         \y[6][1] , \y[6][0] , \y[5][19] , \y[5][18] , \y[5][17] , \y[5][16] ,
         \y[5][15] , \y[5][14] , \y[5][13] , \y[5][12] , \y[5][11] ,
         \y[5][10] , \y[5][9] , \y[5][8] , \y[5][7] , \y[5][6] , \y[5][5] ,
         \y[5][4] , \y[5][3] , \y[5][2] , \y[5][1] , \y[5][0] , \y[4][19] ,
         \y[4][18] , \y[4][17] , \y[4][16] , \y[4][15] , \y[4][14] ,
         \y[4][13] , \y[4][12] , \y[4][11] , \y[4][10] , \y[4][9] , \y[4][8] ,
         \y[4][7] , \y[4][6] , \y[4][5] , \y[4][4] , \y[4][3] , \y[4][2] ,
         \y[4][1] , \y[4][0] , \y[3][19] , \y[3][18] , \y[3][17] , \y[3][16] ,
         \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] ,
         \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] ,
         \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] , \y[2][19] ,
         \y[2][18] , \y[2][17] , \y[2][16] , \y[2][15] , \y[2][14] ,
         \y[2][13] , \y[2][12] , \y[2][11] , \y[2][10] , \y[2][9] , \y[2][8] ,
         \y[2][7] , \y[2][6] , \y[2][5] , \y[2][4] , \y[2][3] , \y[2][2] ,
         \y[2][1] , \y[2][0] , \y[1][19] , \y[1][18] , \y[1][17] , \y[1][16] ,
         \y[1][15] , \y[1][14] , \y[1][13] , \y[1][12] , \y[1][11] ,
         \y[1][10] , \y[1][9] , \y[1][8] , \y[1][7] , \y[1][6] , \y[1][5] ,
         \y[1][4] , \y[1][3] , \y[1][2] , \y[1][1] , \y[1][0] , \y[0][19] ,
         \y[0][18] , \y[0][17] , \y[0][16] , \y[0][15] , \y[0][14] ,
         \y[0][13] , \y[0][12] , \y[0][11] , \y[0][10] , \y[0][9] , \y[0][8] ,
         \y[0][7] , \y[0][6] , \y[0][5] , \y[0][4] , \y[0][3] , \y[0][2] ,
         \y[0][1] , \y[0][0] , input_ready, output_taken;
  wire   done, \reg_yHat[14][19] , \reg_yHat[14][18] , \reg_yHat[14][17] ,
         \reg_yHat[14][16] , \reg_yHat[14][15] , \reg_yHat[14][14] ,
         \reg_yHat[14][13] , \reg_yHat[14][12] , \reg_yHat[14][11] ,
         \reg_yHat[14][10] , \reg_yHat[14][9] , \reg_yHat[14][8] ,
         \reg_yHat[14][7] , \reg_yHat[14][6] , \reg_yHat[14][5] ,
         \reg_yHat[14][4] , \reg_yHat[14][3] , \reg_yHat[14][2] ,
         \reg_yHat[14][1] , \reg_yHat[14][0] , \reg_yHat[13][19] ,
         \reg_yHat[13][18] , \reg_yHat[13][17] , \reg_yHat[13][16] ,
         \reg_yHat[13][15] , \reg_yHat[13][14] , \reg_yHat[13][13] ,
         \reg_yHat[13][12] , \reg_yHat[13][11] , \reg_yHat[13][10] ,
         \reg_yHat[13][9] , \reg_yHat[13][8] , \reg_yHat[13][7] ,
         \reg_yHat[13][6] , \reg_yHat[13][5] , \reg_yHat[13][4] ,
         \reg_yHat[13][3] , \reg_yHat[13][2] , \reg_yHat[13][1] ,
         \reg_yHat[13][0] , \reg_yHat[12][19] , \reg_yHat[12][18] ,
         \reg_yHat[12][17] , \reg_yHat[12][16] , \reg_yHat[12][15] ,
         \reg_yHat[12][14] , \reg_yHat[12][13] , \reg_yHat[12][12] ,
         \reg_yHat[12][11] , \reg_yHat[12][10] , \reg_yHat[12][9] ,
         \reg_yHat[12][8] , \reg_yHat[12][7] , \reg_yHat[12][6] ,
         \reg_yHat[12][5] , \reg_yHat[12][4] , \reg_yHat[12][3] ,
         \reg_yHat[12][2] , \reg_yHat[12][1] , \reg_yHat[12][0] ,
         \reg_yHat[11][19] , \reg_yHat[11][18] , \reg_yHat[11][17] ,
         \reg_yHat[11][16] , \reg_yHat[11][15] , \reg_yHat[11][14] ,
         \reg_yHat[11][13] , \reg_yHat[11][12] , \reg_yHat[11][11] ,
         \reg_yHat[11][10] , \reg_yHat[11][9] , \reg_yHat[11][8] ,
         \reg_yHat[11][7] , \reg_yHat[11][6] , \reg_yHat[11][5] ,
         \reg_yHat[11][4] , \reg_yHat[11][3] , \reg_yHat[11][2] ,
         \reg_yHat[11][1] , \reg_yHat[11][0] , \reg_yHat[10][19] ,
         \reg_yHat[10][18] , \reg_yHat[10][17] , \reg_yHat[10][16] ,
         \reg_yHat[10][15] , \reg_yHat[10][14] , \reg_yHat[10][13] ,
         \reg_yHat[10][12] , \reg_yHat[10][11] , \reg_yHat[10][10] ,
         \reg_yHat[10][9] , \reg_yHat[10][8] , \reg_yHat[10][7] ,
         \reg_yHat[10][6] , \reg_yHat[10][5] , \reg_yHat[10][4] ,
         \reg_yHat[10][3] , \reg_yHat[10][2] , \reg_yHat[10][1] ,
         \reg_yHat[10][0] , \reg_yHat[9][19] , \reg_yHat[9][18] ,
         \reg_yHat[9][17] , \reg_yHat[9][16] , \reg_yHat[9][15] ,
         \reg_yHat[9][14] , \reg_yHat[9][13] , \reg_yHat[9][12] ,
         \reg_yHat[9][11] , \reg_yHat[9][10] , \reg_yHat[9][9] ,
         \reg_yHat[9][8] , \reg_yHat[9][7] , \reg_yHat[9][6] ,
         \reg_yHat[9][5] , \reg_yHat[9][4] , \reg_yHat[9][3] ,
         \reg_yHat[9][2] , \reg_yHat[9][1] , \reg_yHat[9][0] ,
         \reg_yHat[8][19] , \reg_yHat[8][18] , \reg_yHat[8][17] ,
         \reg_yHat[8][16] , \reg_yHat[8][15] , \reg_yHat[8][14] ,
         \reg_yHat[8][13] , \reg_yHat[8][12] , \reg_yHat[8][11] ,
         \reg_yHat[8][10] , \reg_yHat[8][9] , \reg_yHat[8][8] ,
         \reg_yHat[8][7] , \reg_yHat[8][6] , \reg_yHat[8][5] ,
         \reg_yHat[8][4] , \reg_yHat[8][3] , \reg_yHat[8][2] ,
         \reg_yHat[8][1] , \reg_yHat[8][0] , \reg_yHat[7][19] ,
         \reg_yHat[7][18] , \reg_yHat[7][17] , \reg_yHat[7][16] ,
         \reg_yHat[7][15] , \reg_yHat[7][14] , \reg_yHat[7][13] ,
         \reg_yHat[7][12] , \reg_yHat[7][11] , \reg_yHat[7][10] ,
         \reg_yHat[7][9] , \reg_yHat[7][8] , \reg_yHat[7][7] ,
         \reg_yHat[7][6] , \reg_yHat[7][5] , \reg_yHat[7][4] ,
         \reg_yHat[7][3] , \reg_yHat[7][2] , \reg_yHat[7][1] ,
         \reg_yHat[7][0] , \reg_yHat[6][19] , \reg_yHat[6][18] ,
         \reg_yHat[6][17] , \reg_yHat[6][16] , \reg_yHat[6][15] ,
         \reg_yHat[6][14] , \reg_yHat[6][13] , \reg_yHat[6][12] ,
         \reg_yHat[6][11] , \reg_yHat[6][10] , \reg_yHat[6][9] ,
         \reg_yHat[6][8] , \reg_yHat[6][7] , \reg_yHat[6][6] ,
         \reg_yHat[6][5] , \reg_yHat[6][4] , \reg_yHat[6][3] ,
         \reg_yHat[6][2] , \reg_yHat[6][1] , \reg_yHat[6][0] ,
         \reg_yHat[5][19] , \reg_yHat[5][18] , \reg_yHat[5][17] ,
         \reg_yHat[5][16] , \reg_yHat[5][15] , \reg_yHat[5][14] ,
         \reg_yHat[5][13] , \reg_yHat[5][12] , \reg_yHat[5][11] ,
         \reg_yHat[5][10] , \reg_yHat[5][9] , \reg_yHat[5][8] ,
         \reg_yHat[5][7] , \reg_yHat[5][6] , \reg_yHat[5][5] ,
         \reg_yHat[5][4] , \reg_yHat[5][3] , \reg_yHat[5][2] ,
         \reg_yHat[5][1] , \reg_yHat[5][0] , \reg_yHat[4][19] ,
         \reg_yHat[4][18] , \reg_yHat[4][17] , \reg_yHat[4][16] ,
         \reg_yHat[4][15] , \reg_yHat[4][14] , \reg_yHat[4][13] ,
         \reg_yHat[4][12] , \reg_yHat[4][11] , \reg_yHat[4][10] ,
         \reg_yHat[4][9] , \reg_yHat[4][8] , \reg_yHat[4][7] ,
         \reg_yHat[4][6] , \reg_yHat[4][5] , \reg_yHat[4][4] ,
         \reg_yHat[4][3] , \reg_yHat[4][2] , \reg_yHat[4][1] ,
         \reg_yHat[4][0] , \reg_yHat[3][19] , \reg_yHat[3][18] ,
         \reg_yHat[3][17] , \reg_yHat[3][16] , \reg_yHat[3][15] ,
         \reg_yHat[3][14] , \reg_yHat[3][13] , \reg_yHat[3][12] ,
         \reg_yHat[3][11] , \reg_yHat[3][10] , \reg_yHat[3][9] ,
         \reg_yHat[3][8] , \reg_yHat[3][7] , \reg_yHat[3][6] ,
         \reg_yHat[3][5] , \reg_yHat[3][4] , \reg_yHat[3][3] ,
         \reg_yHat[3][2] , \reg_yHat[3][1] , \reg_yHat[3][0] ,
         \reg_yHat[2][19] , \reg_yHat[2][18] , \reg_yHat[2][17] ,
         \reg_yHat[2][16] , \reg_yHat[2][15] , \reg_yHat[2][14] ,
         \reg_yHat[2][13] , \reg_yHat[2][12] , \reg_yHat[2][11] ,
         \reg_yHat[2][10] , \reg_yHat[2][9] , \reg_yHat[2][8] ,
         \reg_yHat[2][7] , \reg_yHat[2][6] , \reg_yHat[2][5] ,
         \reg_yHat[2][4] , \reg_yHat[2][3] , \reg_yHat[2][2] ,
         \reg_yHat[2][1] , \reg_yHat[2][0] , \reg_yHat[1][19] ,
         \reg_yHat[1][18] , \reg_yHat[1][17] , \reg_yHat[1][16] ,
         \reg_yHat[1][15] , \reg_yHat[1][14] , \reg_yHat[1][13] ,
         \reg_yHat[1][12] , \reg_yHat[1][11] , \reg_yHat[1][10] ,
         \reg_yHat[1][9] , \reg_yHat[1][8] , \reg_yHat[1][7] ,
         \reg_yHat[1][6] , \reg_yHat[1][5] , \reg_yHat[1][4] ,
         \reg_yHat[1][3] , \reg_yHat[1][2] , \reg_yHat[1][1] ,
         \reg_yHat[1][0] , \reg_yHat[0][19] , \reg_yHat[0][18] ,
         \reg_yHat[0][17] , \reg_yHat[0][16] , \reg_yHat[0][15] ,
         \reg_yHat[0][14] , \reg_yHat[0][13] , \reg_yHat[0][12] ,
         \reg_yHat[0][11] , \reg_yHat[0][10] , \reg_yHat[0][9] ,
         \reg_yHat[0][8] , \reg_yHat[0][7] , \reg_yHat[0][6] ,
         \reg_yHat[0][5] , \reg_yHat[0][4] , \reg_yHat[0][3] ,
         \reg_yHat[0][2] , \reg_yHat[0][1] , \reg_yHat[0][0] , \reg_y[14][19] ,
         \reg_y[14][18] , \reg_y[14][17] , \reg_y[14][16] , \reg_y[14][15] ,
         \reg_y[14][14] , \reg_y[14][13] , \reg_y[14][12] , \reg_y[14][11] ,
         \reg_y[14][10] , \reg_y[14][9] , \reg_y[14][8] , \reg_y[14][7] ,
         \reg_y[14][6] , \reg_y[14][5] , \reg_y[14][4] , \reg_y[14][3] ,
         \reg_y[14][2] , \reg_y[14][1] , \reg_y[14][0] , \reg_y[13][19] ,
         \reg_y[13][18] , \reg_y[13][17] , \reg_y[13][16] , \reg_y[13][15] ,
         \reg_y[13][14] , \reg_y[13][13] , \reg_y[13][12] , \reg_y[13][11] ,
         \reg_y[13][10] , \reg_y[13][9] , \reg_y[13][8] , \reg_y[13][7] ,
         \reg_y[13][6] , \reg_y[13][5] , \reg_y[13][4] , \reg_y[13][3] ,
         \reg_y[13][2] , \reg_y[13][1] , \reg_y[13][0] , \reg_y[12][19] ,
         \reg_y[12][18] , \reg_y[12][17] , \reg_y[12][16] , \reg_y[12][15] ,
         \reg_y[12][14] , \reg_y[12][13] , \reg_y[12][12] , \reg_y[12][11] ,
         \reg_y[12][10] , \reg_y[12][9] , \reg_y[12][8] , \reg_y[12][7] ,
         \reg_y[12][6] , \reg_y[12][5] , \reg_y[12][4] , \reg_y[12][3] ,
         \reg_y[12][2] , \reg_y[12][1] , \reg_y[12][0] , \reg_y[11][19] ,
         \reg_y[11][18] , \reg_y[11][17] , \reg_y[11][16] , \reg_y[11][15] ,
         \reg_y[11][14] , \reg_y[11][13] , \reg_y[11][12] , \reg_y[11][11] ,
         \reg_y[11][10] , \reg_y[11][9] , \reg_y[11][8] , \reg_y[11][7] ,
         \reg_y[11][6] , \reg_y[11][5] , \reg_y[11][4] , \reg_y[11][3] ,
         \reg_y[11][2] , \reg_y[11][1] , \reg_y[11][0] , \reg_y[10][19] ,
         \reg_y[10][18] , \reg_y[10][17] , \reg_y[10][16] , \reg_y[10][15] ,
         \reg_y[10][14] , \reg_y[10][13] , \reg_y[10][12] , \reg_y[10][11] ,
         \reg_y[10][10] , \reg_y[10][9] , \reg_y[10][8] , \reg_y[10][7] ,
         \reg_y[10][6] , \reg_y[10][5] , \reg_y[10][4] , \reg_y[10][3] ,
         \reg_y[10][2] , \reg_y[10][1] , \reg_y[10][0] , \reg_y[9][19] ,
         \reg_y[9][18] , \reg_y[9][17] , \reg_y[9][16] , \reg_y[9][15] ,
         \reg_y[9][14] , \reg_y[9][13] , \reg_y[9][12] , \reg_y[9][11] ,
         \reg_y[9][10] , \reg_y[9][9] , \reg_y[9][8] , \reg_y[9][7] ,
         \reg_y[9][6] , \reg_y[9][5] , \reg_y[9][4] , \reg_y[9][3] ,
         \reg_y[9][2] , \reg_y[9][1] , \reg_y[9][0] , \reg_y[8][19] ,
         \reg_y[8][18] , \reg_y[8][17] , \reg_y[8][16] , \reg_y[8][15] ,
         \reg_y[8][14] , \reg_y[8][13] , \reg_y[8][12] , \reg_y[8][11] ,
         \reg_y[8][10] , \reg_y[8][9] , \reg_y[8][8] , \reg_y[8][7] ,
         \reg_y[8][6] , \reg_y[8][5] , \reg_y[8][4] , \reg_y[8][3] ,
         \reg_y[8][2] , \reg_y[8][1] , \reg_y[8][0] , \reg_y[7][19] ,
         \reg_y[7][18] , \reg_y[7][17] , \reg_y[7][16] , \reg_y[7][15] ,
         \reg_y[7][14] , \reg_y[7][13] , \reg_y[7][12] , \reg_y[7][11] ,
         \reg_y[7][10] , \reg_y[7][9] , \reg_y[7][8] , \reg_y[7][7] ,
         \reg_y[7][6] , \reg_y[7][5] , \reg_y[7][4] , \reg_y[7][3] ,
         \reg_y[7][2] , \reg_y[7][1] , \reg_y[7][0] , \reg_y[6][19] ,
         \reg_y[6][18] , \reg_y[6][17] , \reg_y[6][16] , \reg_y[6][15] ,
         \reg_y[6][14] , \reg_y[6][13] , \reg_y[6][12] , \reg_y[6][11] ,
         \reg_y[6][10] , \reg_y[6][9] , \reg_y[6][8] , \reg_y[6][7] ,
         \reg_y[6][6] , \reg_y[6][5] , \reg_y[6][4] , \reg_y[6][3] ,
         \reg_y[6][2] , \reg_y[6][1] , \reg_y[6][0] , \reg_y[5][19] ,
         \reg_y[5][18] , \reg_y[5][17] , \reg_y[5][16] , \reg_y[5][15] ,
         \reg_y[5][14] , \reg_y[5][13] , \reg_y[5][12] , \reg_y[5][11] ,
         \reg_y[5][10] , \reg_y[5][9] , \reg_y[5][8] , \reg_y[5][7] ,
         \reg_y[5][6] , \reg_y[5][5] , \reg_y[5][4] , \reg_y[5][3] ,
         \reg_y[5][2] , \reg_y[5][1] , \reg_y[5][0] , \reg_y[4][19] ,
         \reg_y[4][18] , \reg_y[4][17] , \reg_y[4][16] , \reg_y[4][15] ,
         \reg_y[4][14] , \reg_y[4][13] , \reg_y[4][12] , \reg_y[4][11] ,
         \reg_y[4][10] , \reg_y[4][9] , \reg_y[4][8] , \reg_y[4][7] ,
         \reg_y[4][6] , \reg_y[4][5] , \reg_y[4][4] , \reg_y[4][3] ,
         \reg_y[4][2] , \reg_y[4][1] , \reg_y[4][0] , \reg_y[3][19] ,
         \reg_y[3][18] , \reg_y[3][17] , \reg_y[3][16] , \reg_y[3][15] ,
         \reg_y[3][14] , \reg_y[3][13] , \reg_y[3][12] , \reg_y[3][11] ,
         \reg_y[3][10] , \reg_y[3][9] , \reg_y[3][8] , \reg_y[3][7] ,
         \reg_y[3][6] , \reg_y[3][5] , \reg_y[3][4] , \reg_y[3][3] ,
         \reg_y[3][2] , \reg_y[3][1] , \reg_y[3][0] , \reg_y[2][19] ,
         \reg_y[2][18] , \reg_y[2][17] , \reg_y[2][16] , \reg_y[2][15] ,
         \reg_y[2][14] , \reg_y[2][13] , \reg_y[2][12] , \reg_y[2][11] ,
         \reg_y[2][10] , \reg_y[2][9] , \reg_y[2][8] , \reg_y[2][7] ,
         \reg_y[2][6] , \reg_y[2][5] , \reg_y[2][4] , \reg_y[2][3] ,
         \reg_y[2][2] , \reg_y[2][1] , \reg_y[2][0] , \reg_y[1][19] ,
         \reg_y[1][18] , \reg_y[1][17] , \reg_y[1][16] , \reg_y[1][15] ,
         \reg_y[1][14] , \reg_y[1][13] , \reg_y[1][12] , \reg_y[1][11] ,
         \reg_y[1][10] , \reg_y[1][9] , \reg_y[1][8] , \reg_y[1][7] ,
         \reg_y[1][6] , \reg_y[1][5] , \reg_y[1][4] , \reg_y[1][3] ,
         \reg_y[1][2] , \reg_y[1][1] , \reg_y[1][0] , \reg_y[0][19] ,
         \reg_y[0][18] , \reg_y[0][17] , \reg_y[0][16] , \reg_y[0][15] ,
         \reg_y[0][14] , \reg_y[0][13] , \reg_y[0][12] , \reg_y[0][11] ,
         \reg_y[0][10] , \reg_y[0][9] , \reg_y[0][8] , \reg_y[0][7] ,
         \reg_y[0][6] , \reg_y[0][5] , \reg_y[0][4] , \reg_y[0][3] ,
         \reg_y[0][2] , \reg_y[0][1] , \reg_y[0][0] , reg_model, n1358, n1359,
         n1360, n1361, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n55799, n55798, n39253, n39254, n39255, n39256,
         n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
         n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272,
         n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280,
         n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288,
         n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
         n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
         n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312,
         n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
         n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
         n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336,
         n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
         n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
         n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360,
         n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368,
         n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
         n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384,
         n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
         n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400,
         n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408,
         n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
         n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424,
         n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432,
         n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440,
         n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
         n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456,
         n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
         n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472,
         n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480,
         n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
         n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496,
         n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504,
         n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
         n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
         n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
         n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
         n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
         n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552,
         n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
         n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568,
         n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576,
         n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584,
         n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
         n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600,
         n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
         n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616,
         n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624,
         n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632,
         n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640,
         n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
         n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656,
         n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
         n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672,
         n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
         n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688,
         n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696,
         n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
         n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712,
         n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
         n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728,
         n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
         n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744,
         n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
         n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
         n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
         n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
         n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
         n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
         n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800,
         n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
         n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816,
         n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
         n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832,
         n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840,
         n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848,
         n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856,
         n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
         n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872,
         n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
         n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888,
         n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
         n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904,
         n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
         n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920,
         n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928,
         n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936,
         n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944,
         n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
         n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960,
         n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
         n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
         n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984,
         n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992,
         n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000,
         n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008,
         n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016,
         n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
         n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032,
         n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
         n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
         n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056,
         n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064,
         n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072,
         n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080,
         n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088,
         n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
         n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
         n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
         n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
         n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128,
         n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
         n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144,
         n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152,
         n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
         n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
         n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
         n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
         n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
         n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200,
         n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
         n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216,
         n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
         n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
         n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
         n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248,
         n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
         n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
         n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
         n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
         n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288,
         n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296,
         n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304,
         n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
         n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320,
         n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
         n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
         n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
         n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
         n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360,
         n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368,
         n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376,
         n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
         n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392,
         n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
         n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
         n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
         n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424,
         n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432,
         n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440,
         n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448,
         n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
         n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464,
         n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
         n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480,
         n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488,
         n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496,
         n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504,
         n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512,
         n40513, n40514, n40515, n40516, n40517, n40518, n9999, n9998, n9997,
         n9996, n9995, n9994, n9993, n9992, n9991, n9990, n9989, n9988, n9987,
         n9986, n9985, n9984, n9983, n9982, n9981, n9980, n9979, n9978, n9977,
         n9976, n9975, n9974, n9973, n9972, n9971, n9970, n9969, n9968, n9967,
         n9966, n9965, n9964, n9963, n9962, n9961, n9960, n9959, n9958, n9957,
         n9956, n9955, n9954, n9953, n9952, n9951, n9950, n9949, n9948, n9947,
         n9946, n9945, n9944, n9943, n9942, n9941, n9940, n9939, n9938, n9937,
         n9936, n9935, n9934, n9933, n9932, n9931, n9930, n9929, n9928, n9927,
         n9926, n9925, n9924, n9923, n9922, n9921, n9920, n9919, n9918, n9917,
         n9916, n9915, n9914, n9913, n9912, n9911, n9910, n9909, n9908, n9907,
         n9906, n9905, n9904, n9903, n9902, n9901, n9900, n9899, n9898, n9897,
         n9896, n9895, n9894, n9893, n9892, n9891, n9890, n9889, n9888, n9887,
         n9886, n9885, n9884, n9883, n9882, n9881, n9880, n9879, n9878, n9877,
         n9876, n9875, n9874, n9873, n9872, n9871, n9870, n9869, n9868, n9867,
         n9866, n9865, n9864, n9863, n9862, n9861, n9860, n9859, n9858, n9857,
         n9856, n9855, n9854, n9853, n9852, n9851, n9850, n9849, n9848, n9847,
         n9846, n9845, n9844, n9843, n9842, n9841, n9840, n9839, n9838, n9837,
         n9836, n9835, n9834, n9833, n9832, n9831, n9830, n9829, n9828, n9827,
         n9826, n9825, n9824, n9823, n9822, n9821, n9820, n9819, n9818, n9817,
         n9816, n9815, n9814, n9813, n9812, n9811, n9810, n9809, n9808, n9807,
         n9806, n9805, n9804, n9803, n9802, n9801, n9800, n9799, n9798, n9797,
         n9796, n9795, n9794, n9793, n9792, n9791, n9790, n9789, n9788, n9787,
         n9786, n9785, n9784, n9783, n9782, n9781, n9780, n9779, n9778, n9777,
         n9776, n9775, n9774, n9773, n9772, n9771, n9770, n9769, n9768, n9767,
         n9766, n9765, n9764, n9763, n9762, n9761, n9760, n9759, n9758, n9757,
         n9756, n9755, n9754, n9753, n9752, n9751, n9750, n9749, n9748, n9747,
         n9746, n9745, n9744, n9743, n9742, n9741, n9740, n9739, n9738, n9737,
         n9736, n9735, n9734, n9733, n9732, n9731, n9730, n9729, n9728, n9727,
         n9726, n9725, n9724, n9723, n9722, n9721, n9720, n9719, n9718, n9717,
         n9716, n9715, n9714, n9713, n9712, n9711, n9710, n9709, n9708, n9707,
         n9706, n9705, n9704, n9703, n9702, n9701, n9700, n9699, n9698, n9697,
         n9696, n9695, n9694, n9693, n9692, n9691, n9690, n9689, n9688, n9687,
         n9686, n9685, n9684, n9683, n9682, n9681, n9680, n9679, n9678, n9677,
         n9676, n9675, n9674, n9673, n9672, n9671, n9670, n9669, n9668, n9667,
         n9666, n9665, n9664, n9663, n9662, n9661, n9660, n9659, n9658, n9657,
         n9656, n9655, n9654, n9653, n9652, n9651, n9650, n9649, n9648, n9647,
         n9646, n9645, n9644, n9643, n9642, n9641, n9640, n9639, n9638, n9637,
         n9636, n9635, n9634, n9633, n9632, n9631, n9630, n9629, n9628, n9627,
         n9626, n9625, n9624, n9623, n9622, n9621, n9620, n9619, n9618, n9617,
         n9616, n9615, n9614, n9613, n9612, n9611, n9610, n9609, n9608, n9607,
         n9606, n9605, n9604, n9603, n9602, n9601, n9600, n9599, n9598, n9597,
         n9596, n9595, n9594, n9593, n9592, n9591, n9590, n9589, n9588, n9587,
         n9586, n9585, n9584, n9583, n9582, n9581, n9580, n9579, n9578, n9577,
         n9576, n9575, n9574, n9573, n9572, n9571, n9570, n9569, n9568, n9567,
         n9566, n9565, n9564, n9563, n9562, n9561, n9560, n9559, n9558, n9557,
         n9556, n9555, n9554, n9553, n9552, n9551, n9550, n9549, n9548, n9547,
         n9546, n9545, n9544, n9543, n9542, n9541, n9540, n9539, n9538, n9537,
         n9536, n9535, n9534, n9533, n9532, n9531, n9530, n9529, n9528, n9527,
         n9526, n9525, n9524, n9523, n9522, n9521, n9520, n9519, n9518, n9517,
         n9516, n9515, n9514, n9513, n9512, n9511, n9510, n9509, n9508, n9507,
         n9506, n9505, n9504, n9503, n9502, n9501, n9500, n9499, n9498, n9497,
         n9496, n9495, n9494, n9493, n9492, n9491, n9490, n9489, n9488, n9487,
         n9486, n9485, n9484, n9483, n9482, n9481, n9480, n9479, n9478, n9477,
         n9476, n9475, n9474, n9473, n9472, n9471, n9470, n9469, n9468, n9467,
         n9466, n9465, n9464, n9463, n9462, n9461, n9460, n9459, n9458, n9457,
         n9456, n9455, n9454, n9453, n9452, n9451, n9450, n9449, n9448, n9447,
         n9446, n9445, n9444, n9443, n9442, n9441, n9440, n9439, n9438, n9437,
         n9436, n9435, n9434, n9433, n9432, n9431, n9430, n9429, n9428, n9427,
         n9426, n9425, n9424, n9423, n9422, n9421, n9420, n9419, n9418, n9417,
         n9416, n9415, n9414, n9413, n9412, n9411, n9410, n9409, n9408, n9407,
         n9406, n9405, n9404, n9403, n9402, n9401, n9400, n9399, n9398, n9397,
         n9396, n9395, n9394, n9393, n9392, n9391, n9390, n9389, n9388, n9387,
         n9386, n9385, n9384, n9383, n9382, n9381, n9380, n9379, n9378, n9377,
         n9376, n9375, n9374, n9373, n9372, n9371, n9370, n9369, n9368, n9367,
         n9366, n9365, n9364, n9363, n9362, n9361, n9360, n9359, n9358, n9357,
         n9356, n9355, n9354, n9353, n9352, n9351, n9350, n9349, n9348, n9347,
         n9346, n9345, n9344, n9343, n9342, n9341, n9340, n9339, n9338, n9337,
         n9336, n9335, n9334, n9333, n9332, n9331, n9330, n9329, n9328, n9327,
         n9326, n9325, n9324, n9323, n9322, n9321, n9320, n9319, n9318, n9317,
         n9316, n9315, n9314, n9313, n9312, n9311, n9310, n9309, n9308, n9307,
         n9306, n9305, n9304, n9303, n9302, n9301, n9300, n9299, n9298, n9297,
         n9296, n9295, n9294, n9293, n9292, n9291, n9290, n9289, n9288, n9287,
         n9286, n9285, n9284, n9283, n9282, n9281, n9280, n9279, n9278, n9277,
         n9276, n9275, n9274, n9273, n9272, n9271, n9270, n9269, n9268, n9267,
         n9266, n9265, n9264, n9263, n9262, n9261, n9260, n9259, n9258, n9257,
         n9256, n9255, n9254, n9253, n9252, n9251, n9250, n9249, n9248, n9247,
         n9246, n9245, n9244, n9243, n9242, n9241, n9240, n9239, n9238, n9237,
         n9236, n9235, n9234, n9233, n9232, n9231, n9230, n9229, n9228, n9227,
         n9226, n9225, n9224, n9223, n9222, n9221, n9220, n9219, n9218, n9217,
         n9216, n9215, n9214, n9213, n9212, n9211, n9210, n9209, n9208, n9207,
         n9206, n9205, n9204, n9203, n9202, n9201, n9200, n9199, n9198, n9197,
         n9196, n9195, n9194, n9193, n9192, n9191, n9190, n9189, n9188, n9187,
         n9186, n9185, n9184, n9183, n9182, n9181, n9180, n9179, n9178, n9177,
         n9176, n9175, n9174, n9173, n9172, n9171, n9170, n9169, n9168, n9167,
         n9166, n9165, n9164, n9163, n9162, n9161, n9160, n9159, n9158, n9157,
         n9156, n9155, n9154, n9153, n9152, n9151, n9150, n9149, n9148, n9147,
         n9146, n9145, n9144, n9143, n9142, n9141, n9140, n9139, n9138, n9137,
         n9136, n9135, n9134, n9133, n9132, n9131, n9130, n9129, n9128, n9127,
         n9126, n9125, n9124, n9123, n9122, n9121, n9120, n9119, n9118, n9117,
         n9116, n9115, n9114, n9113, n9112, n9111, n9110, n9109, n9108, n9107,
         n9106, n9105, n9104, n9103, n9102, n9101, n9100, n9099, n9098, n9097,
         n9096, n9095, n9094, n9093, n9092, n9091, n9090, n9089, n9088, n9087,
         n9086, n9085, n9084, n9083, n9082, n9081, n9080, n9079, n9078, n9077,
         n9076, n9075, n9074, n9073, n9072, n9071, n9070, n9069, n9068, n9067,
         n9066, n9065, n9064, n9063, n9062, n9061, n9060, n9059, n9058, n9057,
         n9056, n9055, n9054, n9053, n9052, n9051, n9050, n9049, n9048, n9047,
         n9046, n9045, n9044, n9043, n9042, n9041, n9040, n9039, n9038, n9037,
         n9036, n9035, n9034, n9033, n9032, n9031, n9030, n9029, n9028, n9027,
         n9026, n9025, n9024, n9023, n9022, n9021, n9020, n9019, n9018, n9017,
         n9016, n9015, n9014, n9013, n9012, n9011, n9010, n9009, n9008, n9007,
         n9006, n9005, n9004, n9003, n9002, n9001, n9000, n8999, n8998, n8997,
         n8996, n8995, n8994, n8993, n8992, n8991, n8990, n8989, n8988, n8987,
         n8986, n8985, n8984, n8983, n8982, n8981, n8980, n8979, n8978, n8977,
         n8976, n8975, n8974, n8973, n8972, n8971, n8970, n8969, n8968, n8967,
         n8966, n8965, n8964, n8963, n8962, n8961, n8960, n8959, n8958, n8957,
         n8956, n8955, n8954, n8953, n8952, n8951, n8950, n8949, n8948, n8947,
         n8946, n8945, n8944, n8943, n8942, n8941, n8940, n8939, n8938, n8937,
         n8936, n8935, n8934, n8933, n8932, n8931, n8930, n8929, n8928, n8927,
         n8926, n8925, n8924, n8923, n8922, n8921, n8920, n8919, n8918, n8917,
         n8916, n8915, n8914, n8913, n8912, n8911, n8910, n8909, n8908, n8907,
         n8906, n8905, n8904, n8903, n8902, n8901, n8900, n8899, n8898, n8897,
         n8896, n8895, n8894, n8893, n8892, n8891, n8890, n8889, n8888, n8887,
         n8886, n8885, n8884, n8883, n8882, n8881, n8880, n8879, n8878, n8877,
         n8876, n8875, n8874, n8873, n8872, n8871, n8870, n8869, n8868, n8867,
         n8866, n8865, n8864, n8863, n8862, n8861, n8860, n8859, n8858, n8857,
         n8856, n8855, n8854, n8853, n8852, n8851, n8850, n8849, n8848, n8847,
         n8846, n8845, n8844, n8843, n8842, n8841, n8840, n8839, n8838, n8837,
         n8836, n8835, n8834, n8833, n8832, n8831, n8830, n8829, n8828, n8827,
         n8826, n8825, n8824, n8823, n8822, n8821, n8820, n8819, n8818, n8817,
         n8816, n8815, n8814, n8813, n8812, n8811, n8810, n8809, n8808, n8807,
         n8806, n8805, n8804, n8803, n8802, n8801, n8800, n8799, n8798, n8797,
         n8796, n8795, n8794, n8793, n8792, n8791, n8790, n8789, n8788, n8787,
         n8786, n8785, n8784, n8783, n8782, n8781, n8780, n8779, n8778, n8777,
         n8776, n8775, n8774, n8773, n8772, n8771, n8770, n8769, n8768, n8767,
         n8766, n8765, n8764, n8763, n8762, n8761, n8760, n8759, n8758, n8757,
         n8756, n8755, n8754, n8753, n8752, n8751, n8750, n8749, n8748, n8747,
         n8746, n8745, n8744, n8743, n8742, n8741, n8740, n8739, n8738, n8737,
         n8736, n8735, n8734, n8733, n8732, n8731, n8730, n8729, n8728, n8727,
         n8726, n8725, n8724, n8723, n8722, n8721, n8720, n8719, n8718, n8717,
         n8716, n8715, n8714, n8713, n8712, n8711, n8710, n8709, n8708, n8707,
         n8706, n8705, n8704, n8703, n8702, n8701, n8700, n8699, n8698, n8697,
         n8696, n8695, n8694, n8693, n8692, n8691, n8690, n8689, n8688, n8687,
         n8686, n8685, n8684, n8683, n8682, n8681, n8680, n8679, n8678, n8677,
         n8676, n8675, n8674, n8673, n8672, n8671, n8670, n8669, n8668, n8667,
         n8666, n8665, n8664, n8663, n8662, n8661, n8660, n8659, n8658, n8657,
         n8656, n8655, n8654, n8653, n8652, n8651, n8650, n8649, n8648, n8647,
         n8646, n8645, n8644, n8643, n8642, n8641, n8640, n8639, n8638, n8637,
         n8636, n8635, n8634, n8633, n8632, n8631, n8630, n8629, n8628, n8627,
         n8626, n8625, n8624, n8623, n8622, n8621, n8620, n8619, n8618, n8617,
         n8616, n8615, n8614, n8613, n8612, n8611, n8610, n8609, n8608, n8607,
         n8606, n8605, n8604, n8603, n8602, n8601, n8600, n8599, n8598, n8597,
         n8596, n8595, n8594, n8593, n8592, n8591, n8590, n8589, n8588, n8587,
         n8586, n8585, n8584, n8583, n8582, n8581, n8580, n8579, n8578, n8577,
         n8576, n8575, n8574, n8573, n8572, n8571, n8570, n8569, n8568, n8567,
         n8566, n8565, n8564, n8563, n8562, n8561, n8560, n8559, n8558, n8557,
         n8556, n8555, n8554, n8553, n8552, n8551, n8550, n8549, n8548, n8547,
         n8546, n8545, n8544, n8543, n8542, n8541, n8540, n8539, n8538, n8537,
         n8536, n8535, n8534, n8533, n8532, n8531, n8530, n8529, n8528, n8527,
         n8526, n8525, n8524, n8523, n8522, n8521, n8520, n8519, n8518, n8517,
         n8516, n8515, n8514, n8513, n8512, n8511, n8510, n8509, n8508, n8507,
         n8506, n8505, n8504, n8503, n8502, n8501, n8500, n8499, n8498, n8497,
         n8496, n8495, n8494, n8493, n8492, n8491, n8490, n8489, n8488, n8487,
         n8486, n8485, n8484, n8483, n8482, n8481, n8480, n8479, n8478, n8477,
         n8476, n8475, n8474, n8473, n8472, n8471, n8470, n8469, n8468, n8467,
         n8466, n8465, n8464, n8463, n8462, n8461, n8460, n8459, n8458, n8457,
         n8456, n8455, n8454, n8453, n8452, n8451, n8450, n8449, n8448, n8447,
         n8446, n8445, n8444, n8443, n8442, n8441, n8440, n8439, n8438, n8437,
         n8436, n8435, n8434, n8433, n8432, n8431, n8430, n8429, n8428, n8427,
         n8426, n8425, n8424, n8423, n8422, n8421, n8420, n8419, n8418, n8417,
         n8416, n8415, n8414, n8413, n8412, n8411, n8410, n8409, n8408, n8407,
         n8406, n8405, n8404, n8403, n8402, n8401, n8400, n8399, n8398, n8397,
         n8396, n8395, n8394, n8393, n8392, n8391, n8390, n8389, n8388, n8387,
         n8386, n8385, n8384, n8383, n8382, n8381, n8380, n8379, n8378, n8377,
         n8376, n8375, n8374, n8373, n8372, n8371, n8370, n8369, n8368, n8367,
         n8366, n8365, n8364, n8363, n8362, n8361, n8360, n8359, n8358, n8357,
         n8356, n8355, n8354, n8353, n8352, n8351, n8350, n8349, n8348, n8347,
         n8346, n8345, n8344, n8343, n8342, n8341, n8340, n8339, n8338, n8337,
         n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328, n8327,
         n8326, n8325, n8324, n8323, n8322, n8321, n8320, n8319, n8318, n8317,
         n8316, n8315, n8314, n8313, n8312, n8311, n8310, n8309, n8308, n8307,
         n8306, n8305, n8304, n8303, n8302, n8301, n8300, n8299, n8298, n8297,
         n8296, n8295, n8294, n8293, n8292, n8291, n8290, n8289, n8288, n8287,
         n8286, n8285, n8284, n8283, n8282, n8281, n8280, n8279, n8278, n8277,
         n8276, n8275, n8274, n8273, n8272, n8271, n8270, n8269, n8268, n8267,
         n8266, n8265, n8264, n8263, n8262, n8261, n8260, n8259, n8258, n8257,
         n8256, n8255, n8254, n8253, n8252, n8251, n8250, n8249, n8248, n8247,
         n8246, n8245, n8244, n8243, n8242, n8241, n8240, n8239, n8238, n8237,
         n8236, n8235, n8234, n8233, n8232, n8231, n8230, n8229, n8228, n8227,
         n8226, n8225, n8224, n8223, n8222, n8221, n8220, n8219, n8218, n8217,
         n8216, n8215, n8214, n8213, n8212, n8211, n8210, n8209, n8208, n8207,
         n8206, n8205, n8204, n8203, n8202, n8201, n8200, n8199, n8198, n8197,
         n8196, n8195, n8194, n8193, n8192, n8191, n8190, n8189, n8188, n8187,
         n8186, n8185, n8184, n8183, n8182, n8181, n8180, n8179, n8178, n8177,
         n8176, n8175, n8174, n8173, n8172, n8171, n8170, n8169, n8168, n8167,
         n8166, n8165, n8164, n8163, n8162, n8161, n8160, n8159, n8158, n8157,
         n8156, n8155, n8154, n8153, n8152, n8151, n8150, n8149, n8148, n8147,
         n8146, n8145, n8144, n8143, n8142, n8141, n8140, n8139, n8138, n8137,
         n8136, n8135, n8134, n8133, n8132, n8131, n8130, n8129, n8128, n8127,
         n8126, n8125, n8124, n8123, n8122, n8121, n8120, n8119, n8118, n8117,
         n8116, n8115, n8114, n8113, n8112, n8111, n8110, n8109, n8108, n8107,
         n8106, n8105, n8104, n8103, n8102, n8101, n8100, n8099, n8098, n8097,
         n8096, n8095, n8094, n8093, n8092, n8091, n8090, n8089, n8088, n8087,
         n8086, n8085, n8084, n8083, n8082, n8081, n8080, n8079, n8078, n8077,
         n8076, n8075, n8074, n8073, n8072, n8071, n8070, n8069, n8068, n8067,
         n8066, n8065, n8064, n8063, n8062, n8061, n8060, n8059, n8058, n8057,
         n8056, n8055, n8054, n8053, n8052, n8051, n8050, n8049, n8048, n8047,
         n8046, n8045, n8044, n8043, n8042, n8041, n8040, n8039, n8038, n8037,
         n8036, n8035, n8034, n8033, n8032, n8031, n8030, n8029, n8028, n8027,
         n8026, n8025, n8024, n8023, n8022, n8021, n8020, n8019, n8018, n8017,
         n8016, n8015, n8014, n8013, n8012, n8011, n8010, n8009, n8008, n8007,
         n8006, n8005, n8004, n8003, n8002, n8001, n8000, n7999, n7998, n7997,
         n7996, n7995, n7994, n7993, n7992, n7991, n7990, n7989, n7988, n7987,
         n7986, n7985, n7984, n7983, n7982, n7981, n7980, n7979, n7978, n7977,
         n7976, n7975, n7974, n7973, n7972, n7971, n7970, n7969, n7968, n7967,
         n7966, n7965, n7964, n7963, n7962, n7961, n7960, n7959, n7958, n7957,
         n7956, n7955, n7954, n7953, n7952, n7951, n7950, n7949, n7948, n7947,
         n7946, n7945, n7944, n7943, n7942, n7941, n7940, n7939, n7938, n7937,
         n7936, n7935, n7934, n7933, n7932, n7931, n7930, n7929, n7928, n7927,
         n7926, n7925, n7924, n7923, n7922, n7921, n7920, n7919, n7918, n7917,
         n7916, n7915, n7914, n7913, n7912, n7911, n7910, n7909, n7908, n7907,
         n7906, n7905, n7904, n7903, n7902, n7901, n7900, n7899, n7898, n7897,
         n7896, n7895, n7894, n7893, n7892, n32139, n32138, n32137, n32136,
         n32135, n32134, n32133, n32132, n32131, n32130, n32129, n32128,
         n32127, n32126, n32125, n32124, n32123, n32122, n32121, n32120,
         n32119, n32118, n32117, n32116, n32115, n32114, n32113, n32112,
         n32111, n32110, n32109, n32108, n32107, n32106, n32105, n32104,
         n32103, n32102, n32101, n32100, n32099, n32098, n32097, n32096,
         n32095, n32094, n32093, n32092, n32091, n32090, n32089, n32088,
         n32087, n32086, n32085, n32084, n32083, n32082, n32081, n32080,
         n32079, n32078, n32077, n32076, n32075, n32074, n32073, n32072,
         n32071, n32070, n32069, n32068, n32067, n32066, n32065, n32064,
         n32063, n32062, n32061, n32060, n32059, n32058, n32057, n32056,
         n32055, n32054, n32053, n32052, n32051, n32050, n32049, n32048,
         n32047, n32046, n32045, n32044, n32043, n32042, n32041, n32040,
         n32039, n32038, n32037, n32036, n32035, n32034, n32033, n32032,
         n32031, n32030, n32029, n32028, n32027, n32026, n32025, n32024,
         n32023, n32022, n32021, n32020, n32019, n32018, n32017, n32016,
         n32015, n32014, n32013, n32012, n32011, n32010, n32009, n32008,
         n32007, n32006, n32005, n32004, n32003, n32002, n32001, n32000,
         n31999, n31998, n31997, n31995, n31994, n31993, n31992, n31991,
         n31990, n31989, n31988, n31987, n31986, n31985, n31984, n31983,
         n31982, n31981, n31980, n31979, n31978, n31977, n31976, n31975,
         n31974, n31973, n31972, n31971, n31970, n31969, n31968, n31967,
         n31966, n31965, n31964, n31963, n31962, n31961, n31960, n31959,
         n31958, n31957, n31956, n31955, n31954, n31953, n31952, n31951,
         n31950, n31949, n31948, n31947, n31946, n31945, n31944, n31943,
         n31942, n31941, n31940, n31939, n31938, n31937, n31936, n31935,
         n31934, n31933, n31932, n31931, n31930, n31929, n31928, n31927,
         n31926, n31925, n31924, n31923, n31922, n31921, n31920, n31919,
         n31918, n31917, n31916, n31915, n31914, n31913, n31912, n31911,
         n31910, n31909, n31908, n31907, n31906, n31905, n31904, n31903,
         n31902, n31901, n31900, n31899, n31898, n31897, n31896, n31895,
         n31894, n31893, n31892, n31891, n31890, n31889, n31888, n31887,
         n31886, n31885, n31884, n31883, n31882, n31881, n31880, n31879,
         n31878, n31877, n31876, n31875, n31874, n31873, n31872, n31871,
         n31870, n31869, n31868, n31867, n31866, n31865, n31864, n31863,
         n31862, n31861, n31860, n31859, n31858, n31857, n31856, n31855,
         n31854, n31853, n31852, n31851, n31850, n31849, n31848, n31847,
         n31846, n31845, n31844, n31843, n31842, n31841, n31840, n31839,
         n31838, n31837, n31836, n31835, n31834, n31833, n31832, n31831,
         n31830, n31829, n31828, n31827, n31826, n31825, n31824, n31823,
         n31822, n31821, n31820, n31819, n31818, n31817, n31816, n31815,
         n31814, n31813, n31812, n31811, n31810, n31809, n31808, n31807,
         n31806, n31805, n31804, n31803, n31802, n31801, n31800, n31799,
         n31798, n31797, n31796, n31795, n31794, n31793, n31792, n31791,
         n31790, n31789, n31788, n31787, n31786, n31785, n31784, n31783,
         n31782, n31781, n31780, n31779, n31778, n31777, n31776, n31775,
         n31774, n31773, n31772, n31771, n31770, n31769, n31768, n31767,
         n31766, n31765, n31764, n31763, n31762, n31761, n31760, n31759,
         n31758, n31757, n31756, n31755, n31754, n31753, n31752, n31751,
         n31750, n31749, n31748, n31747, n31746, n31745, n31744, n31743,
         n31742, n31741, n31740, n31739, n31738, n31737, n31736, n31735,
         n31734, n31733, n31732, n31731, n31730, n31729, n31728, n31727,
         n31726, n31725, n31724, n31723, n31722, n31721, n31720, n31719,
         n31718, n31717, n31716, n31715, n31714, n31713, n31712, n31711,
         n31710, n31709, n31708, n31707, n31706, n31705, n31704, n31703,
         n31702, n31701, n31700, n31699, n31698, n31697, n31696, n31695,
         n31694, n31693, n31692, n31691, n31690, n31689, n31688, n31687,
         n31686, n31685, n31684, n31683, n31682, n31681, n31680, n31679,
         n31678, n31677, n31676, n31675, n31674, n31673, n31672, n31671,
         n31670, n31669, n31668, n31667, n31666, n31665, n31664, n31663,
         n31662, n31661, n31660, n31659, n31658, n31657, n31656, n31655,
         n31654, n31653, n31652, n31651, n31650, n31649, n31648, n31647,
         n31646, n31645, n31644, n31643, n31642, n31641, n31640, n31639,
         n31638, n31637, n31636, n31635, n31634, n31633, n31632, n31631,
         n31630, n31629, n31628, n31627, n31626, n31625, n31624, n31623,
         n31622, n31621, n31620, n31619, n31618, n31617, n31616, n31615,
         n31614, n31613, n31612, n31611, n31610, n31609, n31608, n31607,
         n31606, n31605, n31604, n31603, n31602, n31601, n31600, n31599,
         n31598, n31597, n31596, n31595, n31594, n31593, n31592, n31591,
         n31590, n31589, n31588, n31587, n31586, n31585, n31584, n31583,
         n31582, n31581, n31580, n31579, n31578, n31577, n31576, n31575,
         n31574, n31573, n31572, n31571, n31570, n31569, n31568, n31567,
         n31566, n31565, n31564, n31563, n31562, n31561, n31560, n31559,
         n31558, n31557, n31556, n31555, n31554, n31553, n31552, n31551,
         n31550, n31549, n31548, n31547, n31546, n31545, n31544, n31543,
         n31542, n31541, n31540, n31539, n31538, n31537, n31536, n31535,
         n31534, n31533, n31532, n31531, n31530, n31529, n31528, n31527,
         n31526, n31525, n31524, n31523, n31522, n31521, n31520, n31519,
         n31518, n31517, n31516, n31515, n31514, n31513, n31512, n31511,
         n31510, n31509, n31508, n31507, n31506, n31505, n31504, n31503,
         n31502, n31501, n31500, n31499, n31498, n31497, n31496, n31495,
         n31494, n31493, n31492, n31491, n31490, n31489, n31488, n31487,
         n31486, n31485, n31484, n31483, n31482, n31481, n31480, n31479,
         n31478, n31477, n31476, n31475, n31474, n31473, n31472, n31471,
         n31470, n31469, n31468, n31467, n31466, n31465, n31464, n31463,
         n31462, n31461, n31460, n31459, n31458, n31457, n31456, n31455,
         n31454, n31453, n31452, n31451, n31450, n31449, n31448, n31447,
         n31446, n31445, n31444, n31443, n31442, n31441, n31440, n31439,
         n31438, n31437, n31436, n31435, n31434, n31433, n31432, n31431,
         n31430, n31429, n31428, n31427, n31426, n31425, n31424, n31423,
         n31422, n31421, n31420, n31419, n31418, n31417, n31416, n31415,
         n31414, n31413, n31412, n31411, n31410, n31409, n31408, n31407,
         n31406, n31405, n31404, n31403, n31402, n31401, n31400, n31399,
         n31398, n31397, n31396, n31395, n31394, n31393, n31392, n31391,
         n31390, n31389, n31388, n31387, n31386, n31385, n31384, n31383,
         n31382, n31381, n31380, n31379, n31378, n31377, n31376, n31375,
         n31374, n31373, n31372, n31371, n31370, n31369, n31368, n31367,
         n31366, n31365, n31364, n31363, n31362, n31361, n31360, n31359,
         n31358, n31357, n31356, n31355, n31354, n31353, n31352, n31351,
         n31350, n31349, n31348, n31347, n31346, n31345, n31344, n31343,
         n31342, n31341, n31340, n31339, n31338, n31337, n31336, n31335,
         n31334, n31333, n31332, n31331, n31330, n31329, n31328, n31327,
         n31326, n31325, n31324, n31323, n31322, n31321, n31320, n31319,
         n31318, n31317, n31316, n31315, n31314, n31313, n31312, n31311,
         n31310, n31309, n31308, n31307, n31306, n31305, n31304, n31303,
         n31302, n31301, n31300, n31299, n31298, n31297, n31296, n31295,
         n31294, n31293, n31292, n31291, n31290, n31289, n31288, n31287,
         n31286, n31285, n31284, n31283, n31282, n31281, n31280, n31279,
         n31278, n31277, n31276, n31275, n31274, n31273, n31272, n31271,
         n31270, n31269, n31268, n31267, n31266, n31265, n31264, n31263,
         n31262, n31261, n31260, n31259, n31258, n31257, n31256, n31255,
         n31254, n31253, n31252, n31251, n31250, n31249, n31248, n31247,
         n31246, n31245, n31244, n31243, n31242, n31241, n31240, n31239,
         n31238, n31237, n31236, n31235, n31234, n31233, n31232, n31231,
         n31230, n31229, n31228, n31227, n31226, n31225, n31224, n31223,
         n31222, n31221, n31220, n31219, n31218, n31217, n31216, n31215,
         n31214, n31213, n31212, n31211, n31210, n31209, n31208, n31207,
         n31206, n31205, n31204, n31203, n31202, n31201, n31200, n31199,
         n31198, n31197, n31196, n31195, n31194, n31193, n31192, n31191,
         n31190, n31189, n31188, n31187, n31186, n31185, n31184, n31183,
         n31182, n31181, n31180, n31179, n31178, n31177, n31176, n31175,
         n31174, n31173, n31172, n31171, n31170, n31169, n31168, n31167,
         n31166, n31165, n31164, n31163, n31162, n31161, n31160, n31159,
         n31158, n31157, n31156, n31155, n31154, n31153, n31152, n31151,
         n31150, n31149, n31148, n31147, n31146, n31145, n31144, n31143,
         n31142, n31141, n31140, n31139, n31138, n31137, n31136, n31135,
         n31134, n31133, n31132, n31131, n31130, n31129, n31128, n31127,
         n31126, n31125, n31124, n31123, n31122, n31121, n31120, n31119,
         n31118, n31117, n31116, n31115, n31114, n31113, n31112, n31111,
         n31110, n31109, n31108, n31107, n31106, n31105, n31104, n31103,
         n31102, n31101, n31100, n31099, n31098, n31097, n31096, n31095,
         n31094, n31093, n31092, n31091, n31090, n31089, n31088, n31087,
         n31086, n31085, n31084, n31083, n31082, n31081, n31080, n31079,
         n31078, n31077, n31076, n31075, n31074, n31073, n31072, n31071,
         n31070, n31069, n31068, n31067, n31066, n31065, n31064, n31063,
         n31062, n31061, n31060, n31059, n31058, n31057, n31056, n31055,
         n31054, n31053, n31052, n31051, n31050, n31049, n31048, n31047,
         n31046, n31045, n31044, n31043, n31042, n31041, n31040, n31039,
         n31038, n31037, n31036, n31035, n31034, n31033, n31032, n31031,
         n31030, n31029, n31028, n31027, n31026, n31025, n31024, n31023,
         n31022, n31021, n31020, n31019, n31018, n31017, n31016, n31015,
         n31014, n31013, n31012, n31011, n31010, n31009, n31008, n31007,
         n31006, n31005, n31004, n31003, n31002, n31001, n31000, n30999,
         n30998, n30997, n30996, n30995, n30994, n30993, n30992, n30991,
         n30990, n30989, n30988, n30987, n30986, n30985, n30984, n30983,
         n30982, n30981, n30980, n30979, n30978, n30977, n30976, n30975,
         n30974, n30973, n30972, n30971, n30970, n30969, n30968, n30967,
         n30966, n30965, n30964, n30963, n30962, n30961, n30960, n30959,
         n30958, n30957, n30956, n30955, n30954, n30953, n30952, n30951,
         n30950, n30949, n30948, n30947, n30946, n30945, n30944, n30943,
         n30942, n30941, n30940, n30939, n30938, n30937, n30936, n30935,
         n30934, n30933, n30932, n30931, n30930, n30929, n30928, n30927,
         n30926, n30925, n30924, n30923, n30922, n30921, n30920, n30919,
         n30918, n30917, n30916, n30915, n30914, n30913, n30912, n30911,
         n30910, n30909, n30908, n30907, n30906, n30905, n30904, n30903,
         n30902, n30901, n30900, n30899, n30898, n30897, n30896, n30895,
         n30894, n30893, n30892, n30891, n30890, n30889, n30888, n30887,
         n30886, n30885, n30884, n30883, n30882, n30881, n30880, n30879,
         n30878, n30877, n30876, n30875, n30874, n30873, n30872, n30871,
         n30870, n30869, n30868, n30867, n30866, n30865, n30864, n30863,
         n30862, n30861, n30860, n30859, n30858, n30857, n30856, n30855,
         n30854, n30853, n30852, n30851, n30850, n30849, n30848, n30847,
         n30846, n30845, n30844, n30843, n30842, n30841, n30840, n30839,
         n30838, n30837, n30836, n30835, n30834, n30833, n30832, n30831,
         n30830, n30829, n30828, n30827, n30826, n30825, n30824, n30823,
         n30822, n30821, n30820, n30819, n30818, n30817, n30816, n30815,
         n30814, n30813, n30812, n30811, n30810, n30809, n30808, n30807,
         n30806, n30805, n30804, n30803, n30802, n30801, n30800, n30799,
         n30798, n30797, n30796, n30795, n30794, n30793, n30792, n30791,
         n30790, n30789, n30788, n30787, n30786, n30785, n30784, n30783,
         n30782, n30781, n30780, n30779, n30778, n30777, n30776, n30775,
         n30774, n30773, n30772, n30771, n30770, n30769, n30768, n30767,
         n30766, n30765, n30764, n30763, n30762, n30761, n30760, n30759,
         n30758, n30757, n30756, n30755, n30754, n30753, n30752, n30751,
         n30750, n30749, n30748, n30747, n30746, n30745, n30744, n30743,
         n30742, n30741, n30740, n30739, n30738, n30737, n30736, n30735,
         n30734, n30733, n30732, n30731, n30730, n30729, n30728, n30727,
         n30726, n30725, n30724, n30723, n30722, n30721, n30720, n30719,
         n30718, n30717, n30716, n30715, n30714, n30713, n30712, n30711,
         n30710, n30709, n30708, n30707, n30706, n30705, n30704, n30703,
         n30702, n30701, n30700, n30699, n30698, n30697, n30696, n30695,
         n30694, n30693, n30692, n30691, n30690, n30689, n30688, n30687,
         n30686, n30685, n30684, n30683, n30682, n30681, n30680, n30679,
         n30678, n30677, n30676, n30675, n30674, n30673, n30672, n30671,
         n30670, n30669, n30668, n30667, n30666, n30665, n30664, n30663,
         n30662, n30661, n30660, n30659, n30658, n30657, n30656, n30655,
         n30654, n30653, n30652, n30651, n30650, n30649, n30648, n30647,
         n30646, n30645, n30644, n30643, n30642, n30641, n30640, n30639,
         n30638, n30637, n30636, n30635, n30634, n30633, n30632, n30631,
         n30630, n30629, n30628, n30627, n30626, n30625, n30624, n30623,
         n30622, n30621, n30620, n30619, n30618, n30617, n30616, n30615,
         n30614, n30613, n30612, n30611, n30610, n30609, n30608, n30607,
         n30606, n30605, n30604, n30603, n30602, n30601, n30600, n30599,
         n30598, n30597, n30596, n30595, n30594, n30593, n30592, n30591,
         n30590, n30589, n30588, n30587, n30586, n30585, n30584, n30583,
         n30582, n30581, n30580, n30579, n30578, n30577, n30576, n30575,
         n30574, n30573, n30572, n30571, n30570, n30569, n30568, n30567,
         n30566, n30565, n30564, n30563, n30562, n30561, n30560, n30559,
         n30558, n30557, n30556, n30555, n30554, n30553, n30552, n30551,
         n30550, n30549, n30548, n30547, n30546, n30545, n30544, n30543,
         n30542, n30541, n30540, n30539, n30538, n30537, n30536, n30535,
         n30534, n30533, n30532, n30531, n30530, n30529, n30528, n30527,
         n30526, n30525, n30524, n30523, n30522, n30521, n30520, n30519,
         n30518, n30517, n30516, n30515, n30514, n30513, n30512, n30511,
         n30510, n30509, n30508, n30507, n30506, n30505, n30504, n30503,
         n30502, n30501, n30500, n30499, n30498, n30497, n30496, n30495,
         n30494, n30493, n30492, n30491, n30490, n30489, n30488, n30487,
         n30486, n30485, n30484, n30483, n30482, n30481, n30480, n30479,
         n30478, n30477, n30476, n30475, n30474, n30473, n30472, n30471,
         n30470, n30469, n30468, n30467, n30466, n30465, n30464, n30463,
         n30462, n30461, n30460, n30459, n30458, n30457, n30456, n30455,
         n30454, n30453, n30452, n30451, n30450, n30449, n30448, n30447,
         n30446, n30445, n30444, n30443, n30442, n30441, n30440, n30439,
         n30438, n30437, n30436, n30435, n30434, n30433, n30432, n30431,
         n30430, n30429, n30428, n30427, n30426, n30425, n30424, n30423,
         n30422, n30421, n30420, n30419, n30418, n30417, n30416, n30415,
         n30414, n30413, n30412, n30411, n30410, n30409, n30408, n30407,
         n30406, n30405, n30404, n30403, n30402, n30401, n30400, n30399,
         n30398, n30397, n30396, n30395, n30394, n30393, n30392, n30391,
         n30390, n30389, n30388, n30387, n30386, n30385, n30384, n30383,
         n30382, n30381, n30380, n30379, n30378, n30377, n30376, n30375,
         n30374, n30373, n30372, n30371, n30370, n30369, n30368, n30367,
         n30366, n30365, n30364, n30363, n30362, n30361, n30360, n30359,
         n30358, n30357, n30356, n30355, n30354, n30353, n30352, n30351,
         n30350, n30349, n30348, n30347, n30346, n30345, n30344, n30343,
         n30342, n30341, n30340, n30339, n30338, n30337, n30336, n30335,
         n30334, n30333, n30332, n30331, n30330, n30329, n30328, n30327,
         n30326, n30325, n30324, n30323, n30322, n30321, n30320, n30319,
         n30318, n30317, n30316, n30315, n30314, n30313, n30312, n30311,
         n30310, n30309, n30308, n30307, n30306, n30305, n30304, n30303,
         n30302, n30301, n30300, n30299, n30298, n30297, n30296, n30295,
         n30294, n30293, n30292, n30291, n30290, n30289, n30288, n30287,
         n30286, n30285, n30284, n30283, n30282, n30281, n30280, n30279,
         n30278, n30277, n30276, n30275, n30274, n30273, n30272, n30271,
         n30270, n30269, n30268, n30267, n30266, n30265, n30264, n30263,
         n30262, n30261, n30260, n30259, n30258, n30257, n30256, n30255,
         n30254, n30253, n30252, n30251, n30250, n30249, n30248, n30247,
         n30246, n30245, n30244, n30243, n30242, n30241, n30240, n30239,
         n30238, n30237, n30236, n30235, n30234, n30233, n30232, n30231,
         n30230, n30229, n30228, n30227, n30226, n30225, n30224, n30223,
         n30222, n30221, n30220, n30219, n30218, n30217, n30216, n30215,
         n30214, n30213, n30212, n30211, n30210, n30209, n30208, n30207,
         n30206, n30205, n30204, n30203, n30202, n30201, n30200, n30199,
         n30198, n30197, n30196, n30195, n30194, n30193, n30192, n30191,
         n30190, n30189, n30188, n30187, n30186, n30185, n30184, n30183,
         n30182, n30181, n30180, n30179, n30178, n30177, n30176, n30175,
         n30174, n30173, n30172, n30171, n30170, n30169, n30168, n30167,
         n30166, n30165, n30164, n30163, n30162, n30161, n30160, n30159,
         n30158, n30157, n30156, n30155, n30154, n30153, n30152, n30151,
         n30150, n30149, n30148, n30147, n30146, n30145, n30144, n30143,
         n30142, n30141, n30140, n30139, n30138, n30137, n30136, n30135,
         n30134, n30133, n30132, n30131, n30130, n30129, n30128, n30127,
         n30126, n30125, n30124, n30123, n30122, n30121, n30120, n30119,
         n30118, n30117, n30116, n30115, n30114, n30113, n30112, n30111,
         n30110, n30109, n30108, n30107, n30106, n30105, n30104, n30103,
         n30102, n30101, n30100, n30099, n30098, n30097, n30096, n30095,
         n30094, n30093, n30092, n30091, n30090, n30089, n30088, n30087,
         n30086, n30085, n30084, n30083, n30082, n30081, n30080, n30079,
         n30078, n30077, n30076, n30075, n30074, n30073, n30072, n30071,
         n30070, n30069, n30068, n30067, n30066, n30065, n30064, n30063,
         n30062, n30061, n30060, n30059, n30058, n30057, n30056, n30055,
         n30054, n30053, n30052, n30051, n30050, n30049, n30048, n30047,
         n30046, n30045, n30044, n30043, n30042, n30041, n30040, n30039,
         n30038, n30037, n30036, n30035, n30034, n30033, n30032, n30031,
         n30030, n30029, n30028, n30027, n30026, n30025, n30024, n30023,
         n30022, n30021, n30020, n30019, n30018, n30017, n30016, n30015,
         n30014, n30013, n30012, n30011, n30010, n30009, n30008, n30007,
         n30006, n30005, n30004, n30003, n30002, n30001, n30000, n29999,
         n29998, n29997, n29996, n29995, n29994, n29993, n29992, n29991,
         n29990, n29989, n29988, n29987, n29986, n29985, n29984, n29983,
         n29982, n29981, n29980, n29979, n29978, n29977, n29976, n29975,
         n29974, n29973, n29972, n29971, n29970, n29969, n29968, n29967,
         n29966, n29965, n29964, n29963, n29962, n29961, n29960, n29959,
         n29958, n29957, n29956, n29955, n29954, n29953, n29952, n29951,
         n29950, n29949, n29948, n29947, n29946, n29945, n29944, n29943,
         n29942, n29941, n29940, n29939, n29938, n29937, n29936, n29935,
         n29934, n29933, n29932, n29931, n29930, n29929, n29928, n29927,
         n29926, n29925, n29924, n29923, n29922, n29921, n29920, n29919,
         n29918, n29917, n29916, n29915, n29914, n29913, n29912, n29911,
         n29910, n29909, n29908, n29907, n29906, n29905, n29904, n29903,
         n29902, n29901, n29900, n29899, n29898, n29897, n29896, n29895,
         n29894, n29893, n29892, n29891, n29890, n29889, n29888, n29887,
         n29886, n29885, n29884, n29883, n29882, n29881, n29880, n29879,
         n29878, n29877, n29876, n29875, n29874, n29873, n29872, n29871,
         n29870, n29869, n29868, n29867, n29866, n29865, n29864, n29863,
         n29862, n29861, n29860, n29859, n29858, n29857, n29856, n29855,
         n29854, n29853, n29852, n29851, n29850, n29849, n29848, n29847,
         n29846, n29845, n29844, n29843, n29842, n29841, n29840, n29839,
         n29838, n29837, n29836, n29835, n29834, n29833, n29832, n29831,
         n29830, n29829, n29828, n29827, n29826, n29825, n29824, n29823,
         n29822, n29821, n29820, n29819, n29818, n29817, n29816, n29815,
         n29814, n29813, n29812, n29811, n29810, n29809, n29808, n29807,
         n29806, n29805, n29804, n29803, n29802, n29801, n29800, n29799,
         n29798, n29797, n29796, n29795, n29794, n29793, n29792, n29791,
         n29790, n29789, n29788, n29787, n29786, n29785, n29784, n29783,
         n29782, n29781, n29780, n29779, n29778, n29777, n29776, n29775,
         n29774, n29773, n29772, n29771, n29770, n29769, n29768, n29767,
         n29766, n29765, n29764, n29763, n29762, n29761, n29760, n29759,
         n29758, n29757, n29756, n29755, n29754, n29753, n29752, n29751,
         n29750, n29749, n29748, n29747, n29746, n29745, n29744, n29743,
         n29742, n29741, n29740, n29739, n29738, n29737, n29736, n29735,
         n29734, n29733, n29732, n29731, n29730, n29729, n29728, n29727,
         n29726, n29725, n29724, n29723, n29722, n29721, n29720, n29719,
         n29718, n29717, n29716, n29715, n29714, n29713, n29712, n29711,
         n29710, n29709, n29708, n29707, n29706, n29705, n29704, n29703,
         n29702, n29701, n29700, n29699, n29698, n29697, n29696, n29695,
         n29694, n29693, n29692, n29691, n29690, n29689, n29688, n29687,
         n29686, n29685, n29684, n29683, n29682, n29681, n29680, n29679,
         n29678, n29677, n29676, n29675, n29674, n29673, n29672, n29671,
         n29670, n29669, n29668, n29667, n29666, n29665, n29664, n29663,
         n29662, n29661, n29660, n29659, n29658, n29657, n29656, n29655,
         n29654, n29653, n29652, n29651, n29650, n29649, n29648, n29647,
         n29646, n29645, n29644, n29643, n29642, n29641, n29640, n29639,
         n29638, n29637, n29636, n29635, n29634, n29633, n29632, n29631,
         n29630, n29629, n29628, n29627, n29626, n29625, n29624, n29623,
         n29622, n29621, n29620, n29619, n29618, n29617, n29616, n29615,
         n29614, n29613, n29612, n29611, n29610, n29609, n29608, n29607,
         n29606, n29605, n29604, n29603, n29602, n29601, n29600, n29599,
         n29598, n29597, n29596, n29595, n29594, n29593, n29592, n29591,
         n29590, n29589, n29588, n29587, n29586, n29585, n29584, n29583,
         n29582, n29581, n29580, n29579, n29578, n29577, n29576, n29575,
         n29574, n29573, n29572, n29571, n29570, n29569, n29568, n29567,
         n29566, n29565, n29564, n29563, n29562, n29561, n29560, n29559,
         n29558, n29557, n29556, n29555, n29554, n29553, n29552, n29551,
         n29550, n29549, n29548, n29547, n29546, n29545, n29544, n29543,
         n29542, n29541, n29540, n29539, n29538, n29537, n29536, n29535,
         n29534, n29533, n29532, n29531, n29530, n29529, n29528, n29527,
         n29526, n29525, n29524, n29523, n29522, n29521, n29520, n29519,
         n29518, n29517, n29516, n29515, n29514, n29513, n29512, n29511,
         n29510, n29509, n29508, n29507, n29506, n29505, n29504, n29503,
         n29502, n29501, n29500, n29499, n29498, n29497, n29496, n29495,
         n29494, n29493, n29492, n29491, n29490, n29489, n29488, n29487,
         n29486, n29485, n29484, n29483, n29482, n29481, n29480, n29479,
         n29478, n29477, n29476, n29475, n29474, n29473, n29472, n29471,
         n29470, n29469, n29468, n29467, n29466, n29465, n29464, n29463,
         n29462, n29461, n29460, n29459, n29458, n29457, n29456, n29455,
         n29454, n29453, n29452, n29451, n29450, n29449, n29448, n29447,
         n29446, n29445, n29444, n29443, n29442, n29441, n29440, n29439,
         n29438, n29437, n29436, n29435, n29434, n29433, n29432, n29431,
         n29430, n29429, n29428, n29427, n29426, n29425, n29424, n29423,
         n29422, n29421, n29420, n29419, n29418, n29417, n29416, n29415,
         n29414, n29413, n29412, n29411, n29410, n29409, n29408, n29407,
         n29406, n29405, n29404, n29403, n29402, n29401, n29400, n29399,
         n29398, n29397, n29396, n29395, n29394, n29393, n29392, n29391,
         n29390, n29389, n29388, n29387, n29386, n29385, n29384, n29383,
         n29382, n29381, n29380, n29379, n29378, n29377, n29376, n29375,
         n29374, n29373, n29372, n29371, n29370, n29369, n29368, n29367,
         n29366, n29365, n29364, n29363, n29362, n29361, n29360, n29359,
         n29358, n29357, n29356, n29355, n29354, n29353, n29352, n29351,
         n29350, n29349, n29348, n29347, n29346, n29345, n29344, n29343,
         n29342, n29341, n29340, n29339, n29338, n29337, n29336, n29335,
         n29334, n29333, n29332, n29331, n29330, n29329, n29328, n29327,
         n29326, n29325, n29324, n29323, n29322, n29321, n29320, n29319,
         n29318, n29317, n29316, n29315, n29314, n29313, n29312, n29311,
         n29310, n29309, n29308, n29307, n29306, n29305, n29304, n29303,
         n29302, n29301, n29300, n29299, n29298, n29297, n29296, n29295,
         n29294, n29293, n29292, n29291, n29290, n29289, n29288, n29287,
         n29286, n29285, n29284, n29283, n29282, n29281, n29280, n29279,
         n29278, n29277, n29276, n29275, n29274, n29273, n29272, n29271,
         n29270, n29269, n29268, n29267, n29266, n29265, n29264, n29263,
         n29262, n29261, n29260, n29259, n29258, n29257, n29256, n29255,
         n29254, n29253, n29252, n29251, n29250, n29249, n29248, n29247,
         n29246, n29245, n29244, n29243, n29242, n29241, n29240, n29239,
         n29238, n29237, n29236, n29235, n29234, n29233, n29232, n29231,
         n29230, n29229, n29228, n29227, n29226, n29225, n29224, n29223,
         n29222, n29221, n29220, n29219, n29218, n29217, n29216, n29215,
         n29214, n29213, n29212, n29211, n29210, n29209, n29208, n29207,
         n29206, n29205, n29204, n29203, n29202, n29201, n29200, n29199,
         n29198, n29197, n29196, n29195, n29194, n29193, n29192, n29191,
         n29190, n29189, n29188, n29187, n29186, n29185, n29184, n29183,
         n29182, n29181, n29180, n29179, n29178, n29177, n29176, n29175,
         n29174, n29173, n29172, n29171, n29170, n29169, n29168, n29167,
         n29166, n29165, n29164, n29163, n29162, n29161, n29160, n29159,
         n29158, n29157, n29156, n29155, n29154, n29153, n29152, n29151,
         n29150, n29149, n29148, n29147, n29146, n29145, n29144, n29143,
         n29142, n29141, n29140, n29139, n29138, n29137, n29136, n29135,
         n29134, n29133, n29132, n29131, n29130, n29129, n29128, n29127,
         n29126, n29125, n29124, n29123, n29122, n29121, n29120, n29119,
         n29118, n29117, n29116, n29115, n29114, n29113, n29112, n29111,
         n29110, n29109, n29108, n29107, n29106, n29105, n29104, n29103,
         n29102, n29101, n29100, n29099, n29098, n29097, n29096, n29095,
         n29094, n29093, n29092, n29091, n29090, n29089, n29088, n29087,
         n29086, n29085, n29084, n29083, n29082, n29081, n29080, n29079,
         n29078, n29077, n29076, n29075, n29074, n29073, n29072, n29071,
         n29070, n29069, n29068, n29067, n29066, n29065, n29064, n29063,
         n29062, n29061, n29060, n29059, n29058, n29057, n29056, n29055,
         n29054, n29053, n29052, n29051, n29050, n29049, n29048, n29047,
         n29046, n29045, n29044, n29043, n29042, n29041, n29040, n29039,
         n29038, n29037, n29036, n29035, n29034, n29033, n29032, n29031,
         n29030, n29029, n29028, n29027, n29026, n29025, n29024, n29023,
         n29022, n29021, n29020, n29019, n29018, n29017, n29016, n29015,
         n29014, n29013, n29012, n29011, n29010, n29009, n29008, n29007,
         n29006, n29005, n29004, n29003, n29002, n29001, n29000, n28999,
         n28998, n28997, n28996, n28995, n28994, n28993, n28992, n28991,
         n28990, n28989, n28988, n28987, n28986, n28985, n28984, n28983,
         n28982, n28981, n28980, n28979, n28978, n28977, n28976, n28975,
         n28974, n28973, n28972, n28971, n28970, n28969, n28968, n28967,
         n28966, n28965, n28964, n28963, n28962, n28961, n28960, n28959,
         n28958, n28957, n28956, n28955, n28954, n28953, n28952, n28951,
         n28950, n28949, n28948, n28947, n28946, n28945, n28944, n28943,
         n28942, n28941, n28940, n28939, n28938, n28937, n28936, n28935,
         n28934, n28933, n28932, n28931, n28930, n28929, n28928, n28927,
         n28926, n28925, n28924, n28923, n28922, n28921, n28920, n28919,
         n28918, n28917, n28916, n28915, n28914, n28913, n28912, n28911,
         n28910, n28909, n28908, n28907, n28906, n28905, n28904, n28903,
         n28902, n28901, n28900, n28899, n28898, n28897, n28896, n28895,
         n28894, n28893, n28892, n28891, n28890, n28889, n28888, n28887,
         n28886, n28885, n28884, n28883, n28882, n28881, n28880, n28879,
         n28878, n28877, n28876, n28875, n28874, n28873, n28872, n28871,
         n28870, n28869, n28868, n28867, n28866, n28865, n28864, n28863,
         n28862, n28861, n28860, n28859, n28858, n28857, n28856, n28855,
         n28854, n28853, n28852, n28851, n28850, n28849, n28848, n28847,
         n28846, n28845, n28844, n28843, n28842, n28841, n28840, n28839,
         n28838, n28837, n28836, n28835, n28834, n28833, n28832, n28831,
         n28830, n28829, n28828, n28827, n28826, n28825, n28824, n28823,
         n28822, n28821, n28820, n28819, n28818, n28817, n28816, n28815,
         n28814, n28813, n28812, n28811, n28810, n28809, n28808, n28807,
         n28806, n28805, n28804, n28803, n28802, n28801, n28800, n28799,
         n28798, n28797, n28796, n28795, n28794, n28793, n28792, n28791,
         n28790, n28789, n28788, n28787, n28786, n28785, n28784, n28783,
         n28782, n28781, n28780, n28779, n28778, n28777, n28776, n28775,
         n28774, n28773, n28772, n28771, n28770, n28769, n28768, n28767,
         n28766, n28765, n28764, n28763, n28762, n28761, n28760, n28759,
         n28758, n28757, n28756, n28755, n28754, n28753, n28752, n28751,
         n28750, n28749, n28748, n28747, n28746, n28745, n28744, n28743,
         n28742, n28741, n28740, n28739, n28738, n28737, n28736, n28735,
         n28734, n28733, n28732, n28731, n28730, n28729, n28728, n28727,
         n28726, n28725, n28724, n28723, n28722, n28721, n28720, n28719,
         n28718, n28717, n28716, n28715, n28714, n28713, n28712, n28711,
         n28710, n28709, n28708, n28707, n28706, n28705, n28704, n28703,
         n28702, n28701, n28700, n28699, n28698, n28697, n28696, n28695,
         n28694, n28693, n28692, n28691, n28690, n28689, n28688, n28687,
         n28686, n28685, n28684, n28683, n28682, n28681, n28680, n28679,
         n28678, n28677, n28676, n28675, n28674, n28673, n28672, n28671,
         n28670, n28669, n28668, n28667, n28666, n28665, n28664, n28663,
         n28662, n28661, n28660, n28659, n28658, n28657, n28656, n28655,
         n28654, n28653, n28652, n28651, n28650, n28649, n28648, n28647,
         n28646, n28645, n28644, n28643, n28642, n28641, n28640, n28639,
         n28638, n28637, n28636, n28635, n28634, n28633, n28632, n28631,
         n28630, n28629, n28628, n28627, n28626, n28625, n28624, n28623,
         n28622, n28621, n28620, n28619, n28618, n28617, n28616, n28615,
         n28614, n28613, n28612, n28611, n28610, n28609, n28608, n28607,
         n28606, n28605, n28604, n28603, n28602, n28601, n28600, n28599,
         n28598, n28597, n28596, n28595, n28594, n28593, n28592, n28591,
         n28590, n28589, n28588, n28587, n28586, n28585, n28584, n28583,
         n28582, n28581, n28580, n28579, n28578, n28577, n28576, n28575,
         n28574, n28573, n28572, n28571, n28570, n28569, n28568, n28567,
         n28566, n28565, n28564, n28563, n28562, n28561, n28560, n28559,
         n28558, n28557, n28556, n28555, n28554, n28553, n28552, n28551,
         n28550, n28549, n28548, n28547, n28546, n28545, n28544, n28543,
         n28542, n28541, n28540, n28539, n28538, n28537, n28536, n28535,
         n28534, n28533, n28532, n28531, n28530, n28529, n28528, n28527,
         n28526, n28525, n28524, n28523, n28522, n28521, n28520, n28519,
         n28518, n28517, n28516, n28515, n28514, n28513, n28512, n28511,
         n28510, n28509, n28508, n28507, n28506, n28505, n28504, n28503,
         n28502, n28501, n28500, n28499, n28498, n28497, n28496, n28495,
         n28494, n28493, n28492, n28491, n28490, n28489, n28488, n28487,
         n28486, n28485, n28484, n28483, n28482, n28481, n28480, n28479,
         n28478, n28477, n28476, n28475, n28474, n28473, n28472, n28471,
         n28470, n28469, n28468, n28467, n28466, n28465, n28464, n28463,
         n28462, n28461, n28460, n28459, n28458, n28457, n28456, n28455,
         n28454, n28453, n28452, n28451, n28450, n28449, n28448, n28447,
         n28446, n28445, n28444, n28443, n28442, n28441, n28440, n28439,
         n28438, n28437, n28436, n28435, n28434, n28433, n28432, n28431,
         n28430, n28429, n28428, n28427, n28426, n28425, n28424, n28423,
         n28422, n28421, n28420, n28419, n28418, n28417, n28416, n28415,
         n28414, n28413, n28412, n28411, n28410, n28409, n28408, n28407,
         n28406, n28405, n28404, n28403, n28402, n28401, n28400, n28399,
         n28398, n28397, n28396, n28395, n28394, n28393, n28392, n28391,
         n28390, n28389, n28388, n28387, n28386, n28385, n28384, n28383,
         n28382, n28381, n28380, n28379, n28378, n28377, n28376, n28375,
         n28374, n28373, n28372, n28371, n28370, n28369, n28368, n28367,
         n28366, n28365, n28364, n28363, n28362, n28361, n28360, n28359,
         n28358, n28357, n28356, n28355, n28354, n28353, n28352, n28351,
         n28350, n28349, n28348, n28347, n28346, n28345, n28344, n28343,
         n28342, n28341, n28340, n28339, n28338, n28337, n28336, n28335,
         n28334, n28333, n28332, n28331, n28330, n28329, n28328, n28327,
         n28326, n28325, n28324, n28323, n28322, n28321, n28320, n28319,
         n28318, n28317, n28316, n28315, n28314, n28313, n28312, n28311,
         n28310, n28309, n28308, n28307, n28306, n28305, n28304, n28303,
         n28302, n28301, n28300, n28299, n28298, n28297, n28296, n28295,
         n28294, n28293, n28292, n28291, n28290, n28289, n28288, n28287,
         n28286, n28285, n28284, n28283, n28282, n28281, n28280, n28279,
         n28278, n28277, n28276, n28275, n28274, n28273, n28272, n28271,
         n28270, n28269, n28268, n28267, n28266, n28265, n28264, n28263,
         n28262, n28261, n28260, n28259, n28258, n28257, n28256, n28255,
         n28254, n28253, n28252, n28251, n28250, n28249, n28248, n28247,
         n28246, n28245, n28244, n28243, n28242, n28241, n28240, n28239,
         n28238, n28237, n28236, n28235, n28234, n28233, n28232, n28231,
         n28230, n28229, n28228, n28227, n28226, n28225, n28224, n28223,
         n28222, n28221, n28220, n28219, n28218, n28217, n28216, n28215,
         n28214, n28213, n28212, n28211, n28210, n28209, n28208, n28207,
         n28206, n28205, n28204, n28203, n28202, n28201, n28200, n28199,
         n28198, n28197, n28196, n28195, n28194, n28193, n28192, n28191,
         n28190, n28189, n28188, n28187, n28186, n28185, n28184, n28183,
         n28182, n28181, n28180, n28179, n28178, n28177, n28176, n28175,
         n28174, n28173, n28172, n28171, n28170, n28169, n28168, n28167,
         n28166, n28165, n28164, n28163, n28162, n28161, n28160, n28159,
         n28158, n28157, n28156, n28155, n28154, n28153, n28152, n28151,
         n28150, n28149, n28148, n28147, n28146, n28145, n28144, n28143,
         n28142, n28141, n28140, n28139, n28138, n28137, n28136, n28135,
         n28134, n28133, n28132, n28131, n28130, n28129, n28128, n28127,
         n28126, n28125, n28124, n28123, n28122, n28121, n28120, n28119,
         n28118, n28117, n28116, n28115, n28114, n28113, n28112, n28111,
         n28110, n28109, n28108, n28107, n28106, n28105, n28104, n28103,
         n28102, n28101, n28100, n28099, n28098, n28097, n28096, n28095,
         n28094, n28093, n28092, n28091, n28090, n28089, n28088, n28087,
         n28086, n28085, n28084, n28083, n28082, n28081, n28080, n28079,
         n28078, n28077, n28076, n28075, n28074, n28073, n28072, n28071,
         n28070, n28069, n28068, n28067, n28066, n28065, n28064, n28063,
         n28062, n28061, n28060, n28059, n28058, n28057, n28056, n28055,
         n28054, n28053, n28052, n28051, n28050, n28049, n28048, n28047,
         n28046, n28045, n28044, n28043, n28042, n28041, n28040, n28039,
         n28038, n28037, n28036, n28035, n28034, n28033, n28032, n28031,
         n28030, n28029, n28028, n28027, n28026, n28025, n28024, n28023,
         n28022, n28021, n28020, n28019, n28018, n28017, n28016, n28015,
         n28014, n28013, n28012, n28011, n28010, n28009, n28008, n28007,
         n28006, n28005, n28004, n28003, n28002, n28001, n28000, n27999,
         n27998, n27997, n27996, n27995, n27994, n27993, n27992, n27991,
         n27990, n27989, n27988, n27987, n27986, n27985, n27984, n27983,
         n27982, n27981, n27980, n27979, n27978, n27977, n27976, n27975,
         n27974, n27973, n27972, n27971, n27970, n27969, n27968, n27967,
         n27966, n27965, n27964, n27963, n27962, n27961, n27960, n27959,
         n27958, n27957, n27956, n27955, n27954, n27953, n27952, n27951,
         n27950, n27949, n27948, n27947, n27946, n27945, n27944, n27943,
         n27942, n27941, n27940, n27939, n27938, n27937, n27936, n27935,
         n27934, n27933, n27932, n27931, n27930, n27929, n27928, n27927,
         n27926, n27925, n27924, n27923, n27922, n27921, n27920, n27919,
         n27918, n27917, n27916, n27915, n27914, n27913, n27912, n27911,
         n27910, n27909, n27908, n27907, n27906, n27905, n27904, n27903,
         n27902, n27901, n27900, n27899, n27898, n27897, n27896, n27895,
         n27894, n27893, n27892, n27891, n27890, n27889, n27888, n27887,
         n27886, n27885, n27884, n27883, n27882, n27881, n27880, n27879,
         n27878, n27877, n27876, n27875, n27874, n27873, n27872, n27871,
         n27870, n27869, n27868, n27867, n27866, n27865, n27864, n27863,
         n27862, n27861, n27860, n27859, n27858, n27857, n27856, n27855,
         n27854, n27853, n27852, n27851, n27850, n27849, n27848, n27847,
         n27846, n27845, n27844, n27843, n27842, n27841, n27840, n27839,
         n27838, n27837, n27836, n27835, n27834, n27833, n27832, n27831,
         n27830, n27829, n27828, n27827, n27826, n27825, n27824, n27823,
         n27822, n27821, n27820, n27819, n27818, n27817, n27816, n27815,
         n27814, n27813, n27812, n27811, n27810, n27809, n27808, n27807,
         n27806, n27805, n27804, n27803, n27802, n27801, n27800, n27799,
         n27798, n27797, n27796, n27795, n27794, n27793, n27792, n27791,
         n27790, n27789, n27788, n27787, n27786, n27785, n27784, n27783,
         n27782, n27781, n27780, n27779, n27778, n27777, n27776, n27775,
         n27774, n27773, n27772, n27771, n27770, n27769, n27768, n27767,
         n27766, n27765, n27764, n27763, n27762, n27761, n27760, n27759,
         n27758, n27757, n27756, n27755, n27754, n27753, n27752, n27751,
         n27750, n27749, n27748, n27747, n27746, n27745, n27744, n27743,
         n27742, n27741, n27740, n27739, n27738, n27737, n27736, n27735,
         n27734, n27733, n27732, n27731, n27730, n27729, n27728, n27727,
         n27726, n27725, n27724, n27723, n27722, n27721, n27720, n27719,
         n27718, n27717, n27716, n27715, n27714, n27713, n27712, n27711,
         n27710, n27709, n27708, n27707, n27706, n27705, n27704, n27703,
         n27702, n27701, n27700, n27699, n27698, n27697, n27696, n27695,
         n27694, n27693, n27692, n27691, n27690, n27689, n27688, n27687,
         n27686, n27685, n27684, n27683, n27682, n27681, n27680, n27679,
         n27678, n27677, n27676, n27675, n27674, n27673, n27672, n27671,
         n27670, n27669, n27668, n27667, n27666, n27665, n27664, n27663,
         n27662, n27661, n27660, n27659, n27658, n27657, n27656, n27655,
         n27654, n27653, n27652, n27651, n27650, n27649, n27648, n27647,
         n27646, n27645, n27644, n27643, n27642, n27641, n27640, n27639,
         n27638, n27637, n27636, n27635, n27634, n27633, n27632, n27631,
         n27630, n27629, n27628, n27627, n27626, n27625, n27624, n27623,
         n27622, n27621, n27620, n27619, n27618, n27617, n27616, n27615,
         n27614, n27613, n27612, n27611, n27610, n27609, n27608, n27607,
         n27606, n27605, n27604, n27603, n27602, n27601, n27600, n27599,
         n27598, n27597, n27596, n27595, n27594, n27593, n27592, n27591,
         n27590, n27589, n27588, n27587, n27586, n27585, n27584, n27583,
         n27582, n27581, n27580, n27579, n27578, n27577, n27576, n27575,
         n27574, n27573, n27572, n27571, n27570, n27569, n27568, n27567,
         n27566, n27565, n27564, n27563, n27562, n27561, n27560, n27559,
         n27558, n27557, n27556, n27555, n27554, n27553, n27552, n27551,
         n27550, n27549, n27548, n27547, n27546, n27545, n27544, n27543,
         n27542, n27541, n27540, n27539, n27538, n27537, n27536, n27535,
         n27534, n27533, n27532, n27531, n27530, n27529, n27528, n27527,
         n27526, n27525, n27524, n27523, n27522, n27521, n27520, n27519,
         n27518, n27517, n27516, n27515, n27514, n27513, n27512, n27511,
         n27510, n27509, n27508, n27507, n27506, n27505, n27504, n27503,
         n27502, n27501, n27500, n27499, n27498, n27497, n27496, n27495,
         n27494, n27493, n27492, n27491, n27490, n27489, n27488, n27487,
         n27486, n27485, n27484, n27483, n27482, n27481, n27480, n27479,
         n27478, n27477, n27476, n27475, n27474, n27473, n27472, n27471,
         n27470, n27469, n27468, n27467, n27466, n27465, n27464, n27463,
         n27462, n27461, n27460, n27459, n27458, n27457, n27456, n27455,
         n27454, n27453, n27452, n27451, n27450, n27449, n27448, n27447,
         n27446, n27445, n27444, n27443, n27442, n27441, n27440, n27439,
         n27438, n27437, n27436, n27435, n27434, n27433, n27432, n27431,
         n27430, n27429, n27428, n27427, n27426, n27425, n27424, n27423,
         n27422, n27421, n27420, n27419, n27418, n27417, n27416, n27415,
         n27414, n27413, n27412, n27411, n27410, n27409, n27408, n27407,
         n27406, n27405, n27404, n27403, n27402, n27401, n27400, n27399,
         n27398, n27397, n27396, n27395, n27394, n27393, n27392, n27391,
         n27390, n27389, n27388, n27387, n27386, n27385, n27384, n27383,
         n27382, n27381, n27380, n27379, n27378, n27377, n27376, n27375,
         n27374, n27373, n27372, n27371, n27370, n27369, n27368, n27367,
         n27366, n27365, n27364, n27363, n27362, n27361, n27360, n27359,
         n27358, n27357, n27356, n27355, n27354, n27353, n27352, n27351,
         n27350, n27349, n27348, n27347, n27346, n27345, n27344, n27343,
         n27342, n27341, n27340, n27339, n27338, n27337, n27336, n27335,
         n27334, n27333, n27332, n27331, n27330, n27329, n27328, n27327,
         n27326, n27325, n27324, n27323, n27322, n27321, n27320, n27319,
         n27318, n27317, n27316, n27315, n27314, n27313, n27312, n27311,
         n27310, n27309, n27308, n27307, n27306, n27305, n27304, n27303,
         n27302, n27301, n27300, n27299, n27298, n27297, n27296, n27295,
         n27294, n27293, n27292, n27291, n27290, n27289, n27288, n27287,
         n27286, n27285, n27284, n27283, n27282, n27281, n27280, n27279,
         n27278, n27277, n27276, n27275, n27274, n27273, n27272, n27271,
         n27270, n27269, n27268, n27267, n27266, n27265, n27264, n27263,
         n27262, n27261, n27260, n27259, n27258, n27257, n27256, n27255,
         n27254, n27253, n27252, n27251, n27250, n27249, n27248, n27247,
         n27246, n27245, n27244, n27243, n27242, n27241, n27240, n27239,
         n27238, n27237, n27236, n27235, n27234, n27233, n27232, n27231,
         n27230, n27229, n27228, n27227, n27226, n27225, n27224, n27223,
         n27222, n27221, n27220, n27219, n27218, n27217, n27216, n27215,
         n27214, n27213, n27212, n27211, n27210, n27209, n27208, n27207,
         n27206, n27205, n27204, n27203, n27202, n27201, n27200, n27199,
         n27198, n27197, n27196, n27195, n27194, n27193, n27192, n27191,
         n27190, n27189, n27188, n27187, n27186, n27185, n27184, n27183,
         n27182, n27181, n27180, n27179, n27178, n27177, n27176, n27175,
         n27174, n27173, n27172, n27171, n27170, n27169, n27168, n27167,
         n27166, n27165, n27164, n27163, n27162, n27161, n27160, n27159,
         n27158, n27157, n27156, n27155, n27154, n27153, n27152, n27151,
         n27150, n27149, n27148, n27147, n27146, n27145, n27144, n27143,
         n27142, n27141, n27140, n27139, n27138, n27137, n27136, n27135,
         n27134, n27133, n27132, n27131, n27130, n27129, n27128, n27127,
         n27126, n27125, n27124, n27123, n27122, n27121, n27120, n27119,
         n27118, n27117, n27116, n27115, n27114, n27113, n27112, n27111,
         n27110, n27109, n27108, n27107, n27106, n27105, n27104, n27103,
         n27102, n27101, n27100, n27099, n27098, n27097, n27096, n27095,
         n27094, n27093, n27092, n27091, n27090, n27089, n27088, n27087,
         n27086, n27085, n27084, n27083, n27082, n27081, n27080, n27079,
         n27078, n27077, n27076, n27075, n27074, n27073, n27072, n27071,
         n27070, n27069, n27068, n27067, n27066, n27065, n27064, n27063,
         n27062, n27061, n27060, n27059, n27058, n27057, n27056, n27055,
         n27054, n27053, n27052, n27051, n27050, n27049, n27048, n27047,
         n27046, n27045, n27044, n27043, n27042, n27041, n27040, n27039,
         n27038, n27037, n27036, n27035, n27034, n27033, n27032, n27031,
         n27030, n27029, n27028, n27027, n27026, n27025, n27024, n27023,
         n27022, n27021, n27020, n27019, n27018, n27017, n27016, n27015,
         n27014, n27013, n27012, n27011, n27010, n27009, n27008, n27007,
         n27006, n27005, n27004, n27003, n27002, n27001, n27000, n26999,
         n26998, n26997, n26996, n26995, n26994, n26993, n26992, n26991,
         n26990, n26989, n26988, n26987, n26986, n26985, n26984, n26983,
         n26982, n26981, n26980, n26979, n26978, n26977, n26976, n26975,
         n26974, n26973, n26972, n26971, n26970, n26969, n26968, n26967,
         n26966, n26965, n26964, n26963, n26962, n26961, n26960, n26959,
         n26958, n26957, n26956, n26955, n26954, n26953, n26952, n26951,
         n26950, n26949, n26948, n26947, n26946, n26945, n26944, n26943,
         n26942, n26941, n26940, n26939, n26938, n26937, n26936, n26935,
         n26934, n26933, n26932, n26931, n26930, n26929, n26928, n26927,
         n26926, n26925, n26924, n26923, n26922, n26921, n26920, n26919,
         n26918, n26917, n26916, n26915, n26914, n26913, n26912, n26911,
         n26910, n26909, n26908, n26907, n26906, n26905, n26904, n26903,
         n26902, n26901, n26900, n26899, n26898, n26897, n26896, n26895,
         n26894, n26893, n26892, n26891, n26890, n26889, n26888, n26887,
         n26886, n26885, n26884, n26883, n26882, n26881, n26880, n26879,
         n26878, n26877, n26876, n26875, n26874, n26873, n26872, n26871,
         n26870, n26869, n26868, n26867, n26866, n26865, n26864, n26863,
         n26862, n26861, n26860, n26859, n26858, n26857, n26856, n26855,
         n26854, n26853, n26852, n26851, n26850, n26849, n26848, n26847,
         n26846, n26845, n26844, n26843, n26842, n26841, n26840, n26839,
         n26838, n26837, n26836, n26835, n26834, n26833, n26832, n26831,
         n26830, n26829, n26828, n26827, n26826, n26825, n26824, n26823,
         n26822, n26821, n26820, n26819, n26818, n26817, n26816, n26815,
         n26814, n26813, n26812, n26811, n26810, n26809, n26808, n26807,
         n26806, n26805, n26804, n26803, n26802, n26801, n26800, n26799,
         n26798, n26797, n26796, n26795, n26794, n26793, n26792, n26791,
         n26790, n26789, n26788, n26787, n26786, n26785, n26784, n26783,
         n26782, n26781, n26780, n26779, n26778, n26777, n26776, n26775,
         n26774, n26773, n26772, n26771, n26770, n26769, n26768, n26767,
         n26766, n26765, n26764, n26763, n26762, n26761, n26760, n26759,
         n26758, n26757, n26756, n26755, n26754, n26753, n26752, n26751,
         n26750, n26749, n26748, n26747, n26746, n26745, n26744, n26743,
         n26742, n26741, n26740, n26739, n26738, n26737, n26736, n26735,
         n26734, n26733, n26732, n26731, n26730, n26729, n26728, n26727,
         n26726, n26725, n26724, n26723, n26722, n26721, n26720, n26719,
         n26718, n26717, n26716, n26715, n26714, n26713, n26712, n26711,
         n26710, n26709, n26708, n26707, n26706, n26705, n26704, n26703,
         n26702, n26701, n26700, n26699, n26698, n26697, n26696, n26695,
         n26694, n26693, n26692, n26691, n26690, n26689, n26688, n26687,
         n26686, n26685, n26684, n26683, n26682, n26681, n26680, n26679,
         n26678, n26677, n26676, n26675, n26674, n26673, n26672, n26671,
         n26670, n26669, n26668, n26667, n26666, n26665, n26664, n26663,
         n26662, n26661, n26660, n26659, n26658, n26657, n26656, n26655,
         n26654, n26653, n26652, n26651, n26650, n26649, n26648, n26647,
         n26646, n26645, n26644, n26643, n26642, n26641, n26640, n26639,
         n26638, n26637, n26636, n26635, n26634, n26633, n26632, n26631,
         n26630, n26629, n26628, n26627, n26626, n26625, n26624, n26623,
         n26622, n26621, n26620, n26619, n26618, n26617, n26616, n26615,
         n26614, n26613, n26612, n26611, n26610, n26609, n26608, n26607,
         n26606, n26605, n26604, n26603, n26602, n26601, n26600, n26599,
         n26598, n26597, n26596, n26595, n26594, n26593, n26592, n26591,
         n26590, n26589, n26588, n26587, n26586, n26585, n26584, n26583,
         n26582, n26581, n26580, n26579, n26578, n26577, n26576, n26575,
         n26574, n26573, n26572, n26571, n26570, n26569, n26568, n26567,
         n26566, n26565, n26564, n26563, n26562, n26561, n26560, n26559,
         n26558, n26557, n26556, n26555, n26554, n26553, n26552, n26551,
         n26550, n26549, n26548, n26547, n26546, n26545, n26544, n26543,
         n26542, n26541, n26540, n26539, n26538, n26537, n26536, n26535,
         n26534, n26533, n26532, n26531, n26530, n26529, n26528, n26527,
         n26526, n26525, n26524, n26523, n26522, n26521, n26520, n26519,
         n26518, n26517, n26516, n26515, n26514, n26513, n26512, n26511,
         n26510, n26509, n26508, n26507, n26506, n26505, n26504, n26503,
         n26502, n26501, n26500, n26499, n26498, n26497, n26496, n26495,
         n26494, n26493, n26492, n26491, n26490, n26489, n26488, n26487,
         n26486, n26485, n26484, n26483, n26482, n26481, n26480, n26479,
         n26478, n26477, n26476, n26475, n26474, n26473, n26472, n26471,
         n26470, n26469, n26468, n26467, n26466, n26465, n26464, n26463,
         n26462, n26461, n26460, n26459, n26458, n26457, n26456, n26455,
         n26454, n26453, n26452, n26451, n26450, n26449, n26448, n26447,
         n26446, n26445, n26444, n26443, n26442, n26441, n26440, n26439,
         n26438, n26437, n26436, n26435, n26434, n26433, n26432, n26431,
         n26430, n26429, n26428, n26427, n26426, n26425, n26424, n26423,
         n26422, n26421, n26420, n26419, n26418, n26417, n26416, n26415,
         n26414, n26413, n26412, n26411, n26410, n26409, n26408, n26407,
         n26406, n26405, n26404, n26403, n26402, n26401, n26400, n26399,
         n26398, n26397, n26396, n26395, n26394, n26393, n26392, n26391,
         n26390, n26389, n26388, n26387, n26386, n26385, n26384, n26383,
         n26382, n26381, n26380, n26379, n26378, n26377, n26376, n26375,
         n26374, n26373, n26372, n26371, n26370, n26369, n26368, n26367,
         n26366, n26365, n26364, n26363, n26362, n26361, n26360, n26359,
         n26358, n26357, n26356, n26355, n26354, n26353, n26352, n26351,
         n26350, n26349, n26348, n26347, n26346, n26345, n26344, n26343,
         n26342, n26341, n26340, n26339, n26338, n26337, n26336, n26335,
         n26334, n26333, n26332, n26331, n26330, n26329, n26328, n26327,
         n26326, n26325, n26324, n26323, n26322, n26321, n26320, n26319,
         n26318, n26317, n26316, n26315, n26314, n26313, n26312, n26311,
         n26310, n26309, n26308, n26307, n26306, n26305, n26304, n26303,
         n26302, n26301, n26300, n26299, n26298, n26297, n26296, n26295,
         n26294, n26293, n26292, n26291, n26290, n26289, n26288, n26287,
         n26286, n26285, n26284, n26283, n26282, n26281, n26280, n26279,
         n26278, n26277, n26276, n26275, n26274, n26273, n26272, n26271,
         n26270, n26269, n26268, n26267, n26266, n26265, n26264, n26263,
         n26262, n26261, n26260, n26259, n26258, n26257, n26256, n26255,
         n26254, n26253, n26252, n26251, n26250, n26249, n26248, n26247,
         n26246, n26245, n26244, n26243, n26242, n26241, n26240, n26239,
         n26238, n26237, n26236, n26235, n26234, n26233, n26232, n26231,
         n26230, n26229, n26228, n26227, n26226, n26225, n26224, n26223,
         n26222, n26221, n26220, n26219, n26218, n26217, n26216, n26215,
         n26214, n26213, n26212, n26211, n26210, n26209, n26208, n26207,
         n26206, n26205, n26204, n26203, n26202, n26201, n26200, n26199,
         n26198, n26197, n26196, n26195, n26194, n26193, n26192, n26191,
         n26190, n26189, n26188, n26187, n26186, n26185, n26184, n26183,
         n26182, n26181, n26180, n26179, n26178, n26177, n26176, n26175,
         n26174, n26173, n26172, n26171, n26170, n26169, n26168, n26167,
         n26166, n26165, n26164, n26163, n26162, n26161, n26160, n26159,
         n26158, n26157, n26156, n26155, n26154, n26153, n26152, n26151,
         n26150, n26149, n26148, n26147, n26146, n26145, n26144, n26143,
         n26142, n26141, n26140, n26139, n26138, n26137, n26136, n26135,
         n26134, n26133, n26132, n26131, n26130, n26129, n26128, n26127,
         n26126, n26125, n26124, n26123, n26122, n26121, n26120, n26119,
         n26118, n26117, n26116, n26115, n26114, n26113, n26112, n26111,
         n26110, n26109, n26108, n26107, n26106, n26105, n26104, n26103,
         n26102, n26101, n26100, n26099, n26098, n26097, n26096, n26095,
         n26094, n26093, n26092, n26091, n26090, n26089, n26088, n26087,
         n26086, n26085, n26084, n26083, n26082, n26081, n26080, n26079,
         n26078, n26077, n26076, n26075, n26074, n26073, n26072, n26071,
         n26070, n26069, n26068, n26067, n26066, n26065, n26064, n26063,
         n26062, n26061, n26060, n26059, n26058, n26057, n26056, n26055,
         n26054, n26053, n26052, n26051, n26050, n26049, n26048, n26047,
         n26046, n26045, n26044, n26043, n26042, n26041, n26040, n26039,
         n26038, n26037, n26036, n26035, n26034, n26033, n26032, n26031,
         n26030, n26029, n26028, n26027, n26026, n26025, n26024, n26023,
         n26022, n26021, n26020, n26019, n26018, n26017, n26016, n26015,
         n26014, n26013, n26012, n26011, n26010, n26009, n26008, n26007,
         n26006, n26005, n26004, n26003, n26002, n26001, n26000, n25999,
         n25998, n25997, n25996, n25995, n25994, n25993, n25992, n25991,
         n25990, n25989, n25988, n25987, n25986, n25985, n25984, n25983,
         n25982, n25981, n25980, n25979, n25978, n25977, n25976, n25975,
         n25974, n25973, n25972, n25971, n25970, n25969, n25968, n25967,
         n25966, n25965, n25964, n25963, n25962, n25961, n25960, n25959,
         n25958, n25957, n25956, n25955, n25954, n25953, n25952, n25951,
         n25950, n25949, n25948, n25947, n25946, n25945, n25944, n25943,
         n25942, n25941, n25940, n25939, n25938, n25937, n25936, n25935,
         n25934, n25933, n25932, n25931, n25930, n25929, n25928, n25927,
         n25926, n25925, n25924, n25923, n25922, n25921, n25920, n25919,
         n25918, n25917, n25916, n25915, n25914, n25913, n25912, n25911,
         n25910, n25909, n25908, n25907, n25906, n25905, n25904, n25903,
         n25902, n25901, n25900, n25899, n25898, n25897, n25896, n25895,
         n25894, n25893, n25892, n25891, n25890, n25889, n25888, n25887,
         n25886, n25885, n25884, n25883, n25882, n25881, n25880, n25879,
         n25878, n25877, n25876, n25875, n25874, n25873, n25872, n25871,
         n25870, n25869, n25868, n25867, n25866, n25865, n25864, n25863,
         n25862, n25861, n25860, n25859, n25858, n25857, n25856, n25855,
         n25854, n25853, n25852, n25851, n25850, n25849, n25848, n25847,
         n25846, n25845, n25844, n25843, n25842, n25841, n25840, n25839,
         n25838, n25837, n25836, n25835, n25834, n25833, n25832, n25831,
         n25830, n25829, n25828, n25827, n25826, n25825, n25824, n25823,
         n25822, n25821, n25820, n25819, n25818, n25817, n25816, n25815,
         n25814, n25813, n25812, n25811, n25810, n25809, n25808, n25807,
         n25806, n25805, n25804, n25803, n25802, n25801, n25800, n25799,
         n25798, n25797, n25796, n25795, n25794, n25793, n25792, n25791,
         n25790, n25789, n25788, n25787, n25786, n25785, n25784, n25783,
         n25782, n25781, n25780, n25779, n25778, n25777, n25776, n25775,
         n25774, n25773, n25772, n25771, n25770, n25769, n25768, n25767,
         n25766, n25765, n25764, n25763, n25762, n25761, n25760, n25759,
         n25758, n25757, n25756, n25755, n25754, n25753, n25752, n25751,
         n25750, n25749, n25748, n25747, n25746, n25745, n25744, n25743,
         n25742, n25741, n25740, n25739, n25738, n25737, n25736, n25735,
         n25734, n25733, n25732, n25731, n25730, n25729, n25728, n25727,
         n25726, n25725, n25724, n25723, n25722, n25721, n25720, n25719,
         n25718, n25717, n25716, n25715, n25714, n25713, n25712, n25711,
         n25710, n25709, n25708, n25707, n25706, n25705, n25704, n25703,
         n25702, n25701, n25700, n25699, n25698, n25697, n25696, n25695,
         n25694, n25693, n25692, n25691, n25690, n25689, n25688, n25687,
         n25686, n25685, n25684, n25683, n25682, n25681, n25680, n25679,
         n25678, n25677, n25676, n25675, n25674, n25673, n25672, n25671,
         n25670, n25669, n25668, n25667, n25666, n25665, n25664, n25663,
         n25662, n25661, n25660, n25659, n25658, n25657, n25656, n25655,
         n25654, n25653, n25652, n25651, n25650, n25649, n25648, n25647,
         n25646, n25645, n25644, n25643, n25642, n25641, n25640, n25639,
         n25638, n25637, n25636, n25635, n25634, n25633, n25632, n25631,
         n25630, n25629, n25628, n25627, n25626, n25625, n25624, n25623,
         n25622, n25621, n25620, n25619, n25618, n25617, n25616, n25615,
         n25614, n25613, n25612, n25611, n25610, n25609, n25608, n25607,
         n25606, n25605, n25604, n25603, n25602, n25601, n25600, n25599,
         n25598, n25597, n25596, n25595, n25594, n25593, n25592, n25591,
         n25590, n25589, n25588, n25587, n25586, n25585, n25584, n25583,
         n25582, n25581, n25580, n25579, n25578, n25577, n25576, n25575,
         n25574, n25573, n25572, n25571, n25570, n25569, n25568, n25567,
         n25566, n25565, n25564, n25563, n25562, n25561, n25560, n25559,
         n25558, n25557, n25556, n25555, n25554, n25553, n25552, n25551,
         n25550, n25549, n25548, n25547, n25546, n25545, n25544, n25543,
         n25542, n25541, n25540, n25539, n25538, n25537, n25536, n25535,
         n25534, n25533, n25532, n25531, n25530, n25529, n25528, n25527,
         n25526, n25525, n25524, n25523, n25522, n25521, n25520, n25519,
         n25518, n25517, n25516, n25515, n25514, n25513, n25512, n25511,
         n25510, n25509, n25508, n25507, n25506, n25505, n25504, n25503,
         n25502, n25501, n25500, n25499, n25498, n25497, n25496, n25495,
         n25494, n25493, n25492, n25491, n25490, n25489, n25488, n25487,
         n25486, n25485, n25484, n25483, n25482, n25481, n25480, n25479,
         n25478, n25477, n25476, n25475, n25474, n25473, n25472, n25471,
         n25470, n25469, n25468, n25467, n25466, n25465, n25464, n25463,
         n25462, n25461, n25460, n25459, n25458, n25457, n25456, n25455,
         n25454, n25453, n25452, n25451, n25450, n25449, n25448, n25447,
         n25446, n25445, n25444, n25443, n25442, n25441, n25440, n25439,
         n25438, n25437, n25436, n25435, n25434, n25433, n25432, n25431,
         n25430, n25429, n25428, n25427, n25426, n25425, n25424, n25423,
         n25422, n25421, n25420, n25419, n25418, n25417, n25416, n25415,
         n25414, n25413, n25412, n25411, n25410, n25409, n25408, n25407,
         n25406, n25405, n25404, n25403, n25402, n25401, n25400, n25399,
         n25398, n25397, n25396, n25395, n25394, n25393, n25392, n25391,
         n25390, n25389, n25388, n25387, n25386, n25385, n25384, n25383,
         n25382, n25381, n25380, n25379, n25378, n25377, n25376, n25375,
         n25374, n25373, n25372, n25371, n25370, n25369, n25368, n25367,
         n25366, n25365, n25364, n25363, n25362, n25361, n25360, n25359,
         n25358, n25357, n25356, n25355, n25354, n25353, n25352, n25351,
         n25350, n25349, n25348, n25347, n25346, n25345, n25344, n25343,
         n25342, n25341, n25340, n25339, n25338, n25337, n25336, n25335,
         n25334, n25333, n25332, n25331, n25330, n25329, n25328, n25327,
         n25326, n25325, n25324, n25323, n25322, n25321, n25320, n25319,
         n25318, n25317, n25316, n25315, n25314, n25313, n25312, n25311,
         n25310, n25309, n25308, n25307, n25306, n25305, n25304, n25303,
         n25302, n25301, n25300, n25299, n25298, n25297, n25296, n25295,
         n25294, n25293, n25292, n25291, n25290, n25289, n25288, n25287,
         n25286, n25285, n25284, n25283, n25282, n25281, n25280, n25279,
         n25278, n25277, n25276, n25275, n25274, n25273, n25272, n25271,
         n25270, n25269, n25268, n25267, n25266, n25265, n25264, n25263,
         n25262, n25261, n25260, n25259, n25258, n25257, n25256, n25255,
         n25254, n25253, n25252, n25251, n25250, n25249, n25248, n25247,
         n25246, n25245, n25244, n25243, n25242, n25241, n25240, n25239,
         n25238, n25237, n25236, n25235, n25234, n25233, n25232, n25231,
         n25230, n25229, n25228, n25227, n25226, n25225, n25224, n25223,
         n25222, n25221, n25220, n25219, n25218, n25217, n25216, n25215,
         n25214, n25213, n25212, n25211, n25210, n25209, n25208, n25207,
         n25206, n25205, n25204, n25203, n25202, n25201, n25200, n25199,
         n25198, n25197, n25196, n25195, n25194, n25193, n25192, n25191,
         n25190, n25189, n25188, n25187, n25186, n25185, n25184, n25183,
         n25182, n25181, n25180, n25179, n25178, n25177, n25176, n25175,
         n25174, n25173, n25172, n25171, n25170, n25169, n25168, n25167,
         n25166, n25165, n25164, n25163, n25162, n25161, n25160, n25159,
         n25158, n25157, n25156, n25155, n25154, n25153, n25152, n25151,
         n25150, n25149, n25148, n25147, n25146, n25145, n25144, n25143,
         n25142, n25141, n25140, n25139, n25138, n25137, n25136, n25135,
         n25134, n25133, n25132, n25131, n25130, n25129, n25128, n25127,
         n25126, n25125, n25124, n25123, n25122, n25121, n25120, n25119,
         n25118, n25117, n25116, n25115, n25114, n25113, n25112, n25111,
         n25110, n25109, n25108, n25107, n25106, n25105, n25104, n25103,
         n25102, n25101, n25100, n25099, n25098, n25097, n25096, n25095,
         n25094, n25093, n25092, n25091, n25090, n25089, n25088, n25087,
         n25086, n25085, n25084, n25083, n25082, n25081, n25080, n25079,
         n25078, n25077, n25076, n25075, n25074, n25073, n25072, n25071,
         n25070, n25069, n25068, n25067, n25066, n25065, n25064, n25063,
         n25062, n25061, n25060, n25059, n25058, n25057, n25056, n25055,
         n25054, n25053, n25052, n25051, n25050, n25049, n25048, n25047,
         n25046, n25045, n25044, n25043, n25042, n25041, n25040, n25039,
         n25038, n25037, n25036, n25035, n25034, n25033, n25032, n25031,
         n25030, n25029, n25028, n25027, n25026, n25025, n25024, n25023,
         n25022, n25021, n25020, n25019, n25018, n25017, n25016, n25015,
         n25014, n25013, n25012, n25011, n25010, n25009, n25008, n25007,
         n25006, n25005, n25004, n25003, n25002, n25001, n25000, n24999,
         n24998, n24997, n24996, n24995, n24994, n24993, n24992, n24991,
         n24990, n24989, n24988, n24987, n24986, n24985, n24984, n24983,
         n24982, n24981, n24980, n24979, n24978, n24977, n24976, n24975,
         n24974, n24973, n24972, n24971, n24970, n24969, n24968, n24967,
         n24966, n24965, n24964, n24963, n24962, n24961, n24960, n24959,
         n24958, n24957, n24956, n24955, n24954, n24953, n24952, n24951,
         n24950, n24949, n24948, n24947, n24946, n24945, n24944, n24943,
         n24942, n24941, n24940, n24939, n24938, n24937, n24936, n24935,
         n24934, n24933, n24932, n24931, n24930, n24929, n24928, n24927,
         n24926, n24925, n24924, n24923, n24922, n24921, n24920, n24919,
         n24918, n24917, n24916, n24915, n24914, n24913, n24912, n24911,
         n24910, n24909, n24908, n24907, n24906, n24905, n24904, n24903,
         n24902, n24901, n24900, n24899, n24898, n24897, n24896, n24895,
         n24894, n24893, n24892, n24891, n24890, n24889, n24888, n24887,
         n24886, n24885, n24884, n24883, n24882, n24881, n24880, n24879,
         n24878, n24877, n24876, n24875, n24874, n24873, n24872, n24871,
         n24870, n24869, n24868, n24867, n24866, n24865, n24864, n24863,
         n24862, n24861, n24860, n24859, n24858, n24857, n24856, n24855,
         n24854, n24853, n24852, n24851, n24850, n24849, n24848, n24847,
         n24846, n24845, n24844, n24843, n24842, n24841, n24840, n24839,
         n24838, n24837, n24836, n24835, n24834, n24833, n24832, n24831,
         n24830, n24829, n24828, n24827, n24826, n24825, n24824, n24823,
         n24822, n24821, n24820, n24819, n24818, n24817, n24816, n24815,
         n24814, n24813, n24812, n24811, n24810, n24809, n24808, n24807,
         n24806, n24805, n24804, n24803, n24802, n24801, n24800, n24799,
         n24798, n24797, n24796, n24795, n24794, n24793, n24792, n24791,
         n24790, n24789, n24788, n24787, n24786, n24785, n24784, n24783,
         n24782, n24781, n24780, n24779, n24778, n24777, n24776, n24775,
         n24774, n24773, n24772, n24771, n24770, n24769, n24768, n24767,
         n24766, n24765, n24764, n24763, n24762, n24761, n24760, n24759,
         n24758, n24757, n24756, n24755, n24754, n24753, n24752, n24751,
         n24750, n24749, n24748, n24747, n24746, n24745, n24744, n24743,
         n24742, n24741, n24740, n24739, n24738, n24737, n24736, n24735,
         n24734, n24733, n24732, n24731, n24730, n24729, n24728, n24727,
         n24726, n24725, n24724, n24723, n24722, n24721, n24720, n24719,
         n24718, n24717, n24716, n24715, n24714, n24713, n24712, n24711,
         n24710, n24709, n24708, n24707, n24706, n24705, n24704, n24703,
         n24702, n24701, n24700, n24699, n24698, n24697, n24696, n24695,
         n24694, n24693, n24692, n24691, n24690, n24689, n24688, n24687,
         n24686, n24685, n24684, n24683, n24682, n24681, n24680, n24679,
         n24678, n24677, n24676, n24675, n24674, n24673, n24672, n24671,
         n24670, n24669, n24668, n24667, n24666, n24665, n24664, n24663,
         n24662, n24661, n24660, n24659, n24658, n24657, n24656, n24655,
         n24654, n24653, n24652, n24651, n24650, n24649, n24648, n24647,
         n24646, n24645, n24644, n24643, n24642, n24641, n24640, n24639,
         n24638, n24637, n24636, n24635, n24634, n24633, n24632, n24631,
         n24630, n24629, n24628, n24627, n24626, n24625, n24624, n24623,
         n24622, n24621, n24620, n24619, n24618, n24617, n24616, n24615,
         n24614, n24613, n24612, n24611, n24610, n24609, n24608, n24607,
         n24606, n24605, n24604, n24603, n24602, n24601, n24600, n24599,
         n24598, n24597, n24596, n24595, n24594, n24593, n24592, n24591,
         n24590, n24589, n24588, n24587, n24586, n24585, n24584, n24583,
         n24582, n24581, n24580, n24579, n24578, n24577, n24576, n24575,
         n24574, n24573, n24572, n24571, n24570, n24569, n24568, n24567,
         n24566, n24565, n24564, n24563, n24562, n24561, n24560, n24559,
         n24558, n24557, n24556, n24555, n24554, n24553, n24552, n24551,
         n24550, n24549, n24548, n24547, n24546, n24545, n24544, n24543,
         n24542, n24541, n24540, n24539, n24538, n24537, n24536, n24535,
         n24534, n24533, n24532, n24531, n24530, n24529, n24528, n24527,
         n24526, n24525, n24524, n24523, n24522, n24521, n24520, n24519,
         n24518, n24517, n24516, n24515, n24514, n24513, n24512, n24511,
         n24510, n24509, n24508, n24507, n24506, n24505, n24504, n24503,
         n24502, n24501, n24500, n24499, n24498, n24497, n24496, n24495,
         n24494, n24493, n24492, n24491, n24490, n24489, n24488, n24487,
         n24486, n24485, n24484, n24483, n24482, n24481, n24480, n24479,
         n24478, n24477, n24476, n24475, n24474, n24473, n24472, n24471,
         n24470, n24469, n24468, n24467, n24466, n24465, n24464, n24463,
         n24462, n24461, n24460, n24459, n24458, n24457, n24456, n24455,
         n24454, n24453, n24452, n24451, n24450, n24449, n24448, n24447,
         n24446, n24445, n24444, n24443, n24442, n24441, n24440, n24439,
         n24438, n24437, n24436, n24435, n24434, n24433, n24432, n24431,
         n24430, n24429, n24428, n24427, n24426, n24425, n24424, n24423,
         n24422, n24421, n24420, n24419, n24418, n24417, n24416, n24415,
         n24414, n24413, n24412, n24411, n24410, n24409, n24408, n24407,
         n24406, n24405, n24404, n24403, n24402, n24401, n24400, n24399,
         n24398, n24397, n24396, n24395, n24394, n24393, n24392, n24391,
         n24390, n24389, n24388, n24387, n24386, n24385, n24384, n24383,
         n24382, n24381, n24380, n24379, n24378, n24377, n24376, n24375,
         n24374, n24373, n24372, n24371, n24370, n24369, n24368, n24367,
         n24366, n24365, n24364, n24363, n24362, n24361, n24360, n24359,
         n24358, n24357, n24356, n24355, n24354, n24353, n24352, n24351,
         n24350, n24349, n24348, n24347, n24346, n24345, n24344, n24343,
         n24342, n24341, n24340, n24339, n24338, n24337, n24336, n24335,
         n24334, n24333, n24332, n24331, n24329, n24328, n24327, n24326,
         n24325, n24324, n24323, n24322, n24321, n24320, n24319, n24318,
         n24317, n24316, n24315, n24314, n24313, n24312, n24311, n24310,
         n24309, n24308, n24307, n24306, n24305, n24304, n24303, n24302,
         n24301, n24300, n24299, n24298, n24297, n24296, n24295, n24294,
         n24293, n24292, n24291, n24290, n24289, n24288, n24287, n24286,
         n24285, n24284, n24283, n24282, n24281, n24280, n24279, n24278,
         n24277, n24276, n24275, n24274, n24273, n24272, n24271, n24270,
         n24269, n24268, n24267, n24266, n24265, n24264, n24263, n24262,
         n24261, n24260, n24259, n24258, n24257, n24256, n24255, n24254,
         n24253, n24252, n24251, n24250, n24249, n24248, n24247, n24246,
         n24245, n24244, n24243, n24242, n24241, n24240, n24239, n24238,
         n24237, n24236, n24235, n24234, n24233, n24232, n24231, n24230,
         n24229, n24228, n24227, n24226, n24225, n24224, n24223, n24222,
         n24221, n24220, n24219, n24218, n24217, n24216, n24215, n24214,
         n24213, n24212, n24211, n24210, n24209, n24208, n24207, n24206,
         n24205, n24204, n24203, n24202, n24201, n24200, n24199, n24198,
         n24197, n24196, n24195, n24194, n24193, n24192, n24191, n24190,
         n24189, n24188, n24187, n24186, n24185, n24184, n24183, n24182,
         n24181, n24180, n24179, n24178, n24177, n24176, n24175, n24174,
         n24173, n24172, n24171, n24170, n24169, n24168, n24167, n24166,
         n24165, n24164, n24163, n24162, n24161, n24160, n24159, n24158,
         n24157, n24156, n24155, n24154, n24153, n24152, n24151, n24150,
         n24149, n24148, n24147, n24146, n24145, n24144, n24143, n24142,
         n24141, n24140, n24139, n24138, n24137, n24136, n24135, n24134,
         n24133, n24132, n24131, n24130, n24129, n24128, n24127, n24126,
         n24125, n24124, n24123, n24122, n24121, n24120, n24119, n24118,
         n24117, n24116, n24115, n24114, n24113, n24112, n24111, n24110,
         n24109, n24108, n24107, n24106, n24105, n24104, n24103, n24102,
         n24101, n24100, n24099, n24098, n24097, n24096, n24095, n24094,
         n24093, n24092, n24091, n24090, n24089, n24088, n24087, n24086,
         n24085, n24084, n24083, n24082, n24081, n24080, n24079, n24078,
         n24077, n24076, n24075, n24074, n24073, n24072, n24071, n24070,
         n24069, n24068, n24067, n24066, n24065, n24064, n24063, n24062,
         n24061, n24060, n24059, n24058, n24057, n24056, n24055, n24054,
         n24053, n24052, n24051, n24050, n24049, n24048, n24047, n24046,
         n24045, n24044, n24043, n24042, n24041, n24040, n24039, n24038,
         n24037, n24036, n24035, n24034, n24033, n24032, n24031, n24030,
         n24029, n24028, n24027, n24026, n24025, n24024, n24023, n24022,
         n24021, n24020, n24019, n24018, n24017, n24016, n24015, n24014,
         n24013, n24012, n24011, n24010, n24009, n24008, n24007, n24006,
         n24005, n24004, n24003, n24002, n24001, n24000, n23999, n23998,
         n23997, n23996, n23995, n23994, n23993, n23992, n23991, n23990,
         n23989, n23988, n23987, n23986, n23985, n23984, n23983, n23982,
         n23981, n23980, n23979, n23978, n23977, n23976, n23975, n23974,
         n23973, n23972, n23971, n23970, n23969, n23968, n23967, n23966,
         n23965, n23964, n23963, n23962, n23961, n23960, n23959, n23958,
         n23957, n23956, n23955, n23954, n23953, n23952, n23951, n23950,
         n23949, n23948, n23947, n23946, n23945, n23944, n23943, n23942,
         n23941, n23940, n23939, n23938, n23937, n23936, n23935, n23934,
         n23933, n23932, n23931, n23930, n23929, n23928, n23927, n23926,
         n23925, n23924, n23923, n23922, n23921, n23920, n23919, n23918,
         n23917, n23916, n23915, n23914, n23913, n23912, n23911, n23910,
         n23909, n23908, n23907, n23906, n23905, n23904, n23903, n23902,
         n23901, n23900, n23899, n23898, n23897, n23896, n23895, n23894,
         n23893, n23892, n23891, n23890, n23889, n23888, n23887, n23886,
         n23885, n23884, n23883, n23882, n23881, n23880, n23879, n23878,
         n23877, n23876, n23875, n23874, n23873, n23872, n23871, n23870,
         n23869, n23868, n23867, n23866, n23865, n23864, n23863, n23862,
         n23861, n23860, n23859, n23858, n23857, n23856, n23855, n23854,
         n23853, n23852, n23851, n23850, n23849, n23848, n23847, n23846,
         n23845, n23844, n23843, n23842, n23841, n23840, n23839, n23838,
         n23837, n23836, n23835, n23834, n23833, n23832, n23831, n23830,
         n23829, n23828, n23827, n23826, n23825, n23824, n23823, n23822,
         n23821, n23820, n23819, n23818, n23817, n23816, n23815, n23814,
         n23813, n23812, n23811, n23810, n23809, n23808, n23807, n23806,
         n23805, n23804, n23803, n23802, n23801, n23800, n23799, n23798,
         n23797, n23796, n23795, n23794, n23793, n23792, n23791, n23790,
         n23789, n23788, n23787, n23786, n23785, n23784, n23783, n23782,
         n23781, n23780, n23779, n23778, n23777, n23776, n23775, n23774,
         n23773, n23772, n23771, n23770, n23769, n23768, n23767, n23766,
         n23765, n23764, n23763, n23762, n23761, n23760, n23759, n23758,
         n23757, n23756, n23755, n23754, n23753, n23752, n23751, n23750,
         n23749, n23748, n23747, n23746, n23745, n23744, n23743, n23742,
         n23741, n23740, n23739, n23738, n23737, n23736, n23735, n23734,
         n23733, n23732, n23731, n23730, n23729, n23728, n23727, n23726,
         n23725, n23724, n23723, n23722, n23721, n23720, n23719, n23718,
         n23717, n23716, n23715, n23714, n23713, n23712, n23711, n23710,
         n23709, n23708, n23707, n23706, n23705, n23704, n23703, n23702,
         n23701, n23700, n23699, n23698, n23697, n23696, n23695, n23694,
         n23693, n23692, n23691, n23690, n23689, n23688, n23687, n23686,
         n23685, n23684, n23683, n23682, n23681, n23680, n23679, n23678,
         n23677, n23676, n23675, n23674, n23673, n23672, n23671, n23670,
         n23669, n23668, n23667, n23666, n23665, n23664, n23663, n23662,
         n23661, n23660, n23659, n23658, n23657, n23656, n23655, n23654,
         n23653, n23652, n23651, n23650, n23649, n23648, n23647, n23646,
         n23645, n23644, n23643, n23642, n23641, n23640, n23639, n23638,
         n23637, n23636, n23635, n23634, n23633, n23632, n23631, n23630,
         n23629, n23628, n23627, n23626, n23625, n23624, n23623, n23622,
         n23621, n23620, n23619, n23618, n23617, n23616, n23615, n23614,
         n23613, n23612, n23611, n23610, n23609, n23608, n23607, n23606,
         n23605, n23604, n23603, n23602, n23601, n23600, n23599, n23598,
         n23597, n23596, n23595, n23594, n23593, n23592, n23591, n23590,
         n23589, n23588, n23587, n23586, n23585, n23584, n23583, n23582,
         n23581, n23580, n23579, n23578, n23577, n23576, n23575, n23574,
         n23573, n23572, n23571, n23570, n23569, n23568, n23567, n23566,
         n23565, n23564, n23563, n23562, n23561, n23560, n23559, n23558,
         n23557, n23556, n23555, n23554, n23553, n23552, n23551, n23550,
         n23549, n23548, n23547, n23546, n23545, n23544, n23543, n23542,
         n23541, n23540, n23539, n23538, n23537, n23536, n23535, n23534,
         n23533, n23532, n23531, n23530, n23529, n23528, n23527, n23526,
         n23525, n23524, n23523, n23522, n23521, n23520, n23519, n23518,
         n23517, n23516, n23515, n23514, n23513, n23512, n23511, n23510,
         n23509, n23508, n23507, n23506, n23505, n23504, n23503, n23502,
         n23501, n23500, n23499, n23498, n23497, n23496, n23495, n23494,
         n23493, n23492, n23491, n23490, n23489, n23488, n23487, n23486,
         n23485, n23484, n23483, n23482, n23481, n23480, n23479, n23478,
         n23477, n23476, n23475, n23474, n23473, n23472, n23471, n23470,
         n23469, n23468, n23467, n23466, n23465, n23464, n23463, n23462,
         n23461, n23460, n23459, n23458, n23457, n23456, n23455, n23454,
         n23453, n23452, n23451, n23450, n23449, n23448, n23447, n23446,
         n23445, n23444, n23443, n23442, n23441, n23440, n23439, n23438,
         n23437, n23436, n23435, n23434, n23433, n23432, n23431, n23430,
         n23429, n23428, n23427, n23426, n23425, n23424, n23423, n23422,
         n23421, n23420, n23419, n23418, n23417, n23416, n23415, n23414,
         n23413, n23412, n23411, n23410, n23409, n23408, n23407, n23406,
         n23405, n23404, n23403, n23402, n23401, n23400, n23399, n23398,
         n23397, n23396, n23395, n23394, n23393, n23392, n23391, n23390,
         n23389, n23388, n23387, n23386, n23385, n23384, n23383, n23382,
         n23381, n23380, n23379, n23378, n23377, n23376, n23375, n23374,
         n23373, n23372, n23371, n23370, n23369, n23368, n23367, n23366,
         n23365, n23364, n23363, n23362, n23361, n23360, n23359, n23358,
         n23357, n23356, n23355, n23354, n23353, n23352, n23351, n23350,
         n23349, n23348, n23347, n23346, n23345, n23344, n23343, n23342,
         n23341, n23340, n23339, n23338, n23337, n23336, n23335, n23334,
         n23333, n23332, n23331, n23330, n23329, n23328, n23327, n23326,
         n23325, n23324, n23323, n23322, n23321, n23320, n23319, n23318,
         n23317, n23316, n23315, n23314, n23313, n23312, n23311, n23310,
         n23309, n23308, n23307, n23306, n23305, n23304, n23303, n23302,
         n23301, n23300, n23299, n23298, n23297, n23296, n23295, n23294,
         n23293, n23292, n23291, n23290, n23289, n23288, n23287, n23286,
         n23285, n23284, n23283, n23282, n23281, n23280, n23279, n23278,
         n23277, n23276, n23275, n23274, n23273, n23272, n23271, n23270,
         n23269, n23268, n23267, n23266, n23265, n23264, n23263, n23262,
         n23261, n23260, n23259, n23258, n23257, n23256, n23255, n23254,
         n23253, n23252, n23251, n23250, n23249, n23248, n23247, n23246,
         n23245, n23244, n23243, n23242, n23241, n23240, n23239, n23238,
         n23237, n23236, n23235, n23234, n23233, n23232, n23231, n23230,
         n23229, n23228, n23227, n23226, n23225, n23224, n23223, n23222,
         n23221, n23220, n23219, n23218, n23217, n23216, n23215, n23214,
         n23213, n23212, n23211, n23210, n23209, n23208, n23207, n23206,
         n23205, n23204, n23203, n23202, n23201, n23200, n23199, n23198,
         n23197, n23196, n23195, n23194, n23193, n23192, n23191, n23190,
         n23189, n23188, n23187, n23186, n23185, n23184, n23183, n23182,
         n23181, n23180, n23179, n23178, n23177, n23176, n23175, n23174,
         n23173, n23172, n23171, n23170, n23169, n23168, n23167, n23166,
         n23165, n23164, n23163, n23162, n23161, n23160, n23159, n23158,
         n23157, n23156, n23155, n23154, n23153, n23152, n23151, n23150,
         n23149, n23148, n23147, n23146, n23145, n23144, n23143, n23142,
         n23141, n23140, n23139, n23138, n23137, n23136, n23135, n23134,
         n23133, n23132, n23131, n23130, n23129, n23128, n23127, n23126,
         n23125, n23124, n23123, n23122, n23121, n23120, n23119, n23118,
         n23117, n23116, n23115, n23114, n23113, n23112, n23111, n23110,
         n23109, n23108, n23107, n23106, n23105, n23104, n23103, n23102,
         n23101, n23100, n23099, n23098, n23097, n23096, n23095, n23094,
         n23093, n23092, n23091, n23090, n23089, n23088, n23087, n23086,
         n23085, n23084, n23083, n23082, n23081, n23080, n23079, n23078,
         n23077, n23076, n23075, n23074, n23073, n23072, n23071, n23070,
         n23069, n23068, n23067, n23066, n23065, n23064, n23063, n23062,
         n23061, n23060, n23059, n23058, n23057, n23056, n23055, n23054,
         n23053, n23052, n23051, n23050, n23049, n23048, n23047, n23046,
         n23045, n23044, n23043, n23042, n23041, n23040, n23039, n23038,
         n23037, n23036, n23035, n23034, n23033, n23032, n23031, n23030,
         n23029, n23028, n23027, n23026, n23025, n23024, n23023, n23022,
         n23021, n23020, n23019, n23018, n23017, n23016, n23015, n23014,
         n23013, n23012, n23011, n23010, n23009, n23008, n23007, n23006,
         n23005, n23004, n23003, n23002, n23001, n23000, n22999, n22998,
         n22997, n22996, n22995, n22994, n22993, n22992, n22991, n22990,
         n22989, n22988, n22987, n22986, n22985, n22984, n22983, n22982,
         n22981, n22980, n22979, n22978, n22977, n22976, n22975, n22974,
         n22973, n22972, n22971, n22970, n22969, n22968, n22967, n22966,
         n22965, n22964, n22963, n22962, n22961, n22960, n22959, n22958,
         n22957, n22956, n22955, n22954, n22953, n22952, n22951, n22950,
         n22949, n22948, n22947, n22946, n22945, n22944, n22943, n22942,
         n22941, n22940, n22939, n22938, n22937, n22936, n22935, n22934,
         n22933, n22932, n22931, n22930, n22929, n22928, n22927, n22926,
         n22925, n22924, n22923, n22922, n22921, n22920, n22919, n22918,
         n22917, n22916, n22915, n22914, n22913, n22912, n22911, n22910,
         n22909, n22908, n22907, n22906, n22905, n22904, n22903, n22902,
         n22901, n22900, n22899, n22898, n22897, n22896, n22895, n22894,
         n22893, n22892, n22891, n22890, n22889, n22888, n22887, n22886,
         n22885, n22884, n22883, n22882, n22881, n22880, n22879, n22878,
         n22877, n22876, n22875, n22874, n22873, n22872, n22871, n22870,
         n22869, n22868, n22867, n22866, n22865, n22864, n22863, n22862,
         n22861, n22860, n22859, n22858, n22857, n22856, n22855, n22854,
         n22853, n22852, n22851, n22850, n22849, n22848, n22847, n22846,
         n22845, n22844, n22843, n22842, n22841, n22840, n22839, n22838,
         n22837, n22836, n22835, n22834, n22833, n22832, n22831, n22830,
         n22829, n22828, n22827, n22826, n22825, n22824, n22823, n22822,
         n22821, n22820, n22819, n22818, n22817, n22816, n22815, n22814,
         n22813, n22812, n22811, n22810, n22809, n22808, n22807, n22806,
         n22805, n22804, n22803, n22802, n22801, n22800, n22799, n22798,
         n22797, n22796, n22795, n22794, n22793, n22792, n22791, n22790,
         n22789, n22788, n22787, n22786, n22785, n22784, n22783, n22782,
         n22781, n22780, n22779, n22778, n22777, n22776, n22775, n22774,
         n22773, n22772, n22771, n22770, n22769, n22768, n22767, n22766,
         n22765, n22764, n22763, n22762, n22761, n22760, n22759, n22758,
         n22757, n22756, n22755, n22754, n22753, n22752, n22751, n22750,
         n22749, n22748, n22747, n22746, n22745, n22744, n22743, n22742,
         n22741, n22740, n22739, n22738, n22737, n22736, n22735, n22734,
         n22733, n22732, n22731, n22730, n22729, n22728, n22727, n22726,
         n22725, n22724, n22723, n22722, n22721, n22720, n22719, n22718,
         n22717, n22716, n22715, n22714, n22713, n22712, n22711, n22710,
         n22709, n22708, n22707, n22706, n22705, n22704, n22703, n22702,
         n22701, n22700, n22699, n22698, n22697, n22696, n22695, n22694,
         n22693, n22692, n22691, n22690, n22689, n22688, n22687, n22686,
         n22685, n22684, n22683, n22682, n22681, n22680, n22679, n22678,
         n22677, n22676, n22675, n22674, n22673, n22672, n22671, n22670,
         n22669, n22668, n22667, n22666, n22665, n22664, n22663, n22662,
         n22661, n22660, n22659, n22658, n22657, n22656, n22655, n22654,
         n22653, n22652, n22651, n22650, n22649, n22648, n22647, n22646,
         n22645, n22644, n22643, n22642, n22641, n22640, n22639, n22638,
         n22637, n22636, n22635, n22634, n22633, n22632, n22631, n22630,
         n22629, n22628, n22627, n22626, n22625, n22624, n22623, n22622,
         n22621, n22620, n22619, n22618, n22617, n22616, n22615, n22614,
         n22613, n22612, n22611, n22610, n22609, n22608, n22607, n22606,
         n22605, n22604, n22603, n22602, n22601, n22600, n22599, n22598,
         n22597, n22596, n22595, n22594, n22593, n22592, n22591, n22590,
         n22589, n22588, n22587, n22586, n22585, n22584, n22583, n22582,
         n22581, n22580, n22579, n22578, n22577, n22576, n22575, n22574,
         n22573, n22572, n22571, n22570, n22569, n22568, n22567, n22566,
         n22565, n22564, n22563, n22562, n22561, n22560, n22559, n22558,
         n22557, n22556, n22555, n22554, n22553, n22552, n22551, n22550,
         n22549, n22548, n22547, n22546, n22545, n22544, n22543, n22542,
         n22541, n22540, n22539, n22538, n22537, n22536, n22535, n22534,
         n22533, n22532, n22531, n22530, n22529, n22528, n22527, n22526,
         n22525, n22524, n22523, n22522, n22521, n22520, n22519, n22518,
         n22517, n22516, n22515, n22514, n22513, n22512, n22511, n22510,
         n22509, n22508, n22507, n22506, n22505, n22504, n22503, n22502,
         n22501, n22500, n22499, n22498, n22497, n22496, n22495, n22494,
         n22493, n22492, n22491, n22490, n22489, n22488, n22487, n22486,
         n22485, n22484, n22483, n22482, n22481, n22480, n22479, n22478,
         n22477, n22476, n22475, n22474, n22473, n22472, n22471, n22470,
         n22469, n22468, n22467, n22466, n22465, n22464, n22463, n22462,
         n22461, n22460, n22459, n22458, n22457, n22456, n22455, n22454,
         n22453, n22452, n22451, n22450, n22449, n22448, n22447, n22446,
         n22445, n22444, n22443, n22442, n22441, n22440, n22439, n22438,
         n22437, n22436, n22435, n22434, n22433, n22432, n22431, n22430,
         n22429, n22428, n22427, n22426, n22425, n22424, n22423, n22422,
         n22421, n22420, n22419, n22418, n22417, n22416, n22415, n22414,
         n22413, n22412, n22411, n22410, n22409, n22408, n22407, n22406,
         n22405, n22404, n22403, n22402, n22401, n22400, n22399, n22398,
         n22397, n22396, n22395, n22394, n22393, n22392, n22391, n22390,
         n22389, n22388, n22387, n22386, n22385, n22384, n22383, n22382,
         n22381, n22380, n22379, n22378, n22377, n22376, n22375, n22374,
         n22373, n22372, n22371, n22370, n22369, n22368, n22367, n22366,
         n22365, n22364, n22363, n22362, n22361, n22360, n22359, n22358,
         n22357, n22356, n22355, n22354, n22353, n22352, n22351, n22350,
         n22349, n22348, n22347, n22346, n22345, n22344, n22343, n22342,
         n22341, n22340, n22339, n22338, n22337, n22336, n22335, n22334,
         n22333, n22332, n22331, n22330, n22329, n22328, n22327, n22326,
         n22325, n22324, n22323, n22322, n22321, n22320, n22319, n22318,
         n22317, n22316, n22315, n22314, n22313, n22312, n22311, n22310,
         n22309, n22308, n22307, n22306, n22305, n22304, n22303, n22302,
         n22301, n22300, n22299, n22298, n22297, n22296, n22295, n22294,
         n22293, n22292, n22291, n22290, n22289, n22288, n22287, n22286,
         n22285, n22284, n22283, n22282, n22281, n22280, n22279, n22278,
         n22277, n22276, n22275, n22274, n22273, n22272, n22271, n22270,
         n22269, n22268, n22267, n22266, n22265, n22264, n22263, n22262,
         n22261, n22260, n22259, n22258, n22257, n22256, n22255, n22254,
         n22253, n22252, n22251, n22250, n22249, n22248, n22247, n22246,
         n22245, n22244, n22243, n22242, n22241, n22240, n22239, n22238,
         n22237, n22236, n22235, n22234, n22233, n22232, n22231, n22230,
         n22229, n22228, n22227, n22226, n22225, n22224, n22223, n22222,
         n22221, n22220, n22219, n22218, n22217, n22216, n22215, n22214,
         n22213, n22212, n22211, n22210, n22209, n22208, n22207, n22206,
         n22205, n22204, n22203, n22202, n22201, n22200, n22199, n22198,
         n22197, n22196, n22195, n22194, n22193, n22192, n22191, n22190,
         n22189, n22188, n22187, n22186, n22185, n22184, n22183, n22182,
         n22181, n22180, n22179, n22178, n22177, n22176, n22175, n22174,
         n22173, n22172, n22171, n22170, n22169, n22168, n22167, n22166,
         n22165, n22164, n22163, n22162, n22161, n22160, n22159, n22158,
         n22157, n22156, n22155, n22154, n22153, n22152, n22151, n22150,
         n22149, n22148, n22147, n22146, n22145, n22144, n22143, n22142,
         n22141, n22140, n22139, n22138, n22137, n22136, n22135, n22134,
         n22133, n22132, n22131, n22130, n22129, n22128, n22127, n22126,
         n22125, n22124, n22123, n22122, n22121, n22120, n22119, n22118,
         n22117, n22116, n22115, n22114, n22113, n22112, n22111, n22110,
         n22109, n22108, n22107, n22106, n22105, n22104, n22103, n22102,
         n22101, n22100, n22099, n22098, n22097, n22096, n22095, n22094,
         n22093, n22092, n22091, n22090, n22089, n22088, n22087, n22086,
         n22085, n22084, n22083, n22082, n22081, n22080, n22079, n22078,
         n22077, n22076, n22075, n22074, n22073, n22072, n22071, n22070,
         n22069, n22068, n22067, n22066, n22065, n22064, n22063, n22062,
         n22061, n22060, n22059, n22058, n22057, n22056, n22055, n22054,
         n22053, n22052, n22051, n22050, n22049, n22048, n22047, n22046,
         n22045, n22044, n22043, n22042, n22041, n22040, n22039, n22038,
         n22037, n22036, n22035, n22034, n22033, n22032, n22031, n22030,
         n22029, n22028, n22027, n22026, n22025, n22024, n22023, n22022,
         n22021, n22020, n22019, n22018, n22017, n22016, n22015, n22014,
         n22013, n22012, n22011, n22010, n22009, n22008, n22007, n22006,
         n22005, n22004, n22003, n22002, n22001, n22000, n21999, n21998,
         n21997, n21996, n21995, n21994, n21993, n21992, n21991, n21990,
         n21989, n21988, n21987, n21986, n21985, n21984, n21983, n21982,
         n21981, n21980, n21979, n21978, n21977, n21976, n21975, n21974,
         n21973, n21972, n21971, n21970, n21969, n21968, n21967, n21966,
         n21965, n21964, n21963, n21962, n21961, n21960, n21959, n21958,
         n21957, n21956, n21955, n21954, n21953, n21952, n21951, n21950,
         n21949, n21948, n21947, n21946, n21945, n21944, n21943, n21942,
         n21941, n21940, n21939, n21938, n21937, n21936, n21935, n21934,
         n21933, n21932, n21931, n21930, n21929, n21928, n21927, n21926,
         n21925, n21924, n21923, n21922, n21921, n21920, n21919, n21918,
         n21917, n21916, n21915, n21914, n21913, n21912, n21911, n21910,
         n21909, n21908, n21907, n21906, n21905, n21904, n21903, n21902,
         n21901, n21900, n21899, n21898, n21897, n21896, n21895, n21894,
         n21893, n21892, n21891, n21890, n21889, n21888, n21887, n21886,
         n21885, n21884, n21883, n21882, n21881, n21880, n21879, n21878,
         n21877, n21876, n21875, n21874, n21873, n21872, n21871, n21870,
         n21869, n21868, n21867, n21866, n21865, n21864, n21863, n21862,
         n21861, n21860, n21859, n21858, n21857, n21856, n21855, n21854,
         n21853, n21852, n21851, n21850, n21849, n21848, n21847, n21846,
         n21845, n21844, n21843, n21842, n21841, n21840, n21839, n21838,
         n21837, n21836, n21835, n21834, n21833, n21832, n21831, n21830,
         n21829, n21828, n21827, n21826, n21825, n21824, n21823, n21822,
         n21821, n21820, n21819, n21818, n21817, n21816, n21815, n21814,
         n21813, n21812, n21811, n21810, n21809, n21808, n21807, n21806,
         n21805, n21804, n21803, n21802, n21801, n21800, n21799, n21798,
         n21797, n21796, n21795, n21794, n21793, n21792, n21791, n21790,
         n21789, n21788, n21787, n21786, n21785, n21784, n21783, n21782,
         n21781, n21780, n21779, n21778, n21777, n21776, n21775, n21774,
         n21773, n21772, n21771, n21770, n21769, n21768, n21767, n21766,
         n21765, n21764, n21763, n21762, n21761, n21760, n21759, n21758,
         n21757, n21756, n21755, n21754, n21753, n21752, n21751, n21750,
         n21749, n21748, n21747, n21746, n21745, n21744, n21743, n21742,
         n21741, n21740, n21739, n21738, n21737, n21736, n21735, n21734,
         n21733, n21732, n21731, n21730, n21729, n21728, n21727, n21726,
         n21725, n21724, n21723, n21722, n21721, n21720, n21719, n21718,
         n21717, n21716, n21715, n21714, n21713, n21712, n21711, n21710,
         n21709, n21708, n21707, n21706, n21705, n21704, n21703, n21702,
         n21701, n21700, n21699, n21698, n21697, n21696, n21695, n21694,
         n21693, n21692, n21691, n21690, n21689, n21688, n21687, n21686,
         n21685, n21684, n21683, n21682, n21681, n21680, n21679, n21678,
         n21677, n21676, n21675, n21674, n21673, n21672, n21671, n21670,
         n21669, n21668, n21667, n21666, n21665, n21664, n21663, n21662,
         n21661, n21660, n21659, n21658, n21657, n21656, n21655, n21654,
         n21653, n21652, n21651, n21650, n21649, n21648, n21647, n21646,
         n21645, n21644, n21643, n21642, n21641, n21639, n21638, n21637,
         n21636, n21635, n21634, n21633, n21632, n21631, n21630, n21629,
         n21628, n21627, n21626, n21625, n21624, n21623, n21622, n21621,
         n21620, n21619, n21618, n21617, n21616, n21615, n21614, n21613,
         n21612, n21611, n21610, n21609, n21608, n21607, n21606, n21605,
         n21604, n21603, n21602, n21601, n21600, n21599, n21598, n21597,
         n21596, n21595, n21594, n21593, n21592, n21591, n21590, n21589,
         n21588, n21587, n21586, n21585, n21584, n21583, n21582, n21581,
         n21580, n21579, n21578, n21577, n21576, n21575, n21574, n21573,
         n21572, n21571, n21570, n21569, n21568, n21567, n21566, n21565,
         n21564, n21563, n21562, n21561, n21560, n21559, n21558, n21557,
         n21556, n21555, n21554, n21553, n21552, n21551, n21550, n21549,
         n21548, n21547, n21546, n21545, n21544, n21543, n21542, n21541,
         n21540, n21539, n21538, n21537, n21536, n21535, n21534, n21533,
         n21532, n21531, n21530, n21529, n21528, n21527, n21526, n21525,
         n21524, n21523, n21522, n21521, n21520, n21519, n21518, n21517,
         n21516, n21515, n21514, n21513, n21512, n21511, n21510, n21509,
         n21508, n21507, n21506, n21505, n21504, n21503, n21502, n21501,
         n21500, n21499, n21498, n21497, n21496, n21495, n21494, n21493,
         n21492, n21491, n21490, n21489, n21488, n21487, n21486, n21485,
         n21484, n21483, n21482, n21481, n21480, n21479, n21478, n21477,
         n21476, n21475, n21474, n21473, n21472, n21471, n21470, n21469,
         n21468, n21467, n21466, n21465, n21464, n21463, n21462, n21461,
         n21460, n21459, n21458, n21457, n21456, n21455, n21454, n21453,
         n21452, n21451, n21450, n21449, n21448, n21447, n21446, n21445,
         n21444, n21443, n21442, n21441, n21440, n21439, n21438, n21437,
         n21436, n21435, n21434, n21433, n21432, n21431, n21430, n21429,
         n21428, n21427, n21426, n21425, n21424, n21423, n21422, n21421,
         n21420, n21419, n21418, n21417, n21416, n21415, n21414, n21413,
         n21412, n21411, n21410, n21409, n21408, n21407, n21406, n21405,
         n21404, n21403, n21402, n21401, n21400, n21399, n21398, n21397,
         n21396, n21395, n21394, n21393, n21392, n21391, n21390, n21389,
         n21388, n21387, n21386, n21385, n21384, n21383, n21382, n21381,
         n21380, n21379, n21378, n21377, n21376, n21375, n21374, n21373,
         n21372, n21371, n21370, n21369, n21368, n21367, n21366, n21365,
         n21364, n21363, n21362, n21361, n21360, n21359, n21358, n21357,
         n21356, n21355, n21354, n21353, n21352, n21351, n21350, n21349,
         n21348, n21347, n21346, n21345, n21344, n21343, n21342, n21341,
         n21340, n21339, n21338, n21337, n21336, n21335, n21334, n21333,
         n21332, n21331, n21330, n21329, n21328, n21327, n21326, n21325,
         n21324, n21323, n21322, n21321, n21320, n21319, n21318, n21317,
         n21316, n21315, n21314, n21313, n21312, n21311, n21310, n21309,
         n21308, n21307, n21306, n21305, n21304, n21303, n21302, n21301,
         n21300, n21299, n21298, n21297, n21296, n21295, n21294, n21293,
         n21292, n21291, n21290, n21289, n21288, n21287, n21286, n21285,
         n21284, n21283, n21282, n21281, n21280, n21279, n21278, n21277,
         n21276, n21275, n21274, n21273, n21272, n21271, n21270, n21269,
         n21268, n21267, n21266, n21265, n21264, n21263, n21262, n21261,
         n21260, n21259, n21258, n21257, n21256, n21255, n21254, n21253,
         n21252, n21251, n21250, n21249, n21248, n21247, n21246, n21245,
         n21244, n21243, n21242, n21241, n21240, n21239, n21238, n21237,
         n21236, n21235, n21234, n21233, n21232, n21231, n21230, n21229,
         n21228, n21227, n21226, n21225, n21224, n21223, n21222, n21221,
         n21220, n21219, n21218, n21217, n21216, n21215, n21214, n21213,
         n21212, n21211, n21210, n21209, n21208, n21207, n21206, n21205,
         n21204, n21203, n21202, n21201, n21200, n21199, n21198, n21197,
         n21196, n21195, n21194, n21193, n21192, n21191, n21190, n21189,
         n21188, n21187, n21186, n21185, n21184, n21183, n21182, n21181,
         n21180, n21179, n21178, n21177, n21176, n21175, n21174, n21173,
         n21172, n21171, n21170, n21169, n21168, n21167, n21166, n21165,
         n21164, n21163, n21162, n21161, n21160, n21159, n21158, n21157,
         n21156, n21155, n21154, n21153, n21152, n21151, n21150, n21149,
         n21148, n21147, n21146, n21145, n21144, n21143, n21142, n21141,
         n21140, n21139, n21138, n21137, n21136, n21135, n21134, n21133,
         n21132, n21131, n21130, n21129, n21128, n21127, n21126, n21125,
         n21124, n21123, n21122, n21121, n21120, n21119, n21118, n21117,
         n21116, n21115, n21114, n21113, n21112, n21111, n21110, n21109,
         n21108, n21107, n21106, n21105, n21104, n21103, n21102, n21101,
         n21100, n21099, n21098, n21097, n21096, n21095, n21094, n21093,
         n21092, n21091, n21090, n21089, n21088, n21087, n21086, n21085,
         n21084, n21083, n21082, n21081, n21080, n21079, n21078, n21077,
         n21076, n21075, n21074, n21073, n21072, n21071, n21070, n21069,
         n21068, n21067, n21066, n21065, n21064, n21063, n21062, n21061,
         n21060, n21059, n21058, n21057, n21056, n21055, n21054, n21053,
         n21052, n21051, n21050, n21049, n21048, n21047, n21046, n21045,
         n21044, n21043, n21042, n21041, n21040, n21039, n21038, n21037,
         n21036, n21035, n21034, n21033, n21032, n21031, n21030, n21029,
         n21028, n21027, n21026, n21025, n21024, n21023, n21022, n21021,
         n21020, n21019, n21018, n21017, n21016, n21015, n21014, n21013,
         n21012, n21011, n21010, n21009, n21008, n21007, n21006, n21005,
         n21004, n21003, n21002, n21001, n21000, n20999, n20998, n20997,
         n20996, n20995, n20994, n20993, n20992, n20991, n20990, n20989,
         n20988, n20987, n20986, n20985, n20984, n20983, n20982, n20981,
         n20980, n20979, n20978, n20977, n20976, n20975, n20974, n20973,
         n20972, n20971, n20970, n20969, n20968, n20967, n20966, n20965,
         n20964, n20963, n20962, n20961, n20960, n20959, n20958, n20957,
         n20956, n20955, n20954, n20953, n20952, n20951, n20950, n20949,
         n20948, n20947, n20946, n20945, n20944, n20943, n20942, n20941,
         n20940, n20939, n20938, n20937, n20936, n20935, n20934, n20933,
         n20932, n20931, n20930, n20929, n20928, n20927, n20926, n20925,
         n20924, n20923, n20922, n20921, n20920, n20919, n20918, n20917,
         n20916, n20915, n20914, n20913, n20912, n20911, n20910, n20909,
         n20908, n20907, n20906, n20905, n20904, n20903, n20902, n20901,
         n20900, n20899, n20898, n20897, n20896, n20895, n20894, n20893,
         n20892, n20891, n20890, n20889, n20888, n20887, n20886, n20885,
         n20884, n20883, n20882, n20881, n20880, n20879, n20878, n20877,
         n20876, n20875, n20874, n20873, n20872, n20870, n20869, n20868,
         n20867, n20866, n20865, n20864, n20863, n20862, n20861, n20860,
         n20858, n20857, n20856, n20855, n20854, n20853, n20852, n20851,
         n20850, n20849, n20848, n20847, n20846, n20845, n20844, n20843,
         n20842, n20841, n20840, n20839, n20838, n20837, n20836, n20835,
         n20834, n20833, n20832, n20831, n20830, n20829, n20828, n20827,
         n20826, n20825, n20824, n20823, n20822, n20821, n20820, n20819,
         n20818, n20817, n20816, n20815, n20814, n20813, n20812, n20811,
         n20810, n20809, n20808, n20807, n20806, n20805, n20804, n20803,
         n20802, n20801, n20800, n20799, n20798, n20797, n20796, n20795,
         n20794, n20793, n20792, n20791, n20790, n20789, n20788, n20787,
         n20786, n20785, n20784, n20783, n20782, n20781, n20780, n20779,
         n20778, n20777, n20776, n20775, n20774, n20773, n20772, n20771,
         n20770, n20769, n20768, n20767, n20766, n20765, n20764, n20763,
         n20762, n20761, n20760, n20759, n20758, n20757, n20756, n20755,
         n20754, n20753, n20752, n20751, n20750, n20749, n20748, n20747,
         n20746, n20745, n20744, n20743, n20742, n20741, n20740, n20739,
         n20738, n20737, n20736, n20735, n20734, n20733, n20732, n20731,
         n20730, n20729, n20728, n20727, n20726, n20725, n20724, n20723,
         n20722, n20721, n20720, n20719, n20718, n20717, n20716, n20715,
         n20714, n20713, n20712, n20711, n20710, n20709, n20708, n20707,
         n20706, n20705, n20704, n20703, n20702, n20701, n20700, n20699,
         n20698, n20697, n20696, n20695, n20694, n20693, n20692, n20691,
         n20690, n20689, n20688, n20687, n20686, n20685, n20684, n20683,
         n20682, n20681, n20680, n20679, n20678, n20677, n20676, n20675,
         n20674, n20673, n20672, n20671, n20670, n20669, n20668, n20667,
         n20666, n20665, n20664, n20663, n20662, n20661, n20660, n20659,
         n20658, n20657, n20656, n20655, n20654, n20653, n20652, n20651,
         n20650, n20649, n20648, n20647, n20646, n20645, n20644, n20643,
         n20642, n20641, n20640, n20639, n20638, n20637, n20636, n20635,
         n20634, n20633, n20632, n20631, n20630, n20629, n20628, n20627,
         n20626, n20625, n20624, n20623, n20622, n20621, n20620, n20619,
         n20618, n20617, n20616, n20615, n20614, n20613, n20612, n20611,
         n20610, n20609, n20608, n20607, n20606, n20605, n20604, n20603,
         n20602, n20601, n20600, n20599, n20598, n20597, n20596, n20595,
         n20594, n20593, n20592, n20591, n20590, n20589, n20588, n20587,
         n20586, n20585, n20584, n20583, n20582, n20581, n20580, n20579,
         n20578, n20577, n20576, n20575, n20574, n20573, n20572, n20571,
         n20570, n20569, n20568, n20567, n20566, n20565, n20564, n20563,
         n20562, n20561, n20560, n20559, n20558, n20557, n20556, n20555,
         n20554, n20553, n20552, n20551, n20550, n20549, n20548, n20547,
         n20546, n20545, n20544, n20543, n20542, n20541, n20540, n20539,
         n20538, n20537, n20536, n20535, n20534, n20533, n20532, n20531,
         n20530, n20529, n20528, n20527, n20526, n20525, n20524, n20523,
         n20522, n20521, n20520, n20519, n20518, n20517, n20516, n20515,
         n20514, n20513, n20512, n20511, n20510, n20509, n20508, n20507,
         n20506, n20505, n20504, n20503, n20502, n20501, n20500, n20499,
         n20498, n20497, n20496, n20495, n20494, n20493, n20492, n20491,
         n20490, n20489, n20488, n20487, n20486, n20485, n20484, n20483,
         n20482, n20481, n20480, n20479, n20478, n20477, n20476, n20475,
         n20474, n20473, n20472, n20471, n20470, n20469, n20468, n20467,
         n20466, n20465, n20464, n20463, n20462, n20461, n20460, n20459,
         n20458, n20457, n20456, n20455, n20454, n20453, n20452, n20451,
         n20450, n20449, n20448, n20447, n20446, n20445, n20444, n20443,
         n20442, n20441, n20440, n20439, n20438, n20437, n20436, n20435,
         n20434, n20433, n20432, n20431, n20430, n20429, n20428, n20427,
         n20426, n20425, n20424, n20423, n20422, n20421, n20420, n20419,
         n20418, n20417, n20416, n20415, n20414, n20413, n20412, n20411,
         n20410, n20409, n20408, n20407, n20406, n20405, n20404, n20403,
         n20402, n20401, n20400, n20399, n20398, n20397, n20396, n20395,
         n20394, n20393, n20392, n20391, n20390, n20389, n20388, n20387,
         n20386, n20385, n20384, n20383, n20382, n20381, n20380, n20379,
         n20378, n20377, n20376, n20375, n20374, n20373, n20372, n20371,
         n20370, n20369, n20368, n20367, n20366, n20365, n20364, n20363,
         n20362, n20361, n20360, n20359, n20358, n20357, n20356, n20355,
         n20354, n20353, n20352, n20351, n20350, n20349, n20348, n20347,
         n20346, n20345, n20344, n20343, n20342, n20341, n20340, n20339,
         n20338, n20337, n20336, n20335, n20334, n20333, n20332, n20331,
         n20330, n20329, n20328, n20327, n20326, n20325, n20324, n20323,
         n20322, n20321, n20320, n20319, n20318, n20317, n20316, n20315,
         n20314, n20313, n20312, n20311, n20310, n20309, n20308, n20307,
         n20306, n20305, n20304, n20303, n20302, n20301, n20300, n20299,
         n20298, n20297, n20296, n20295, n20294, n20293, n20292, n20291,
         n20290, n20289, n20288, n20287, n20286, n20285, n20284, n20283,
         n20282, n20281, n20280, n20279, n20278, n20277, n20276, n20275,
         n20274, n20273, n20272, n20271, n20270, n20269, n20268, n20267,
         n20266, n20265, n20264, n20263, n20262, n20261, n20260, n20259,
         n20258, n20257, n20256, n20255, n20254, n20253, n20252, n20251,
         n20250, n20249, n20248, n20247, n20246, n20245, n20244, n20243,
         n20242, n20241, n20240, n20239, n20238, n20237, n20236, n20235,
         n20234, n20233, n20232, n20231, n20230, n20229, n20228, n20227,
         n20226, n20225, n20224, n20223, n20222, n20221, n20220, n20219,
         n20218, n20217, n20216, n20215, n20214, n20213, n20212, n20211,
         n20210, n20209, n20208, n20207, n20206, n20205, n20204, n20203,
         n20202, n20201, n20200, n20199, n20198, n20197, n20196, n20195,
         n20194, n20193, n20192, n20191, n20190, n20189, n20188, n20187,
         n20186, n20185, n20184, n20183, n20182, n20181, n20180, n20179,
         n20178, n20177, n20176, n20175, n20174, n20173, n20172, n20171,
         n20170, n20169, n20168, n20167, n20166, n20165, n20164, n20163,
         n20162, n20161, n20160, n20159, n20158, n20157, n20156, n20155,
         n20154, n20153, n20152, n20151, n20150, n20149, n20148, n20147,
         n20146, n20145, n20144, n20143, n20142, n20141, n20140, n20139,
         n20138, n20137, n20136, n20135, n20134, n20133, n20132, n20131,
         n20130, n20129, n20128, n20127, n20126, n20125, n20124, n20123,
         n20122, n20121, n20120, n20119, n20118, n20117, n20116, n20115,
         n20114, n20113, n20112, n20111, n20110, n20109, n20108, n20107,
         n20106, n20105, n20104, n20103, n20102, n20101, n20100, n20099,
         n20098, n20097, n20096, n20094, n20093, n20092, n20091, n20090,
         n20089, n20088, n20087, n20086, n20085, n20084, n20083, n20082,
         n20081, n20080, n20079, n20078, n20077, n20076, n20075, n20074,
         n20073, n20072, n20071, n20070, n20069, n20068, n20067, n20066,
         n20065, n20064, n20063, n20062, n20061, n20060, n20059, n20058,
         n20057, n20056, n20055, n20054, n20053, n20052, n20051, n20050,
         n20049, n20048, n20047, n20046, n20045, n20044, n20043, n20042,
         n20041, n20040, n20039, n20038, n20037, n20036, n20035, n20034,
         n20033, n20032, n20031, n20030, n20029, n20028, n20027, n20026,
         n20025, n20024, n20023, n20022, n20021, n20020, n20019, n20018,
         n20017, n20016, n20015, n20014, n20013, n20012, n20011, n20010,
         n20009, n20008, n20007, n20006, n20005, n20004, n20003, n20002,
         n20001, n20000, n19999, n19998, n19997, n19996, n19995, n19994,
         n19993, n19992, n19991, n19990, n19989, n19988, n19987, n19986,
         n19985, n19984, n19983, n19982, n19981, n19980, n19979, n19978,
         n19977, n19976, n19975, n19974, n19973, n19972, n19971, n19970,
         n19969, n19968, n19967, n19966, n19965, n19964, n19963, n19962,
         n19961, n19960, n19959, n19958, n19957, n19956, n19955, n19954,
         n19953, n19952, n19951, n19950, n19949, n19948, n19947, n19946,
         n19945, n19944, n19943, n19942, n19941, n19940, n19939, n19938,
         n19937, n19936, n19935, n19934, n19933, n19932, n19931, n19930,
         n19929, n19928, n19927, n19926, n19925, n19924, n19923, n19922,
         n19921, n19920, n19919, n19918, n19917, n19916, n19915, n19914,
         n19913, n19912, n19911, n19910, n19909, n19908, n19907, n19906,
         n19905, n19904, n19903, n19902, n19901, n19900, n19899, n19898,
         n19897, n19896, n19895, n19894, n19893, n19892, n19891, n19890,
         n19889, n19888, n19887, n19886, n19885, n19884, n19883, n19882,
         n19881, n19880, n19879, n19878, n19877, n19876, n19875, n19874,
         n19873, n19872, n19871, n19870, n19869, n19868, n19867, n19866,
         n19865, n19864, n19863, n19862, n19861, n19860, n19859, n19858,
         n19857, n19856, n19855, n19854, n19853, n19852, n19851, n19850,
         n19849, n19848, n19847, n19846, n19845, n19844, n19843, n19842,
         n19841, n19840, n19839, n19838, n19837, n19836, n19835, n19834,
         n19833, n19832, n19831, n19830, n19829, n19828, n19827, n19826,
         n19825, n19824, n19823, n19822, n19821, n19820, n19819, n19818,
         n19817, n19816, n19815, n19814, n19813, n19812, n19811, n19810,
         n19809, n19808, n19807, n19806, n19805, n19804, n19803, n19802,
         n19801, n19800, n19799, n19798, n19797, n19796, n19795, n19794,
         n19793, n19792, n19791, n19790, n19789, n19788, n19787, n19786,
         n19785, n19784, n19783, n19782, n19781, n19780, n19779, n19778,
         n19777, n19776, n19775, n19774, n19773, n19772, n19771, n19770,
         n19769, n19768, n19767, n19766, n19765, n19764, n19763, n19762,
         n19761, n19760, n19759, n19758, n19757, n19756, n19755, n19754,
         n19753, n19752, n19751, n19750, n19749, n19748, n19747, n19746,
         n19745, n19744, n19743, n19742, n19741, n19740, n19739, n19738,
         n19737, n19736, n19735, n19734, n19733, n19732, n19731, n19730,
         n19729, n19728, n19727, n19726, n19725, n19724, n19723, n19722,
         n19721, n19720, n19719, n19718, n19717, n19716, n19715, n19714,
         n19713, n19712, n19711, n19710, n19709, n19708, n19707, n19706,
         n19705, n19704, n19703, n19702, n19701, n19700, n19699, n19698,
         n19697, n19696, n19695, n19694, n19693, n19692, n19691, n19690,
         n19689, n19688, n19687, n19686, n19685, n19684, n19683, n19682,
         n19681, n19680, n19679, n19678, n19677, n19676, n19675, n19674,
         n19673, n19672, n19671, n19670, n19669, n19668, n19667, n19666,
         n19665, n19664, n19663, n19662, n19661, n19660, n19659, n19658,
         n19657, n19656, n19655, n19654, n19653, n19652, n19651, n19650,
         n19649, n19648, n19647, n19646, n19645, n19644, n19643, n19642,
         n19641, n19640, n19639, n19638, n19637, n19636, n19635, n19634,
         n19633, n19632, n19631, n19630, n19629, n19628, n19627, n19626,
         n19625, n19624, n19623, n19622, n19621, n19620, n19619, n19618,
         n19617, n19616, n19615, n19614, n19613, n19612, n19611, n19610,
         n19609, n19608, n19607, n19606, n19605, n19604, n19603, n19602,
         n19601, n19600, n19599, n19598, n19597, n19596, n19595, n19594,
         n19593, n19592, n19591, n19590, n19589, n19588, n19587, n19586,
         n19585, n19584, n19583, n19582, n19581, n19580, n19579, n19578,
         n19577, n19576, n19575, n19574, n19573, n19572, n19571, n19570,
         n19569, n19568, n19567, n19566, n19565, n19564, n19563, n19562,
         n19561, n19560, n19559, n19558, n19557, n19556, n19555, n19554,
         n19553, n19552, n19551, n19550, n19549, n19548, n19547, n19546,
         n19545, n19544, n19543, n19542, n19541, n19540, n19539, n19538,
         n19537, n19536, n19535, n19534, n19533, n19532, n19531, n19530,
         n19529, n19528, n19527, n19526, n19525, n19524, n19523, n19522,
         n19521, n19520, n19519, n19518, n19517, n19516, n19515, n19514,
         n19513, n19512, n19511, n19510, n19509, n19508, n19507, n19506,
         n19505, n19504, n19503, n19502, n19501, n19500, n19499, n19498,
         n19497, n19496, n19495, n19494, n19493, n19492, n19491, n19490,
         n19489, n19488, n19487, n19486, n19485, n19484, n19483, n19482,
         n19481, n19480, n19479, n19478, n19477, n19476, n19475, n19474,
         n19473, n19472, n19471, n19470, n19469, n19468, n19467, n19466,
         n19465, n19464, n19463, n19462, n19461, n19460, n19459, n19458,
         n19457, n19456, n19455, n19454, n19453, n19452, n19451, n19450,
         n19449, n19448, n19447, n19446, n19445, n19444, n19443, n19442,
         n19441, n19440, n19439, n19438, n19437, n19436, n19435, n19434,
         n19433, n19432, n19431, n19430, n19429, n19428, n19427, n19426,
         n19425, n19424, n19423, n19422, n19421, n19420, n19419, n19418,
         n19417, n19416, n19415, n19414, n19413, n19412, n19411, n19410,
         n19409, n19408, n19407, n19406, n19405, n19404, n19403, n19402,
         n19401, n19400, n19399, n19398, n19397, n19396, n19395, n19394,
         n19393, n19392, n19391, n19390, n19389, n19388, n19387, n19386,
         n19385, n19384, n19383, n19382, n19381, n19380, n19379, n19378,
         n19377, n19376, n19375, n19374, n19373, n19372, n19371, n19370,
         n19369, n19368, n19367, n19366, n19365, n19364, n19363, n19362,
         n19361, n19360, n19359, n19358, n19357, n19356, n19355, n19354,
         n19353, n19352, n19351, n19350, n19349, n19348, n19347, n19346,
         n19345, n19344, n19343, n19342, n19341, n19340, n19339, n19338,
         n19337, n19336, n19335, n19334, n19333, n19332, n19331, n19330,
         n19329, n19328, n19326, n19325, n19324, n19323, n19322, n19321,
         n19320, n19319, n19318, n19317, n19316, n19314, n19313, n19312,
         n19311, n19310, n19309, n19308, n19307, n19306, n19305, n19304,
         n19303, n19302, n19301, n19300, n19299, n19298, n19297, n19296,
         n19295, n19294, n19293, n19292, n19291, n19290, n19289, n19288,
         n19287, n19286, n19285, n19284, n19283, n19282, n19281, n19280,
         n19279, n19278, n19277, n19276, n19275, n19274, n19273, n19272,
         n19271, n19270, n19269, n19268, n19267, n19266, n19265, n19264,
         n19263, n19262, n19261, n19260, n19259, n19258, n19257, n19256,
         n19255, n19254, n19253, n19252, n19251, n19250, n19249, n19248,
         n19247, n19246, n19245, n19244, n19243, n19242, n19241, n19240,
         n19239, n19238, n19237, n19236, n19235, n19234, n19233, n19232,
         n19231, n19230, n19229, n19228, n19227, n19226, n19225, n19224,
         n19223, n19222, n19221, n19220, n19219, n19218, n19217, n19216,
         n19215, n19214, n19213, n19212, n19211, n19210, n19209, n19208,
         n19207, n19206, n19205, n19204, n19203, n19202, n19201, n19200,
         n19199, n19198, n19197, n19196, n19195, n19194, n19193, n19192,
         n19191, n19190, n19189, n19188, n19187, n19186, n19185, n19184,
         n19183, n19182, n19181, n19180, n19179, n19178, n19177, n19176,
         n19175, n19174, n19173, n19172, n19171, n19170, n19169, n19168,
         n19167, n19166, n19165, n19164, n19163, n19162, n19161, n19160,
         n19159, n19158, n19157, n19156, n19155, n19154, n19153, n19152,
         n19151, n19150, n19149, n19148, n19147, n19146, n19145, n19144,
         n19143, n19142, n19141, n19140, n19139, n19138, n19137, n19136,
         n19135, n19134, n19133, n19132, n19131, n19130, n19129, n19128,
         n19127, n19126, n19125, n19124, n19123, n19122, n19121, n19120,
         n19119, n19118, n19117, n19116, n19115, n19114, n19113, n19112,
         n19111, n19110, n19109, n19108, n19107, n19106, n19105, n19104,
         n19103, n19102, n19101, n19100, n19099, n19098, n19097, n19096,
         n19095, n19094, n19093, n19092, n19091, n19090, n19089, n19088,
         n19087, n19086, n19085, n19084, n19083, n19082, n19081, n19080,
         n19079, n19078, n19077, n19076, n19075, n19074, n19073, n19072,
         n19071, n19070, n19069, n19068, n19067, n19066, n19065, n19064,
         n19063, n19062, n19061, n19060, n19059, n19058, n19057, n19056,
         n19055, n19054, n19053, n19052, n19051, n19050, n19049, n19048,
         n19047, n19046, n19045, n19044, n19043, n19042, n19041, n19040,
         n19039, n19038, n19037, n19036, n19035, n19034, n19033, n19032,
         n19031, n19030, n19029, n19028, n19027, n19026, n19025, n19024,
         n19023, n19022, n19021, n19020, n19019, n19018, n19017, n19016,
         n19015, n19014, n19013, n19012, n19011, n19010, n19009, n19008,
         n19007, n19006, n19005, n19004, n19003, n19002, n19001, n19000,
         n18999, n18998, n18997, n18996, n18995, n18994, n18993, n18992,
         n18991, n18990, n18989, n18988, n18987, n18986, n18985, n18984,
         n18983, n18982, n18981, n18980, n18979, n18978, n18977, n18976,
         n18975, n18974, n18973, n18972, n18971, n18970, n18969, n18968,
         n18967, n18966, n18965, n18964, n18963, n18962, n18961, n18960,
         n18959, n18958, n18957, n18956, n18955, n18954, n18953, n18952,
         n18951, n18950, n18949, n18948, n18947, n18946, n18945, n18944,
         n18943, n18942, n18941, n18940, n18939, n18938, n18937, n18936,
         n18935, n18934, n18933, n18932, n18931, n18930, n18929, n18928,
         n18927, n18926, n18925, n18924, n18923, n18922, n18921, n18920,
         n18919, n18918, n18917, n18916, n18915, n18914, n18913, n18912,
         n18911, n18910, n18909, n18908, n18907, n18906, n18905, n18904,
         n18903, n18902, n18901, n18900, n18899, n18898, n18897, n18896,
         n18895, n18894, n18893, n18892, n18891, n18890, n18889, n18888,
         n18887, n18886, n18885, n18884, n18883, n18882, n18881, n18880,
         n18879, n18878, n18877, n18876, n18875, n18874, n18873, n18872,
         n18871, n18870, n18869, n18868, n18867, n18866, n18865, n18864,
         n18863, n18862, n18861, n18860, n18859, n18858, n18857, n18856,
         n18855, n18854, n18853, n18852, n18851, n18850, n18849, n18848,
         n18847, n18846, n18845, n18844, n18843, n18842, n18841, n18840,
         n18839, n18838, n18837, n18836, n18835, n18834, n18833, n18832,
         n18831, n18830, n18829, n18828, n18827, n18826, n18825, n18824,
         n18823, n18822, n18821, n18820, n18819, n18818, n18817, n18816,
         n18815, n18814, n18813, n18812, n18811, n18810, n18809, n18808,
         n18807, n18806, n18805, n18804, n18803, n18802, n18801, n18800,
         n18799, n18798, n18797, n18796, n18795, n18794, n18793, n18792,
         n18791, n18790, n18789, n18788, n18787, n18786, n18785, n18784,
         n18783, n18782, n18781, n18780, n18779, n18778, n18777, n18776,
         n18775, n18774, n18773, n18772, n18771, n18770, n18769, n18768,
         n18767, n18766, n18765, n18764, n18763, n18762, n18761, n18760,
         n18759, n18758, n18757, n18756, n18755, n18754, n18753, n18752,
         n18751, n18750, n18749, n18748, n18747, n18746, n18745, n18744,
         n18743, n18742, n18741, n18740, n18739, n18738, n18737, n18736,
         n18735, n18734, n18733, n18732, n18731, n18730, n18729, n18728,
         n18727, n18726, n18725, n18724, n18723, n18722, n18721, n18720,
         n18719, n18718, n18717, n18716, n18715, n18714, n18713, n18712,
         n18711, n18710, n18709, n18708, n18707, n18706, n18705, n18704,
         n18703, n18702, n18701, n18700, n18699, n18698, n18697, n18696,
         n18695, n18694, n18693, n18692, n18691, n18690, n18689, n18688,
         n18687, n18686, n18685, n18684, n18683, n18682, n18681, n18680,
         n18679, n18678, n18677, n18676, n18675, n18674, n18673, n18672,
         n18671, n18670, n18669, n18668, n18667, n18666, n18665, n18664,
         n18663, n18662, n18661, n18660, n18659, n18658, n18657, n18656,
         n18655, n18654, n18653, n18652, n18651, n18650, n18648, n18647,
         n18646, n18645, n18644, n18643, n18642, n18641, n18640, n18639,
         n18638, n18637, n18636, n18635, n18634, n18633, n18632, n18631,
         n18630, n18629, n18628, n18627, n18626, n18625, n18624, n18623,
         n18622, n18621, n18620, n18619, n18618, n18617, n18616, n18615,
         n18614, n18613, n18612, n18611, n18610, n18609, n18608, n18607,
         n18606, n18605, n18604, n18603, n18602, n18601, n18600, n18599,
         n18597, n18596, n18595, n18594, n18593, n18592, n18591, n18590,
         n18589, n18588, n18587, n18586, n18585, n18584, n18583, n18582,
         n18581, n18580, n18579, n18578, n18577, n18576, n18575, n18574,
         n18573, n18572, n18571, n18570, n18569, n18568, n18567, n18566,
         n18565, n18564, n18563, n18562, n18561, n18560, n18559, n18558,
         n18557, n18556, n18555, n18554, n18553, n18552, n18551, n18549,
         n18548, n18547, n18546, n18545, n18544, n18543, n18542, n18541,
         n18540, n18539, n18538, n18537, n18536, n18535, n18534, n18533,
         n18532, n18531, n18530, n18529, n18528, n18527, n18526, n18525,
         n18524, n18523, n18522, n18521, n18520, n18519, n18518, n18517,
         n18516, n18515, n18514, n18513, n18512, n18511, n18510, n18509,
         n18508, n18507, n18506, n18505, n18504, n18503, n18502, n18501,
         n18500, n18499, n18498, n18497, n18496, n18495, n18494, n18493,
         n18492, n18491, n18490, n18489, n18488, n18487, n18486, n18485,
         n18484, n18483, n18482, n18481, n18480, n18479, n18478, n18477,
         n18476, n18475, n18474, n18473, n18472, n18471, n18470, n18469,
         n18468, n18467, n18466, n18465, n18464, n18463, n18462, n18461,
         n18460, n18459, n18458, n18457, n18456, n18455, n18454, n18453,
         n18452, n18451, n18450, n18449, n18448, n18447, n18446, n18445,
         n18444, n18443, n18442, n18441, n18440, n18439, n18438, n18437,
         n18436, n18435, n18434, n18433, n18432, n18431, n18430, n18429,
         n18428, n18427, n18426, n18425, n18424, n18423, n18422, n18421,
         n18420, n18419, n18418, n18417, n18416, n18415, n18414, n18413,
         n18412, n18411, n18410, n18409, n18408, n18407, n18406, n18405,
         n18404, n18403, n18402, n18401, n18400, n18399, n18398, n18397,
         n18396, n18395, n18394, n18393, n18392, n18391, n18390, n18389,
         n18388, n18387, n18386, n18385, n18384, n18383, n18382, n18381,
         n18380, n18379, n18378, n18377, n18376, n18375, n18374, n18373,
         n18372, n18371, n18370, n18369, n18368, n18367, n18366, n18365,
         n18364, n18363, n18362, n18361, n18360, n18359, n18358, n18357,
         n18356, n18355, n18354, n18353, n18352, n18351, n18350, n18349,
         n18348, n18347, n18346, n18345, n18344, n18343, n18342, n18341,
         n18340, n18339, n18338, n18337, n18336, n18335, n18334, n18333,
         n18332, n18331, n18330, n18329, n18328, n18327, n18326, n18325,
         n18324, n18323, n18322, n18321, n18320, n18319, n18318, n18317,
         n18316, n18315, n18314, n18313, n18312, n18311, n18310, n18309,
         n18308, n18307, n18306, n18305, n18304, n18303, n18302, n18301,
         n18300, n18299, n18298, n18297, n18296, n18295, n18294, n18293,
         n18292, n18291, n18290, n18289, n18288, n18287, n18286, n18285,
         n18284, n18283, n18282, n18281, n18280, n18279, n18278, n18277,
         n18276, n18275, n18274, n18273, n18272, n18271, n18270, n18269,
         n18268, n18267, n18266, n18265, n18264, n18263, n18262, n18261,
         n18260, n18259, n18258, n18257, n18256, n18255, n18254, n18253,
         n18252, n18251, n18250, n18249, n18248, n18247, n18246, n18245,
         n18244, n18243, n18242, n18241, n18240, n18239, n18238, n18237,
         n18236, n18235, n18234, n18233, n18232, n18231, n18230, n18229,
         n18228, n18227, n18226, n18225, n18224, n18223, n18222, n18221,
         n18220, n18219, n18218, n18217, n18216, n18215, n18214, n18213,
         n18212, n18211, n18210, n18209, n18208, n18207, n18206, n18205,
         n18204, n18203, n18201, n18200, n18199, n18198, n18197, n18196,
         n18195, n18194, n18193, n18192, n18191, n18190, n18189, n18188,
         n18187, n18186, n18185, n18184, n18183, n18182, n18181, n18180,
         n18179, n18178, n18177, n18176, n18175, n18174, n18173, n18172,
         n18171, n18170, n18169, n18168, n18167, n18166, n18165, n18164,
         n18163, n18162, n18161, n18160, n18159, n18158, n18157, n18156,
         n18155, n18154, n18153, n18152, n18151, n18150, n18149, n18148,
         n18147, n18146, n18145, n18144, n18143, n18142, n18141, n18140,
         n18139, n18138, n18137, n18136, n18135, n18134, n18133, n18132,
         n18131, n18130, n18129, n18128, n18127, n18126, n18125, n18124,
         n18123, n18122, n18121, n18120, n18119, n18118, n18117, n18116,
         n18115, n18114, n18113, n18112, n18111, n18110, n18109, n18108,
         n18107, n18106, n18105, n18104, n18103, n18102, n18101, n18100,
         n18099, n18098, n18097, n18096, n18095, n18094, n18093, n18092,
         n18091, n18090, n18089, n18088, n18087, n18086, n18085, n18084,
         n18083, n18082, n18081, n18080, n18079, n18078, n18077, n18076,
         n18075, n18074, n18073, n18072, n18071, n18070, n18069, n18068,
         n18067, n18066, n18065, n18064, n18063, n18062, n18061, n18060,
         n18059, n18058, n18057, n18056, n18055, n18054, n18053, n18052,
         n18051, n18050, n18049, n18048, n18047, n18046, n18045, n18044,
         n18043, n18042, n18041, n18040, n18039, n18038, n18037, n18036,
         n18035, n18034, n18033, n18032, n18031, n18030, n18029, n18028,
         n18027, n18026, n18025, n18024, n18023, n18022, n18021, n18020,
         n18019, n18018, n18017, n18016, n18015, n18014, n18013, n18012,
         n18011, n18010, n18009, n18008, n18007, n18006, n18005, n18004,
         n18003, n18002, n18001, n18000, n17999, n17998, n17997, n17996,
         n17995, n17994, n17993, n17992, n17991, n17990, n17989, n17988,
         n17987, n17986, n17985, n17984, n17983, n17982, n17981, n17980,
         n17979, n17978, n17977, n17976, n17975, n17974, n17973, n17972,
         n17971, n17970, n17969, n17968, n17967, n17966, n17965, n17964,
         n17963, n17962, n17961, n17960, n17959, n17958, n17957, n17956,
         n17955, n17954, n17953, n17952, n17951, n17950, n17949, n17948,
         n17947, n17946, n17945, n17944, n17943, n17942, n17941, n17940,
         n17939, n17938, n17937, n17936, n17935, n17934, n17933, n17932,
         n17931, n17930, n17929, n17928, n17927, n17926, n17925, n17924,
         n17923, n17922, n17921, n17920, n17919, n17918, n17917, n17916,
         n17915, n17914, n17913, n17912, n17911, n17910, n17909, n17908,
         n17907, n17906, n17905, n17904, n17903, n17902, n17901, n17900,
         n17899, n17898, n17897, n17896, n17895, n17894, n17893, n17892,
         n17891, n17890, n17889, n17888, n17887, n17886, n17885, n17884,
         n17883, n17882, n17881, n17880, n17879, n17878, n17877, n17876,
         n17875, n17874, n17873, n17872, n17871, n17870, n17869, n17868,
         n17867, n17866, n17865, n17864, n17863, n17862, n17861, n17860,
         n17859, n17858, n17857, n17856, n17855, n17854, n17853, n17852,
         n17851, n17850, n17849, n17848, n17847, n17846, n17845, n17844,
         n17843, n17842, n17841, n17840, n17839, n17838, n17837, n17836,
         n17835, n17834, n17833, n17832, n17831, n17830, n17829, n17828,
         n17827, n17826, n17825, n17824, n17823, n17822, n17821, n17820,
         n17819, n17818, n17817, n17816, n17815, n17814, n17813, n17812,
         n17811, n17810, n17809, n17808, n17807, n17806, n17805, n17804,
         n17803, n17802, n17801, n17800, n17799, n17798, n17797, n17796,
         n17795, n17794, n17793, n17792, n17791, n17790, n17789, n17788,
         n17787, n17786, n17785, n17784, n17783, n17781, n17780, n17779,
         n17778, n17777, n17776, n17775, n17774, n17773, n17772, n17771,
         n17769, n17768, n17767, n17766, n17765, n17764, n17763, n17762,
         n17761, n17760, n17759, n17758, n17757, n17756, n17755, n17754,
         n17753, n17752, n17751, n17750, n17749, n17748, n17747, n17746,
         n17745, n17744, n17743, n17742, n17741, n17740, n17739, n17738,
         n17737, n17736, n17735, n17734, n17733, n17732, n17731, n17730,
         n17729, n17728, n17727, n17726, n17725, n17724, n17723, n17722,
         n17721, n17720, n17719, n17718, n17717, n17716, n17715, n17714,
         n17713, n17712, n17711, n17710, n17709, n17708, n17707, n17706,
         n17705, n17704, n17703, n17702, n17701, n17700, n17699, n17698,
         n17697, n17696, n17695, n17694, n17693, n17692, n17691, n17690,
         n17689, n17688, n17687, n17686, n17685, n17684, n17683, n17682,
         n17681, n17680, n17679, n17678, n17677, n17676, n17675, n17674,
         n17673, n17672, n17671, n17670, n17669, n17668, n17667, n17666,
         n17665, n17664, n17663, n17662, n17661, n17660, n17659, n17658,
         n17657, n17656, n17655, n17654, n17653, n17652, n17651, n17650,
         n17649, n17648, n17647, n17646, n17645, n17644, n17643, n17642,
         n17641, n17640, n17639, n17638, n17637, n17636, n17635, n17634,
         n17633, n17632, n17631, n17630, n17629, n17628, n17627, n17626,
         n17625, n17624, n17623, n17622, n17621, n17620, n17619, n17618,
         n17617, n17616, n17615, n17614, n17613, n17612, n17611, n17610,
         n17609, n17608, n17607, n17606, n17605, n17604, n17603, n17602,
         n17601, n17600, n17599, n17598, n17597, n17596, n17595, n17594,
         n17593, n17592, n17591, n17590, n17589, n17588, n17587, n17586,
         n17585, n17584, n17583, n17582, n17581, n17580, n17579, n17578,
         n17577, n17576, n17575, n17574, n17573, n17572, n17571, n17570,
         n17569, n17568, n17567, n17566, n17565, n17564, n17563, n17562,
         n17561, n17560, n17559, n17558, n17557, n17556, n17555, n17554,
         n17553, n17552, n17551, n17550, n17549, n17548, n17547, n17546,
         n17545, n17544, n17543, n17542, n17541, n17540, n17539, n17538,
         n17537, n17536, n17535, n17534, n17533, n17532, n17531, n17530,
         n17529, n17528, n17527, n17526, n17525, n17524, n17523, n17522,
         n17521, n17520, n17519, n17518, n17517, n17516, n17515, n17514,
         n17513, n17512, n17511, n17510, n17509, n17508, n17507, n17506,
         n17505, n17504, n17503, n17502, n17501, n17500, n17499, n17498,
         n17497, n17496, n17495, n17494, n17493, n17492, n17491, n17490,
         n17489, n17488, n17487, n17486, n17485, n17484, n17483, n17482,
         n17481, n17480, n17479, n17478, n17477, n17476, n17475, n17474,
         n17473, n17472, n17471, n17470, n17469, n17468, n17467, n17466,
         n17465, n17464, n17463, n17462, n17461, n17460, n17459, n17458,
         n17457, n17456, n17455, n17454, n17453, n17452, n17451, n17450,
         n17449, n17448, n17447, n17446, n17445, n17444, n17443, n17442,
         n17441, n17440, n17439, n17438, n17437, n17436, n17435, n17434,
         n17433, n17432, n17431, n17430, n17429, n17428, n17427, n17426,
         n17425, n17424, n17423, n17422, n17421, n17420, n17419, n17418,
         n17417, n17416, n17415, n17414, n17413, n17412, n17411, n17410,
         n17409, n17408, n17407, n17406, n17405, n17404, n17403, n17402,
         n17401, n17400, n17399, n17398, n17397, n17396, n17395, n17394,
         n17393, n17392, n17391, n17390, n17389, n17388, n17387, n17386,
         n17385, n17384, n17383, n17382, n17381, n17380, n17379, n17378,
         n17377, n17376, n17375, n17374, n17373, n17372, n17371, n17370,
         n17369, n17368, n17367, n17366, n17365, n17364, n17363, n17362,
         n17361, n17360, n17359, n17358, n17357, n17356, n17355, n17354,
         n17353, n17352, n17351, n17350, n17349, n17348, n17347, n17346,
         n17345, n17344, n17343, n17342, n17341, n17340, n17339, n17338,
         n17337, n17336, n17335, n17334, n17333, n17332, n17331, n17330,
         n17329, n17328, n17327, n17326, n17325, n17324, n17323, n17322,
         n17321, n17320, n17319, n17318, n17317, n17316, n17315, n17314,
         n17313, n17312, n17311, n17310, n17309, n17308, n17307, n17306,
         n17305, n17304, n17303, n17302, n17301, n17300, n17299, n17298,
         n17297, n17296, n17295, n17294, n17293, n17292, n17291, n17290,
         n17289, n17288, n17287, n17286, n17285, n17284, n17283, n17282,
         n17281, n17280, n17279, n17278, n17277, n17276, n17275, n17274,
         n17273, n17272, n17271, n17270, n17269, n17268, n17267, n17266,
         n17265, n17264, n17263, n17262, n17261, n17260, n17259, n17258,
         n17257, n17256, n17255, n17254, n17253, n17252, n17251, n17250,
         n17249, n17248, n17247, n17246, n17245, n17244, n17243, n17242,
         n17241, n17240, n17239, n17238, n17237, n17236, n17235, n17234,
         n17233, n17232, n17231, n17230, n17229, n17228, n17227, n17226,
         n17225, n17224, n17223, n17222, n17221, n17220, n17219, n17218,
         n17217, n17216, n17215, n17214, n17213, n17212, n17211, n17210,
         n17209, n17208, n17207, n17206, n17205, n17204, n17203, n17202,
         n17201, n17200, n17199, n17198, n17197, n17196, n17195, n17194,
         n17193, n17192, n17191, n17190, n17189, n17188, n17187, n17186,
         n17185, n17184, n17183, n17182, n17181, n17180, n17179, n17178,
         n17177, n17176, n17175, n17174, n17173, n17172, n17171, n17170,
         n17169, n17168, n17167, n17166, n17165, n17164, n17163, n17162,
         n17161, n17160, n17159, n17158, n17157, n17156, n17155, n17154,
         n17153, n17152, n17151, n17150, n17149, n17148, n17147, n17146,
         n17145, n17144, n17143, n17142, n17141, n17140, n17139, n17138,
         n17137, n17136, n17135, n17134, n17133, n17132, n17131, n17130,
         n17129, n17128, n17127, n17126, n17125, n17124, n17123, n17122,
         n17121, n17120, n17118, n17117, n17116, n17115, n17114, n17113,
         n17112, n17111, n17110, n17109, n17108, n17107, n17106, n17105,
         n17104, n17103, n17102, n17101, n17100, n17099, n17098, n17097,
         n17096, n17095, n17094, n17093, n17092, n17091, n17090, n17089,
         n17088, n17087, n17086, n17085, n17084, n17083, n17082, n17081,
         n17080, n17079, n17078, n17077, n17076, n17075, n17074, n17073,
         n17072, n17071, n17070, n17069, n17068, n17067, n17066, n17065,
         n17064, n17063, n17062, n17061, n17060, n17059, n17057, n17056,
         n17055, n17054, n17053, n17052, n17051, n17050, n17049, n17048,
         n17047, n17046, n17045, n17044, n17043, n17042, n17041, n17040,
         n17039, n17038, n17037, n17036, n17035, n17034, n17033, n17032,
         n17031, n17030, n17029, n17028, n17027, n17026, n17025, n17024,
         n17023, n17022, n17021, n17020, n17019, n17018, n17017, n17016,
         n17015, n17014, n17013, n17012, n17011, n17010, n17009, n17008,
         n17007, n17006, n17005, n17004, n17003, n17002, n17001, n17000,
         n16998, n16997, n16996, n16995, n16994, n16993, n16992, n16991,
         n16990, n16989, n16988, n16987, n16986, n16985, n16984, n16983,
         n16982, n16981, n16980, n16979, n16978, n16977, n16976, n16975,
         n16974, n16973, n16972, n16971, n16970, n16969, n16968, n16967,
         n16966, n16965, n16964, n16963, n16962, n16961, n16960, n16959,
         n16958, n16957, n16956, n16955, n16954, n16953, n16952, n16951,
         n16950, n16949, n16948, n16947, n16946, n16945, n16944, n16943,
         n16942, n16941, n16940, n16939, n16938, n16937, n16936, n16935,
         n16934, n16933, n16932, n16931, n16930, n16929, n16928, n16927,
         n16926, n16925, n16924, n16923, n16922, n16921, n16920, n16919,
         n16918, n16917, n16916, n16915, n16914, n16913, n16912, n16911,
         n16910, n16909, n16908, n16907, n16906, n16905, n16904, n16903,
         n16902, n16901, n16900, n16899, n16898, n16897, n16896, n16895,
         n16894, n16893, n16892, n16891, n16890, n16889, n16888, n16887,
         n16886, n16885, n16884, n16883, n16882, n16881, n16880, n16879,
         n16878, n16877, n16876, n16875, n16874, n16873, n16872, n16871,
         n16870, n16869, n16868, n16867, n16866, n16865, n16864, n16863,
         n16862, n16861, n16860, n16859, n16858, n16857, n16856, n16855,
         n16854, n16853, n16852, n16851, n16850, n16849, n16848, n16847,
         n16846, n16845, n16844, n16843, n16842, n16841, n16840, n16839,
         n16838, n16837, n16836, n16835, n16834, n16833, n16832, n16831,
         n16830, n16829, n16828, n16827, n16826, n16825, n16824, n16823,
         n16822, n16821, n16820, n16819, n16818, n16817, n16816, n16815,
         n16814, n16813, n16812, n16811, n16810, n16809, n16808, n16807,
         n16806, n16805, n16804, n16803, n16802, n16801, n16800, n16799,
         n16798, n16797, n16796, n16795, n16794, n16793, n16792, n16791,
         n16790, n16789, n16788, n16787, n16786, n16785, n16784, n16783,
         n16782, n16781, n16780, n16779, n16778, n16777, n16776, n16775,
         n16774, n16773, n16772, n16771, n16770, n16769, n16768, n16767,
         n16766, n16765, n16764, n16763, n16762, n16761, n16760, n16759,
         n16758, n16757, n16756, n16755, n16754, n16753, n16752, n16751,
         n16750, n16749, n16748, n16747, n16746, n16745, n16744, n16743,
         n16742, n16741, n16740, n16739, n16738, n16737, n16736, n16735,
         n16734, n16733, n16732, n16731, n16730, n16729, n16728, n16727,
         n16726, n16725, n16724, n16723, n16722, n16721, n16720, n16719,
         n16718, n16717, n16716, n16715, n16714, n16713, n16712, n16711,
         n16710, n16709, n16708, n16707, n16706, n16705, n16704, n16703,
         n16702, n16701, n16700, n16699, n16698, n16697, n16696, n16695,
         n16694, n16693, n16692, n16691, n16690, n16689, n16688, n16687,
         n16686, n16685, n16684, n16683, n16682, n16681, n16680, n16679,
         n16678, n16677, n16676, n16675, n16674, n16673, n16672, n16671,
         n16670, n16669, n16668, n16667, n16666, n16665, n16664, n16663,
         n16662, n16661, n16660, n16659, n16658, n16657, n16656, n16655,
         n16654, n16653, n16652, n16651, n16650, n16649, n16648, n16647,
         n16646, n16645, n16644, n16643, n16642, n16641, n16640, n16639,
         n16638, n16637, n16636, n16635, n16634, n16633, n16632, n16631,
         n16630, n16629, n16628, n16627, n16626, n16625, n16624, n16623,
         n16622, n16621, n16620, n16619, n16618, n16617, n16616, n16615,
         n16614, n16613, n16612, n16611, n16610, n16609, n16608, n16607,
         n16606, n16605, n16604, n16603, n16602, n16601, n16600, n16599,
         n16598, n16597, n16596, n16595, n16594, n16593, n16592, n16590,
         n16589, n16588, n16587, n16586, n16585, n16584, n16583, n16582,
         n16581, n16580, n16579, n16578, n16577, n16576, n16575, n16574,
         n16573, n16572, n16571, n16570, n16569, n16568, n16567, n16566,
         n16565, n16564, n16563, n16562, n16561, n16560, n16559, n16558,
         n16557, n16556, n16555, n16554, n16553, n16552, n16551, n16550,
         n16549, n16548, n16547, n16546, n16545, n16544, n16543, n16542,
         n16541, n16540, n16539, n16538, n16537, n16536, n16535, n16534,
         n16533, n16532, n16531, n16530, n16529, n16528, n16527, n16526,
         n16525, n16524, n16523, n16522, n16521, n16520, n16519, n16518,
         n16517, n16516, n16515, n16514, n16513, n16512, n16511, n16510,
         n16509, n16508, n16507, n16506, n16505, n16504, n16503, n16502,
         n16501, n16500, n16499, n16498, n16497, n16496, n16495, n16494,
         n16493, n16492, n16491, n16490, n16489, n16488, n16487, n16486,
         n16485, n16484, n16483, n16482, n16481, n16480, n16479, n16478,
         n16477, n16476, n16475, n16474, n16473, n16472, n16471, n16470,
         n16469, n16468, n16467, n16466, n16465, n16464, n16463, n16462,
         n16461, n16460, n16459, n16458, n16457, n16456, n16455, n16454,
         n16453, n16452, n16451, n16450, n16449, n16448, n16447, n16446,
         n16445, n16444, n16443, n16442, n16441, n16440, n16439, n16438,
         n16437, n16436, n16435, n16434, n16433, n16432, n16431, n16430,
         n16429, n16428, n16427, n16426, n16425, n16424, n16423, n16422,
         n16421, n16420, n16419, n16418, n16417, n16416, n16415, n16414,
         n16413, n16412, n16411, n16410, n16409, n16408, n16407, n16406,
         n16405, n16404, n16403, n16402, n16401, n16400, n16399, n16398,
         n16397, n16396, n16395, n16394, n16393, n16392, n16391, n16390,
         n16389, n16388, n16387, n16386, n16385, n16384, n16383, n16382,
         n16381, n16380, n16379, n16378, n16377, n16376, n16375, n16374,
         n16373, n16372, n16371, n16370, n16369, n16368, n16367, n16366,
         n16365, n16364, n16363, n16362, n16361, n16360, n16359, n16358,
         n16357, n16356, n16355, n16354, n16353, n16352, n16351, n16350,
         n16349, n16348, n16347, n16346, n16345, n16344, n16343, n16342,
         n16341, n16340, n16339, n16338, n16337, n16336, n16335, n16334,
         n16333, n16332, n16331, n16330, n16329, n16328, n16327, n16326,
         n16325, n16324, n16323, n16322, n16321, n16320, n16319, n16318,
         n16317, n16316, n16315, n16314, n16313, n16312, n16311, n16310,
         n16309, n16308, n16307, n16306, n16305, n16304, n16303, n16302,
         n16301, n16300, n16299, n16298, n16297, n16296, n16295, n16294,
         n16293, n16292, n16291, n16290, n16289, n16288, n16287, n16286,
         n16285, n16284, n16283, n16282, n16281, n16280, n16279, n16278,
         n16277, n16276, n16275, n16274, n16273, n16272, n16271, n16270,
         n16269, n16268, n16267, n16266, n16265, n16264, n16263, n16262,
         n16261, n16260, n16259, n16258, n16257, n16256, n16255, n16254,
         n16253, n16252, n16251, n16250, n16249, n16248, n16247, n16246,
         n16245, n16244, n16243, n16242, n16241, n16240, n16239, n16238,
         n16237, n16236, n16235, n16234, n16233, n16232, n16231, n16230,
         n16228, n16227, n16226, n16225, n16224, n16223, n16222, n16221,
         n16220, n16219, n16218, n16217, n16216, n16215, n16213, n16212,
         n16211, n16210, n16209, n16208, n16207, n16206, n16205, n16204,
         n16203, n16202, n16201, n16200, n16199, n16198, n16197, n16196,
         n16195, n16194, n16193, n16192, n16191, n16190, n16189, n16188,
         n16187, n16186, n16185, n16184, n16183, n16182, n16181, n16180,
         n16179, n16178, n16177, n16176, n16175, n16174, n16173, n16172,
         n16171, n16170, n16169, n16168, n16167, n16166, n16165, n16164,
         n16163, n16162, n16161, n16160, n16159, n16158, n16157, n16156,
         n16155, n16154, n16153, n16152, n16151, n16150, n16149, n16148,
         n16147, n16146, n16145, n16144, n16143, n16142, n16141, n16140,
         n16139, n16138, n16137, n16136, n16135, n16134, n16133, n16132,
         n16131, n16130, n16129, n16128, n16127, n16126, n16125, n16124,
         n16123, n16122, n16121, n16120, n16119, n16118, n16117, n16116,
         n16115, n16114, n16113, n16112, n16111, n16110, n16109, n16108,
         n16107, n16106, n16105, n16104, n16103, n16102, n16101, n16100,
         n16099, n16098, n16097, n16096, n16095, n16094, n16093, n16092,
         n16091, n16090, n16089, n16088, n16087, n16086, n16085, n16084,
         n16083, n16082, n16081, n16080, n16079, n16078, n16077, n16076,
         n16075, n16074, n16073, n16072, n16071, n16070, n16069, n16068,
         n16067, n16066, n16065, n16064, n16063, n16062, n16061, n16060,
         n16059, n16058, n16057, n16056, n16055, n16054, n16053, n16052,
         n16051, n16050, n16049, n16048, n16047, n16046, n16045, n16044,
         n16043, n16042, n16041, n16040, n16039, n16038, n16037, n16036,
         n16035, n16034, n16033, n16032, n16031, n16030, n16029, n16028,
         n16027, n16026, n16025, n16024, n16023, n16022, n16021, n16020,
         n16019, n16018, n16017, n16016, n16015, n16014, n16013, n16012,
         n16011, n16010, n16009, n16008, n16007, n16006, n16005, n16004,
         n16003, n16002, n16001, n16000, n15999, n15998, n15997, n15996,
         n15995, n15994, n15993, n15992, n15991, n15990, n15989, n15988,
         n15987, n15986, n15985, n15984, n15983, n15982, n15981, n15980,
         n15979, n15978, n15977, n15976, n15975, n15974, n15973, n15972,
         n15971, n15970, n15969, n15968, n15967, n15966, n15965, n15964,
         n15963, n15962, n15961, n15960, n15959, n15958, n15957, n15956,
         n15955, n15954, n15953, n15952, n15951, n15950, n15949, n15948,
         n15947, n15946, n15945, n15944, n15943, n15942, n15941, n15940,
         n15939, n15938, n15937, n15936, n15935, n15934, n15933, n15932,
         n15931, n15930, n15929, n15928, n15927, n15926, n15925, n15924,
         n15923, n15922, n15921, n15920, n15919, n15918, n15917, n15916,
         n15915, n15914, n15913, n15912, n15911, n15910, n15909, n15908,
         n15907, n15906, n15905, n15904, n15903, n15902, n15901, n15900,
         n15899, n15898, n15897, n15896, n15895, n15894, n15893, n15892,
         n15891, n15890, n15889, n15888, n15887, n15886, n15885, n15884,
         n15883, n15882, n15881, n15880, n15879, n15878, n15877, n15876,
         n15875, n15874, n15873, n15872, n15871, n15870, n15869, n15868,
         n15867, n15866, n15865, n15864, n15863, n15862, n15861, n15860,
         n15859, n15858, n15857, n15856, n15855, n15854, n15853, n15852,
         n15851, n15850, n15849, n15848, n15847, n15846, n15845, n15844,
         n15843, n15842, n15841, n15840, n15839, n15838, n15837, n15836,
         n15835, n15834, n15833, n15832, n15831, n15830, n15829, n15828,
         n15827, n15826, n15825, n15824, n15823, n15822, n15821, n15820,
         n15819, n15818, n15817, n15816, n15815, n15814, n15813, n15812,
         n15811, n15810, n15809, n15808, n15807, n15806, n15805, n15804,
         n15803, n15802, n15801, n15800, n15799, n15798, n15797, n15796,
         n15795, n15794, n15793, n15792, n15791, n15790, n15789, n15788,
         n15787, n15786, n15785, n15784, n15783, n15782, n15781, n15780,
         n15779, n15778, n15777, n15776, n15775, n15774, n15773, n15772,
         n15771, n15770, n15769, n15768, n15767, n15766, n15765, n15764,
         n15763, n15762, n15761, n15760, n15759, n15758, n15757, n15756,
         n15755, n15754, n15753, n15752, n15751, n15750, n15749, n15748,
         n15747, n15746, n15745, n15744, n15743, n15742, n15741, n15740,
         n15739, n15738, n15737, n15736, n15735, n15734, n15733, n15732,
         n15731, n15730, n15729, n15728, n15727, n15726, n15725, n15724,
         n15723, n15722, n15721, n15720, n15719, n15718, n15717, n15716,
         n15715, n15714, n15713, n15712, n15711, n15710, n15709, n15708,
         n15707, n15706, n15705, n15704, n15703, n15702, n15701, n15700,
         n15699, n15698, n15697, n15696, n15695, n15694, n15693, n15692,
         n15691, n15690, n15689, n15688, n15687, n15686, n15685, n15684,
         n15683, n15682, n15681, n15680, n15679, n15678, n15677, n15676,
         n15675, n15674, n15673, n15672, n15671, n15670, n15669, n15668,
         n15667, n15666, n15665, n15664, n15663, n15662, n15661, n15660,
         n15659, n15658, n15657, n15656, n15655, n15654, n15653, n15652,
         n15651, n15650, n15649, n15648, n15647, n15646, n15645, n15644,
         n15643, n15642, n15641, n15640, n15639, n15638, n15637, n15636,
         n15635, n15634, n15633, n15632, n15631, n15630, n15629, n15628,
         n15627, n15626, n15625, n15624, n15623, n15622, n15621, n15620,
         n15619, n15618, n15617, n15616, n15615, n15614, n15613, n15612,
         n15611, n15610, n15609, n15608, n15607, n15606, n15605, n15604,
         n15603, n15602, n15601, n15600, n15599, n15598, n15597, n15596,
         n15595, n15594, n15593, n15592, n15591, n15590, n15589, n15588,
         n15587, n15586, n15585, n15584, n15583, n15582, n15581, n15580,
         n15579, n15578, n15577, n15576, n15575, n15574, n15573, n15572,
         n15571, n15570, n15569, n15568, n15567, n15566, n15565, n15564,
         n15563, n15562, n15561, n15560, n15559, n15558, n15557, n15556,
         n15555, n15554, n15552, n15551, n15550, n15549, n15548, n15547,
         n15546, n15545, n15544, n15543, n15542, n15541, n15540, n15539,
         n15538, n15537, n15536, n15535, n15534, n15533, n15532, n15531,
         n15530, n15529, n15528, n15527, n15526, n15525, n15524, n15523,
         n15522, n15521, n15520, n15519, n15518, n15517, n15516, n15515,
         n15514, n15513, n15512, n15511, n15510, n15509, n15508, n15507,
         n15506, n15505, n15504, n15503, n15502, n15501, n15500, n15499,
         n15498, n15497, n15496, n15495, n15494, n15493, n15491, n15490,
         n15489, n15488, n15487, n15486, n15485, n15484, n15483, n15482,
         n15481, n15480, n15479, n15478, n15477, n15476, n15475, n15474,
         n15473, n15472, n15471, n15470, n15469, n15468, n15467, n15466,
         n15465, n15464, n15463, n15462, n15461, n15460, n15459, n15458,
         n15457, n15456, n15455, n15454, n15453, n15452, n15451, n15450,
         n15449, n15448, n15447, n15446, n15445, n15444, n15443, n15442,
         n15441, n15440, n15439, n15438, n15437, n15436, n15435, n15434,
         n15432, n15431, n15430, n15429, n15428, n15427, n15426, n15425,
         n15424, n15423, n15422, n15421, n15420, n15419, n15418, n15417,
         n15416, n15415, n15414, n15413, n15412, n15411, n15410, n15409,
         n15408, n15407, n15406, n15405, n15404, n15403, n15402, n15401,
         n15400, n15399, n15398, n15397, n15396, n15395, n15394, n15393,
         n15392, n15391, n15390, n15389, n15388, n15387, n15386, n15385,
         n15384, n15383, n15382, n15381, n15380, n15379, n15378, n15377,
         n15376, n15375, n15374, n15373, n15372, n15371, n15370, n15369,
         n15368, n15367, n15366, n15365, n15364, n15363, n15362, n15361,
         n15360, n15359, n15358, n15357, n15356, n15355, n15354, n15353,
         n15352, n15351, n15350, n15349, n15348, n15347, n15346, n15345,
         n15344, n15343, n15342, n15341, n15340, n15339, n15338, n15337,
         n15336, n15335, n15334, n15333, n15332, n15331, n15330, n15329,
         n15328, n15327, n15326, n15325, n15324, n15323, n15322, n15321,
         n15320, n15319, n15318, n15317, n15316, n15315, n15314, n15313,
         n15312, n15311, n15310, n15309, n15308, n15307, n15306, n15305,
         n15304, n15303, n15302, n15301, n15300, n15299, n15298, n15297,
         n15296, n15295, n15294, n15293, n15292, n15291, n15290, n15289,
         n15288, n15287, n15286, n15285, n15284, n15283, n15282, n15281,
         n15280, n15279, n15278, n15277, n15276, n15275, n15274, n15273,
         n15272, n15271, n15270, n15269, n15268, n15267, n15266, n15265,
         n15264, n15263, n15262, n15261, n15260, n15259, n15258, n15257,
         n15256, n15255, n15254, n15253, n15252, n15251, n15250, n15249,
         n15248, n15247, n15246, n15245, n15244, n15243, n15242, n15241,
         n15240, n15239, n15238, n15237, n15236, n15235, n15234, n15233,
         n15232, n15231, n15230, n15229, n15228, n15227, n15226, n15225,
         n15224, n15223, n15222, n15221, n15220, n15219, n15218, n15217,
         n15216, n15215, n15214, n15213, n15212, n15211, n15210, n15209,
         n15208, n15207, n15206, n15205, n15204, n15203, n15202, n15201,
         n15200, n15199, n15198, n15197, n15196, n15195, n15194, n15193,
         n15192, n15191, n15190, n15189, n15188, n15187, n15186, n15185,
         n15184, n15183, n15182, n15181, n15180, n15179, n15178, n15177,
         n15176, n15175, n15174, n15173, n15172, n15171, n15170, n15169,
         n15168, n15167, n15166, n15165, n15164, n15163, n15162, n15161,
         n15160, n15159, n15158, n15157, n15156, n15155, n15154, n15153,
         n15152, n15151, n15150, n15149, n15148, n15147, n15146, n15145,
         n15144, n15143, n15142, n15141, n15140, n15139, n15138, n15137,
         n15136, n15135, n15134, n15133, n15132, n15131, n15130, n15129,
         n15128, n15127, n15126, n15125, n15124, n15123, n15122, n15121,
         n15120, n15119, n15118, n15117, n15116, n15115, n15114, n15113,
         n15112, n15111, n15110, n15109, n15108, n15107, n15106, n15105,
         n15104, n15103, n15102, n15101, n15100, n15099, n15098, n15097,
         n15096, n15095, n15094, n15093, n15092, n15091, n15090, n15089,
         n15088, n15087, n15086, n15085, n15084, n15083, n15082, n15081,
         n15080, n15079, n15078, n15077, n15076, n15075, n15074, n15073,
         n15072, n15071, n15070, n15069, n15068, n15067, n15066, n15065,
         n15064, n15063, n15062, n15061, n15060, n15059, n15058, n15057,
         n15056, n15055, n15054, n15053, n15052, n15051, n15050, n15049,
         n15048, n15047, n15046, n15045, n15044, n15043, n15042, n15041,
         n15040, n15039, n15038, n15037, n15036, n15035, n15034, n15033,
         n15032, n15031, n15030, n15029, n15028, n15027, n15026, n15024,
         n15023, n15022, n15021, n15020, n15019, n15018, n15017, n15016,
         n15015, n15014, n15013, n15012, n15011, n15010, n15009, n15008,
         n15007, n15006, n15005, n15004, n15003, n15002, n15001, n15000,
         n14999, n14998, n14997, n14996, n14995, n14994, n14993, n14992,
         n14991, n14990, n14989, n14988, n14987, n14986, n14985, n14984,
         n14983, n14982, n14981, n14980, n14979, n14978, n14977, n14976,
         n14975, n14974, n14973, n14972, n14971, n14970, n14969, n14968,
         n14967, n14966, n14965, n14964, n14963, n14962, n14961, n14960,
         n14959, n14958, n14957, n14956, n14955, n14954, n14953, n14952,
         n14951, n14950, n14949, n14948, n14947, n14946, n14945, n14944,
         n14943, n14942, n14941, n14940, n14939, n14938, n14937, n14936,
         n14935, n14934, n14933, n14932, n14931, n14930, n14929, n14928,
         n14927, n14926, n14925, n14924, n14923, n14922, n14921, n14920,
         n14919, n14918, n14917, n14916, n14915, n14914, n14913, n14912,
         n14911, n14910, n14909, n14908, n14907, n14906, n14905, n14904,
         n14903, n14902, n14901, n14900, n14899, n14898, n14897, n14896,
         n14895, n14894, n14893, n14892, n14891, n14890, n14889, n14888,
         n14887, n14886, n14885, n14884, n14883, n14882, n14881, n14880,
         n14879, n14878, n14877, n14876, n14875, n14874, n14873, n14872,
         n14871, n14870, n14869, n14868, n14867, n14866, n14865, n14864,
         n14863, n14862, n14861, n14860, n14859, n14858, n14857, n14856,
         n14855, n14854, n14853, n14852, n14851, n14850, n14849, n14848,
         n14847, n14846, n14845, n14844, n14843, n14842, n14841, n14840,
         n14839, n14838, n14837, n14836, n14835, n14834, n14833, n14832,
         n14831, n14830, n14829, n14828, n14827, n14826, n14825, n14824,
         n14823, n14822, n14821, n14820, n14819, n14818, n14817, n14816,
         n14815, n14814, n14813, n14812, n14811, n14810, n14809, n14808,
         n14807, n14806, n14805, n14804, n14803, n14802, n14801, n14800,
         n14799, n14798, n14797, n14796, n14795, n14794, n14793, n14792,
         n14791, n14790, n14789, n14788, n14787, n14786, n14785, n14784,
         n14783, n14782, n14781, n14780, n14779, n14778, n14777, n14776,
         n14775, n14774, n14773, n14772, n14771, n14770, n14769, n14768,
         n14767, n14766, n14765, n14764, n14763, n14762, n14761, n14760,
         n14759, n14758, n14757, n14756, n14755, n14754, n14753, n14752,
         n14751, n14750, n14749, n14748, n14747, n14746, n14745, n14744,
         n14743, n14742, n14741, n14740, n14739, n14738, n14737, n14736,
         n14735, n14734, n14733, n14732, n14731, n14730, n14729, n14728,
         n14727, n14726, n14725, n14724, n14723, n14722, n14721, n14720,
         n14719, n14718, n14717, n14716, n14715, n14714, n14713, n14712,
         n14711, n14710, n14709, n14708, n14707, n14706, n14705, n14704,
         n14703, n14702, n14701, n14700, n14699, n14698, n14697, n14696,
         n14695, n14694, n14693, n14692, n14691, n14690, n14689, n14688,
         n14687, n14686, n14685, n14684, n14683, n14682, n14681, n14680,
         n14679, n14678, n14677, n14676, n14675, n14674, n14673, n14672,
         n14671, n14670, n14669, n14668, n14667, n14666, n14665, n14664,
         n14663, n14662, n14660, n14659, n14658, n14657, n14656, n14655,
         n14654, n14653, n14652, n14651, n14650, n14648, n14647, n14646,
         n14645, n14644, n14643, n14642, n14641, n14640, n14639, n14638,
         n14637, n14636, n14635, n14634, n14633, n14632, n14631, n14630,
         n14629, n14628, n14627, n14626, n14625, n14624, n14623, n14622,
         n14621, n14620, n14619, n14618, n14617, n14616, n14615, n14614,
         n14613, n14612, n14611, n14610, n14609, n14608, n14607, n14606,
         n14605, n14604, n14603, n14602, n14601, n14600, n14599, n14598,
         n14597, n14596, n14595, n14594, n14593, n14592, n14591, n14590,
         n14589, n14588, n14587, n14586, n14585, n14584, n14583, n14582,
         n14581, n14580, n14579, n14578, n14577, n14576, n14575, n14574,
         n14573, n14572, n14571, n14570, n14569, n14568, n14567, n14566,
         n14565, n14564, n14563, n14562, n14561, n14560, n14559, n14558,
         n14557, n14556, n14555, n14554, n14553, n14552, n14551, n14550,
         n14549, n14548, n14547, n14546, n14545, n14544, n14543, n14542,
         n14541, n14540, n14539, n14538, n14537, n14536, n14535, n14534,
         n14533, n14532, n14531, n14530, n14529, n14528, n14527, n14526,
         n14525, n14524, n14523, n14522, n14521, n14520, n14519, n14518,
         n14517, n14516, n14515, n14514, n14513, n14512, n14511, n14510,
         n14509, n14508, n14507, n14506, n14505, n14504, n14503, n14502,
         n14501, n14500, n14499, n14498, n14497, n14496, n14495, n14494,
         n14493, n14492, n14491, n14490, n14489, n14488, n14487, n14486,
         n14485, n14484, n14483, n14482, n14481, n14480, n14479, n14478,
         n14477, n14476, n14475, n14474, n14473, n14472, n14471, n14470,
         n14469, n14468, n14467, n14466, n14465, n14464, n14463, n14462,
         n14461, n14460, n14459, n14458, n14457, n14456, n14455, n14454,
         n14453, n14452, n14451, n14450, n14449, n14448, n14447, n14446,
         n14445, n14444, n14443, n14442, n14441, n14440, n14439, n14438,
         n14437, n14436, n14435, n14434, n14433, n14432, n14431, n14430,
         n14429, n14428, n14427, n14426, n14425, n14424, n14423, n14422,
         n14421, n14420, n14419, n14418, n14417, n14416, n14415, n14414,
         n14413, n14412, n14411, n14410, n14409, n14408, n14407, n14406,
         n14405, n14404, n14403, n14402, n14401, n14400, n14399, n14398,
         n14397, n14396, n14395, n14394, n14393, n14392, n14391, n14390,
         n14389, n14388, n14387, n14386, n14385, n14384, n14383, n14382,
         n14381, n14380, n14379, n14378, n14377, n14376, n14375, n14374,
         n14373, n14372, n14371, n14370, n14369, n14368, n14367, n14366,
         n14365, n14364, n14363, n14362, n14361, n14360, n14359, n14358,
         n14357, n14356, n14355, n14354, n14353, n14352, n14351, n14350,
         n14349, n14348, n14347, n14346, n14345, n14344, n14343, n14342,
         n14341, n14340, n14339, n14338, n14337, n14336, n14335, n14334,
         n14333, n14332, n14331, n14330, n14329, n14328, n14327, n14326,
         n14325, n14324, n14323, n14322, n14321, n14320, n14319, n14318,
         n14317, n14316, n14315, n14314, n14313, n14312, n14311, n14310,
         n14309, n14308, n14307, n14306, n14305, n14304, n14303, n14302,
         n14301, n14300, n14299, n14298, n14297, n14296, n14295, n14294,
         n14293, n14292, n14291, n14290, n14289, n14288, n14287, n14286,
         n14285, n14284, n14283, n14282, n14281, n14280, n14279, n14278,
         n14277, n14276, n14275, n14274, n14273, n14272, n14271, n14270,
         n14269, n14268, n14267, n14266, n14265, n14264, n14263, n14262,
         n14261, n14260, n14259, n14258, n14257, n14256, n14255, n14254,
         n14253, n14252, n14251, n14250, n14249, n14248, n14247, n14246,
         n14245, n14244, n14243, n14242, n14241, n14240, n14239, n14238,
         n14237, n14236, n14235, n14234, n14233, n14232, n14231, n14230,
         n14229, n14228, n14227, n14226, n14225, n14224, n14223, n14222,
         n14221, n14220, n14219, n14218, n14217, n14216, n14215, n14214,
         n14213, n14212, n14211, n14210, n14209, n14208, n14207, n14206,
         n14205, n14204, n14203, n14202, n14201, n14200, n14199, n14198,
         n14197, n14196, n14195, n14194, n14193, n14192, n14191, n14190,
         n14189, n14188, n14187, n14186, n14185, n14184, n14183, n14182,
         n14181, n14180, n14179, n14178, n14177, n14176, n14175, n14174,
         n14173, n14172, n14171, n14170, n14169, n14168, n14167, n14166,
         n14165, n14164, n14163, n14162, n14161, n14160, n14159, n14158,
         n14157, n14156, n14155, n14154, n14153, n14152, n14151, n14150,
         n14149, n14148, n14147, n14146, n14145, n14144, n14143, n14142,
         n14141, n14140, n14139, n14138, n14137, n14136, n14135, n14134,
         n14133, n14132, n14131, n14130, n14129, n14128, n14127, n14126,
         n14125, n14124, n14123, n14122, n14121, n14120, n14119, n14118,
         n14117, n14116, n14115, n14114, n14113, n14112, n14111, n14110,
         n14109, n14108, n14107, n14106, n14105, n14104, n14103, n14102,
         n14101, n14100, n14099, n14098, n14097, n14096, n14095, n14094,
         n14093, n14092, n14091, n14090, n14089, n14088, n14087, n14086,
         n14085, n14084, n14083, n14082, n14081, n14080, n14079, n14078,
         n14077, n14076, n14075, n14074, n14073, n14072, n14071, n14070,
         n14069, n14068, n14067, n14066, n14065, n14064, n14063, n14062,
         n14061, n14060, n14059, n14058, n14057, n14056, n14055, n14054,
         n14053, n14052, n14051, n14050, n14049, n14048, n14047, n14046,
         n14045, n14044, n14043, n14042, n14041, n14040, n14039, n14038,
         n14037, n14036, n14035, n14034, n14033, n14032, n14031, n14030,
         n14029, n14028, n14027, n14026, n14025, n14024, n14023, n14022,
         n14021, n14020, n14019, n14018, n14017, n14016, n14015, n14014,
         n14013, n14012, n14011, n14010, n14009, n14008, n14007, n14006,
         n14005, n14004, n14003, n14002, n14001, n13999, n13998, n13997,
         n13996, n13995, n13994, n13993, n13992, n13991, n13990, n13988,
         n13987, n13986, n13985, n13984, n13983, n13982, n13981, n13980,
         n13979, n13978, n13977, n13976, n13975, n13974, n13973, n13972,
         n13971, n13970, n13969, n13968, n13967, n13966, n13965, n13964,
         n13963, n13962, n13961, n13960, n13959, n13958, n13957, n13956,
         n13955, n13954, n13953, n13952, n13951, n13950, n13949, n13948,
         n13947, n13946, n13945, n13944, n13943, n13942, n13941, n13940,
         n13938, n13937, n13936, n13935, n13934, n13933, n13932, n13931,
         n13930, n13929, n13928, n13927, n13926, n13925, n13924, n13923,
         n13922, n13921, n13920, n13919, n13918, n13917, n13916, n13915,
         n13914, n13913, n13912, n13911, n13910, n13909, n13908, n13907,
         n13906, n13905, n13904, n13903, n13902, n13901, n13900, n13899,
         n13898, n13897, n13896, n13895, n13894, n13893, n13892, n13891,
         n13890, n13889, n13888, n13887, n13886, n13885, n13884, n13883,
         n13882, n13881, n13879, n13878, n13877, n13876, n13875, n13874,
         n13873, n13872, n13871, n13870, n13869, n13868, n13867, n13866,
         n13865, n13864, n13863, n13862, n13861, n13860, n13859, n13858,
         n13857, n13856, n13855, n13854, n13853, n13852, n13851, n13850,
         n13849, n13848, n13847, n13846, n13845, n13844, n13843, n13842,
         n13841, n13840, n13839, n13838, n13837, n13836, n13835, n13834,
         n13833, n13832, n13831, n13830, n13829, n13828, n13827, n13826,
         n13825, n13824, n13823, n13822, n13821, n13820, n13819, n13818,
         n13817, n13816, n13815, n13814, n13813, n13812, n13811, n13810,
         n13809, n13808, n13807, n13806, n13805, n13804, n13803, n13802,
         n13801, n13800, n13799, n13798, n13797, n13796, n13795, n13794,
         n13793, n13792, n13791, n13790, n13789, n13788, n13787, n13786,
         n13785, n13784, n13783, n13782, n13781, n13780, n13779, n13778,
         n13777, n13776, n13775, n13774, n13773, n13772, n13771, n13770,
         n13769, n13768, n13767, n13766, n13765, n13764, n13763, n13762,
         n13761, n13760, n13759, n13758, n13757, n13756, n13755, n13754,
         n13753, n13752, n13751, n13750, n13749, n13748, n13747, n13746,
         n13745, n13744, n13743, n13742, n13741, n13740, n13739, n13738,
         n13737, n13736, n13735, n13734, n13733, n13732, n13731, n13730,
         n13729, n13728, n13727, n13726, n13725, n13724, n13723, n13722,
         n13721, n13720, n13719, n13718, n13717, n13716, n13715, n13714,
         n13713, n13712, n13711, n13710, n13709, n13708, n13707, n13706,
         n13705, n13704, n13703, n13702, n13701, n13700, n13699, n13698,
         n13697, n13696, n13695, n13694, n13693, n13692, n13691, n13690,
         n13689, n13688, n13687, n13686, n13685, n13684, n13683, n13682,
         n13681, n13680, n13679, n13678, n13677, n13676, n13675, n13674,
         n13673, n13672, n13671, n13670, n13669, n13668, n13667, n13666,
         n13665, n13664, n13663, n13662, n13661, n13660, n13659, n13658,
         n13657, n13656, n13655, n13654, n13653, n13652, n13651, n13650,
         n13649, n13648, n13647, n13646, n13645, n13644, n13643, n13642,
         n13641, n13640, n13639, n13638, n13637, n13636, n13635, n13634,
         n13633, n13632, n13631, n13630, n13629, n13628, n13627, n13626,
         n13625, n13624, n13623, n13622, n13621, n13620, n13619, n13618,
         n13617, n13616, n13615, n13614, n13613, n13612, n13611, n13610,
         n13609, n13608, n13607, n13606, n13605, n13604, n13603, n13602,
         n13601, n13600, n13599, n13598, n13597, n13596, n13595, n13594,
         n13593, n13592, n13591, n13590, n13589, n13588, n13587, n13586,
         n13585, n13584, n13583, n13582, n13581, n13580, n13579, n13578,
         n13577, n13576, n13575, n13574, n13573, n13572, n13571, n13570,
         n13569, n13568, n13567, n13566, n13565, n13564, n13563, n13562,
         n13561, n13560, n13559, n13558, n13557, n13556, n13555, n13554,
         n13553, n13552, n13551, n13550, n13549, n13548, n13547, n13546,
         n13545, n13544, n13543, n13542, n13541, n13540, n13539, n13538,
         n13537, n13536, n13535, n13534, n13533, n13532, n13531, n13530,
         n13529, n13528, n13527, n13526, n13525, n13524, n13523, n13522,
         n13521, n13520, n13519, n13518, n13517, n13516, n13515, n13514,
         n13513, n13512, n13511, n13510, n13509, n13508, n13507, n13506,
         n13505, n13504, n13503, n13502, n13501, n13500, n13499, n13498,
         n13497, n13496, n13495, n13494, n13493, n13492, n13491, n13490,
         n13489, n13488, n13487, n13486, n13485, n13484, n13483, n13482,
         n13481, n13480, n13479, n13478, n13477, n13475, n13474, n13473,
         n13472, n13471, n13470, n13469, n13468, n13467, n13466, n13465,
         n13464, n13463, n13462, n13461, n13460, n13459, n13458, n13457,
         n13456, n13455, n13454, n13453, n13452, n13451, n13450, n13449,
         n13448, n13447, n13446, n13445, n13444, n13443, n13442, n13441,
         n13440, n13439, n13438, n13437, n13436, n13435, n13434, n13433,
         n13432, n13431, n13430, n13429, n13428, n13427, n13426, n13425,
         n13424, n13423, n13422, n13421, n13420, n13419, n13418, n13417,
         n13416, n13415, n13414, n13413, n13412, n13411, n13410, n13409,
         n13408, n13407, n13406, n13405, n13404, n13403, n13402, n13401,
         n13400, n13399, n13398, n13397, n13396, n13395, n13394, n13393,
         n13392, n13391, n13390, n13389, n13388, n13387, n13386, n13385,
         n13384, n13383, n13382, n13381, n13380, n13379, n13378, n13377,
         n13376, n13375, n13374, n13373, n13372, n13371, n13370, n13369,
         n13368, n13367, n13366, n13365, n13364, n13363, n13362, n13361,
         n13360, n13359, n13358, n13357, n13356, n13355, n13354, n13353,
         n13352, n13351, n13350, n13349, n13348, n13347, n13346, n13345,
         n13344, n13343, n13342, n13341, n13340, n13339, n13338, n13337,
         n13336, n13335, n13334, n13333, n13332, n13331, n13330, n13329,
         n13328, n13327, n13326, n13325, n13324, n13323, n13322, n13321,
         n13320, n13319, n13318, n13317, n13316, n13315, n13314, n13313,
         n13312, n13311, n13310, n13309, n13308, n13307, n13306, n13305,
         n13304, n13303, n13302, n13301, n13300, n13299, n13298, n13297,
         n13296, n13295, n13294, n13293, n13292, n13291, n13290, n13289,
         n13288, n13287, n13286, n13285, n13284, n13283, n13282, n13281,
         n13280, n13279, n13278, n13277, n13276, n13275, n13274, n13273,
         n13272, n13271, n13270, n13269, n13268, n13267, n13266, n13265,
         n13264, n13263, n13262, n13261, n13260, n13259, n13258, n13257,
         n13256, n13255, n13254, n13253, n13252, n13251, n13250, n13249,
         n13248, n13247, n13246, n13245, n13244, n13243, n13242, n13241,
         n13240, n13239, n13238, n13237, n13236, n13235, n13234, n13233,
         n13232, n13231, n13230, n13229, n13228, n13227, n13226, n13225,
         n13224, n13223, n13222, n13221, n13219, n13218, n13217, n13216,
         n13215, n13214, n13213, n13212, n13211, n13210, n13209, n13208,
         n13207, n13206, n13205, n13204, n13203, n13202, n13201, n13200,
         n13199, n13198, n13197, n13196, n13195, n13194, n13193, n13192,
         n13191, n13190, n13189, n13188, n13187, n13186, n13185, n13184,
         n13183, n13182, n13181, n13180, n13179, n13178, n13177, n13176,
         n13175, n13174, n13173, n13172, n13171, n13170, n13169, n13168,
         n13167, n13166, n13165, n13164, n13163, n13162, n13161, n13160,
         n13158, n13157, n13156, n13155, n13154, n13153, n13152, n13151,
         n13150, n13149, n13148, n13147, n13146, n13145, n13144, n13143,
         n13142, n13141, n13140, n13139, n13138, n13137, n13136, n13135,
         n13134, n13133, n13132, n13131, n13130, n13129, n13128, n13127,
         n13126, n13125, n13124, n13123, n13122, n13121, n13120, n13119,
         n13118, n13117, n13116, n13115, n13114, n13113, n13112, n13111,
         n13110, n13109, n13108, n13107, n13106, n13105, n13104, n13103,
         n13102, n13101, n13099, n13098, n13097, n13096, n13095, n13094,
         n13093, n13092, n13091, n13090, n13089, n13088, n13087, n13086,
         n13085, n13084, n13083, n13082, n13081, n13080, n13079, n13078,
         n13077, n13076, n13075, n13074, n13073, n13072, n13071, n13070,
         n13069, n13068, n13067, n13066, n13065, n13064, n13063, n13062,
         n13061, n13060, n13059, n13058, n13057, n13056, n13055, n13054,
         n13053, n13052, n13051, n13050, n13049, n13048, n13047, n13046,
         n13045, n13044, n13043, n13042, n13041, n13040, n13039, n13038,
         n13037, n13036, n13035, n13034, n13033, n13032, n13031, n13030,
         n13029, n13028, n13027, n13026, n13025, n13024, n13023, n13022,
         n13021, n13020, n13019, n13018, n13017, n13016, n13015, n13014,
         n13013, n13012, n13011, n13010, n13009, n13008, n13007, n13006,
         n13005, n13004, n13003, n13002, n13001, n13000, n12999, n12998,
         n12997, n12996, n12995, n12994, n12993, n12992, n12991, n12990,
         n12989, n12988, n12987, n12986, n12985, n12984, n12983, n12982,
         n12981, n12980, n12979, n12978, n12977, n12976, n12975, n12974,
         n12973, n12972, n12971, n12970, n12969, n12968, n12967, n12966,
         n12965, n12964, n12963, n12962, n12961, n12960, n12959, n12958,
         n12957, n12956, n12955, n12954, n12953, n12952, n12951, n12950,
         n12949, n12948, n12947, n12946, n12945, n12944, n12943, n12942,
         n12941, n12940, n12939, n12938, n12937, n12936, n12935, n12934,
         n12933, n12932, n12931, n12930, n12929, n12928, n12927, n12926,
         n12925, n12924, n12923, n12922, n12921, n12920, n12919, n12918,
         n12917, n12916, n12915, n12914, n12913, n12912, n12911, n12910,
         n12909, n12908, n12907, n12906, n12905, n12904, n12903, n12902,
         n12901, n12900, n12899, n12898, n12897, n12896, n12895, n12894,
         n12893, n12892, n12891, n12890, n12889, n12888, n12887, n12886,
         n12885, n12884, n12883, n12882, n12881, n12880, n12879, n12878,
         n12877, n12876, n12875, n12874, n12873, n12872, n12871, n12870,
         n12869, n12868, n12867, n12866, n12865, n12864, n12863, n12862,
         n12861, n12860, n12859, n12858, n12857, n12856, n12855, n12854,
         n12853, n12852, n12851, n12850, n12849, n12848, n12847, n12846,
         n12845, n12844, n12843, n12842, n12841, n12840, n12839, n12838,
         n12837, n12836, n12835, n12834, n12833, n12832, n12831, n12830,
         n12829, n12828, n12827, n12826, n12825, n12824, n12823, n12822,
         n12821, n12820, n12819, n12818, n12817, n12816, n12815, n12814,
         n12813, n12812, n12811, n12810, n12809, n12808, n12807, n12806,
         n12805, n12804, n12803, n12802, n12801, n12800, n12799, n12798,
         n12797, n12796, n12795, n12794, n12793, n12792, n12791, n12790,
         n12789, n12788, n12787, n12786, n12785, n12784, n12783, n12782,
         n12781, n12780, n12779, n12778, n12777, n12776, n12775, n12774,
         n12773, n12772, n12771, n12770, n12769, n12768, n12767, n12766,
         n12765, n12764, n12763, n12762, n12761, n12760, n12759, n12758,
         n12757, n12756, n12755, n12754, n12753, n12752, n12751, n12750,
         n12749, n12748, n12747, n12746, n12745, n12744, n12743, n12742,
         n12741, n12740, n12739, n12738, n12737, n12736, n12735, n12734,
         n12733, n12732, n12731, n12730, n12729, n12728, n12727, n12726,
         n12725, n12724, n12723, n12722, n12721, n12720, n12719, n12718,
         n12717, n12716, n12715, n12714, n12713, n12712, n12711, n12710,
         n12709, n12708, n12707, n12706, n12705, n12704, n12703, n12702,
         n12701, n12700, n12699, n12698, n12697, n12696, n12695, n12694,
         n12693, n12691, n12690, n12689, n12688, n12687, n12686, n12685,
         n12684, n12683, n12682, n12681, n12680, n12679, n12678, n12677,
         n12676, n12675, n12674, n12673, n12672, n12671, n12670, n12669,
         n12668, n12667, n12666, n12665, n12664, n12663, n12662, n12661,
         n12660, n12659, n12658, n12657, n12656, n12655, n12654, n12653,
         n12652, n12651, n12650, n12649, n12648, n12647, n12646, n12645,
         n12644, n12643, n12642, n12641, n12640, n12639, n12638, n12637,
         n12636, n12635, n12634, n12633, n12632, n12631, n12630, n12629,
         n12628, n12627, n12626, n12625, n12624, n12623, n12622, n12621,
         n12620, n12619, n12618, n12617, n12616, n12615, n12614, n12613,
         n12612, n12611, n12610, n12609, n12608, n12607, n12606, n12605,
         n12604, n12603, n12602, n12601, n12600, n12599, n12598, n12597,
         n12596, n12595, n12594, n12593, n12592, n12591, n12590, n12589,
         n12588, n12587, n12586, n12585, n12584, n12583, n12582, n12581,
         n12580, n12579, n12578, n12577, n12576, n12575, n12574, n12573,
         n12572, n12571, n12570, n12569, n12568, n12567, n12566, n12565,
         n12564, n12563, n12562, n12561, n12560, n12559, n12558, n12557,
         n12556, n12555, n12554, n12553, n12552, n12551, n12550, n12549,
         n12548, n12547, n12546, n12545, n12544, n12543, n12542, n12541,
         n12540, n12539, n12538, n12537, n12536, n12535, n12534, n12533,
         n12532, n12531, n12530, n12529, n12528, n12527, n12526, n12525,
         n12524, n12523, n12522, n12521, n12520, n12519, n12518, n12517,
         n12516, n12515, n12514, n12513, n12512, n12511, n12510, n12509,
         n12508, n12507, n12506, n12505, n12504, n12503, n12502, n12501,
         n12500, n12499, n12498, n12497, n12496, n12495, n12494, n12493,
         n12492, n12491, n12490, n12489, n12488, n12487, n12486, n12485,
         n12484, n12483, n12482, n12481, n12480, n12479, n12478, n12477,
         n12476, n12475, n12474, n12473, n12472, n12471, n12470, n12469,
         n12468, n12467, n12466, n12465, n12464, n12463, n12462, n12461,
         n12460, n12459, n12458, n12457, n12456, n12455, n12454, n12453,
         n12452, n12451, n12450, n12449, n12448, n12447, n12446, n12445,
         n12444, n12443, n12442, n12441, n12440, n12438, n12437, n12436,
         n12435, n12434, n12433, n12432, n12431, n12430, n12429, n12428,
         n12427, n12426, n12425, n12424, n12423, n12422, n12421, n12420,
         n12419, n12418, n12417, n12416, n12415, n12414, n12413, n12412,
         n12411, n12410, n12409, n12408, n12407, n12406, n12405, n12404,
         n12403, n12402, n12401, n12400, n12399, n12398, n12397, n12396,
         n12395, n12394, n12393, n12392, n12391, n12390, n12389, n12388,
         n12387, n12386, n12385, n12384, n12383, n12382, n12381, n12380,
         n12378, n12377, n12376, n12375, n12374, n12373, n12372, n12371,
         n12370, n12369, n12368, n12367, n12366, n12365, n12364, n12363,
         n12362, n12361, n12360, n12359, n12358, n12357, n12356, n12355,
         n12354, n12353, n12352, n12351, n12350, n12349, n12348, n12347,
         n12346, n12345, n12344, n12343, n12342, n12341, n12340, n12339,
         n12338, n12337, n12336, n12335, n12334, n12333, n12332, n12331,
         n12330, n12329, n12328, n12327, n12326, n12325, n12324, n12323,
         n12322, n12321, n12320, n12318, n12317, n12316, n12315, n12314,
         n12313, n12312, n12311, n12310, n12309, n12308, n12307, n12306,
         n12305, n12304, n12303, n12302, n12301, n12300, n12299, n12298,
         n12297, n12296, n12295, n12294, n12293, n12292, n12291, n12290,
         n12289, n12288, n12287, n12286, n12285, n12284, n12283, n12282,
         n12281, n12280, n12279, n12278, n12277, n12276, n12275, n12274,
         n12273, n12272, n12271, n12270, n12269, n12268, n12267, n12266,
         n12265, n12264, n12263, n12262, n12261, n12260, n12259, n12258,
         n12257, n12256, n12255, n12254, n12253, n12252, n12251, n12250,
         n12249, n12248, n12247, n12246, n12245, n12244, n12243, n12242,
         n12241, n12240, n12239, n12238, n12237, n12236, n12235, n12234,
         n12233, n12232, n12231, n12230, n12229, n12228, n12227, n12226,
         n12225, n12224, n12223, n12222, n12221, n12220, n12219, n12218,
         n12217, n12216, n12215, n12214, n12213, n12212, n12211, n12210,
         n12209, n12208, n12207, n12206, n12205, n12204, n12203, n12202,
         n12201, n12200, n12199, n12198, n12197, n12196, n12195, n12194,
         n12193, n12192, n12191, n12190, n12189, n12188, n12187, n12186,
         n12185, n12184, n12183, n12182, n12181, n12180, n12179, n12178,
         n12177, n12176, n12175, n12174, n12173, n12172, n12171, n12170,
         n12169, n12168, n12167, n12166, n12165, n12164, n12163, n12162,
         n12161, n12160, n12159, n12158, n12157, n12156, n12155, n12154,
         n12153, n12152, n12151, n12150, n12149, n12148, n12147, n12146,
         n12145, n12144, n12143, n12142, n12141, n12140, n12139, n12138,
         n12137, n12136, n12135, n12134, n12133, n12132, n12131, n12130,
         n12129, n12128, n12127, n12126, n12125, n12124, n12123, n12122,
         n12121, n12120, n12119, n12118, n12117, n12116, n12115, n12114,
         n12113, n12112, n12111, n12110, n12109, n12108, n12107, n12106,
         n12105, n12104, n12103, n12102, n12101, n12100, n12099, n12098,
         n12097, n12096, n12095, n12094, n12093, n12092, n12091, n12090,
         n12089, n12088, n12087, n12086, n12085, n12084, n12083, n12082,
         n12081, n12080, n12079, n12078, n12077, n12076, n12075, n12074,
         n12073, n12072, n12071, n12070, n12069, n12068, n12067, n12066,
         n12065, n12064, n12063, n12062, n12061, n12060, n12059, n12058,
         n12057, n12056, n12055, n12054, n12053, n12052, n12051, n12050,
         n12049, n12048, n12047, n12046, n12045, n12044, n12043, n12042,
         n12041, n12040, n12039, n12038, n12037, n12036, n12035, n12034,
         n12033, n12032, n12031, n12030, n12029, n12028, n12027, n12026,
         n12025, n12024, n12023, n12022, n12021, n12020, n12019, n12018,
         n12017, n12016, n12015, n12014, n12013, n12012, n12011, n12010,
         n12009, n12008, n12007, n12006, n12005, n12004, n12003, n12002,
         n12001, n12000, n11999, n11998, n11997, n11996, n11995, n11994,
         n11993, n11992, n11991, n11990, n11989, n11988, n11987, n11986,
         n11985, n11984, n11983, n11982, n11981, n11980, n11979, n11978,
         n11977, n11976, n11975, n11974, n11973, n11972, n11971, n11970,
         n11969, n11968, n11967, n11966, n11965, n11964, n11963, n11962,
         n11961, n11960, n11959, n11958, n11957, n11956, n11955, n11954,
         n11953, n11952, n11951, n11950, n11949, n11948, n11947, n11946,
         n11945, n11944, n11943, n11942, n11941, n11940, n11939, n11938,
         n11937, n11936, n11935, n11934, n11933, n11932, n11931, n11930,
         n11929, n11928, n11927, n11926, n11925, n11924, n11923, n11922,
         n11921, n11920, n11919, n11918, n11917, n11916, n11915, n11913,
         n11912, n11911, n11910, n11909, n11908, n11907, n11906, n11905,
         n11904, n11903, n11902, n11901, n11900, n11899, n11898, n11897,
         n11896, n11895, n11894, n11893, n11892, n11891, n11890, n11889,
         n11888, n11887, n11886, n11885, n11884, n11883, n11882, n11881,
         n11880, n11879, n11878, n11877, n11876, n11875, n11874, n11873,
         n11872, n11871, n11870, n11869, n11868, n11867, n11866, n11865,
         n11864, n11863, n11862, n11861, n11860, n11859, n11858, n11857,
         n11856, n11855, n11854, n11853, n11852, n11851, n11850, n11849,
         n11848, n11847, n11846, n11845, n11844, n11843, n11842, n11841,
         n11840, n11839, n11838, n11837, n11836, n11835, n11834, n11833,
         n11832, n11831, n11830, n11829, n11828, n11827, n11826, n11825,
         n11824, n11823, n11822, n11821, n11820, n11819, n11818, n11817,
         n11816, n11815, n11814, n11813, n11812, n11811, n11810, n11809,
         n11808, n11807, n11806, n11805, n11804, n11803, n11802, n11801,
         n11800, n11799, n11798, n11797, n11796, n11795, n11794, n11793,
         n11792, n11791, n11790, n11789, n11788, n11787, n11786, n11785,
         n11784, n11783, n11782, n11781, n11780, n11779, n11778, n11777,
         n11776, n11775, n11774, n11773, n11772, n11771, n11770, n11769,
         n11768, n11767, n11766, n11765, n11764, n11763, n11762, n11761,
         n11760, n11759, n11758, n11757, n11756, n11755, n11754, n11753,
         n11752, n11751, n11750, n11749, n11748, n11747, n11746, n11745,
         n11744, n11743, n11742, n11741, n11740, n11739, n11738, n11737,
         n11736, n11735, n11734, n11733, n11732, n11731, n11730, n11729,
         n11728, n11727, n11726, n11725, n11724, n11723, n11722, n11721,
         n11720, n11719, n11718, n11717, n11716, n11715, n11714, n11713,
         n11712, n11711, n11710, n11709, n11708, n11707, n11706, n11705,
         n11704, n11703, n11702, n11701, n11700, n11699, n11698, n11697,
         n11696, n11695, n11694, n11693, n11692, n11691, n11690, n11689,
         n11688, n11687, n11686, n11685, n11684, n11683, n11682, n11681,
         n11680, n11679, n11678, n11677, n11676, n11675, n11674, n11673,
         n11672, n11671, n11670, n11669, n11668, n11667, n11666, n11665,
         n11664, n11663, n11662, n11661, n11660, n11659, n11658, n11657,
         n11656, n11655, n11654, n11653, n11652, n11651, n11650, n11649,
         n11648, n11647, n11646, n11645, n11644, n11643, n11642, n11641,
         n11640, n11639, n11638, n11637, n11636, n11635, n11634, n11633,
         n11632, n11631, n11630, n11629, n11628, n11627, n11626, n11625,
         n11624, n11623, n11622, n11621, n11620, n11619, n11618, n11617,
         n11616, n11615, n11614, n11613, n11612, n11611, n11610, n11609,
         n11608, n11607, n11606, n11605, n11604, n11603, n11602, n11601,
         n11600, n11599, n11597, n11596, n11595, n11594, n11593, n11592,
         n11591, n11590, n11589, n11588, n11587, n11586, n11585, n11584,
         n11583, n11582, n11581, n11580, n11579, n11578, n11577, n11576,
         n11575, n11574, n11573, n11572, n11571, n11570, n11569, n11568,
         n11567, n11566, n11565, n11564, n11563, n11562, n11561, n11560,
         n11559, n11558, n11557, n11556, n11555, n11554, n11553, n11552,
         n11550, n11549, n11548, n11547, n11546, n11545, n11544, n11543,
         n11542, n11541, n11540, n11538, n11537, n11536, n11535, n11534,
         n11533, n11532, n11531, n11530, n11529, n11528, n11527, n11526,
         n11525, n11524, n11523, n11522, n11521, n11520, n11519, n11518,
         n11517, n11516, n11515, n11514, n11513, n11512, n11511, n11510,
         n11509, n11508, n11507, n11506, n11505, n11504, n11503, n11502,
         n11501, n11500, n11499, n11498, n11497, n11496, n11495, n11494,
         n11493, n11492, n11491, n11490, n11489, n11488, n11487, n11486,
         n11485, n11484, n11483, n11482, n11481, n11480, n11479, n11478,
         n11477, n11476, n11475, n11474, n11473, n11472, n11471, n11470,
         n11469, n11468, n11467, n11466, n11465, n11464, n11463, n11462,
         n11461, n11460, n11459, n11458, n11457, n11456, n11455, n11454,
         n11453, n11452, n11451, n11450, n11449, n11448, n11447, n11446,
         n11445, n11444, n11443, n11442, n11441, n11440, n11439, n11438,
         n11437, n11436, n11435, n11434, n11433, n11432, n11431, n11430,
         n11429, n11428, n11427, n11426, n11425, n11424, n11423, n11422,
         n11421, n11420, n11419, n11418, n11417, n11416, n11415, n11414,
         n11413, n11412, n11411, n11410, n11409, n11408, n11407, n11406,
         n11405, n11404, n11403, n11402, n11401, n11400, n11399, n11398,
         n11397, n11396, n11395, n11394, n11393, n11392, n11391, n11390,
         n11389, n11388, n11387, n11386, n11385, n11384, n11383, n11382,
         n11381, n11380, n11379, n11378, n11377, n11376, n11375, n11374,
         n11373, n11372, n11371, n11370, n11369, n11368, n11367, n11366,
         n11365, n11364, n11363, n11362, n11361, n11360, n11359, n11358,
         n11357, n11356, n11355, n11354, n11353, n11352, n11351, n11350,
         n11349, n11348, n11347, n11346, n11345, n11344, n11343, n11342,
         n11341, n11340, n11339, n11338, n11337, n11336, n11335, n11334,
         n11333, n11332, n11331, n11330, n11329, n11328, n11327, n11326,
         n11325, n11324, n11323, n11322, n11321, n11320, n11319, n11318,
         n11317, n11316, n11315, n11314, n11313, n11312, n11311, n11310,
         n11309, n11308, n11307, n11306, n11305, n11304, n11303, n11302,
         n11301, n11300, n11299, n11298, n11297, n11296, n11295, n11294,
         n11293, n11292, n11291, n11290, n11289, n11288, n11287, n11286,
         n11285, n11284, n11283, n11282, n11281, n11280, n11279, n11278,
         n11277, n11276, n11275, n11274, n11273, n11272, n11271, n11270,
         n11269, n11268, n11267, n11266, n11265, n11264, n11263, n11262,
         n11261, n11260, n11259, n11258, n11257, n11256, n11255, n11254,
         n11253, n11252, n11251, n11250, n11249, n11248, n11247, n11246,
         n11245, n11244, n11243, n11242, n11241, n11240, n11239, n11238,
         n11237, n11236, n11235, n11234, n11233, n11232, n11231, n11230,
         n11229, n11228, n11227, n11226, n11225, n11224, n11223, n11222,
         n11221, n11220, n11219, n11218, n11217, n11216, n11215, n11214,
         n11213, n11212, n11211, n11210, n11209, n11208, n11207, n11206,
         n11205, n11204, n11203, n11202, n11201, n11200, n11199, n11198,
         n11197, n11196, n11195, n11194, n11193, n11192, n11191, n11190,
         n11189, n11188, n11187, n11186, n11185, n11184, n11183, n11182,
         n11181, n11180, n11179, n11178, n11177, n11176, n11175, n11174,
         n11173, n11172, n11171, n11170, n11169, n11168, n11167, n11166,
         n11165, n11164, n11163, n11162, n11161, n11160, n11159, n11158,
         n11157, n11156, n11155, n11154, n11153, n11152, n11151, n11150,
         n11149, n11148, n11147, n11146, n11145, n11144, n11143, n11142,
         n11141, n11140, n11139, n11138, n11137, n11136, n11135, n11134,
         n11133, n11132, n11131, n11130, n11129, n11128, n11127, n11126,
         n11125, n11124, n11123, n11122, n11121, n11120, n11119, n11118,
         n11117, n11116, n11115, n11114, n11113, n11112, n11111, n11110,
         n11109, n11108, n11107, n11106, n11105, n11104, n11103, n11102,
         n11101, n11100, n11099, n11098, n11097, n11096, n11095, n11094,
         n11093, n11092, n11091, n11090, n11089, n11088, n11087, n11086,
         n11085, n11084, n11083, n11082, n11081, n11080, n11079, n11078,
         n11077, n11076, n11075, n11074, n11073, n11072, n11071, n11070,
         n11069, n11068, n11067, n11066, n11065, n11064, n11063, n11062,
         n11061, n11060, n11059, n11058, n11057, n11056, n11055, n11054,
         n11053, n11052, n11051, n11050, n11049, n11048, n11047, n11046,
         n11045, n11044, n11043, n11042, n11041, n11040, n11039, n11038,
         n11037, n11036, n11035, n11034, n11033, n11032, n11031, n11030,
         n11029, n11028, n11027, n11026, n11025, n11024, n11023, n11022,
         n11021, n11020, n11019, n11018, n11017, n11016, n11015, n11014,
         n11013, n11012, n11011, n11010, n11009, n11008, n11007, n11006,
         n11005, n11004, n11003, n11002, n11001, n11000, n10999, n10998,
         n10997, n10996, n10995, n10994, n10993, n10992, n10991, n10990,
         n10989, n10988, n10987, n10986, n10985, n10984, n10983, n10982,
         n10981, n10980, n10979, n10978, n10977, n10976, n10975, n10974,
         n10973, n10972, n10971, n10970, n10969, n10968, n10967, n10966,
         n10965, n10964, n10963, n10962, n10961, n10960, n10959, n10958,
         n10957, n10956, n10955, n10954, n10953, n10952, n10951, n10950,
         n10949, n10948, n10947, n10946, n10945, n10944, n10943, n10942,
         n10941, n10940, n10939, n10938, n10937, n10936, n10935, n10934,
         n10933, n10932, n10931, n10930, n10929, n10928, n10927, n10926,
         n10925, n10924, n10923, n10922, n10921, n10920, n10919, n10918,
         n10917, n10916, n10915, n10914, n10913, n10912, n10911, n10910,
         n10909, n10908, n10907, n10906, n10905, n10904, n10903, n10902,
         n10901, n10900, n10899, n10898, n10897, n10896, n10895, n10894,
         n10893, n10892, n10891, n10890, n10889, n10888, n10887, n10886,
         n10885, n10884, n10883, n10882, n10881, n10880, n10879, n10878,
         n10877, n10876, n10875, n10874, n10873, n10872, n10871, n10870,
         n10869, n10868, n10867, n10866, n10865, n10864, n10863, n10862,
         n10861, n10860, n10859, n10858, n10857, n10856, n10855, n10854,
         n10853, n10852, n10851, n10850, n10849, n10848, n10847, n10846,
         n10845, n10844, n10843, n10842, n10841, n10840, n10839, n10838,
         n10837, n10836, n10835, n10834, n10833, n10832, n10831, n10830,
         n10829, n10828, n10827, n10826, n10825, n10824, n10823, n10822,
         n10821, n10820, n10819, n10818, n10817, n10816, n10815, n10814,
         n10813, n10812, n10811, n10810, n10809, n10808, n10807, n10806,
         n10805, n10804, n10803, n10802, n10801, n10800, n10799, n10798,
         n10797, n10796, n10795, n10794, n10793, n10792, n10791, n10790,
         n10789, n10788, n10787, n10786, n10785, n10784, n10783, n10782,
         n10781, n10780, n10779, n10778, n10777, n10776, n10775, n10774,
         n10773, n10771, n10770, n10769, n10768, n10767, n10766, n10765,
         n10764, n10763, n10762, n10761, n10760, n10759, n10758, n10757,
         n10756, n10755, n10754, n10753, n10752, n10751, n10750, n10749,
         n10748, n10747, n10746, n10745, n10744, n10743, n10742, n10741,
         n10740, n10739, n10737, n10736, n10735, n10734, n10733, n10732,
         n10731, n10730, n10729, n10728, n10727, n10726, n10725, n10724,
         n10723, n10722, n10721, n10720, n10719, n10718, n10717, n10716,
         n10715, n10714, n10713, n10712, n10711, n10710, n10709, n10707,
         n10706, n10705, n10704, n10703, n10702, n10701, n10700, n10699,
         n10698, n10697, n10696, n10695, n10694, n10693, n10692, n10691,
         n10690, n10689, n10688, n10687, n10686, n10685, n10684, n10683,
         n10682, n10681, n10680, n10679, n10678, n10677, n10676, n10675,
         n10674, n10673, n10672, n10671, n10670, n10669, n10668, n10667,
         n10666, n10665, n10664, n10663, n10662, n10661, n10660, n10659,
         n10658, n10657, n10656, n10655, n10654, n10653, n10652, n10651,
         n10650, n10649, n10648, n10647, n10646, n10645, n10644, n10643,
         n10642, n10641, n10640, n10639, n10638, n10637, n10636, n10635,
         n10634, n10633, n10632, n10631, n10630, n10629, n10628, n10627,
         n10626, n10625, n10624, n10623, n10622, n10621, n10620, n10619,
         n10618, n10617, n10616, n10615, n10614, n10613, n10612, n10611,
         n10610, n10609, n10608, n10607, n10606, n10605, n10604, n10603,
         n10602, n10601, n10600, n10599, n10598, n10597, n10596, n10595,
         n10594, n10593, n10592, n10591, n10590, n10589, n10588, n10587,
         n10586, n10585, n10584, n10583, n10582, n10581, n10580, n10579,
         n10578, n10577, n10576, n10575, n10574, n10573, n10572, n10571,
         n10570, n10569, n10568, n10567, n10566, n10565, n10564, n10563,
         n10562, n10561, n10560, n10559, n10558, n10557, n10556, n10555,
         n10554, n10553, n10552, n10551, n10550, n10549, n10548, n10547,
         n10546, n10545, n10544, n10543, n10542, n10541, n10540, n10539,
         n10538, n10537, n10536, n10535, n10534, n10533, n10532, n10531,
         n10530, n10529, n10528, n10527, n10526, n10525, n10524, n10523,
         n10522, n10521, n10520, n10519, n10518, n10517, n10516, n10515,
         n10514, n10513, n10512, n10511, n10510, n10509, n10508, n10507,
         n10506, n10505, n10504, n10503, n10502, n10501, n10500, n10499,
         n10498, n10497, n10496, n10495, n10494, n10493, n10492, n10491,
         n10490, n10489, n10488, n10487, n10486, n10485, n10484, n10483,
         n10482, n10481, n10480, n10479, n10478, n10477, n10476, n10475,
         n10474, n10473, n10472, n10471, n10470, n10469, n10468, n10467,
         n10466, n10465, n10464, n10463, n10462, n10461, n10460, n10459,
         n10458, n10457, n10456, n10455, n10454, n10453, n10452, n10451,
         n10450, n10449, n10448, n10447, n10446, n10445, n10444, n10443,
         n10442, n10441, n10440, n10439, n10438, n10437, n10436, n10435,
         n10434, n10433, n10432, n10431, n10430, n10429, n10428, n10427,
         n10426, n10425, n10424, n10423, n10422, n10421, n10420, n10419,
         n10418, n10417, n10416, n10415, n10414, n10413, n10412, n10411,
         n10410, n10409, n10408, n10407, n10406, n10405, n10404, n10403,
         n10402, n10401, n10400, n10399, n10398, n10397, n10396, n10395,
         n10394, n10393, n10392, n10391, n10390, n10389, n10388, n10387,
         n10386, n10385, n10384, n10383, n10382, n10381, n10380, n10379,
         n10378, n10377, n10376, n10375, n10374, n10373, n10372, n10371,
         n10370, n10369, n10368, n10367, n10366, n10365, n10364, n10363,
         n10362, n10361, n10360, n10359, n10358, n10357, n10356, n10355,
         n10354, n10353, n10352, n10351, n10350, n10349, n10348, n10347,
         n10346, n10345, n10344, n10343, n10342, n10341, n10340, n10339,
         n10338, n10337, n10336, n10335, n10334, n10333, n10332, n10331,
         n10330, n10329, n10328, n10327, n10326, n10325, n10324, n10323,
         n10322, n10321, n10320, n10319, n10318, n10317, n10316, n10315,
         n10314, n10313, n10312, n10311, n10310, n10309, n10308, n10307,
         n10306, n10305, n10304, n10303, n10302, n10301, n10300, n10299,
         n10298, n10297, n10296, n10295, n10294, n10293, n10292, n10291,
         n10290, n10289, n10288, n10287, n10286, n10285, n10284, n10283,
         n10282, n10281, n10280, n10279, n10278, n10277, n10276, n10275,
         n10274, n10273, n10272, n10271, n10270, n10269, n10268, n10267,
         n10266, n10265, n10264, n10263, n10262, n10261, n10260, n10259,
         n10258, n10257, n10256, n10255, n10254, n10253, n10252, n10251,
         n10250, n10249, n10248, n10247, n10246, n10245, n10244, n10243,
         n10242, n10241, n10240, n10239, n10238, n10237, n10236, n10235,
         n10234, n10233, n10232, n10231, n10230, n10229, n10228, n10227,
         n10226, n10225, n10224, n10223, n10222, n10221, n10220, n10219,
         n10218, n10217, n10216, n10215, n10214, n10213, n10212, n10211,
         n10210, n10209, n10208, n10207, n10206, n10205, n10204, n10203,
         n10202, n10201, n10200, n10199, n10198, n10197, n10196, n10195,
         n10194, n10193, n10192, n10191, n10190, n10189, n10188, n10187,
         n10186, n10185, n10184, n10183, n10182, n10181, n10180, n10179,
         n10178, n10177, n10176, n10175, n10174, n10173, n10172, n10171,
         n10170, n10169, n10168, n10167, n10166, n10165, n10164, n10163,
         n10162, n10161, n10160, n10159, n10158, n10157, n10156, n10155,
         n10154, n10153, n10152, n10151, n10150, n10149, n10148, n10147,
         n10146, n10145, n10144, n10143, n10142, n10141, n10140, n10139,
         n10138, n10137, n10136, n10135, n10134, n10133, n10132, n10131,
         n10130, n10129, n10128, n10127, n10126, n10125, n10124, n10123,
         n10122, n10121, n10120, n10119, n10118, n10117, n10116, n10115,
         n10114, n10113, n10112, n10111, n10110, n10109, n10108, n10107,
         n10106, n10105, n10104, n10103, n10102, n10101, n10100, n10099,
         n10098, n10097, n10096, n10095, n10094, n10093, n10092, n10091,
         n10090, n10089, n10088, n10087, n10086, n10085, n10084, n10083,
         n10082, n10081, n10080, n10079, n10078, n10077, n10076, n10075,
         n10074, n10073, n10072, n10071, n10070, n10069, n10068, n10067,
         n10066, n10065, n10064, n10063, n10062, n10061, n10060, n10059,
         n10058, n10057, n10056, n10055, n10054, n10053, n10052, n10051,
         n10050, n10049, n10048, n10047, n10046, n10045, n10044, n10043,
         n10042, n10041, n10040, n10039, n10038, n10037, n10036, n10035,
         n10034, n10033, n10032, n10031, n10030, n10029, n10028, n10027,
         n10026, n10025, n10024, n10023, n10022, n10021, n10020, n10019,
         n10018, n10017, n10016, n10015, n10014, n10013, n10012, n10011,
         n10010, n10009, n10008, n10007, n10006, n10005, n10004, n10003,
         n10002, n10001, n10000, \L2_0/n4220 , \L2_0/n4219 , \L2_0/n4216 ,
         \L2_0/n4215 , \L2_0/n4212 , \L2_0/n4211 , \L2_0/n4208 , \L2_0/n4207 ,
         \L2_0/n4204 , \L2_0/n4203 , \L2_0/n4200 , \L2_0/n4199 , \L2_0/n4196 ,
         \L2_0/n4195 , \L2_0/n4192 , \L2_0/n4191 , \L2_0/n4188 , \L2_0/n4187 ,
         \L2_0/n4184 , \L2_0/n4183 , \L2_0/n4180 , \L2_0/n4179 , \L2_0/n4176 ,
         \L2_0/n4175 , \L2_0/n4172 , \L2_0/n4171 , \L2_0/n4168 , \L2_0/n4167 ,
         \L2_0/n4164 , \L2_0/n4163 , \L2_0/n4160 , \L2_0/n4159 , \L2_0/n4156 ,
         \L2_0/n4155 , \L2_0/n4152 , \L2_0/n4151 , \L2_0/n4148 , \L2_0/n4147 ,
         \L2_0/n4144 , \L2_0/n4136 , \L2_0/n4132 , \L2_0/n4128 , \L2_0/n4124 ,
         \L2_0/n4120 , \L2_0/n4116 , \L2_0/n4112 , \L2_0/n4108 , \L2_0/n4104 ,
         \L2_0/n4100 , \L2_0/n4096 , \L2_0/n4092 , \L2_0/n4088 , \L2_0/n4084 ,
         \L2_0/n4080 , \L2_0/n4076 , \L2_0/n4072 , \L2_0/n4068 , \L2_0/n4064 ,
         \L2_0/n4056 , \L2_0/n4052 , \L2_0/n4048 , \L2_0/n4044 , \L2_0/n4040 ,
         \L2_0/n4036 , \L2_0/n4032 , \L2_0/n4028 , \L2_0/n4024 , \L2_0/n4020 ,
         \L2_0/n4016 , \L2_0/n4012 , \L2_0/n4008 , \L2_0/n4004 , \L2_0/n4000 ,
         \L2_0/n3996 , \L2_0/n3992 , \L2_0/n3988 , \L2_0/n3984 , \L2_0/n3976 ,
         \L2_0/n3972 , \L2_0/n3968 , \L2_0/n3964 , \L2_0/n3960 , \L2_0/n3956 ,
         \L2_0/n3952 , \L2_0/n3948 , \L2_0/n3944 , \L2_0/n3940 , \L2_0/n3936 ,
         \L2_0/n3932 , \L2_0/n3928 , \L2_0/n3924 , \L2_0/n3920 , \L2_0/n3916 ,
         \L2_0/n3912 , \L2_0/n3908 , \L2_0/n3904 , \L2_0/n3896 , \L2_0/n3892 ,
         \L2_0/n3888 , \L2_0/n3884 , \L2_0/n3880 , \L2_0/n3876 , \L2_0/n3872 ,
         \L2_0/n3868 , \L2_0/n3864 , \L2_0/n3860 , \L2_0/n3856 , \L2_0/n3852 ,
         \L2_0/n3848 , \L2_0/n3844 , \L2_0/n3840 , \L2_0/n3836 , \L2_0/n3832 ,
         \L2_0/n3828 , \L2_0/n3824 , \L2_0/n3816 , \L2_0/n3812 , \L2_0/n3808 ,
         \L2_0/n3804 , \L2_0/n3800 , \L2_0/n3796 , \L2_0/n3792 , \L2_0/n3788 ,
         \L2_0/n3784 , \L2_0/n3780 , \L2_0/n3776 , \L2_0/n3772 , \L2_0/n3768 ,
         \L2_0/n3764 , \L2_0/n3760 , \L2_0/n3756 , \L2_0/n3752 , \L2_0/n3748 ,
         \L2_0/n3744 , \L2_0/n3736 , \L2_0/n3732 , \L2_0/n3728 , \L2_0/n3724 ,
         \L2_0/n3720 , \L2_0/n3716 , \L2_0/n3712 , \L2_0/n3708 , \L2_0/n3704 ,
         \L2_0/n3700 , \L2_0/n3696 , \L2_0/n3692 , \L2_0/n3688 , \L2_0/n3684 ,
         \L2_0/n3680 , \L2_0/n3676 , \L2_0/n3672 , \L2_0/n3668 , \L2_0/n3664 ,
         \L2_0/n3656 , \L2_0/n3652 , \L2_0/n3648 , \L2_0/n3644 , \L2_0/n3640 ,
         \L2_0/n3636 , \L2_0/n3632 , \L2_0/n3628 , \L2_0/n3624 , \L2_0/n3620 ,
         \L2_0/n3616 , \L2_0/n3612 , \L2_0/n3608 , \L2_0/n3604 , \L2_0/n3600 ,
         \L2_0/n3596 , \L2_0/n3592 , \L2_0/n3588 , \L2_0/n3584 , \L2_0/n3576 ,
         \L2_0/n3572 , \L2_0/n3568 , \L2_0/n3564 , \L2_0/n3560 , \L2_0/n3556 ,
         \L2_0/n3552 , \L2_0/n3548 , \L2_0/n3544 , \L2_0/n3540 , \L2_0/n3536 ,
         \L2_0/n3532 , \L2_0/n3528 , \L2_0/n3524 , \L2_0/n3520 , \L2_0/n3516 ,
         \L2_0/n3512 , \L2_0/n3508 , \L2_0/n3504 , \L2_0/n3496 , \L2_0/n3492 ,
         \L2_0/n3488 , \L2_0/n3484 , \L2_0/n3480 , \L2_0/n3476 , \L2_0/n3472 ,
         \L2_0/n3468 , \L2_0/n3464 , \L2_0/n3460 , \L2_0/n3456 , \L2_0/n3452 ,
         \L2_0/n3448 , \L2_0/n3444 , \L2_0/n3440 , \L2_0/n3436 , \L2_0/n3432 ,
         \L2_0/n3428 , \L2_0/n3424 , \L2_0/n3416 , \L2_0/n3412 , \L2_0/n3408 ,
         \L2_0/n3404 , \L2_0/n3400 , \L2_0/n3396 , \L2_0/n3392 , \L2_0/n3388 ,
         \L2_0/n3384 , \L2_0/n3380 , \L2_0/n3376 , \L2_0/n3372 , \L2_0/n3368 ,
         \L2_0/n3364 , \L2_0/n3360 , \L2_0/n3356 , \L2_0/n3352 , \L2_0/n3348 ,
         \L2_0/n3344 , \L2_0/n3336 , \L2_0/n3332 , \L2_0/n3328 , \L2_0/n3324 ,
         \L2_0/n3320 , \L2_0/n3316 , \L2_0/n3312 , \L2_0/n3308 , \L2_0/n3304 ,
         \L2_0/n3300 , \L2_0/n3296 , \L2_0/n3292 , \L2_0/n3288 , \L2_0/n3284 ,
         \L2_0/n3280 , \L2_0/n3276 , \L2_0/n3272 , \L2_0/n3268 , \L2_0/n3264 ,
         \L2_0/n3256 , \L2_0/n3252 , \L2_0/n3248 , \L2_0/n3244 , \L2_0/n3240 ,
         \L2_0/n3236 , \L2_0/n3232 , \L2_0/n3228 , \L2_0/n3224 , \L2_0/n3220 ,
         \L2_0/n3216 , \L2_0/n3212 , \L2_0/n3208 , \L2_0/n3204 , \L2_0/n3200 ,
         \L2_0/n3196 , \L2_0/n3192 , \L2_0/n3188 , \L2_0/n3184 , \L2_0/n3176 ,
         \L2_0/n3172 , \L2_0/n3168 , \L2_0/n3164 , \L2_0/n3160 , \L2_0/n3156 ,
         \L2_0/n3152 , \L2_0/n3148 , \L2_0/n3144 , \L2_0/n3140 , \L2_0/n3136 ,
         \L2_0/n3132 , \L2_0/n3128 , \L2_0/n3124 , \L2_0/n3120 , \L2_0/n3116 ,
         \L2_0/n3112 , \L2_0/n3108 , \L2_0/n3104 , \L2_0/n3096 , \L2_0/n3092 ,
         \L2_0/n3088 , \L2_0/n3084 , \L2_0/n3080 , \L2_0/n3076 , \L2_0/n3072 ,
         \L2_0/n3068 , \L2_0/n3064 , \L2_0/n3060 , \L2_0/n3056 , \L2_0/n3052 ,
         \L2_0/n3048 , \L2_0/n3044 , \L2_0/n3040 , \L2_0/n3036 , \L2_0/n3032 ,
         \L2_0/n3028 , \L2_0/n3024 , \L2_0/n3016 , \L2_0/n3012 , \L2_0/n3008 ,
         \L2_0/n3004 , \L2_0/n3000 , \L2_0/n2996 , \L2_0/n2992 , \L2_0/n2988 ,
         \L2_0/n2984 , \L2_0/n2980 , \L2_0/n2976 , \L2_0/n2972 , \L2_0/n2968 ,
         \L2_0/n2964 , \L2_0/n2960 , \L2_0/n2956 , \L2_0/n2952 , \L2_0/n2948 ,
         \L2_0/n2904 , \L2_0/n2903 , \L1_0/n4823 , \L1_0/n4822 , \L1_0/n4819 ,
         \L1_0/n4818 , \L1_0/n4815 , \L1_0/n4814 , \L1_0/n4811 , \L1_0/n4810 ,
         \L1_0/n4807 , \L1_0/n4806 , \L1_0/n4803 , \L1_0/n4802 , \L1_0/n4799 ,
         \L1_0/n4798 , \L1_0/n4795 , \L1_0/n4794 , \L1_0/n4791 , \L1_0/n4790 ,
         \L1_0/n4787 , \L1_0/n4786 , \L1_0/n4783 , \L1_0/n4782 , \L1_0/n4779 ,
         \L1_0/n4778 , \L1_0/n4775 , \L1_0/n4774 , \L1_0/n4771 , \L1_0/n4770 ,
         \L1_0/n4767 , \L1_0/n4766 , \L1_0/n4763 , \L1_0/n4762 , \L1_0/n4759 ,
         \L1_0/n4758 , \L1_0/n4755 , \L1_0/n4754 , \L1_0/n4751 , \L1_0/n4750 ,
         \L1_0/n4747 , \L1_0/n4746 , \L1_0/n4743 , \L1_0/n4742 , \L1_0/n4739 ,
         \L1_0/n4738 , \L1_0/n4735 , \L1_0/n4734 , \L1_0/n4731 , \L1_0/n4730 ,
         \L1_0/n4727 , \L1_0/n4726 , \L1_0/n4723 , \L1_0/n4722 , \L1_0/n4719 ,
         \L1_0/n4718 , \L1_0/n4715 , \L1_0/n4714 , \L1_0/n4711 , \L1_0/n4710 ,
         \L1_0/n4707 , \L1_0/n4706 , \L1_0/n4703 , \L1_0/n4702 , \L1_0/n4699 ,
         \L1_0/n4698 , \L1_0/n4695 , \L1_0/n4694 , \L1_0/n4691 , \L1_0/n4690 ,
         \L1_0/n4687 , \L1_0/n4686 , \L1_0/n4683 , \L1_0/n4682 , \L1_0/n4679 ,
         \L1_0/n4678 , \L1_0/n4675 , \L1_0/n4674 , \L1_0/n4671 , \L1_0/n4670 ,
         \L1_0/n4667 , \L1_0/n4666 , \L1_0/n4663 , \L1_0/n4662 , \L1_0/n4659 ,
         \L1_0/n4658 , \L1_0/n4655 , \L1_0/n4654 , \L1_0/n4651 , \L1_0/n4650 ,
         \L1_0/n4647 , \L1_0/n4646 , \L1_0/n4643 , \L1_0/n4642 , \L1_0/n4639 ,
         \L1_0/n4638 , \L1_0/n4635 , \L1_0/n4634 , \L1_0/n4631 , \L1_0/n4630 ,
         \L1_0/n4627 , \L1_0/n4626 , \L1_0/n4623 , \L1_0/n4622 , \L1_0/n4619 ,
         \L1_0/n4618 , \L1_0/n4615 , \L1_0/n4614 , \L1_0/n4611 , \L1_0/n4610 ,
         \L1_0/n4607 , \L1_0/n4606 , \L1_0/n4603 , \L1_0/n4602 , \L1_0/n4599 ,
         \L1_0/n4598 , \L1_0/n4595 , \L1_0/n4594 , \L1_0/n4591 , \L1_0/n4590 ,
         \L1_0/n4587 , \L1_0/n4586 , \L1_0/n4583 , \L1_0/n4582 , \L1_0/n4579 ,
         \L1_0/n4578 , \L1_0/n4575 , \L1_0/n4574 , \L1_0/n4571 , \L1_0/n4570 ,
         \L1_0/n4567 , \L1_0/n4566 , \L1_0/n4563 , \L1_0/n4562 , \L1_0/n4559 ,
         \L1_0/n4558 , \L1_0/n4555 , \L1_0/n4554 , \L1_0/n4551 , \L1_0/n4550 ,
         \L1_0/n4547 , \L1_0/n4546 , \L1_0/n4543 , \L1_0/n4542 , \L1_0/n4539 ,
         \L1_0/n4538 , \L1_0/n4535 , \L1_0/n4534 , \L1_0/n4531 , \L1_0/n4530 ,
         \L1_0/n4527 , \L1_0/n4526 , \L1_0/n4523 , \L1_0/n4522 , \L1_0/n4519 ,
         \L1_0/n4518 , \L1_0/n4515 , \L1_0/n4514 , \L1_0/n4511 , \L1_0/n4510 ,
         \L1_0/n4507 , \L1_0/n4506 , \L1_0/n4503 , \L1_0/n4502 , \L1_0/n4499 ,
         \L1_0/n4498 , \L1_0/n4495 , \L1_0/n4494 , \L1_0/n4491 , \L1_0/n4490 ,
         \L1_0/n4487 , \L1_0/n4486 , \L1_0/n4483 , \L1_0/n4482 , \L1_0/n4479 ,
         \L1_0/n4478 , \L1_0/n4475 , \L1_0/n4474 , \L1_0/n4471 , \L1_0/n4470 ,
         \L1_0/n4467 , \L1_0/n4466 , \L1_0/n4463 , \L1_0/n4462 , \L1_0/n4459 ,
         \L1_0/n4458 , \L1_0/n4455 , \L1_0/n4454 , \L1_0/n4451 , \L1_0/n4450 ,
         \L1_0/n4447 , \L1_0/n4446 , \L1_0/n4443 , \L1_0/n4442 , \L1_0/n4439 ,
         \L1_0/n4438 , \L1_0/n4435 , \L1_0/n4434 , \L1_0/n4431 , \L1_0/n4430 ,
         \L1_0/n4427 , \L1_0/n4426 , \L1_0/n4423 , \L1_0/n4422 , \L1_0/n4419 ,
         \L1_0/n4418 , \L1_0/n4415 , \L1_0/n4414 , \L1_0/n4411 , \L1_0/n4410 ,
         \L1_0/n4407 , \L1_0/n4406 , \L1_0/n4403 , \L1_0/n4402 , \L1_0/n4399 ,
         \L1_0/n4398 , \L1_0/n4395 , \L1_0/n4394 , \L1_0/n4391 , \L1_0/n4390 ,
         \L1_0/n4387 , \L1_0/n4386 , \L1_0/n4383 , \L1_0/n4382 , \L1_0/n4379 ,
         \L1_0/n4378 , \L1_0/n4375 , \L1_0/n4374 , \L1_0/n4371 , \L1_0/n4370 ,
         \L1_0/n4367 , \L1_0/n4366 , \L1_0/n4363 , \L1_0/n4362 , \L1_0/n4359 ,
         \L1_0/n4358 , \L1_0/n4355 , \L1_0/n4354 , \L1_0/n4351 , \L1_0/n4350 ,
         \L1_0/n4347 , \L1_0/n4346 , \L1_0/n4343 , \L1_0/n4342 , \L1_0/n4339 ,
         \L1_0/n4338 , \L1_0/n4335 , \L1_0/n4334 , \L1_0/n4331 , \L1_0/n4330 ,
         \L1_0/n4327 , \L1_0/n4326 , \L1_0/n4323 , \L1_0/n4322 , \L1_0/n4319 ,
         \L1_0/n4318 , \L1_0/n4315 , \L1_0/n4314 , \L1_0/n4311 , \L1_0/n4310 ,
         \L1_0/n4307 , \L1_0/n4306 , \L1_0/n4303 , \L1_0/n4302 , \L1_0/n4299 ,
         \L1_0/n4298 , \L1_0/n4295 , \L1_0/n4294 , \L1_0/n4291 , \L1_0/n4290 ,
         \L1_0/n4287 , \L1_0/n4286 , \L1_0/n4283 , \L1_0/n4282 , \L1_0/n4279 ,
         \L1_0/n4278 , \L1_0/n4275 , \L1_0/n4274 , \L1_0/n4271 , \L1_0/n4270 ,
         \L1_0/n4267 , \L1_0/n4266 , \L1_0/n4263 , \L1_0/n4262 , \L1_0/n4259 ,
         \L1_0/n4258 , \L1_0/n4255 , \L1_0/n4254 , \L1_0/n4251 , \L1_0/n4250 ,
         \L1_0/n4247 , \L1_0/n4246 , \L1_0/n4243 , \L1_0/n4242 , \L1_0/n4239 ,
         \L1_0/n4238 , \L1_0/n4235 , \L1_0/n4234 , \L1_0/n4231 , \L1_0/n4230 ,
         \L1_0/n4227 , \L1_0/n4226 , \L1_0/n4223 , \L1_0/n4222 , \L1_0/n4219 ,
         \L1_0/n4218 , \L1_0/n4215 , \L1_0/n4214 , \L1_0/n4211 , \L1_0/n4210 ,
         \L1_0/n4207 , \L1_0/n4206 , \L1_0/n4203 , \L1_0/n4202 , \L1_0/n4199 ,
         \L1_0/n4198 , \L1_0/n4195 , \L1_0/n4194 , \L1_0/n4191 , \L1_0/n4190 ,
         \L1_0/n4187 , \L1_0/n4186 , \L1_0/n4183 , \L1_0/n4182 , \L1_0/n4179 ,
         \L1_0/n4178 , \L1_0/n4175 , \L1_0/n4174 , \L1_0/n4171 , \L1_0/n4170 ,
         \L1_0/n4167 , \L1_0/n4166 , \L1_0/n4163 , \L1_0/n4162 , \L1_0/n4159 ,
         \L1_0/n4158 , \L1_0/n4155 , \L1_0/n4154 , \L1_0/n4151 , \L1_0/n4150 ,
         \L1_0/n4147 , \L1_0/n4146 , \L1_0/n4143 , \L1_0/n4142 , \L1_0/n4139 ,
         \L1_0/n4138 , \L1_0/n4135 , \L1_0/n4134 , \L1_0/n4131 , \L1_0/n4130 ,
         \L1_0/n4127 , \L1_0/n4126 , \L1_0/n4123 , \L1_0/n4122 , \L1_0/n4119 ,
         \L1_0/n4118 , \L1_0/n4115 , \L1_0/n4114 , \L1_0/n4111 , \L1_0/n4110 ,
         \L1_0/n4107 , \L1_0/n4106 , \L1_0/n4103 , \L1_0/n4102 , \L1_0/n4099 ,
         \L1_0/n4098 , \L1_0/n4095 , \L1_0/n4094 , \L1_0/n4091 , \L1_0/n4090 ,
         \L1_0/n4087 , \L1_0/n4086 , \L1_0/n4083 , \L1_0/n4082 , \L1_0/n4079 ,
         \L1_0/n4078 , \L1_0/n4075 , \L1_0/n4074 , \L1_0/n4071 , \L1_0/n4070 ,
         \L1_0/n4067 , \L1_0/n4066 , \L1_0/n4063 , \L1_0/n4062 , \L1_0/n4059 ,
         \L1_0/n4058 , \L1_0/n4055 , \L1_0/n4054 , \L1_0/n4051 , \L1_0/n4050 ,
         \L1_0/n4047 , \L1_0/n4046 , \L1_0/n4043 , \L1_0/n4042 , \L1_0/n4039 ,
         \L1_0/n4038 , \L1_0/n4035 , \L1_0/n4034 , \L1_0/n4031 , \L1_0/n4030 ,
         \L1_0/n4027 , \L1_0/n4026 , \L1_0/n4023 , \L1_0/n4022 , \L1_0/n4019 ,
         \L1_0/n4018 , \L1_0/n4015 , \L1_0/n4014 , \L1_0/n4011 , \L1_0/n4010 ,
         \L1_0/n4007 , \L1_0/n4006 , \L1_0/n4003 , \L1_0/n4002 , \L1_0/n3999 ,
         \L1_0/n3998 , \L1_0/n3995 , \L1_0/n3994 , \L1_0/n3991 , \L1_0/n3990 ,
         \L1_0/n3987 , \L1_0/n3986 , \L1_0/n3983 , \L1_0/n3982 , \L1_0/n3979 ,
         \L1_0/n3978 , \L1_0/n3975 , \L1_0/n3974 , \L1_0/n3971 , \L1_0/n3970 ,
         \L1_0/n3967 , \L1_0/n3966 , \L1_0/n3963 , \L1_0/n3962 , \L1_0/n3959 ,
         \L1_0/n3958 , \L1_0/n3955 , \L1_0/n3954 , \L1_0/n3951 , \L1_0/n3950 ,
         \L1_0/n3947 , \L1_0/n3946 , \L1_0/n3943 , \L1_0/n3942 , \L1_0/n3939 ,
         \L1_0/n3938 , \L1_0/n3935 , \L1_0/n3934 , \L1_0/n3931 , \L1_0/n3930 ,
         \L1_0/n3927 , \L1_0/n3926 , \L1_0/n3923 , \L1_0/n3922 , \L1_0/n3919 ,
         \L1_0/n3918 , \L1_0/n3915 , \L1_0/n3914 , \L1_0/n3911 , \L1_0/n3910 ,
         \L1_0/n3907 , \L1_0/n3906 , \L1_0/n3903 , \L1_0/n3902 , \L1_0/n3899 ,
         \L1_0/n3898 , \L1_0/n3895 , \L1_0/n3894 , \L1_0/n3891 , \L1_0/n3890 ,
         \L1_0/n3887 , \L1_0/n3886 , \L1_0/n3883 , \L1_0/n3882 , \L1_0/n3879 ,
         \L1_0/n3878 , \L1_0/n3875 , \L1_0/n3874 , \L1_0/n3871 , \L1_0/n3870 ,
         \L1_0/n3867 , \L1_0/n3866 , \L1_0/n3863 , \L1_0/n3862 , \L1_0/n3859 ,
         \L1_0/n3858 , \L1_0/n3855 , \L1_0/n3854 , \L1_0/n3851 , \L1_0/n3850 ,
         \L1_0/n3847 , \L1_0/n3846 , \L1_0/n3843 , \L1_0/n3842 , \L1_0/n3839 ,
         \L1_0/n3838 , \L1_0/n3835 , \L1_0/n3834 , \L1_0/n3831 , \L1_0/n3830 ,
         \L1_0/n3827 , \L1_0/n3826 , \L1_0/n3823 , \L1_0/n3822 , \L1_0/n3819 ,
         \L1_0/n3818 , \L1_0/n3815 , \L1_0/n3814 , \L1_0/n3811 , \L1_0/n3810 ,
         \L1_0/n3807 , \L1_0/n3806 , \L1_0/n3803 , \L1_0/n3802 , \L1_0/n3799 ,
         \L1_0/n3798 , \L1_0/n3795 , \L1_0/n3794 , \L1_0/n3791 , \L1_0/n3790 ,
         \L1_0/n3787 , \L1_0/n3786 , \L1_0/n3783 , \L1_0/n3782 , \L1_0/n3779 ,
         \L1_0/n3778 , \L1_0/n3775 , \L1_0/n3774 , \L1_0/n3771 , \L1_0/n3770 ,
         \L1_0/n3767 , \L1_0/n3766 , \L1_0/n3763 , \L1_0/n3762 , \L1_0/n3759 ,
         \L1_0/n3758 , \L1_0/n3755 , \L1_0/n3754 , \L1_0/n3751 , \L1_0/n3750 ,
         \L1_0/n3747 , \L1_0/n3746 , \L1_0/n3743 , \L1_0/n3742 , \L1_0/n3739 ,
         \L1_0/n3738 , \L1_0/n3735 , \L1_0/n3734 , \L1_0/n3731 , \L1_0/n3730 ,
         \L1_0/n3727 , \L1_0/n3726 , \L1_0/n3723 , \L1_0/n3722 , \L1_0/n3719 ,
         \L1_0/n3718 , \L1_0/n3715 , \L1_0/n3714 , \L1_0/n3711 , \L1_0/n3710 ,
         \L1_0/n3707 , \L1_0/n3706 , \L1_0/n3703 , \L1_0/n3702 , \L1_0/n3699 ,
         \L1_0/n3698 , \L1_0/n3695 , \L1_0/n3694 , \L1_0/n3691 , \L1_0/n3690 ,
         \L1_0/n3687 , \L1_0/n3686 , \L1_0/n3683 , \L1_0/n3682 , \L1_0/n3679 ,
         \L1_0/n3678 , \L1_0/n3675 , \L1_0/n3674 , \L1_0/n3671 , \L1_0/n3670 ,
         \L1_0/n3667 , \L1_0/n3666 , \L1_0/n3663 , \L1_0/n3662 , \L1_0/n3659 ,
         \L1_0/n3658 , \L1_0/n3655 , \L1_0/n3654 , \L1_0/n3651 , \L1_0/n3650 ,
         \L1_0/n3647 , \L1_0/n3646 , \L1_0/n3643 , \L1_0/n3642 , \L1_0/n3639 ,
         \L1_0/n3638 , \L1_0/n3635 , \L1_0/n3634 , \L1_0/n3631 , \L1_0/n3630 ,
         \L1_0/n3627 , \L1_0/n3626 , \L1_0/n3623 , \L1_0/n3622 , \L1_0/n3619 ,
         \L1_0/n3618 , \L1_0/n3615 , \L1_0/n3614 , \L1_0/n3611 , \L1_0/n3610 ,
         \L1_0/n3607 , \L1_0/n3606 , \L1_0/n3603 , \L1_0/n3602 , \L1_0/n3599 ,
         \L1_0/n3598 , \L1_0/n3595 , \L1_0/n3594 , \L1_0/n3591 , \L1_0/n3590 ,
         \L1_0/n3587 , \L1_0/n3586 , \L1_0/n3583 , \L1_0/n3582 , \L1_0/n3579 ,
         \L1_0/n3578 , \L1_0/n3575 , \L1_0/n3574 , \L1_0/n3571 , \L1_0/n3570 ,
         \L1_0/n3567 , \L1_0/n3566 , \L1_0/n3563 , \L1_0/n3562 , \L1_0/n3559 ,
         \L1_0/n3558 , \L1_0/n3555 , \L1_0/n3554 , \L1_0/n3551 , \L1_0/n3550 ,
         \L1_0/n3507 , \L1_0/n3506 , n40519, n40520, n40521, n40522, n40523,
         n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531,
         n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539,
         n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547,
         n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
         n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
         n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
         n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
         n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587,
         n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
         n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603,
         n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611,
         n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
         n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
         n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
         n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
         n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
         n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659,
         n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667,
         n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675,
         n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683,
         n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691,
         n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
         n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
         n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
         n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723,
         n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731,
         n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739,
         n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747,
         n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755,
         n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763,
         n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
         n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779,
         n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
         n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795,
         n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803,
         n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
         n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819,
         n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827,
         n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835,
         n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
         n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851,
         n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
         n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867,
         n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875,
         n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
         n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891,
         n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
         n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907,
         n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
         n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923,
         n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
         n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
         n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947,
         n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
         n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963,
         n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971,
         n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979,
         n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
         n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995,
         n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
         n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
         n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019,
         n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027,
         n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035,
         n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043,
         n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051,
         n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
         n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067,
         n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
         n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083,
         n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091,
         n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099,
         n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107,
         n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115,
         n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123,
         n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
         n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139,
         n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
         n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155,
         n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163,
         n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171,
         n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179,
         n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
         n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195,
         n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
         n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211,
         n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
         n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227,
         n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235,
         n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243,
         n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251,
         n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259,
         n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267,
         n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
         n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283,
         n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
         n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299,
         n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307,
         n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
         n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323,
         n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
         n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339,
         n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
         n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355,
         n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
         n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371,
         n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379,
         n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387,
         n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395,
         n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403,
         n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411,
         n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419,
         n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427,
         n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435,
         n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443,
         n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451,
         n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459,
         n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467,
         n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475,
         n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483,
         n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491,
         n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499,
         n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
         n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515,
         n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523,
         n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531,
         n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539,
         n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547,
         n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555,
         n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563,
         n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
         n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579,
         n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587,
         n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595,
         n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603,
         n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611,
         n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619,
         n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627,
         n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
         n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643,
         n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
         n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659,
         n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667,
         n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675,
         n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683,
         n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691,
         n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699,
         n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707,
         n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715,
         n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723,
         n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731,
         n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739,
         n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747,
         n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755,
         n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763,
         n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771,
         n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779,
         n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787,
         n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
         n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
         n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811,
         n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819,
         n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827,
         n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835,
         n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843,
         n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851,
         n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859,
         n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867,
         n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875,
         n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883,
         n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
         n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899,
         n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907,
         n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915,
         n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
         n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931,
         n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
         n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
         n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955,
         n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963,
         n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971,
         n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979,
         n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987,
         n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995,
         n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003,
         n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011,
         n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019,
         n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027,
         n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035,
         n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043,
         n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051,
         n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059,
         n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
         n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075,
         n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083,
         n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091,
         n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099,
         n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107,
         n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115,
         n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123,
         n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131,
         n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139,
         n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147,
         n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
         n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163,
         n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171,
         n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179,
         n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187,
         n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195,
         n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203,
         n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211,
         n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219,
         n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
         n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235,
         n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243,
         n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251,
         n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259,
         n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267,
         n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275,
         n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283,
         n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291,
         n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
         n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
         n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315,
         n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323,
         n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331,
         n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339,
         n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347,
         n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
         n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363,
         n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371,
         n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379,
         n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387,
         n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395,
         n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403,
         n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411,
         n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419,
         n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427,
         n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435,
         n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
         n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451,
         n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459,
         n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467,
         n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475,
         n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483,
         n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491,
         n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
         n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507,
         n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
         n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
         n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531,
         n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539,
         n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547,
         n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555,
         n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563,
         n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
         n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579,
         n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587,
         n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595,
         n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603,
         n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611,
         n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619,
         n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627,
         n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635,
         n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643,
         n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651,
         n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659,
         n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667,
         n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675,
         n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683,
         n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691,
         n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699,
         n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707,
         n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715,
         n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723,
         n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731,
         n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739,
         n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747,
         n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755,
         n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763,
         n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771,
         n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779,
         n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787,
         n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795,
         n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803,
         n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811,
         n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819,
         n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827,
         n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835,
         n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843,
         n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851,
         n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859,
         n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867,
         n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875,
         n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883,
         n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891,
         n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899,
         n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907,
         n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915,
         n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923,
         n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931,
         n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939,
         n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947,
         n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955,
         n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963,
         n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971,
         n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979,
         n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987,
         n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995,
         n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
         n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011,
         n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
         n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027,
         n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035,
         n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043,
         n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051,
         n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059,
         n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067,
         n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
         n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083,
         n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
         n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099,
         n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107,
         n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115,
         n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123,
         n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131,
         n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139,
         n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
         n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155,
         n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
         n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171,
         n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179,
         n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187,
         n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195,
         n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203,
         n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211,
         n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
         n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227,
         n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
         n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
         n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251,
         n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259,
         n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267,
         n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275,
         n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283,
         n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
         n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299,
         n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
         n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315,
         n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323,
         n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
         n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339,
         n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347,
         n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355,
         n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
         n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371,
         n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
         n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387,
         n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395,
         n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
         n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411,
         n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419,
         n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427,
         n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
         n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443,
         n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
         n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459,
         n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467,
         n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475,
         n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483,
         n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491,
         n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499,
         n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
         n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515,
         n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
         n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531,
         n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539,
         n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547,
         n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555,
         n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563,
         n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571,
         n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
         n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
         n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
         n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603,
         n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611,
         n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
         n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
         n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
         n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643,
         n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
         n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659,
         n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
         n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
         n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683,
         n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
         n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699,
         n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707,
         n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
         n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
         n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731,
         n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
         n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747,
         n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
         n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
         n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771,
         n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779,
         n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787,
         n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
         n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803,
         n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
         n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819,
         n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827,
         n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
         n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
         n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851,
         n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859,
         n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
         n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875,
         n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
         n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891,
         n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899,
         n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
         n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915,
         n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923,
         n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931,
         n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
         n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947,
         n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
         n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963,
         n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
         n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
         n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987,
         n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995,
         n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003,
         n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
         n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019,
         n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
         n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035,
         n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043,
         n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
         n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059,
         n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067,
         n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075,
         n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
         n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091,
         n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
         n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107,
         n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115,
         n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
         n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131,
         n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139,
         n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147,
         n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
         n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163,
         n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
         n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179,
         n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187,
         n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
         n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
         n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211,
         n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219,
         n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
         n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235,
         n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
         n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251,
         n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259,
         n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
         n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275,
         n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283,
         n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291,
         n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
         n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307,
         n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
         n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323,
         n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331,
         n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
         n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347,
         n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355,
         n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363,
         n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
         n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379,
         n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
         n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
         n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403,
         n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
         n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419,
         n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427,
         n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435,
         n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
         n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451,
         n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
         n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467,
         n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475,
         n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
         n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491,
         n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499,
         n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507,
         n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
         n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523,
         n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
         n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539,
         n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547,
         n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
         n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563,
         n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571,
         n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579,
         n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
         n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595,
         n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
         n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611,
         n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619,
         n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
         n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635,
         n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643,
         n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651,
         n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
         n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667,
         n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
         n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683,
         n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691,
         n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
         n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707,
         n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715,
         n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723,
         n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
         n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739,
         n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
         n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755,
         n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763,
         n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
         n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779,
         n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787,
         n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795,
         n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
         n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811,
         n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
         n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827,
         n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835,
         n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
         n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851,
         n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859,
         n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867,
         n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
         n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883,
         n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
         n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899,
         n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907,
         n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
         n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923,
         n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931,
         n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939,
         n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
         n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955,
         n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
         n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971,
         n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979,
         n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
         n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995,
         n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003,
         n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011,
         n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
         n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027,
         n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
         n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043,
         n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051,
         n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
         n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067,
         n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075,
         n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083,
         n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
         n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099,
         n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
         n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115,
         n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123,
         n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
         n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139,
         n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147,
         n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155,
         n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
         n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171,
         n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
         n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187,
         n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195,
         n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
         n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211,
         n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219,
         n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227,
         n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
         n45236, n45237, n45238, n45240, n45241, n45242, n45243, n45244,
         n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252,
         n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260,
         n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268,
         n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276,
         n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284,
         n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292,
         n45293, n45294, n45295, n45296, n45297, n45298, n45299, n45300,
         n45301, n45302, n45303, n45304, n45305, n45306, n45307, n45308,
         n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316,
         n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324,
         n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332,
         n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340,
         n45341, n45342, n45343, n45344, n45345, n45346, n45347, n45348,
         n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356,
         n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364,
         n45365, n45366, n45367, n45368, n45369, n45370, n45371, n45372,
         n45373, n45374, n45375, n45376, n45377, n45378, n45379, n45380,
         n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388,
         n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396,
         n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404,
         n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412,
         n45413, n45414, n45415, n45416, n45417, n45418, n45419, n45420,
         n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428,
         n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436,
         n45437, n45438, n45439, n45440, n45441, n45442, n45443, n45444,
         n45445, n45446, n45447, n45448, n45449, n45450, n45451, n45452,
         n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460,
         n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468,
         n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476,
         n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484,
         n45485, n45486, n45487, n45488, n45489, n45490, n45491, n45492,
         n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500,
         n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508,
         n45509, n45510, n45511, n45512, n45513, n45514, n45515, n45516,
         n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524,
         n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532,
         n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540,
         n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548,
         n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556,
         n45557, n45558, n45559, n45560, n45561, n45562, n45563, n45564,
         n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572,
         n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580,
         n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588,
         n45589, n45590, n45591, n45592, n45593, n45594, n45595, n45596,
         n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604,
         n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612,
         n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620,
         n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628,
         n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636,
         n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644,
         n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652,
         n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660,
         n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668,
         n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676,
         n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684,
         n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692,
         n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700,
         n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708,
         n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716,
         n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724,
         n45725, n45726, n45727, n45728, n45729, n45730, n45731, n45732,
         n45733, n45734, n45735, n45736, n45737, n45738, n45739, n45740,
         n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748,
         n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756,
         n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764,
         n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772,
         n45773, n45774, n45775, n45776, n45777, n45778, n45779, n45780,
         n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788,
         n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796,
         n45797, n45798, n45799, n45800, n45801, n45802, n45803, n45804,
         n45805, n45806, n45807, n45808, n45809, n45810, n45811, n45812,
         n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820,
         n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828,
         n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836,
         n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844,
         n45845, n45846, n45847, n45848, n45849, n45850, n45851, n45852,
         n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860,
         n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868,
         n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876,
         n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884,
         n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892,
         n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900,
         n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908,
         n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916,
         n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924,
         n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932,
         n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940,
         n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948,
         n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956,
         n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964,
         n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972,
         n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980,
         n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988,
         n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996,
         n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004,
         n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012,
         n46013, n46014, n46015, n46016, n46017, n46018, n46019, n46020,
         n46021, n46022, n46023, n46024, n46025, n46026, n46027, n46028,
         n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036,
         n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044,
         n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052,
         n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060,
         n46061, n46062, n46063, n46064, n46065, n46066, n46067, n46068,
         n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076,
         n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084,
         n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092,
         n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100,
         n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108,
         n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116,
         n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124,
         n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132,
         n46133, n46134, n46135, n46136, n46137, n46138, n46139, n46140,
         n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148,
         n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156,
         n46157, n46158, n46159, n46160, n46161, n46162, n46163, n46164,
         n46165, n46166, n46167, n46168, n46169, n46170, n46171, n46172,
         n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180,
         n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188,
         n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197,
         n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205,
         n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213,
         n46214, n46215, n46216, n46217, n46218, n46219, n46220, n46221,
         n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229,
         n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237,
         n46238, n46239, n46240, n46241, n46242, n46243, n46244, n46245,
         n46246, n46247, n46248, n46249, n46250, n46251, n46252, n46253,
         n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261,
         n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269,
         n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277,
         n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285,
         n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293,
         n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301,
         n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309,
         n46310, n46311, n46312, n46313, n46314, n46315, n46316, n46317,
         n46318, n46319, n46320, n46321, n46322, n46323, n46324, n46325,
         n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333,
         n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341,
         n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349,
         n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357,
         n46358, n46359, n46360, n46361, n46362, n46363, n46364, n46365,
         n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373,
         n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381,
         n46382, n46383, n46384, n46385, n46386, n46387, n46388, n46389,
         n46390, n46391, n46392, n46393, n46394, n46395, n46396, n46397,
         n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405,
         n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413,
         n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421,
         n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429,
         n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437,
         n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445,
         n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453,
         n46454, n46455, n46456, n46457, n46458, n46459, n46460, n46461,
         n46462, n46463, n46464, n46465, n46466, n46467, n46468, n46469,
         n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477,
         n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485,
         n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493,
         n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501,
         n46502, n46503, n46504, n46505, n46506, n46507, n46508, n46509,
         n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517,
         n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525,
         n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533,
         n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541,
         n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549,
         n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557,
         n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565,
         n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573,
         n46574, n46575, n46576, n46577, n46578, n46579, n46580, n46581,
         n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589,
         n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597,
         n46598, n46599, n46600, n46601, n46602, n46603, n46604, n46605,
         n46606, n46607, n46608, n46609, n46610, n46611, n46612, n46613,
         n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621,
         n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629,
         n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637,
         n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645,
         n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653,
         n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661,
         n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669,
         n46670, n46671, n46672, n46673, n49249, n49250, n49251, n49252,
         n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260,
         n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268,
         n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276,
         n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284,
         n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292,
         n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300,
         n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308,
         n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316,
         n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324,
         n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332,
         n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340,
         n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348,
         n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356,
         n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364,
         n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372,
         n49373, n49374, n49375, n49376, n49377, n49378, n49379, n49380,
         n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388,
         n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396,
         n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404,
         n49405, n49406, n49407, n49408, n49409, n49410, n49411, n49412,
         n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420,
         n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428,
         n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436,
         n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444,
         n49445, n49446, n49447, n49448, n49449, n49450, n49451, n49452,
         n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460,
         n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468,
         n49469, n49470, n49471, n49472, n49473, n49474, n49475, n49476,
         n49477, n49478, n49479, n49480, n49481, n49482, n49483, n49484,
         n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492,
         n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500,
         n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508,
         n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516,
         n49517, n49518, n49519, n49520, n49521, n49522, n49523, n49524,
         n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532,
         n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540,
         n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548,
         n49549, n49550, n49551, n49552, n49553, n49554, n49555, n49556,
         n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564,
         n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572,
         n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580,
         n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588,
         n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596,
         n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604,
         n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612,
         n49613, n49614, n49615, n49616, n49617, n49618, n49619, n49620,
         n49621, n49622, n49623, n49624, n49625, n49626, n49627, n49628,
         n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636,
         n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644,
         n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652,
         n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660,
         n49661, n49662, n49663, n49664, n49665, n49666, n49667, n49668,
         n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676,
         n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684,
         n49685, n49686, n49687, n49688, n49689, n49690, n49691, n49692,
         n49693, n49694, n49695, n49696, n49697, n49698, n49699, n49700,
         n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708,
         n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716,
         n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724,
         n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732,
         n49733, n49734, n49735, n49736, n49737, n49738, n49739, n49740,
         n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748,
         n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756,
         n49757, n49758, n49759, n49760, n49761, n49762, n49763, n49764,
         n49765, n49766, n49767, n49768, n49769, n49770, n49771, n49772,
         n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780,
         n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788,
         n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796,
         n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804,
         n49805, n49806, n49807, n49808, n49809, n49810, n49811, n49812,
         n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820,
         n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828,
         n49829, n49830, n49831, n49832, n49833, n49834, n49835, n49836,
         n49837, n49838, n49839, n49840, n49841, n49842, n49843, n49844,
         n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852,
         n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860,
         n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868,
         n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876,
         n49877, n49878, n49879, n49880, n49881, n49882, n49883, n49884,
         n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892,
         n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900,
         n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908,
         n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916,
         n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924,
         n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932,
         n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940,
         n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948,
         n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956,
         n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964,
         n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972,
         n49973, n49974, n49975, n49976, n49977, n49978, n49979, n49980,
         n49981, n49982, n49983, n49984, n49985, n49986, n49987, n49988,
         n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996,
         n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004,
         n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012,
         n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020,
         n50021, n50022, n50023, n50024, n50025, n50026, n50027, n50028,
         n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036,
         n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044,
         n50045, n50046, n50047, n50048, n50049, n50050, n50051, n50052,
         n50053, n50054, n50055, n50056, n50057, n50058, n50059, n50060,
         n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068,
         n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076,
         n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084,
         n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092,
         n50093, n50094, n50095, n50096, n50097, n50098, n50099, n50100,
         n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108,
         n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116,
         n50117, n50118, n50119, n50120, n50121, n50122, n50123, n50124,
         n50125, n50126, n50127, n50128, n50129, n50130, n50131, n50132,
         n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140,
         n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148,
         n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156,
         n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164,
         n50165, n50166, n50167, n50168, n50169, n50170, n50171, n50172,
         n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180,
         n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188,
         n50189, n50190, n50191, n50192, n50193, n50194, n50195, n50196,
         n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204,
         n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212,
         n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220,
         n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228,
         n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236,
         n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244,
         n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252,
         n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260,
         n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268,
         n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276,
         n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284,
         n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292,
         n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300,
         n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308,
         n50309, n50310, n50311, n50312, n50313, n50314, n50315, n50316,
         n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324,
         n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332,
         n50333, n50334, n50335, n50336, n50337, n50338, n50339, n50340,
         n50341, n50342, n50343, n50344, n50345, n50346, n50347, n50348,
         n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356,
         n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364,
         n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372,
         n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380,
         n50381, n50382, n50383, n50384, n50385, n50386, n50387, n50388,
         n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396,
         n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404,
         n50405, n50406, n50407, n50408, n50409, n50410, n50411, n50412,
         n50413, n50414, n50415, n50416, n50417, n50418, n50419, n50420,
         n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428,
         n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436,
         n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444,
         n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452,
         n50453, n50454, n50455, n50456, n50457, n50458, n50459, n50460,
         n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468,
         n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476,
         n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484,
         n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492,
         n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500,
         n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508,
         n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516,
         n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524,
         n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532,
         n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540,
         n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548,
         n50549, n50550, n50551, n50552, n50553, n50554, n50555, n50556,
         n50557, n50558, n50559, n50560, n50561, n50562, n50563, n50564,
         n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572,
         n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580,
         n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588,
         n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596,
         n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604,
         n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612,
         n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620,
         n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628,
         n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636,
         n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644,
         n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652,
         n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660,
         n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668,
         n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676,
         n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684,
         n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692,
         n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700,
         n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708,
         n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716,
         n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724,
         n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732,
         n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740,
         n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748,
         n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756,
         n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764,
         n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772,
         n50773, n50774, n50775, n50776, n50777, n50778, n50779, n50780,
         n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788,
         n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796,
         n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804,
         n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812,
         n50813, n50814, n50815, n50816, n50817, n50818, n50819, n50820,
         n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828,
         n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836,
         n50837, n50838, n50839, n50840, n50841, n50842, n50843, n50844,
         n50845, n50846, n50847, n50848, n50849, n50850, n50851, n50852,
         n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860,
         n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868,
         n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876,
         n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884,
         n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892,
         n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900,
         n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908,
         n50909, n50910, n50911, n50912, n50913, n50914, n50915, n50916,
         n50917, n50918, n50919, n50920, n50921, n50922, n50923, n50924,
         n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932,
         n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940,
         n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948,
         n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956,
         n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964,
         n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972,
         n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980,
         n50981, n50982, n50983, n50984, n50985, n50986, n50987, n50988,
         n50989, n50990, n50991, n50992, n50993, n50994, n50995, n50996,
         n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004,
         n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012,
         n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020,
         n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028,
         n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036,
         n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044,
         n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052,
         n51053, n51054, n51055, n51056, n51057, n51058, n51059, n51060,
         n51061, n51062, n51063, n51064, n51065, n51066, n51067, n51068,
         n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076,
         n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084,
         n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092,
         n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100,
         n51101, n51102, n51103, n51104, n51105, n51106, n51107, n51108,
         n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116,
         n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124,
         n51125, n51126, n51127, n51128, n51129, n51130, n51131, n51132,
         n51133, n51134, n51135, n51136, n51137, n51138, n51139, n51140,
         n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148,
         n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156,
         n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164,
         n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172,
         n51173, n51174, n51175, n51176, n51177, n51178, n51179, n51180,
         n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188,
         n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196,
         n51197, n51198, n51199, n51200, n51201, n51202, n51203, n51204,
         n51205, n51206, n51207, n51208, n51209, n51210, n51211, n51212,
         n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220,
         n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228,
         n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236,
         n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244,
         n51245, n51246, n51247, n51248, n51249, n51250, n51251, n51252,
         n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260,
         n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268,
         n51269, n51270, n51271, n51272, n51273, n51274, n51275, n51276,
         n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284,
         n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292,
         n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300,
         n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308,
         n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316,
         n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324,
         n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332,
         n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340,
         n51341, n51342, n51343, n51344, n51345, n51346, n51347, n51348,
         n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356,
         n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364,
         n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372,
         n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380,
         n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388,
         n51389, n51390, n51391, n51392, n51393, n51394, n51395, n51396,
         n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404,
         n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412,
         n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420,
         n51421, n51422, n51423, n51424, n51425, n51426, n51427, n51428,
         n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436,
         n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444,
         n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452,
         n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460,
         n51461, n51462, n51463, n51464, n51465, n51466, n51467, n51468,
         n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476,
         n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484,
         n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492,
         n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500,
         n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508,
         n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516,
         n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524,
         n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532,
         n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540,
         n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548,
         n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556,
         n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51564,
         n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572,
         n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580,
         n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588,
         n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596,
         n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604,
         n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612,
         n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620,
         n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628,
         n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636,
         n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644,
         n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652,
         n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660,
         n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668,
         n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676,
         n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684,
         n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692,
         n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700,
         n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708,
         n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716,
         n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724,
         n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732,
         n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740,
         n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748,
         n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756,
         n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764,
         n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772,
         n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780,
         n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788,
         n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796,
         n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804,
         n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812,
         n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820,
         n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828,
         n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836,
         n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844,
         n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852,
         n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860,
         n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868,
         n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876,
         n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884,
         n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892,
         n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900,
         n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908,
         n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916,
         n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924,
         n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932,
         n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940,
         n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948,
         n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956,
         n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964,
         n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972,
         n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980,
         n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988,
         n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996,
         n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004,
         n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012,
         n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020,
         n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028,
         n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036,
         n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044,
         n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052,
         n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060,
         n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068,
         n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076,
         n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084,
         n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092,
         n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100,
         n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108,
         n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116,
         n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124,
         n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132,
         n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140,
         n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148,
         n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156,
         n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164,
         n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172,
         n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180,
         n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188,
         n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196,
         n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204,
         n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212,
         n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220,
         n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228,
         n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236,
         n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244,
         n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252,
         n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260,
         n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268,
         n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276,
         n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284,
         n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292,
         n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
         n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308,
         n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316,
         n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324,
         n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332,
         n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340,
         n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348,
         n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356,
         n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364,
         n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372,
         n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380,
         n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388,
         n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396,
         n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404,
         n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412,
         n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420,
         n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428,
         n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436,
         n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444,
         n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452,
         n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460,
         n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468,
         n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476,
         n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484,
         n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492,
         n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500,
         n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508,
         n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
         n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524,
         n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532,
         n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540,
         n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548,
         n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556,
         n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564,
         n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572,
         n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580,
         n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
         n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596,
         n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604,
         n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612,
         n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620,
         n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628,
         n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636,
         n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644,
         n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652,
         n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660,
         n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668,
         n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676,
         n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684,
         n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692,
         n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700,
         n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708,
         n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716,
         n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724,
         n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732,
         n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740,
         n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748,
         n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756,
         n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764,
         n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772,
         n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780,
         n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788,
         n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796,
         n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804,
         n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812,
         n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820,
         n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828,
         n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836,
         n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844,
         n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852,
         n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860,
         n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868,
         n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876,
         n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884,
         n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892,
         n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900,
         n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908,
         n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916,
         n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924,
         n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932,
         n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940,
         n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948,
         n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956,
         n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964,
         n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972,
         n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980,
         n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988,
         n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996,
         n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004,
         n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012,
         n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020,
         n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028,
         n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036,
         n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044,
         n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052,
         n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060,
         n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068,
         n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076,
         n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084,
         n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
         n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100,
         n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
         n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116,
         n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124,
         n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132,
         n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140,
         n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148,
         n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156,
         n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164,
         n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172,
         n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180,
         n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188,
         n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196,
         n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204,
         n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212,
         n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220,
         n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228,
         n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
         n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244,
         n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252,
         n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260,
         n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268,
         n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276,
         n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284,
         n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292,
         n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300,
         n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308,
         n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316,
         n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324,
         n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332,
         n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340,
         n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348,
         n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356,
         n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364,
         n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372,
         n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380,
         n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388,
         n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396,
         n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404,
         n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412,
         n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420,
         n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428,
         n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436,
         n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444,
         n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452,
         n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460,
         n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468,
         n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476,
         n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484,
         n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492,
         n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500,
         n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508,
         n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516,
         n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524,
         n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532,
         n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540,
         n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548,
         n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556,
         n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564,
         n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572,
         n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580,
         n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588,
         n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596,
         n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604,
         n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612,
         n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620,
         n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628,
         n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636,
         n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644,
         n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652,
         n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660,
         n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668,
         n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676,
         n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684,
         n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692,
         n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700,
         n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708,
         n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716,
         n53717, n53718, n53719, n53720, n53721, n53722, n53723, n53724,
         n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732,
         n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740,
         n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748,
         n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756,
         n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764,
         n53765, n53766, n53767, n53768, n53769, n53770, n53771, n53772,
         n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780,
         n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788,
         n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796,
         n53797, n53798, n53799, n53800, n53801, n53802, n53803, n53804,
         n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812,
         n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820,
         n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828,
         n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836,
         n53837, n53838, n53839, n53840, n53841, n53842, n53843, n53844,
         n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852,
         n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860,
         n53861, n53862, n53863, n53864, n53865, n53866, n53867, n53868,
         n53869, n53870, n53871, n53872, n53873, n53874, n53875, n53876,
         n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884,
         n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892,
         n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900,
         n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908,
         n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916,
         n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924,
         n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932,
         n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940,
         n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948,
         n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956,
         n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964,
         n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972,
         n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980,
         n53981, n53982, n53983, n53984, n53985, n53986, n53987, n53988,
         n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996,
         n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004,
         n54005, n54006, n54007, n54008, n54009, n54010, n54011, n54012,
         n54013, n54014, n54015, n54016, n54017, n54018, n54019, n54020,
         n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028,
         n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036,
         n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044,
         n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052,
         n54053, n54054, n54055, n54056, n54057, n54058, n54059, n54060,
         n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068,
         n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076,
         n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084,
         n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092,
         n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100,
         n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108,
         n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116,
         n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124,
         n54125, n54126, n54127, n54128, n54129, n54130, n54131, n54132,
         n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140,
         n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148,
         n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156,
         n54157, n54158, n54159, n54160, n54161, n54162, n54163, n54164,
         n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172,
         n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180,
         n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188,
         n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196,
         n54197, n54198, n54199, n54200, n54201, n54202, n54203, n54204,
         n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212,
         n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220,
         n54221, n54222, n54223, n54224, n54225, n54226, n54227, n54228,
         n54229, n54230, n54231, n54232, n54233, n54234, n54235, n54236,
         n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244,
         n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252,
         n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260,
         n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268,
         n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276,
         n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284,
         n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292,
         n54293, n54294, n54295, n54296, n54297, n54298, n54299, n54300,
         n54301, n54302, n54303, n54304, n54305, n54306, n54307, n54308,
         n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316,
         n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324,
         n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332,
         n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340,
         n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348,
         n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356,
         n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364,
         n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372,
         n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380,
         n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388,
         n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396,
         n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404,
         n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412,
         n54413, n54414, n54415, n54416, n54417, n54418, n54419, n54420,
         n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428,
         n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436,
         n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444,
         n54445, n54446, n54447, n54448, n54449, n54450, n54451, n54452,
         n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460,
         n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468,
         n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476,
         n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484,
         n54485, n54486, n54487, n54488, n54489, n54490, n54491, n54492,
         n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500,
         n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508,
         n54509, n54510, n54511, n54512, n54513, n54514, n54515, n54516,
         n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524,
         n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532,
         n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540,
         n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548,
         n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556,
         n54557, n54558, n54559, n54560, n54561, n54562, n54563, n54564,
         n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572,
         n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580,
         n54581, n54582, n54583, n54584, n54585, n54586, n54587, n54588,
         n54589, n54590, n54591, n54592, n54593, n54594, n54595, n54596,
         n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604,
         n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612,
         n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620,
         n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628,
         n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636,
         n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644,
         n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652,
         n54653, n54654, n54655, n54656, n54657, n54658, n54659, n54660,
         n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668,
         n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676,
         n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684,
         n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692,
         n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700,
         n54701, n54702, n54703, n54704, n54705, n54706, n54707, n54708,
         n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716,
         n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724,
         n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732,
         n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740,
         n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748,
         n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756,
         n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764,
         n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772,
         n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780,
         n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788,
         n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796,
         n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804,
         n54805, n54806, n54807, n54808, n54809, n54810, n54811, n54812,
         n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820,
         n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828,
         n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836,
         n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844,
         n54845, n54846, n54847, n54848, n54849, n54850, n54851, n54852,
         n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860,
         n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868,
         n54869, n54870, n54871, n54872, n54873, n54874, n54875, n54876,
         n54877, n54878, n54879, n54880, n54881, n54882, n54883, n54884,
         n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892,
         n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900,
         n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908,
         n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916,
         n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924,
         n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932,
         n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940,
         n54941, n54942, n54943, n54944, n54945, n54946, n54947, n54948,
         n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956,
         n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964,
         n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972,
         n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980,
         n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988,
         n54989, n54990, n54991, n54992, n54993, n54994, n54995, n54996,
         n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004,
         n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012,
         n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020,
         n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028,
         n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036,
         n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044,
         n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052,
         n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060,
         n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068,
         n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076,
         n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084,
         n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092,
         n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100,
         n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108,
         n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116,
         n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124,
         n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132,
         n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140,
         n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148,
         n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156,
         n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164,
         n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172,
         n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180,
         n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188,
         n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196,
         n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204,
         n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212,
         n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220,
         n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228,
         n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236,
         n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244,
         n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252,
         n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260,
         n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268,
         n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276,
         n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284,
         n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292,
         n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300,
         n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308,
         n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316,
         n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324,
         n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332,
         n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340,
         n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348,
         n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356,
         n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364,
         n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372,
         n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380,
         n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388,
         n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396,
         n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404,
         n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412,
         n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420,
         n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428,
         n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436,
         n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444,
         n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452,
         n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460,
         n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468,
         n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476,
         n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484,
         n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492,
         n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500,
         n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508,
         n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516,
         n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524,
         n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532,
         n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540,
         n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548,
         n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556,
         n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564,
         n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572,
         n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580,
         n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588,
         n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596,
         n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604,
         n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612,
         n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620,
         n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628,
         n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636,
         n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644,
         n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652,
         n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660,
         n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668,
         n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676,
         n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684,
         n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692,
         n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700,
         n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708,
         n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716,
         n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724,
         n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732,
         n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740,
         n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748,
         n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756,
         n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764,
         n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772,
         n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780,
         n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788,
         n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796,
         n55797;
  wire   [3:0] reg_num;
  wire   [19:0] out_L1;
  wire   [19:0] out_L2;

  dff_sg done_reg ( .D(n55795), .CP(clk), .Q(done) );
  dff_sg \state_reg[1]  ( .D(n40518), .CP(clk), .Q(n55798) );
  dff_sg \state_reg[0]  ( .D(n40517), .CP(clk), .Q(n55799) );
  dff_sg \reg_num_reg[3]  ( .D(n1358), .CP(clk), .Q(reg_num[3]) );
  dff_sg \reg_num_reg[2]  ( .D(n1359), .CP(clk), .Q(reg_num[2]) );
  dff_sg \reg_num_reg[1]  ( .D(n1360), .CP(clk), .Q(reg_num[1]) );
  dff_sg \reg_num_reg[0]  ( .D(n1361), .CP(clk), .Q(reg_num[0]) );
  dff_sg \reg_y_reg[14][19]  ( .D(n1382), .CP(clk), .Q(\reg_y[14][19] ) );
  dff_sg \reg_y_reg[14][18]  ( .D(n1383), .CP(clk), .Q(\reg_y[14][18] ) );
  dff_sg \reg_y_reg[14][17]  ( .D(n1384), .CP(clk), .Q(\reg_y[14][17] ) );
  dff_sg \reg_y_reg[14][16]  ( .D(n1385), .CP(clk), .Q(\reg_y[14][16] ) );
  dff_sg \reg_y_reg[14][15]  ( .D(n1386), .CP(clk), .Q(\reg_y[14][15] ) );
  dff_sg \reg_y_reg[14][14]  ( .D(n1387), .CP(clk), .Q(\reg_y[14][14] ) );
  dff_sg \reg_y_reg[14][13]  ( .D(n1388), .CP(clk), .Q(\reg_y[14][13] ) );
  dff_sg \reg_y_reg[14][12]  ( .D(n1389), .CP(clk), .Q(\reg_y[14][12] ) );
  dff_sg \reg_y_reg[14][11]  ( .D(n1390), .CP(clk), .Q(\reg_y[14][11] ) );
  dff_sg \reg_y_reg[14][10]  ( .D(n1391), .CP(clk), .Q(\reg_y[14][10] ) );
  dff_sg \reg_y_reg[14][9]  ( .D(n1392), .CP(clk), .Q(\reg_y[14][9] ) );
  dff_sg \reg_y_reg[14][8]  ( .D(n1393), .CP(clk), .Q(\reg_y[14][8] ) );
  dff_sg \reg_y_reg[14][7]  ( .D(n1394), .CP(clk), .Q(\reg_y[14][7] ) );
  dff_sg \reg_y_reg[14][6]  ( .D(n1395), .CP(clk), .Q(\reg_y[14][6] ) );
  dff_sg \reg_y_reg[14][5]  ( .D(n1396), .CP(clk), .Q(\reg_y[14][5] ) );
  dff_sg \reg_y_reg[14][4]  ( .D(n1397), .CP(clk), .Q(\reg_y[14][4] ) );
  dff_sg \reg_y_reg[14][3]  ( .D(n1398), .CP(clk), .Q(\reg_y[14][3] ) );
  dff_sg \reg_y_reg[14][2]  ( .D(n1399), .CP(clk), .Q(\reg_y[14][2] ) );
  dff_sg \reg_y_reg[14][1]  ( .D(n1400), .CP(clk), .Q(\reg_y[14][1] ) );
  dff_sg \reg_y_reg[14][0]  ( .D(n1401), .CP(clk), .Q(\reg_y[14][0] ) );
  dff_sg \reg_y_reg[13][19]  ( .D(n1402), .CP(clk), .Q(\reg_y[13][19] ) );
  dff_sg \reg_y_reg[13][18]  ( .D(n1403), .CP(clk), .Q(\reg_y[13][18] ) );
  dff_sg \reg_y_reg[13][17]  ( .D(n1404), .CP(clk), .Q(\reg_y[13][17] ) );
  dff_sg \reg_y_reg[13][16]  ( .D(n1405), .CP(clk), .Q(\reg_y[13][16] ) );
  dff_sg \reg_y_reg[13][15]  ( .D(n1406), .CP(clk), .Q(\reg_y[13][15] ) );
  dff_sg \reg_y_reg[13][14]  ( .D(n1407), .CP(clk), .Q(\reg_y[13][14] ) );
  dff_sg \reg_y_reg[13][13]  ( .D(n1408), .CP(clk), .Q(\reg_y[13][13] ) );
  dff_sg \reg_y_reg[13][12]  ( .D(n1409), .CP(clk), .Q(\reg_y[13][12] ) );
  dff_sg \reg_y_reg[13][11]  ( .D(n1410), .CP(clk), .Q(\reg_y[13][11] ) );
  dff_sg \reg_y_reg[13][10]  ( .D(n1411), .CP(clk), .Q(\reg_y[13][10] ) );
  dff_sg \reg_y_reg[13][9]  ( .D(n1412), .CP(clk), .Q(\reg_y[13][9] ) );
  dff_sg \reg_y_reg[13][8]  ( .D(n1413), .CP(clk), .Q(\reg_y[13][8] ) );
  dff_sg \reg_y_reg[13][7]  ( .D(n1414), .CP(clk), .Q(\reg_y[13][7] ) );
  dff_sg \reg_y_reg[13][6]  ( .D(n1415), .CP(clk), .Q(\reg_y[13][6] ) );
  dff_sg \reg_y_reg[13][5]  ( .D(n1416), .CP(clk), .Q(\reg_y[13][5] ) );
  dff_sg \reg_y_reg[13][4]  ( .D(n1417), .CP(clk), .Q(\reg_y[13][4] ) );
  dff_sg \reg_y_reg[13][3]  ( .D(n1418), .CP(clk), .Q(\reg_y[13][3] ) );
  dff_sg \reg_y_reg[13][2]  ( .D(n1419), .CP(clk), .Q(\reg_y[13][2] ) );
  dff_sg \reg_y_reg[13][1]  ( .D(n1420), .CP(clk), .Q(\reg_y[13][1] ) );
  dff_sg \reg_y_reg[13][0]  ( .D(n1421), .CP(clk), .Q(\reg_y[13][0] ) );
  dff_sg \reg_y_reg[12][19]  ( .D(n1422), .CP(clk), .Q(\reg_y[12][19] ) );
  dff_sg \reg_y_reg[12][18]  ( .D(n1423), .CP(clk), .Q(\reg_y[12][18] ) );
  dff_sg \reg_y_reg[12][17]  ( .D(n1424), .CP(clk), .Q(\reg_y[12][17] ) );
  dff_sg \reg_y_reg[12][16]  ( .D(n1425), .CP(clk), .Q(\reg_y[12][16] ) );
  dff_sg \reg_y_reg[12][15]  ( .D(n1426), .CP(clk), .Q(\reg_y[12][15] ) );
  dff_sg \reg_y_reg[12][14]  ( .D(n1427), .CP(clk), .Q(\reg_y[12][14] ) );
  dff_sg \reg_y_reg[12][13]  ( .D(n1428), .CP(clk), .Q(\reg_y[12][13] ) );
  dff_sg \reg_y_reg[12][12]  ( .D(n1429), .CP(clk), .Q(\reg_y[12][12] ) );
  dff_sg \reg_y_reg[12][11]  ( .D(n1430), .CP(clk), .Q(\reg_y[12][11] ) );
  dff_sg \reg_y_reg[12][10]  ( .D(n1431), .CP(clk), .Q(\reg_y[12][10] ) );
  dff_sg \reg_y_reg[12][9]  ( .D(n1432), .CP(clk), .Q(\reg_y[12][9] ) );
  dff_sg \reg_y_reg[12][8]  ( .D(n1433), .CP(clk), .Q(\reg_y[12][8] ) );
  dff_sg \reg_y_reg[12][7]  ( .D(n1434), .CP(clk), .Q(\reg_y[12][7] ) );
  dff_sg \reg_y_reg[12][6]  ( .D(n1435), .CP(clk), .Q(\reg_y[12][6] ) );
  dff_sg \reg_y_reg[12][5]  ( .D(n1436), .CP(clk), .Q(\reg_y[12][5] ) );
  dff_sg \reg_y_reg[12][4]  ( .D(n1437), .CP(clk), .Q(\reg_y[12][4] ) );
  dff_sg \reg_y_reg[12][3]  ( .D(n1438), .CP(clk), .Q(\reg_y[12][3] ) );
  dff_sg \reg_y_reg[12][2]  ( .D(n1439), .CP(clk), .Q(\reg_y[12][2] ) );
  dff_sg \reg_y_reg[12][1]  ( .D(n1440), .CP(clk), .Q(\reg_y[12][1] ) );
  dff_sg \reg_y_reg[12][0]  ( .D(n1441), .CP(clk), .Q(\reg_y[12][0] ) );
  dff_sg \reg_y_reg[11][19]  ( .D(n1442), .CP(clk), .Q(\reg_y[11][19] ) );
  dff_sg \reg_y_reg[11][18]  ( .D(n1443), .CP(clk), .Q(\reg_y[11][18] ) );
  dff_sg \reg_y_reg[11][17]  ( .D(n1444), .CP(clk), .Q(\reg_y[11][17] ) );
  dff_sg \reg_y_reg[11][16]  ( .D(n1445), .CP(clk), .Q(\reg_y[11][16] ) );
  dff_sg \reg_y_reg[11][15]  ( .D(n1446), .CP(clk), .Q(\reg_y[11][15] ) );
  dff_sg \reg_y_reg[11][14]  ( .D(n1447), .CP(clk), .Q(\reg_y[11][14] ) );
  dff_sg \reg_y_reg[11][13]  ( .D(n1448), .CP(clk), .Q(\reg_y[11][13] ) );
  dff_sg \reg_y_reg[11][12]  ( .D(n1449), .CP(clk), .Q(\reg_y[11][12] ) );
  dff_sg \reg_y_reg[11][11]  ( .D(n1450), .CP(clk), .Q(\reg_y[11][11] ) );
  dff_sg \reg_y_reg[11][10]  ( .D(n1451), .CP(clk), .Q(\reg_y[11][10] ) );
  dff_sg \reg_y_reg[11][9]  ( .D(n1452), .CP(clk), .Q(\reg_y[11][9] ) );
  dff_sg \reg_y_reg[11][8]  ( .D(n1453), .CP(clk), .Q(\reg_y[11][8] ) );
  dff_sg \reg_y_reg[11][7]  ( .D(n1454), .CP(clk), .Q(\reg_y[11][7] ) );
  dff_sg \reg_y_reg[11][6]  ( .D(n1455), .CP(clk), .Q(\reg_y[11][6] ) );
  dff_sg \reg_y_reg[11][5]  ( .D(n1456), .CP(clk), .Q(\reg_y[11][5] ) );
  dff_sg \reg_y_reg[11][4]  ( .D(n1457), .CP(clk), .Q(\reg_y[11][4] ) );
  dff_sg \reg_y_reg[11][3]  ( .D(n1458), .CP(clk), .Q(\reg_y[11][3] ) );
  dff_sg \reg_y_reg[11][2]  ( .D(n1459), .CP(clk), .Q(\reg_y[11][2] ) );
  dff_sg \reg_y_reg[11][1]  ( .D(n1460), .CP(clk), .Q(\reg_y[11][1] ) );
  dff_sg \reg_y_reg[11][0]  ( .D(n1461), .CP(clk), .Q(\reg_y[11][0] ) );
  dff_sg \reg_y_reg[10][19]  ( .D(n1462), .CP(clk), .Q(\reg_y[10][19] ) );
  dff_sg \reg_y_reg[10][18]  ( .D(n1463), .CP(clk), .Q(\reg_y[10][18] ) );
  dff_sg \reg_y_reg[10][17]  ( .D(n1464), .CP(clk), .Q(\reg_y[10][17] ) );
  dff_sg \reg_y_reg[10][16]  ( .D(n1465), .CP(clk), .Q(\reg_y[10][16] ) );
  dff_sg \reg_y_reg[10][15]  ( .D(n1466), .CP(clk), .Q(\reg_y[10][15] ) );
  dff_sg \reg_y_reg[10][14]  ( .D(n1467), .CP(clk), .Q(\reg_y[10][14] ) );
  dff_sg \reg_y_reg[10][13]  ( .D(n1468), .CP(clk), .Q(\reg_y[10][13] ) );
  dff_sg \reg_y_reg[10][12]  ( .D(n1469), .CP(clk), .Q(\reg_y[10][12] ) );
  dff_sg \reg_y_reg[10][11]  ( .D(n1470), .CP(clk), .Q(\reg_y[10][11] ) );
  dff_sg \reg_y_reg[10][10]  ( .D(n1471), .CP(clk), .Q(\reg_y[10][10] ) );
  dff_sg \reg_y_reg[10][9]  ( .D(n1472), .CP(clk), .Q(\reg_y[10][9] ) );
  dff_sg \reg_y_reg[10][8]  ( .D(n1473), .CP(clk), .Q(\reg_y[10][8] ) );
  dff_sg \reg_y_reg[10][7]  ( .D(n1474), .CP(clk), .Q(\reg_y[10][7] ) );
  dff_sg \reg_y_reg[10][6]  ( .D(n1475), .CP(clk), .Q(\reg_y[10][6] ) );
  dff_sg \reg_y_reg[10][5]  ( .D(n1476), .CP(clk), .Q(\reg_y[10][5] ) );
  dff_sg \reg_y_reg[10][4]  ( .D(n1477), .CP(clk), .Q(\reg_y[10][4] ) );
  dff_sg \reg_y_reg[10][3]  ( .D(n1478), .CP(clk), .Q(\reg_y[10][3] ) );
  dff_sg \reg_y_reg[10][2]  ( .D(n1479), .CP(clk), .Q(\reg_y[10][2] ) );
  dff_sg \reg_y_reg[10][1]  ( .D(n1480), .CP(clk), .Q(\reg_y[10][1] ) );
  dff_sg \reg_y_reg[10][0]  ( .D(n1481), .CP(clk), .Q(\reg_y[10][0] ) );
  dff_sg \reg_y_reg[9][19]  ( .D(n1482), .CP(clk), .Q(\reg_y[9][19] ) );
  dff_sg \reg_y_reg[9][18]  ( .D(n1483), .CP(clk), .Q(\reg_y[9][18] ) );
  dff_sg \reg_y_reg[9][17]  ( .D(n1484), .CP(clk), .Q(\reg_y[9][17] ) );
  dff_sg \reg_y_reg[9][16]  ( .D(n1485), .CP(clk), .Q(\reg_y[9][16] ) );
  dff_sg \reg_y_reg[9][15]  ( .D(n1486), .CP(clk), .Q(\reg_y[9][15] ) );
  dff_sg \reg_y_reg[9][14]  ( .D(n1487), .CP(clk), .Q(\reg_y[9][14] ) );
  dff_sg \reg_y_reg[9][13]  ( .D(n1488), .CP(clk), .Q(\reg_y[9][13] ) );
  dff_sg \reg_y_reg[9][12]  ( .D(n1489), .CP(clk), .Q(\reg_y[9][12] ) );
  dff_sg \reg_y_reg[9][11]  ( .D(n1490), .CP(clk), .Q(\reg_y[9][11] ) );
  dff_sg \reg_y_reg[9][10]  ( .D(n1491), .CP(clk), .Q(\reg_y[9][10] ) );
  dff_sg \reg_y_reg[9][9]  ( .D(n1492), .CP(clk), .Q(\reg_y[9][9] ) );
  dff_sg \reg_y_reg[9][8]  ( .D(n1493), .CP(clk), .Q(\reg_y[9][8] ) );
  dff_sg \reg_y_reg[9][7]  ( .D(n1494), .CP(clk), .Q(\reg_y[9][7] ) );
  dff_sg \reg_y_reg[9][6]  ( .D(n1495), .CP(clk), .Q(\reg_y[9][6] ) );
  dff_sg \reg_y_reg[9][5]  ( .D(n1496), .CP(clk), .Q(\reg_y[9][5] ) );
  dff_sg \reg_y_reg[9][4]  ( .D(n1497), .CP(clk), .Q(\reg_y[9][4] ) );
  dff_sg \reg_y_reg[9][3]  ( .D(n1498), .CP(clk), .Q(\reg_y[9][3] ) );
  dff_sg \reg_y_reg[9][2]  ( .D(n1499), .CP(clk), .Q(\reg_y[9][2] ) );
  dff_sg \reg_y_reg[9][1]  ( .D(n1500), .CP(clk), .Q(\reg_y[9][1] ) );
  dff_sg \reg_y_reg[9][0]  ( .D(n1501), .CP(clk), .Q(\reg_y[9][0] ) );
  dff_sg \reg_y_reg[8][19]  ( .D(n1502), .CP(clk), .Q(\reg_y[8][19] ) );
  dff_sg \reg_y_reg[8][18]  ( .D(n1503), .CP(clk), .Q(\reg_y[8][18] ) );
  dff_sg \reg_y_reg[8][17]  ( .D(n1504), .CP(clk), .Q(\reg_y[8][17] ) );
  dff_sg \reg_y_reg[8][16]  ( .D(n1505), .CP(clk), .Q(\reg_y[8][16] ) );
  dff_sg \reg_y_reg[8][15]  ( .D(n1506), .CP(clk), .Q(\reg_y[8][15] ) );
  dff_sg \reg_y_reg[8][14]  ( .D(n1507), .CP(clk), .Q(\reg_y[8][14] ) );
  dff_sg \reg_y_reg[8][13]  ( .D(n1508), .CP(clk), .Q(\reg_y[8][13] ) );
  dff_sg \reg_y_reg[8][12]  ( .D(n1509), .CP(clk), .Q(\reg_y[8][12] ) );
  dff_sg \reg_y_reg[8][11]  ( .D(n1510), .CP(clk), .Q(\reg_y[8][11] ) );
  dff_sg \reg_y_reg[8][10]  ( .D(n1511), .CP(clk), .Q(\reg_y[8][10] ) );
  dff_sg \reg_y_reg[8][9]  ( .D(n1512), .CP(clk), .Q(\reg_y[8][9] ) );
  dff_sg \reg_y_reg[8][8]  ( .D(n1513), .CP(clk), .Q(\reg_y[8][8] ) );
  dff_sg \reg_y_reg[8][7]  ( .D(n1514), .CP(clk), .Q(\reg_y[8][7] ) );
  dff_sg \reg_y_reg[8][6]  ( .D(n1515), .CP(clk), .Q(\reg_y[8][6] ) );
  dff_sg \reg_y_reg[8][5]  ( .D(n1516), .CP(clk), .Q(\reg_y[8][5] ) );
  dff_sg \reg_y_reg[8][4]  ( .D(n1517), .CP(clk), .Q(\reg_y[8][4] ) );
  dff_sg \reg_y_reg[8][3]  ( .D(n1518), .CP(clk), .Q(\reg_y[8][3] ) );
  dff_sg \reg_y_reg[8][2]  ( .D(n1519), .CP(clk), .Q(\reg_y[8][2] ) );
  dff_sg \reg_y_reg[8][1]  ( .D(n1520), .CP(clk), .Q(\reg_y[8][1] ) );
  dff_sg \reg_y_reg[8][0]  ( .D(n1521), .CP(clk), .Q(\reg_y[8][0] ) );
  dff_sg \reg_y_reg[7][19]  ( .D(n1522), .CP(clk), .Q(\reg_y[7][19] ) );
  dff_sg \reg_y_reg[7][18]  ( .D(n1523), .CP(clk), .Q(\reg_y[7][18] ) );
  dff_sg \reg_y_reg[7][17]  ( .D(n1524), .CP(clk), .Q(\reg_y[7][17] ) );
  dff_sg \reg_y_reg[7][16]  ( .D(n1525), .CP(clk), .Q(\reg_y[7][16] ) );
  dff_sg \reg_y_reg[7][15]  ( .D(n1526), .CP(clk), .Q(\reg_y[7][15] ) );
  dff_sg \reg_y_reg[7][14]  ( .D(n1527), .CP(clk), .Q(\reg_y[7][14] ) );
  dff_sg \reg_y_reg[7][13]  ( .D(n1528), .CP(clk), .Q(\reg_y[7][13] ) );
  dff_sg \reg_y_reg[7][12]  ( .D(n1529), .CP(clk), .Q(\reg_y[7][12] ) );
  dff_sg \reg_y_reg[7][11]  ( .D(n1530), .CP(clk), .Q(\reg_y[7][11] ) );
  dff_sg \reg_y_reg[7][10]  ( .D(n1531), .CP(clk), .Q(\reg_y[7][10] ) );
  dff_sg \reg_y_reg[7][9]  ( .D(n1532), .CP(clk), .Q(\reg_y[7][9] ) );
  dff_sg \reg_y_reg[7][8]  ( .D(n1533), .CP(clk), .Q(\reg_y[7][8] ) );
  dff_sg \reg_y_reg[7][7]  ( .D(n1534), .CP(clk), .Q(\reg_y[7][7] ) );
  dff_sg \reg_y_reg[7][6]  ( .D(n1535), .CP(clk), .Q(\reg_y[7][6] ) );
  dff_sg \reg_y_reg[7][5]  ( .D(n1536), .CP(clk), .Q(\reg_y[7][5] ) );
  dff_sg \reg_y_reg[7][4]  ( .D(n1537), .CP(clk), .Q(\reg_y[7][4] ) );
  dff_sg \reg_y_reg[7][3]  ( .D(n1538), .CP(clk), .Q(\reg_y[7][3] ) );
  dff_sg \reg_y_reg[7][2]  ( .D(n1539), .CP(clk), .Q(\reg_y[7][2] ) );
  dff_sg \reg_y_reg[7][1]  ( .D(n1540), .CP(clk), .Q(\reg_y[7][1] ) );
  dff_sg \reg_y_reg[7][0]  ( .D(n1541), .CP(clk), .Q(\reg_y[7][0] ) );
  dff_sg \reg_y_reg[6][19]  ( .D(n1542), .CP(clk), .Q(\reg_y[6][19] ) );
  dff_sg \reg_y_reg[6][18]  ( .D(n1543), .CP(clk), .Q(\reg_y[6][18] ) );
  dff_sg \reg_y_reg[6][17]  ( .D(n1544), .CP(clk), .Q(\reg_y[6][17] ) );
  dff_sg \reg_y_reg[6][16]  ( .D(n1545), .CP(clk), .Q(\reg_y[6][16] ) );
  dff_sg \reg_y_reg[6][15]  ( .D(n1546), .CP(clk), .Q(\reg_y[6][15] ) );
  dff_sg \reg_y_reg[6][14]  ( .D(n1547), .CP(clk), .Q(\reg_y[6][14] ) );
  dff_sg \reg_y_reg[6][13]  ( .D(n1548), .CP(clk), .Q(\reg_y[6][13] ) );
  dff_sg \reg_y_reg[6][12]  ( .D(n1549), .CP(clk), .Q(\reg_y[6][12] ) );
  dff_sg \reg_y_reg[6][11]  ( .D(n1550), .CP(clk), .Q(\reg_y[6][11] ) );
  dff_sg \reg_y_reg[6][10]  ( .D(n1551), .CP(clk), .Q(\reg_y[6][10] ) );
  dff_sg \reg_y_reg[6][9]  ( .D(n1552), .CP(clk), .Q(\reg_y[6][9] ) );
  dff_sg \reg_y_reg[6][8]  ( .D(n1553), .CP(clk), .Q(\reg_y[6][8] ) );
  dff_sg \reg_y_reg[6][7]  ( .D(n1554), .CP(clk), .Q(\reg_y[6][7] ) );
  dff_sg \reg_y_reg[6][6]  ( .D(n1555), .CP(clk), .Q(\reg_y[6][6] ) );
  dff_sg \reg_y_reg[6][5]  ( .D(n1556), .CP(clk), .Q(\reg_y[6][5] ) );
  dff_sg \reg_y_reg[6][4]  ( .D(n1557), .CP(clk), .Q(\reg_y[6][4] ) );
  dff_sg \reg_y_reg[6][3]  ( .D(n1558), .CP(clk), .Q(\reg_y[6][3] ) );
  dff_sg \reg_y_reg[6][2]  ( .D(n1559), .CP(clk), .Q(\reg_y[6][2] ) );
  dff_sg \reg_y_reg[6][1]  ( .D(n1560), .CP(clk), .Q(\reg_y[6][1] ) );
  dff_sg \reg_y_reg[6][0]  ( .D(n1561), .CP(clk), .Q(\reg_y[6][0] ) );
  dff_sg \reg_y_reg[5][19]  ( .D(n1562), .CP(clk), .Q(\reg_y[5][19] ) );
  dff_sg \reg_y_reg[5][18]  ( .D(n1563), .CP(clk), .Q(\reg_y[5][18] ) );
  dff_sg \reg_y_reg[5][17]  ( .D(n1564), .CP(clk), .Q(\reg_y[5][17] ) );
  dff_sg \reg_y_reg[5][16]  ( .D(n1565), .CP(clk), .Q(\reg_y[5][16] ) );
  dff_sg \reg_y_reg[5][15]  ( .D(n1566), .CP(clk), .Q(\reg_y[5][15] ) );
  dff_sg \reg_y_reg[5][14]  ( .D(n1567), .CP(clk), .Q(\reg_y[5][14] ) );
  dff_sg \reg_y_reg[5][13]  ( .D(n1568), .CP(clk), .Q(\reg_y[5][13] ) );
  dff_sg \reg_y_reg[5][12]  ( .D(n1569), .CP(clk), .Q(\reg_y[5][12] ) );
  dff_sg \reg_y_reg[5][11]  ( .D(n1570), .CP(clk), .Q(\reg_y[5][11] ) );
  dff_sg \reg_y_reg[5][10]  ( .D(n1571), .CP(clk), .Q(\reg_y[5][10] ) );
  dff_sg \reg_y_reg[5][9]  ( .D(n1572), .CP(clk), .Q(\reg_y[5][9] ) );
  dff_sg \reg_y_reg[5][8]  ( .D(n1573), .CP(clk), .Q(\reg_y[5][8] ) );
  dff_sg \reg_y_reg[5][7]  ( .D(n1574), .CP(clk), .Q(\reg_y[5][7] ) );
  dff_sg \reg_y_reg[5][6]  ( .D(n1575), .CP(clk), .Q(\reg_y[5][6] ) );
  dff_sg \reg_y_reg[5][5]  ( .D(n1576), .CP(clk), .Q(\reg_y[5][5] ) );
  dff_sg \reg_y_reg[5][4]  ( .D(n1577), .CP(clk), .Q(\reg_y[5][4] ) );
  dff_sg \reg_y_reg[5][3]  ( .D(n1578), .CP(clk), .Q(\reg_y[5][3] ) );
  dff_sg \reg_y_reg[5][2]  ( .D(n1579), .CP(clk), .Q(\reg_y[5][2] ) );
  dff_sg \reg_y_reg[5][1]  ( .D(n1580), .CP(clk), .Q(\reg_y[5][1] ) );
  dff_sg \reg_y_reg[5][0]  ( .D(n1581), .CP(clk), .Q(\reg_y[5][0] ) );
  dff_sg \reg_y_reg[4][19]  ( .D(n1582), .CP(clk), .Q(\reg_y[4][19] ) );
  dff_sg \reg_y_reg[4][18]  ( .D(n1583), .CP(clk), .Q(\reg_y[4][18] ) );
  dff_sg \reg_y_reg[4][17]  ( .D(n1584), .CP(clk), .Q(\reg_y[4][17] ) );
  dff_sg \reg_y_reg[4][16]  ( .D(n1585), .CP(clk), .Q(\reg_y[4][16] ) );
  dff_sg \reg_y_reg[4][15]  ( .D(n1586), .CP(clk), .Q(\reg_y[4][15] ) );
  dff_sg \reg_y_reg[4][14]  ( .D(n1587), .CP(clk), .Q(\reg_y[4][14] ) );
  dff_sg \reg_y_reg[4][13]  ( .D(n1588), .CP(clk), .Q(\reg_y[4][13] ) );
  dff_sg \reg_y_reg[4][12]  ( .D(n1589), .CP(clk), .Q(\reg_y[4][12] ) );
  dff_sg \reg_y_reg[4][11]  ( .D(n1590), .CP(clk), .Q(\reg_y[4][11] ) );
  dff_sg \reg_y_reg[4][10]  ( .D(n1591), .CP(clk), .Q(\reg_y[4][10] ) );
  dff_sg \reg_y_reg[4][9]  ( .D(n1592), .CP(clk), .Q(\reg_y[4][9] ) );
  dff_sg \reg_y_reg[4][8]  ( .D(n1593), .CP(clk), .Q(\reg_y[4][8] ) );
  dff_sg \reg_y_reg[4][7]  ( .D(n1594), .CP(clk), .Q(\reg_y[4][7] ) );
  dff_sg \reg_y_reg[4][6]  ( .D(n1595), .CP(clk), .Q(\reg_y[4][6] ) );
  dff_sg \reg_y_reg[4][5]  ( .D(n1596), .CP(clk), .Q(\reg_y[4][5] ) );
  dff_sg \reg_y_reg[4][4]  ( .D(n1597), .CP(clk), .Q(\reg_y[4][4] ) );
  dff_sg \reg_y_reg[4][3]  ( .D(n1598), .CP(clk), .Q(\reg_y[4][3] ) );
  dff_sg \reg_y_reg[4][2]  ( .D(n1599), .CP(clk), .Q(\reg_y[4][2] ) );
  dff_sg \reg_y_reg[4][1]  ( .D(n1600), .CP(clk), .Q(\reg_y[4][1] ) );
  dff_sg \reg_y_reg[4][0]  ( .D(n1601), .CP(clk), .Q(\reg_y[4][0] ) );
  dff_sg \reg_y_reg[3][19]  ( .D(n1602), .CP(clk), .Q(\reg_y[3][19] ) );
  dff_sg \reg_y_reg[3][18]  ( .D(n1603), .CP(clk), .Q(\reg_y[3][18] ) );
  dff_sg \reg_y_reg[3][17]  ( .D(n1604), .CP(clk), .Q(\reg_y[3][17] ) );
  dff_sg \reg_y_reg[3][16]  ( .D(n1605), .CP(clk), .Q(\reg_y[3][16] ) );
  dff_sg \reg_y_reg[3][15]  ( .D(n1606), .CP(clk), .Q(\reg_y[3][15] ) );
  dff_sg \reg_y_reg[3][14]  ( .D(n1607), .CP(clk), .Q(\reg_y[3][14] ) );
  dff_sg \reg_y_reg[3][13]  ( .D(n1608), .CP(clk), .Q(\reg_y[3][13] ) );
  dff_sg \reg_y_reg[3][12]  ( .D(n1609), .CP(clk), .Q(\reg_y[3][12] ) );
  dff_sg \reg_y_reg[3][11]  ( .D(n1610), .CP(clk), .Q(\reg_y[3][11] ) );
  dff_sg \reg_y_reg[3][10]  ( .D(n1611), .CP(clk), .Q(\reg_y[3][10] ) );
  dff_sg \reg_y_reg[3][9]  ( .D(n1612), .CP(clk), .Q(\reg_y[3][9] ) );
  dff_sg \reg_y_reg[3][8]  ( .D(n1613), .CP(clk), .Q(\reg_y[3][8] ) );
  dff_sg \reg_y_reg[3][7]  ( .D(n1614), .CP(clk), .Q(\reg_y[3][7] ) );
  dff_sg \reg_y_reg[3][6]  ( .D(n1615), .CP(clk), .Q(\reg_y[3][6] ) );
  dff_sg \reg_y_reg[3][5]  ( .D(n1616), .CP(clk), .Q(\reg_y[3][5] ) );
  dff_sg \reg_y_reg[3][4]  ( .D(n1617), .CP(clk), .Q(\reg_y[3][4] ) );
  dff_sg \reg_y_reg[3][3]  ( .D(n1618), .CP(clk), .Q(\reg_y[3][3] ) );
  dff_sg \reg_y_reg[3][2]  ( .D(n1619), .CP(clk), .Q(\reg_y[3][2] ) );
  dff_sg \reg_y_reg[3][1]  ( .D(n1620), .CP(clk), .Q(\reg_y[3][1] ) );
  dff_sg \reg_y_reg[3][0]  ( .D(n1621), .CP(clk), .Q(\reg_y[3][0] ) );
  dff_sg \reg_y_reg[2][19]  ( .D(n1622), .CP(clk), .Q(\reg_y[2][19] ) );
  dff_sg \reg_y_reg[2][18]  ( .D(n1623), .CP(clk), .Q(\reg_y[2][18] ) );
  dff_sg \reg_y_reg[2][17]  ( .D(n1624), .CP(clk), .Q(\reg_y[2][17] ) );
  dff_sg \reg_y_reg[2][16]  ( .D(n1625), .CP(clk), .Q(\reg_y[2][16] ) );
  dff_sg \reg_y_reg[2][15]  ( .D(n1626), .CP(clk), .Q(\reg_y[2][15] ) );
  dff_sg \reg_y_reg[2][14]  ( .D(n1627), .CP(clk), .Q(\reg_y[2][14] ) );
  dff_sg \reg_y_reg[2][13]  ( .D(n1628), .CP(clk), .Q(\reg_y[2][13] ) );
  dff_sg \reg_y_reg[2][12]  ( .D(n1629), .CP(clk), .Q(\reg_y[2][12] ) );
  dff_sg \reg_y_reg[2][11]  ( .D(n1630), .CP(clk), .Q(\reg_y[2][11] ) );
  dff_sg \reg_y_reg[2][10]  ( .D(n1631), .CP(clk), .Q(\reg_y[2][10] ) );
  dff_sg \reg_y_reg[2][9]  ( .D(n1632), .CP(clk), .Q(\reg_y[2][9] ) );
  dff_sg \reg_y_reg[2][8]  ( .D(n1633), .CP(clk), .Q(\reg_y[2][8] ) );
  dff_sg \reg_y_reg[2][7]  ( .D(n1634), .CP(clk), .Q(\reg_y[2][7] ) );
  dff_sg \reg_y_reg[2][6]  ( .D(n1635), .CP(clk), .Q(\reg_y[2][6] ) );
  dff_sg \reg_y_reg[2][5]  ( .D(n1636), .CP(clk), .Q(\reg_y[2][5] ) );
  dff_sg \reg_y_reg[2][4]  ( .D(n1637), .CP(clk), .Q(\reg_y[2][4] ) );
  dff_sg \reg_y_reg[2][3]  ( .D(n1638), .CP(clk), .Q(\reg_y[2][3] ) );
  dff_sg \reg_y_reg[2][2]  ( .D(n1639), .CP(clk), .Q(\reg_y[2][2] ) );
  dff_sg \reg_y_reg[2][1]  ( .D(n1640), .CP(clk), .Q(\reg_y[2][1] ) );
  dff_sg \reg_y_reg[2][0]  ( .D(n1641), .CP(clk), .Q(\reg_y[2][0] ) );
  dff_sg \reg_y_reg[1][19]  ( .D(n1642), .CP(clk), .Q(\reg_y[1][19] ) );
  dff_sg \reg_y_reg[1][18]  ( .D(n1643), .CP(clk), .Q(\reg_y[1][18] ) );
  dff_sg \reg_y_reg[1][17]  ( .D(n1644), .CP(clk), .Q(\reg_y[1][17] ) );
  dff_sg \reg_y_reg[1][16]  ( .D(n1645), .CP(clk), .Q(\reg_y[1][16] ) );
  dff_sg \reg_y_reg[1][15]  ( .D(n1646), .CP(clk), .Q(\reg_y[1][15] ) );
  dff_sg \reg_y_reg[1][14]  ( .D(n1647), .CP(clk), .Q(\reg_y[1][14] ) );
  dff_sg \reg_y_reg[1][13]  ( .D(n1648), .CP(clk), .Q(\reg_y[1][13] ) );
  dff_sg \reg_y_reg[1][12]  ( .D(n1649), .CP(clk), .Q(\reg_y[1][12] ) );
  dff_sg \reg_y_reg[1][11]  ( .D(n1650), .CP(clk), .Q(\reg_y[1][11] ) );
  dff_sg \reg_y_reg[1][10]  ( .D(n1651), .CP(clk), .Q(\reg_y[1][10] ) );
  dff_sg \reg_y_reg[1][9]  ( .D(n1652), .CP(clk), .Q(\reg_y[1][9] ) );
  dff_sg \reg_y_reg[1][8]  ( .D(n1653), .CP(clk), .Q(\reg_y[1][8] ) );
  dff_sg \reg_y_reg[1][7]  ( .D(n1654), .CP(clk), .Q(\reg_y[1][7] ) );
  dff_sg \reg_y_reg[1][6]  ( .D(n1655), .CP(clk), .Q(\reg_y[1][6] ) );
  dff_sg \reg_y_reg[1][5]  ( .D(n1656), .CP(clk), .Q(\reg_y[1][5] ) );
  dff_sg \reg_y_reg[1][4]  ( .D(n1657), .CP(clk), .Q(\reg_y[1][4] ) );
  dff_sg \reg_y_reg[1][3]  ( .D(n1658), .CP(clk), .Q(\reg_y[1][3] ) );
  dff_sg \reg_y_reg[1][2]  ( .D(n1659), .CP(clk), .Q(\reg_y[1][2] ) );
  dff_sg \reg_y_reg[1][1]  ( .D(n1660), .CP(clk), .Q(\reg_y[1][1] ) );
  dff_sg \reg_y_reg[1][0]  ( .D(n1661), .CP(clk), .Q(\reg_y[1][0] ) );
  dff_sg \reg_y_reg[0][19]  ( .D(n1662), .CP(clk), .Q(\reg_y[0][19] ) );
  dff_sg \reg_y_reg[0][18]  ( .D(n1663), .CP(clk), .Q(\reg_y[0][18] ) );
  dff_sg \reg_y_reg[0][17]  ( .D(n1664), .CP(clk), .Q(\reg_y[0][17] ) );
  dff_sg \reg_y_reg[0][16]  ( .D(n1665), .CP(clk), .Q(\reg_y[0][16] ) );
  dff_sg \reg_y_reg[0][15]  ( .D(n1666), .CP(clk), .Q(\reg_y[0][15] ) );
  dff_sg \reg_y_reg[0][14]  ( .D(n1667), .CP(clk), .Q(\reg_y[0][14] ) );
  dff_sg \reg_y_reg[0][13]  ( .D(n1668), .CP(clk), .Q(\reg_y[0][13] ) );
  dff_sg \reg_y_reg[0][12]  ( .D(n1669), .CP(clk), .Q(\reg_y[0][12] ) );
  dff_sg \reg_y_reg[0][11]  ( .D(n1670), .CP(clk), .Q(\reg_y[0][11] ) );
  dff_sg \reg_y_reg[0][10]  ( .D(n1671), .CP(clk), .Q(\reg_y[0][10] ) );
  dff_sg \reg_y_reg[0][9]  ( .D(n1672), .CP(clk), .Q(\reg_y[0][9] ) );
  dff_sg \reg_y_reg[0][8]  ( .D(n1673), .CP(clk), .Q(\reg_y[0][8] ) );
  dff_sg \reg_y_reg[0][7]  ( .D(n1674), .CP(clk), .Q(\reg_y[0][7] ) );
  dff_sg \reg_y_reg[0][6]  ( .D(n1675), .CP(clk), .Q(\reg_y[0][6] ) );
  dff_sg \reg_y_reg[0][5]  ( .D(n1676), .CP(clk), .Q(\reg_y[0][5] ) );
  dff_sg \reg_y_reg[0][4]  ( .D(n1677), .CP(clk), .Q(\reg_y[0][4] ) );
  dff_sg \reg_y_reg[0][3]  ( .D(n1678), .CP(clk), .Q(\reg_y[0][3] ) );
  dff_sg \reg_y_reg[0][2]  ( .D(n1679), .CP(clk), .Q(\reg_y[0][2] ) );
  dff_sg \reg_y_reg[0][1]  ( .D(n1680), .CP(clk), .Q(\reg_y[0][1] ) );
  dff_sg \reg_y_reg[0][0]  ( .D(n1681), .CP(clk), .Q(\reg_y[0][0] ) );
  dff_sg \reg_yHat_reg[14][19]  ( .D(n1702), .CP(clk), .Q(\reg_yHat[14][19] )
         );
  dff_sg \reg_yHat_reg[14][18]  ( .D(n1703), .CP(clk), .Q(\reg_yHat[14][18] )
         );
  dff_sg \reg_yHat_reg[14][17]  ( .D(n1704), .CP(clk), .Q(\reg_yHat[14][17] )
         );
  dff_sg \reg_yHat_reg[14][16]  ( .D(n1705), .CP(clk), .Q(\reg_yHat[14][16] )
         );
  dff_sg \reg_yHat_reg[14][15]  ( .D(n1706), .CP(clk), .Q(\reg_yHat[14][15] )
         );
  dff_sg \reg_yHat_reg[14][14]  ( .D(n1707), .CP(clk), .Q(\reg_yHat[14][14] )
         );
  dff_sg \reg_yHat_reg[14][13]  ( .D(n1708), .CP(clk), .Q(\reg_yHat[14][13] )
         );
  dff_sg \reg_yHat_reg[14][12]  ( .D(n1709), .CP(clk), .Q(\reg_yHat[14][12] )
         );
  dff_sg \reg_yHat_reg[14][11]  ( .D(n1710), .CP(clk), .Q(\reg_yHat[14][11] )
         );
  dff_sg \reg_yHat_reg[14][10]  ( .D(n1711), .CP(clk), .Q(\reg_yHat[14][10] )
         );
  dff_sg \reg_yHat_reg[14][9]  ( .D(n1712), .CP(clk), .Q(\reg_yHat[14][9] ) );
  dff_sg \reg_yHat_reg[14][8]  ( .D(n1713), .CP(clk), .Q(\reg_yHat[14][8] ) );
  dff_sg \reg_yHat_reg[14][7]  ( .D(n1714), .CP(clk), .Q(\reg_yHat[14][7] ) );
  dff_sg \reg_yHat_reg[14][6]  ( .D(n1715), .CP(clk), .Q(\reg_yHat[14][6] ) );
  dff_sg \reg_yHat_reg[14][5]  ( .D(n1716), .CP(clk), .Q(\reg_yHat[14][5] ) );
  dff_sg \reg_yHat_reg[14][4]  ( .D(n1717), .CP(clk), .Q(\reg_yHat[14][4] ) );
  dff_sg \reg_yHat_reg[14][3]  ( .D(n1718), .CP(clk), .Q(\reg_yHat[14][3] ) );
  dff_sg \reg_yHat_reg[14][2]  ( .D(n1719), .CP(clk), .Q(\reg_yHat[14][2] ) );
  dff_sg \reg_yHat_reg[14][1]  ( .D(n1720), .CP(clk), .Q(\reg_yHat[14][1] ) );
  dff_sg \reg_yHat_reg[14][0]  ( .D(n1721), .CP(clk), .Q(\reg_yHat[14][0] ) );
  dff_sg \reg_yHat_reg[13][19]  ( .D(n1722), .CP(clk), .Q(\reg_yHat[13][19] )
         );
  dff_sg \reg_yHat_reg[13][18]  ( .D(n1723), .CP(clk), .Q(\reg_yHat[13][18] )
         );
  dff_sg \reg_yHat_reg[13][17]  ( .D(n1724), .CP(clk), .Q(\reg_yHat[13][17] )
         );
  dff_sg \reg_yHat_reg[13][16]  ( .D(n1725), .CP(clk), .Q(\reg_yHat[13][16] )
         );
  dff_sg \reg_yHat_reg[13][15]  ( .D(n1726), .CP(clk), .Q(\reg_yHat[13][15] )
         );
  dff_sg \reg_yHat_reg[13][14]  ( .D(n1727), .CP(clk), .Q(\reg_yHat[13][14] )
         );
  dff_sg \reg_yHat_reg[13][13]  ( .D(n1728), .CP(clk), .Q(\reg_yHat[13][13] )
         );
  dff_sg \reg_yHat_reg[13][12]  ( .D(n1729), .CP(clk), .Q(\reg_yHat[13][12] )
         );
  dff_sg \reg_yHat_reg[13][11]  ( .D(n1730), .CP(clk), .Q(\reg_yHat[13][11] )
         );
  dff_sg \reg_yHat_reg[13][10]  ( .D(n1731), .CP(clk), .Q(\reg_yHat[13][10] )
         );
  dff_sg \reg_yHat_reg[13][9]  ( .D(n1732), .CP(clk), .Q(\reg_yHat[13][9] ) );
  dff_sg \reg_yHat_reg[13][8]  ( .D(n1733), .CP(clk), .Q(\reg_yHat[13][8] ) );
  dff_sg \reg_yHat_reg[13][7]  ( .D(n1734), .CP(clk), .Q(\reg_yHat[13][7] ) );
  dff_sg \reg_yHat_reg[13][6]  ( .D(n1735), .CP(clk), .Q(\reg_yHat[13][6] ) );
  dff_sg \reg_yHat_reg[13][5]  ( .D(n1736), .CP(clk), .Q(\reg_yHat[13][5] ) );
  dff_sg \reg_yHat_reg[13][4]  ( .D(n1737), .CP(clk), .Q(\reg_yHat[13][4] ) );
  dff_sg \reg_yHat_reg[13][3]  ( .D(n1738), .CP(clk), .Q(\reg_yHat[13][3] ) );
  dff_sg \reg_yHat_reg[13][2]  ( .D(n1739), .CP(clk), .Q(\reg_yHat[13][2] ) );
  dff_sg \reg_yHat_reg[13][1]  ( .D(n1740), .CP(clk), .Q(\reg_yHat[13][1] ) );
  dff_sg \reg_yHat_reg[13][0]  ( .D(n1741), .CP(clk), .Q(\reg_yHat[13][0] ) );
  dff_sg \reg_yHat_reg[12][19]  ( .D(n1742), .CP(clk), .Q(\reg_yHat[12][19] )
         );
  dff_sg \reg_yHat_reg[12][18]  ( .D(n1743), .CP(clk), .Q(\reg_yHat[12][18] )
         );
  dff_sg \reg_yHat_reg[12][17]  ( .D(n1744), .CP(clk), .Q(\reg_yHat[12][17] )
         );
  dff_sg \reg_yHat_reg[12][16]  ( .D(n1745), .CP(clk), .Q(\reg_yHat[12][16] )
         );
  dff_sg \reg_yHat_reg[12][15]  ( .D(n1746), .CP(clk), .Q(\reg_yHat[12][15] )
         );
  dff_sg \reg_yHat_reg[12][14]  ( .D(n1747), .CP(clk), .Q(\reg_yHat[12][14] )
         );
  dff_sg \reg_yHat_reg[12][13]  ( .D(n1748), .CP(clk), .Q(\reg_yHat[12][13] )
         );
  dff_sg \reg_yHat_reg[12][12]  ( .D(n1749), .CP(clk), .Q(\reg_yHat[12][12] )
         );
  dff_sg \reg_yHat_reg[12][11]  ( .D(n1750), .CP(clk), .Q(\reg_yHat[12][11] )
         );
  dff_sg \reg_yHat_reg[12][10]  ( .D(n1751), .CP(clk), .Q(\reg_yHat[12][10] )
         );
  dff_sg \reg_yHat_reg[12][9]  ( .D(n1752), .CP(clk), .Q(\reg_yHat[12][9] ) );
  dff_sg \reg_yHat_reg[12][8]  ( .D(n1753), .CP(clk), .Q(\reg_yHat[12][8] ) );
  dff_sg \reg_yHat_reg[12][7]  ( .D(n1754), .CP(clk), .Q(\reg_yHat[12][7] ) );
  dff_sg \reg_yHat_reg[12][6]  ( .D(n1755), .CP(clk), .Q(\reg_yHat[12][6] ) );
  dff_sg \reg_yHat_reg[12][5]  ( .D(n1756), .CP(clk), .Q(\reg_yHat[12][5] ) );
  dff_sg \reg_yHat_reg[12][4]  ( .D(n1757), .CP(clk), .Q(\reg_yHat[12][4] ) );
  dff_sg \reg_yHat_reg[12][3]  ( .D(n1758), .CP(clk), .Q(\reg_yHat[12][3] ) );
  dff_sg \reg_yHat_reg[12][2]  ( .D(n1759), .CP(clk), .Q(\reg_yHat[12][2] ) );
  dff_sg \reg_yHat_reg[12][1]  ( .D(n1760), .CP(clk), .Q(\reg_yHat[12][1] ) );
  dff_sg \reg_yHat_reg[12][0]  ( .D(n1761), .CP(clk), .Q(\reg_yHat[12][0] ) );
  dff_sg \reg_yHat_reg[11][19]  ( .D(n1762), .CP(clk), .Q(\reg_yHat[11][19] )
         );
  dff_sg \reg_yHat_reg[11][18]  ( .D(n1763), .CP(clk), .Q(\reg_yHat[11][18] )
         );
  dff_sg \reg_yHat_reg[11][17]  ( .D(n1764), .CP(clk), .Q(\reg_yHat[11][17] )
         );
  dff_sg \reg_yHat_reg[11][16]  ( .D(n1765), .CP(clk), .Q(\reg_yHat[11][16] )
         );
  dff_sg \reg_yHat_reg[11][15]  ( .D(n1766), .CP(clk), .Q(\reg_yHat[11][15] )
         );
  dff_sg \reg_yHat_reg[11][14]  ( .D(n1767), .CP(clk), .Q(\reg_yHat[11][14] )
         );
  dff_sg \reg_yHat_reg[11][13]  ( .D(n1768), .CP(clk), .Q(\reg_yHat[11][13] )
         );
  dff_sg \reg_yHat_reg[11][12]  ( .D(n1769), .CP(clk), .Q(\reg_yHat[11][12] )
         );
  dff_sg \reg_yHat_reg[11][11]  ( .D(n1770), .CP(clk), .Q(\reg_yHat[11][11] )
         );
  dff_sg \reg_yHat_reg[11][10]  ( .D(n1771), .CP(clk), .Q(\reg_yHat[11][10] )
         );
  dff_sg \reg_yHat_reg[11][9]  ( .D(n1772), .CP(clk), .Q(\reg_yHat[11][9] ) );
  dff_sg \reg_yHat_reg[11][8]  ( .D(n1773), .CP(clk), .Q(\reg_yHat[11][8] ) );
  dff_sg \reg_yHat_reg[11][7]  ( .D(n1774), .CP(clk), .Q(\reg_yHat[11][7] ) );
  dff_sg \reg_yHat_reg[11][6]  ( .D(n1775), .CP(clk), .Q(\reg_yHat[11][6] ) );
  dff_sg \reg_yHat_reg[11][5]  ( .D(n1776), .CP(clk), .Q(\reg_yHat[11][5] ) );
  dff_sg \reg_yHat_reg[11][4]  ( .D(n1777), .CP(clk), .Q(\reg_yHat[11][4] ) );
  dff_sg \reg_yHat_reg[11][3]  ( .D(n1778), .CP(clk), .Q(\reg_yHat[11][3] ) );
  dff_sg \reg_yHat_reg[11][2]  ( .D(n1779), .CP(clk), .Q(\reg_yHat[11][2] ) );
  dff_sg \reg_yHat_reg[11][1]  ( .D(n1780), .CP(clk), .Q(\reg_yHat[11][1] ) );
  dff_sg \reg_yHat_reg[11][0]  ( .D(n1781), .CP(clk), .Q(\reg_yHat[11][0] ) );
  dff_sg \reg_yHat_reg[10][19]  ( .D(n1782), .CP(clk), .Q(\reg_yHat[10][19] )
         );
  dff_sg \reg_yHat_reg[10][18]  ( .D(n1783), .CP(clk), .Q(\reg_yHat[10][18] )
         );
  dff_sg \reg_yHat_reg[10][17]  ( .D(n1784), .CP(clk), .Q(\reg_yHat[10][17] )
         );
  dff_sg \reg_yHat_reg[10][16]  ( .D(n1785), .CP(clk), .Q(\reg_yHat[10][16] )
         );
  dff_sg \reg_yHat_reg[10][15]  ( .D(n1786), .CP(clk), .Q(\reg_yHat[10][15] )
         );
  dff_sg \reg_yHat_reg[10][14]  ( .D(n1787), .CP(clk), .Q(\reg_yHat[10][14] )
         );
  dff_sg \reg_yHat_reg[10][13]  ( .D(n1788), .CP(clk), .Q(\reg_yHat[10][13] )
         );
  dff_sg \reg_yHat_reg[10][12]  ( .D(n1789), .CP(clk), .Q(\reg_yHat[10][12] )
         );
  dff_sg \reg_yHat_reg[10][11]  ( .D(n1790), .CP(clk), .Q(\reg_yHat[10][11] )
         );
  dff_sg \reg_yHat_reg[10][10]  ( .D(n1791), .CP(clk), .Q(\reg_yHat[10][10] )
         );
  dff_sg \reg_yHat_reg[10][9]  ( .D(n1792), .CP(clk), .Q(\reg_yHat[10][9] ) );
  dff_sg \reg_yHat_reg[10][8]  ( .D(n1793), .CP(clk), .Q(\reg_yHat[10][8] ) );
  dff_sg \reg_yHat_reg[10][7]  ( .D(n1794), .CP(clk), .Q(\reg_yHat[10][7] ) );
  dff_sg \reg_yHat_reg[10][6]  ( .D(n1795), .CP(clk), .Q(\reg_yHat[10][6] ) );
  dff_sg \reg_yHat_reg[10][5]  ( .D(n1796), .CP(clk), .Q(\reg_yHat[10][5] ) );
  dff_sg \reg_yHat_reg[10][4]  ( .D(n1797), .CP(clk), .Q(\reg_yHat[10][4] ) );
  dff_sg \reg_yHat_reg[10][3]  ( .D(n1798), .CP(clk), .Q(\reg_yHat[10][3] ) );
  dff_sg \reg_yHat_reg[10][2]  ( .D(n1799), .CP(clk), .Q(\reg_yHat[10][2] ) );
  dff_sg \reg_yHat_reg[10][1]  ( .D(n1800), .CP(clk), .Q(\reg_yHat[10][1] ) );
  dff_sg \reg_yHat_reg[10][0]  ( .D(n1801), .CP(clk), .Q(\reg_yHat[10][0] ) );
  dff_sg \reg_yHat_reg[9][19]  ( .D(n1802), .CP(clk), .Q(\reg_yHat[9][19] ) );
  dff_sg \reg_yHat_reg[9][18]  ( .D(n1803), .CP(clk), .Q(\reg_yHat[9][18] ) );
  dff_sg \reg_yHat_reg[9][17]  ( .D(n1804), .CP(clk), .Q(\reg_yHat[9][17] ) );
  dff_sg \reg_yHat_reg[9][16]  ( .D(n1805), .CP(clk), .Q(\reg_yHat[9][16] ) );
  dff_sg \reg_yHat_reg[9][15]  ( .D(n1806), .CP(clk), .Q(\reg_yHat[9][15] ) );
  dff_sg \reg_yHat_reg[9][14]  ( .D(n1807), .CP(clk), .Q(\reg_yHat[9][14] ) );
  dff_sg \reg_yHat_reg[9][13]  ( .D(n1808), .CP(clk), .Q(\reg_yHat[9][13] ) );
  dff_sg \reg_yHat_reg[9][12]  ( .D(n1809), .CP(clk), .Q(\reg_yHat[9][12] ) );
  dff_sg \reg_yHat_reg[9][11]  ( .D(n1810), .CP(clk), .Q(\reg_yHat[9][11] ) );
  dff_sg \reg_yHat_reg[9][10]  ( .D(n1811), .CP(clk), .Q(\reg_yHat[9][10] ) );
  dff_sg \reg_yHat_reg[9][9]  ( .D(n1812), .CP(clk), .Q(\reg_yHat[9][9] ) );
  dff_sg \reg_yHat_reg[9][8]  ( .D(n1813), .CP(clk), .Q(\reg_yHat[9][8] ) );
  dff_sg \reg_yHat_reg[9][7]  ( .D(n1814), .CP(clk), .Q(\reg_yHat[9][7] ) );
  dff_sg \reg_yHat_reg[9][6]  ( .D(n1815), .CP(clk), .Q(\reg_yHat[9][6] ) );
  dff_sg \reg_yHat_reg[9][5]  ( .D(n1816), .CP(clk), .Q(\reg_yHat[9][5] ) );
  dff_sg \reg_yHat_reg[9][4]  ( .D(n1817), .CP(clk), .Q(\reg_yHat[9][4] ) );
  dff_sg \reg_yHat_reg[9][3]  ( .D(n1818), .CP(clk), .Q(\reg_yHat[9][3] ) );
  dff_sg \reg_yHat_reg[9][2]  ( .D(n1819), .CP(clk), .Q(\reg_yHat[9][2] ) );
  dff_sg \reg_yHat_reg[9][1]  ( .D(n1820), .CP(clk), .Q(\reg_yHat[9][1] ) );
  dff_sg \reg_yHat_reg[9][0]  ( .D(n1821), .CP(clk), .Q(\reg_yHat[9][0] ) );
  dff_sg \reg_yHat_reg[8][19]  ( .D(n1822), .CP(clk), .Q(\reg_yHat[8][19] ) );
  dff_sg \reg_yHat_reg[8][18]  ( .D(n1823), .CP(clk), .Q(\reg_yHat[8][18] ) );
  dff_sg \reg_yHat_reg[8][17]  ( .D(n1824), .CP(clk), .Q(\reg_yHat[8][17] ) );
  dff_sg \reg_yHat_reg[8][16]  ( .D(n1825), .CP(clk), .Q(\reg_yHat[8][16] ) );
  dff_sg \reg_yHat_reg[8][15]  ( .D(n1826), .CP(clk), .Q(\reg_yHat[8][15] ) );
  dff_sg \reg_yHat_reg[8][14]  ( .D(n1827), .CP(clk), .Q(\reg_yHat[8][14] ) );
  dff_sg \reg_yHat_reg[8][13]  ( .D(n1828), .CP(clk), .Q(\reg_yHat[8][13] ) );
  dff_sg \reg_yHat_reg[8][12]  ( .D(n1829), .CP(clk), .Q(\reg_yHat[8][12] ) );
  dff_sg \reg_yHat_reg[8][11]  ( .D(n1830), .CP(clk), .Q(\reg_yHat[8][11] ) );
  dff_sg \reg_yHat_reg[8][10]  ( .D(n1831), .CP(clk), .Q(\reg_yHat[8][10] ) );
  dff_sg \reg_yHat_reg[8][9]  ( .D(n1832), .CP(clk), .Q(\reg_yHat[8][9] ) );
  dff_sg \reg_yHat_reg[8][8]  ( .D(n1833), .CP(clk), .Q(\reg_yHat[8][8] ) );
  dff_sg \reg_yHat_reg[8][7]  ( .D(n1834), .CP(clk), .Q(\reg_yHat[8][7] ) );
  dff_sg \reg_yHat_reg[8][6]  ( .D(n1835), .CP(clk), .Q(\reg_yHat[8][6] ) );
  dff_sg \reg_yHat_reg[8][5]  ( .D(n1836), .CP(clk), .Q(\reg_yHat[8][5] ) );
  dff_sg \reg_yHat_reg[8][4]  ( .D(n1837), .CP(clk), .Q(\reg_yHat[8][4] ) );
  dff_sg \reg_yHat_reg[8][3]  ( .D(n1838), .CP(clk), .Q(\reg_yHat[8][3] ) );
  dff_sg \reg_yHat_reg[8][2]  ( .D(n1839), .CP(clk), .Q(\reg_yHat[8][2] ) );
  dff_sg \reg_yHat_reg[8][1]  ( .D(n1840), .CP(clk), .Q(\reg_yHat[8][1] ) );
  dff_sg \reg_yHat_reg[8][0]  ( .D(n1841), .CP(clk), .Q(\reg_yHat[8][0] ) );
  dff_sg \reg_yHat_reg[7][19]  ( .D(n1842), .CP(clk), .Q(\reg_yHat[7][19] ) );
  dff_sg \reg_yHat_reg[7][18]  ( .D(n1843), .CP(clk), .Q(\reg_yHat[7][18] ) );
  dff_sg \reg_yHat_reg[7][17]  ( .D(n1844), .CP(clk), .Q(\reg_yHat[7][17] ) );
  dff_sg \reg_yHat_reg[7][16]  ( .D(n1845), .CP(clk), .Q(\reg_yHat[7][16] ) );
  dff_sg \reg_yHat_reg[7][15]  ( .D(n1846), .CP(clk), .Q(\reg_yHat[7][15] ) );
  dff_sg \reg_yHat_reg[7][14]  ( .D(n1847), .CP(clk), .Q(\reg_yHat[7][14] ) );
  dff_sg \reg_yHat_reg[7][13]  ( .D(n1848), .CP(clk), .Q(\reg_yHat[7][13] ) );
  dff_sg \reg_yHat_reg[7][12]  ( .D(n1849), .CP(clk), .Q(\reg_yHat[7][12] ) );
  dff_sg \reg_yHat_reg[7][11]  ( .D(n1850), .CP(clk), .Q(\reg_yHat[7][11] ) );
  dff_sg \reg_yHat_reg[7][10]  ( .D(n1851), .CP(clk), .Q(\reg_yHat[7][10] ) );
  dff_sg \reg_yHat_reg[7][9]  ( .D(n1852), .CP(clk), .Q(\reg_yHat[7][9] ) );
  dff_sg \reg_yHat_reg[7][8]  ( .D(n1853), .CP(clk), .Q(\reg_yHat[7][8] ) );
  dff_sg \reg_yHat_reg[7][7]  ( .D(n1854), .CP(clk), .Q(\reg_yHat[7][7] ) );
  dff_sg \reg_yHat_reg[7][6]  ( .D(n1855), .CP(clk), .Q(\reg_yHat[7][6] ) );
  dff_sg \reg_yHat_reg[7][5]  ( .D(n1856), .CP(clk), .Q(\reg_yHat[7][5] ) );
  dff_sg \reg_yHat_reg[7][4]  ( .D(n1857), .CP(clk), .Q(\reg_yHat[7][4] ) );
  dff_sg \reg_yHat_reg[7][3]  ( .D(n1858), .CP(clk), .Q(\reg_yHat[7][3] ) );
  dff_sg \reg_yHat_reg[7][2]  ( .D(n1859), .CP(clk), .Q(\reg_yHat[7][2] ) );
  dff_sg \reg_yHat_reg[7][1]  ( .D(n1860), .CP(clk), .Q(\reg_yHat[7][1] ) );
  dff_sg \reg_yHat_reg[7][0]  ( .D(n1861), .CP(clk), .Q(\reg_yHat[7][0] ) );
  dff_sg \reg_yHat_reg[6][19]  ( .D(n1862), .CP(clk), .Q(\reg_yHat[6][19] ) );
  dff_sg \reg_yHat_reg[6][18]  ( .D(n1863), .CP(clk), .Q(\reg_yHat[6][18] ) );
  dff_sg \reg_yHat_reg[6][17]  ( .D(n1864), .CP(clk), .Q(\reg_yHat[6][17] ) );
  dff_sg \reg_yHat_reg[6][16]  ( .D(n1865), .CP(clk), .Q(\reg_yHat[6][16] ) );
  dff_sg \reg_yHat_reg[6][15]  ( .D(n1866), .CP(clk), .Q(\reg_yHat[6][15] ) );
  dff_sg \reg_yHat_reg[6][14]  ( .D(n1867), .CP(clk), .Q(\reg_yHat[6][14] ) );
  dff_sg \reg_yHat_reg[6][13]  ( .D(n1868), .CP(clk), .Q(\reg_yHat[6][13] ) );
  dff_sg \reg_yHat_reg[6][12]  ( .D(n1869), .CP(clk), .Q(\reg_yHat[6][12] ) );
  dff_sg \reg_yHat_reg[6][11]  ( .D(n1870), .CP(clk), .Q(\reg_yHat[6][11] ) );
  dff_sg \reg_yHat_reg[6][10]  ( .D(n1871), .CP(clk), .Q(\reg_yHat[6][10] ) );
  dff_sg \reg_yHat_reg[6][9]  ( .D(n1872), .CP(clk), .Q(\reg_yHat[6][9] ) );
  dff_sg \reg_yHat_reg[6][8]  ( .D(n1873), .CP(clk), .Q(\reg_yHat[6][8] ) );
  dff_sg \reg_yHat_reg[6][7]  ( .D(n1874), .CP(clk), .Q(\reg_yHat[6][7] ) );
  dff_sg \reg_yHat_reg[6][6]  ( .D(n1875), .CP(clk), .Q(\reg_yHat[6][6] ) );
  dff_sg \reg_yHat_reg[6][5]  ( .D(n1876), .CP(clk), .Q(\reg_yHat[6][5] ) );
  dff_sg \reg_yHat_reg[6][4]  ( .D(n1877), .CP(clk), .Q(\reg_yHat[6][4] ) );
  dff_sg \reg_yHat_reg[6][3]  ( .D(n1878), .CP(clk), .Q(\reg_yHat[6][3] ) );
  dff_sg \reg_yHat_reg[6][2]  ( .D(n1879), .CP(clk), .Q(\reg_yHat[6][2] ) );
  dff_sg \reg_yHat_reg[6][1]  ( .D(n1880), .CP(clk), .Q(\reg_yHat[6][1] ) );
  dff_sg \reg_yHat_reg[6][0]  ( .D(n1881), .CP(clk), .Q(\reg_yHat[6][0] ) );
  dff_sg \reg_yHat_reg[5][19]  ( .D(n1882), .CP(clk), .Q(\reg_yHat[5][19] ) );
  dff_sg \reg_yHat_reg[5][18]  ( .D(n1883), .CP(clk), .Q(\reg_yHat[5][18] ) );
  dff_sg \reg_yHat_reg[5][17]  ( .D(n1884), .CP(clk), .Q(\reg_yHat[5][17] ) );
  dff_sg \reg_yHat_reg[5][16]  ( .D(n1885), .CP(clk), .Q(\reg_yHat[5][16] ) );
  dff_sg \reg_yHat_reg[5][15]  ( .D(n1886), .CP(clk), .Q(\reg_yHat[5][15] ) );
  dff_sg \reg_yHat_reg[5][14]  ( .D(n1887), .CP(clk), .Q(\reg_yHat[5][14] ) );
  dff_sg \reg_yHat_reg[5][13]  ( .D(n1888), .CP(clk), .Q(\reg_yHat[5][13] ) );
  dff_sg \reg_yHat_reg[5][12]  ( .D(n1889), .CP(clk), .Q(\reg_yHat[5][12] ) );
  dff_sg \reg_yHat_reg[5][11]  ( .D(n1890), .CP(clk), .Q(\reg_yHat[5][11] ) );
  dff_sg \reg_yHat_reg[5][10]  ( .D(n1891), .CP(clk), .Q(\reg_yHat[5][10] ) );
  dff_sg \reg_yHat_reg[5][9]  ( .D(n1892), .CP(clk), .Q(\reg_yHat[5][9] ) );
  dff_sg \reg_yHat_reg[5][8]  ( .D(n1893), .CP(clk), .Q(\reg_yHat[5][8] ) );
  dff_sg \reg_yHat_reg[5][7]  ( .D(n1894), .CP(clk), .Q(\reg_yHat[5][7] ) );
  dff_sg \reg_yHat_reg[5][6]  ( .D(n1895), .CP(clk), .Q(\reg_yHat[5][6] ) );
  dff_sg \reg_yHat_reg[5][5]  ( .D(n1896), .CP(clk), .Q(\reg_yHat[5][5] ) );
  dff_sg \reg_yHat_reg[5][4]  ( .D(n1897), .CP(clk), .Q(\reg_yHat[5][4] ) );
  dff_sg \reg_yHat_reg[5][3]  ( .D(n1898), .CP(clk), .Q(\reg_yHat[5][3] ) );
  dff_sg \reg_yHat_reg[5][2]  ( .D(n1899), .CP(clk), .Q(\reg_yHat[5][2] ) );
  dff_sg \reg_yHat_reg[5][1]  ( .D(n1900), .CP(clk), .Q(\reg_yHat[5][1] ) );
  dff_sg \reg_yHat_reg[5][0]  ( .D(n1901), .CP(clk), .Q(\reg_yHat[5][0] ) );
  dff_sg \reg_yHat_reg[4][19]  ( .D(n1902), .CP(clk), .Q(\reg_yHat[4][19] ) );
  dff_sg \reg_yHat_reg[4][18]  ( .D(n1903), .CP(clk), .Q(\reg_yHat[4][18] ) );
  dff_sg \reg_yHat_reg[4][17]  ( .D(n1904), .CP(clk), .Q(\reg_yHat[4][17] ) );
  dff_sg \reg_yHat_reg[4][16]  ( .D(n1905), .CP(clk), .Q(\reg_yHat[4][16] ) );
  dff_sg \reg_yHat_reg[4][15]  ( .D(n1906), .CP(clk), .Q(\reg_yHat[4][15] ) );
  dff_sg \reg_yHat_reg[4][14]  ( .D(n1907), .CP(clk), .Q(\reg_yHat[4][14] ) );
  dff_sg \reg_yHat_reg[4][13]  ( .D(n1908), .CP(clk), .Q(\reg_yHat[4][13] ) );
  dff_sg \reg_yHat_reg[4][12]  ( .D(n1909), .CP(clk), .Q(\reg_yHat[4][12] ) );
  dff_sg \reg_yHat_reg[4][11]  ( .D(n1910), .CP(clk), .Q(\reg_yHat[4][11] ) );
  dff_sg \reg_yHat_reg[4][10]  ( .D(n1911), .CP(clk), .Q(\reg_yHat[4][10] ) );
  dff_sg \reg_yHat_reg[4][9]  ( .D(n1912), .CP(clk), .Q(\reg_yHat[4][9] ) );
  dff_sg \reg_yHat_reg[4][8]  ( .D(n1913), .CP(clk), .Q(\reg_yHat[4][8] ) );
  dff_sg \reg_yHat_reg[4][7]  ( .D(n1914), .CP(clk), .Q(\reg_yHat[4][7] ) );
  dff_sg \reg_yHat_reg[4][6]  ( .D(n1915), .CP(clk), .Q(\reg_yHat[4][6] ) );
  dff_sg \reg_yHat_reg[4][5]  ( .D(n1916), .CP(clk), .Q(\reg_yHat[4][5] ) );
  dff_sg \reg_yHat_reg[4][4]  ( .D(n1917), .CP(clk), .Q(\reg_yHat[4][4] ) );
  dff_sg \reg_yHat_reg[4][3]  ( .D(n1918), .CP(clk), .Q(\reg_yHat[4][3] ) );
  dff_sg \reg_yHat_reg[4][2]  ( .D(n1919), .CP(clk), .Q(\reg_yHat[4][2] ) );
  dff_sg \reg_yHat_reg[4][1]  ( .D(n1920), .CP(clk), .Q(\reg_yHat[4][1] ) );
  dff_sg \reg_yHat_reg[4][0]  ( .D(n1921), .CP(clk), .Q(\reg_yHat[4][0] ) );
  dff_sg \reg_yHat_reg[3][19]  ( .D(n1922), .CP(clk), .Q(\reg_yHat[3][19] ) );
  dff_sg \reg_yHat_reg[3][18]  ( .D(n1923), .CP(clk), .Q(\reg_yHat[3][18] ) );
  dff_sg \reg_yHat_reg[3][17]  ( .D(n1924), .CP(clk), .Q(\reg_yHat[3][17] ) );
  dff_sg \reg_yHat_reg[3][16]  ( .D(n1925), .CP(clk), .Q(\reg_yHat[3][16] ) );
  dff_sg \reg_yHat_reg[3][15]  ( .D(n1926), .CP(clk), .Q(\reg_yHat[3][15] ) );
  dff_sg \reg_yHat_reg[3][14]  ( .D(n1927), .CP(clk), .Q(\reg_yHat[3][14] ) );
  dff_sg \reg_yHat_reg[3][13]  ( .D(n1928), .CP(clk), .Q(\reg_yHat[3][13] ) );
  dff_sg \reg_yHat_reg[3][12]  ( .D(n1929), .CP(clk), .Q(\reg_yHat[3][12] ) );
  dff_sg \reg_yHat_reg[3][11]  ( .D(n1930), .CP(clk), .Q(\reg_yHat[3][11] ) );
  dff_sg \reg_yHat_reg[3][10]  ( .D(n1931), .CP(clk), .Q(\reg_yHat[3][10] ) );
  dff_sg \reg_yHat_reg[3][9]  ( .D(n1932), .CP(clk), .Q(\reg_yHat[3][9] ) );
  dff_sg \reg_yHat_reg[3][8]  ( .D(n1933), .CP(clk), .Q(\reg_yHat[3][8] ) );
  dff_sg \reg_yHat_reg[3][7]  ( .D(n1934), .CP(clk), .Q(\reg_yHat[3][7] ) );
  dff_sg \reg_yHat_reg[3][6]  ( .D(n1935), .CP(clk), .Q(\reg_yHat[3][6] ) );
  dff_sg \reg_yHat_reg[3][5]  ( .D(n1936), .CP(clk), .Q(\reg_yHat[3][5] ) );
  dff_sg \reg_yHat_reg[3][4]  ( .D(n1937), .CP(clk), .Q(\reg_yHat[3][4] ) );
  dff_sg \reg_yHat_reg[3][3]  ( .D(n1938), .CP(clk), .Q(\reg_yHat[3][3] ) );
  dff_sg \reg_yHat_reg[3][2]  ( .D(n1939), .CP(clk), .Q(\reg_yHat[3][2] ) );
  dff_sg \reg_yHat_reg[3][1]  ( .D(n1940), .CP(clk), .Q(\reg_yHat[3][1] ) );
  dff_sg \reg_yHat_reg[3][0]  ( .D(n1941), .CP(clk), .Q(\reg_yHat[3][0] ) );
  dff_sg \reg_yHat_reg[2][19]  ( .D(n1942), .CP(clk), .Q(\reg_yHat[2][19] ) );
  dff_sg \reg_yHat_reg[2][18]  ( .D(n1943), .CP(clk), .Q(\reg_yHat[2][18] ) );
  dff_sg \reg_yHat_reg[2][17]  ( .D(n1944), .CP(clk), .Q(\reg_yHat[2][17] ) );
  dff_sg \reg_yHat_reg[2][16]  ( .D(n1945), .CP(clk), .Q(\reg_yHat[2][16] ) );
  dff_sg \reg_yHat_reg[2][15]  ( .D(n1946), .CP(clk), .Q(\reg_yHat[2][15] ) );
  dff_sg \reg_yHat_reg[2][14]  ( .D(n1947), .CP(clk), .Q(\reg_yHat[2][14] ) );
  dff_sg \reg_yHat_reg[2][13]  ( .D(n1948), .CP(clk), .Q(\reg_yHat[2][13] ) );
  dff_sg \reg_yHat_reg[2][12]  ( .D(n1949), .CP(clk), .Q(\reg_yHat[2][12] ) );
  dff_sg \reg_yHat_reg[2][11]  ( .D(n1950), .CP(clk), .Q(\reg_yHat[2][11] ) );
  dff_sg \reg_yHat_reg[2][10]  ( .D(n1951), .CP(clk), .Q(\reg_yHat[2][10] ) );
  dff_sg \reg_yHat_reg[2][9]  ( .D(n1952), .CP(clk), .Q(\reg_yHat[2][9] ) );
  dff_sg \reg_yHat_reg[2][8]  ( .D(n1953), .CP(clk), .Q(\reg_yHat[2][8] ) );
  dff_sg \reg_yHat_reg[2][7]  ( .D(n1954), .CP(clk), .Q(\reg_yHat[2][7] ) );
  dff_sg \reg_yHat_reg[2][6]  ( .D(n1955), .CP(clk), .Q(\reg_yHat[2][6] ) );
  dff_sg \reg_yHat_reg[2][5]  ( .D(n1956), .CP(clk), .Q(\reg_yHat[2][5] ) );
  dff_sg \reg_yHat_reg[2][4]  ( .D(n1957), .CP(clk), .Q(\reg_yHat[2][4] ) );
  dff_sg \reg_yHat_reg[2][3]  ( .D(n1958), .CP(clk), .Q(\reg_yHat[2][3] ) );
  dff_sg \reg_yHat_reg[2][2]  ( .D(n1959), .CP(clk), .Q(\reg_yHat[2][2] ) );
  dff_sg \reg_yHat_reg[2][1]  ( .D(n1960), .CP(clk), .Q(\reg_yHat[2][1] ) );
  dff_sg \reg_yHat_reg[2][0]  ( .D(n1961), .CP(clk), .Q(\reg_yHat[2][0] ) );
  dff_sg \reg_yHat_reg[1][19]  ( .D(n1962), .CP(clk), .Q(\reg_yHat[1][19] ) );
  dff_sg \reg_yHat_reg[1][18]  ( .D(n1963), .CP(clk), .Q(\reg_yHat[1][18] ) );
  dff_sg \reg_yHat_reg[1][17]  ( .D(n1964), .CP(clk), .Q(\reg_yHat[1][17] ) );
  dff_sg \reg_yHat_reg[1][16]  ( .D(n1965), .CP(clk), .Q(\reg_yHat[1][16] ) );
  dff_sg \reg_yHat_reg[1][15]  ( .D(n1966), .CP(clk), .Q(\reg_yHat[1][15] ) );
  dff_sg \reg_yHat_reg[1][14]  ( .D(n1967), .CP(clk), .Q(\reg_yHat[1][14] ) );
  dff_sg \reg_yHat_reg[1][13]  ( .D(n1968), .CP(clk), .Q(\reg_yHat[1][13] ) );
  dff_sg \reg_yHat_reg[1][12]  ( .D(n1969), .CP(clk), .Q(\reg_yHat[1][12] ) );
  dff_sg \reg_yHat_reg[1][11]  ( .D(n1970), .CP(clk), .Q(\reg_yHat[1][11] ) );
  dff_sg \reg_yHat_reg[1][10]  ( .D(n1971), .CP(clk), .Q(\reg_yHat[1][10] ) );
  dff_sg \reg_yHat_reg[1][9]  ( .D(n1972), .CP(clk), .Q(\reg_yHat[1][9] ) );
  dff_sg \reg_yHat_reg[1][8]  ( .D(n1973), .CP(clk), .Q(\reg_yHat[1][8] ) );
  dff_sg \reg_yHat_reg[1][7]  ( .D(n1974), .CP(clk), .Q(\reg_yHat[1][7] ) );
  dff_sg \reg_yHat_reg[1][6]  ( .D(n1975), .CP(clk), .Q(\reg_yHat[1][6] ) );
  dff_sg \reg_yHat_reg[1][5]  ( .D(n1976), .CP(clk), .Q(\reg_yHat[1][5] ) );
  dff_sg \reg_yHat_reg[1][4]  ( .D(n1977), .CP(clk), .Q(\reg_yHat[1][4] ) );
  dff_sg \reg_yHat_reg[1][3]  ( .D(n1978), .CP(clk), .Q(\reg_yHat[1][3] ) );
  dff_sg \reg_yHat_reg[1][2]  ( .D(n1979), .CP(clk), .Q(\reg_yHat[1][2] ) );
  dff_sg \reg_yHat_reg[1][1]  ( .D(n1980), .CP(clk), .Q(\reg_yHat[1][1] ) );
  dff_sg \reg_yHat_reg[1][0]  ( .D(n1981), .CP(clk), .Q(\reg_yHat[1][0] ) );
  dff_sg \reg_yHat_reg[0][19]  ( .D(n1982), .CP(clk), .Q(\reg_yHat[0][19] ) );
  dff_sg \reg_yHat_reg[0][18]  ( .D(n1983), .CP(clk), .Q(\reg_yHat[0][18] ) );
  dff_sg \reg_yHat_reg[0][17]  ( .D(n1984), .CP(clk), .Q(\reg_yHat[0][17] ) );
  dff_sg \reg_yHat_reg[0][16]  ( .D(n1985), .CP(clk), .Q(\reg_yHat[0][16] ) );
  dff_sg \reg_yHat_reg[0][15]  ( .D(n1986), .CP(clk), .Q(\reg_yHat[0][15] ) );
  dff_sg \reg_yHat_reg[0][14]  ( .D(n1987), .CP(clk), .Q(\reg_yHat[0][14] ) );
  dff_sg \reg_yHat_reg[0][13]  ( .D(n1988), .CP(clk), .Q(\reg_yHat[0][13] ) );
  dff_sg \reg_yHat_reg[0][12]  ( .D(n1989), .CP(clk), .Q(\reg_yHat[0][12] ) );
  dff_sg \reg_yHat_reg[0][11]  ( .D(n1990), .CP(clk), .Q(\reg_yHat[0][11] ) );
  dff_sg \reg_yHat_reg[0][10]  ( .D(n1991), .CP(clk), .Q(\reg_yHat[0][10] ) );
  dff_sg \reg_yHat_reg[0][9]  ( .D(n1992), .CP(clk), .Q(\reg_yHat[0][9] ) );
  dff_sg \reg_yHat_reg[0][8]  ( .D(n1993), .CP(clk), .Q(\reg_yHat[0][8] ) );
  dff_sg \reg_yHat_reg[0][7]  ( .D(n1994), .CP(clk), .Q(\reg_yHat[0][7] ) );
  dff_sg \reg_yHat_reg[0][6]  ( .D(n1995), .CP(clk), .Q(\reg_yHat[0][6] ) );
  dff_sg \reg_yHat_reg[0][5]  ( .D(n1996), .CP(clk), .Q(\reg_yHat[0][5] ) );
  dff_sg \reg_yHat_reg[0][4]  ( .D(n1997), .CP(clk), .Q(\reg_yHat[0][4] ) );
  dff_sg \reg_yHat_reg[0][3]  ( .D(n1998), .CP(clk), .Q(\reg_yHat[0][3] ) );
  dff_sg \reg_yHat_reg[0][2]  ( .D(n1999), .CP(clk), .Q(\reg_yHat[0][2] ) );
  dff_sg \reg_yHat_reg[0][1]  ( .D(n2000), .CP(clk), .Q(\reg_yHat[0][1] ) );
  dff_sg \reg_yHat_reg[0][0]  ( .D(n2001), .CP(clk), .Q(\reg_yHat[0][0] ) );
  dff_sg reg_model_reg ( .D(n2002), .CP(clk), .Q(reg_model) );
  \**FFGEN**  \L1_0/abs_reg[14][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3550 ), .force_10(\L1_0/n3551 ), 
        .force_11(1'b0), .QN(n8183) );
  \**FFGEN**  \L1_0/abs_reg[14][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3554 ), .force_10(\L1_0/n3555 ), 
        .force_11(1'b0), .QN(n8184) );
  \**FFGEN**  \L1_0/abs_reg[14][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3558 ), .force_10(\L1_0/n3559 ), 
        .force_11(1'b0), .QN(n8185) );
  \**FFGEN**  \L1_0/abs_reg[14][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3562 ), .force_10(\L1_0/n3563 ), 
        .force_11(1'b0), .QN(n8186) );
  \**FFGEN**  \L1_0/abs_reg[14][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3566 ), .force_10(\L1_0/n3567 ), 
        .force_11(1'b0), .QN(n8187) );
  \**FFGEN**  \L1_0/abs_reg[14][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3570 ), .force_10(\L1_0/n3571 ), 
        .force_11(1'b0), .QN(n8188) );
  \**FFGEN**  \L1_0/abs_reg[14][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3574 ), .force_10(\L1_0/n3575 ), 
        .force_11(1'b0), .QN(n8189) );
  \**FFGEN**  \L1_0/abs_reg[14][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3578 ), .force_10(\L1_0/n3579 ), 
        .force_11(1'b0), .QN(n8190) );
  \**FFGEN**  \L1_0/abs_reg[14][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3582 ), .force_10(\L1_0/n3583 ), 
        .force_11(1'b0), .QN(n8191) );
  \**FFGEN**  \L1_0/abs_reg[14][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3586 ), .force_10(\L1_0/n3587 ), 
        .force_11(1'b0), .QN(n8192) );
  \**FFGEN**  \L1_0/abs_reg[14][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3590 ), .force_10(\L1_0/n3591 ), 
        .force_11(1'b0), .QN(n8193) );
  \**FFGEN**  \L1_0/abs_reg[14][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3594 ), .force_10(\L1_0/n3595 ), 
        .force_11(1'b0), .QN(n8194) );
  \**FFGEN**  \L1_0/abs_reg[14][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3598 ), .force_10(\L1_0/n3599 ), 
        .force_11(1'b0), .QN(n8195) );
  \**FFGEN**  \L1_0/abs_reg[14][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3602 ), .force_10(\L1_0/n3603 ), 
        .force_11(1'b0), .QN(n8196) );
  \**FFGEN**  \L1_0/abs_reg[14][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3606 ), .force_10(\L1_0/n3607 ), 
        .force_11(1'b0), .QN(n8197) );
  \**FFGEN**  \L1_0/abs_reg[14][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3610 ), .force_10(\L1_0/n3611 ), 
        .force_11(1'b0), .QN(n8198) );
  \**FFGEN**  \L1_0/abs_reg[14][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3614 ), .force_10(\L1_0/n3615 ), 
        .force_11(1'b0), .QN(n8199) );
  \**FFGEN**  \L1_0/abs_reg[14][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3618 ), .force_10(\L1_0/n3619 ), 
        .force_11(1'b0), .QN(n8200) );
  \**FFGEN**  \L1_0/abs_reg[14][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3622 ), .force_10(\L1_0/n3623 ), 
        .force_11(1'b0), .Q(n40840), .QN(n8201) );
  \**FFGEN**  \L1_0/abs_reg[14][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3626 ), .force_10(\L1_0/n3627 ), 
        .force_11(1'b0), .Q(n40790), .QN(n8202) );
  \**FFGEN**  \L1_0/abs_reg[13][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3630 ), .force_10(\L1_0/n3631 ), 
        .force_11(1'b0), .QN(n8203) );
  \**FFGEN**  \L1_0/abs_reg[13][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3634 ), .force_10(\L1_0/n3635 ), 
        .force_11(1'b0), .QN(n8204) );
  \**FFGEN**  \L1_0/abs_reg[13][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3638 ), .force_10(\L1_0/n3639 ), 
        .force_11(1'b0), .QN(n8205) );
  \**FFGEN**  \L1_0/abs_reg[13][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3642 ), .force_10(\L1_0/n3643 ), 
        .force_11(1'b0), .QN(n8206) );
  \**FFGEN**  \L1_0/abs_reg[13][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3646 ), .force_10(\L1_0/n3647 ), 
        .force_11(1'b0), .QN(n8207) );
  \**FFGEN**  \L1_0/abs_reg[13][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3650 ), .force_10(\L1_0/n3651 ), 
        .force_11(1'b0), .QN(n8208) );
  \**FFGEN**  \L1_0/abs_reg[13][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3654 ), .force_10(\L1_0/n3655 ), 
        .force_11(1'b0), .QN(n8209) );
  \**FFGEN**  \L1_0/abs_reg[13][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3658 ), .force_10(\L1_0/n3659 ), 
        .force_11(1'b0), .QN(n8210) );
  \**FFGEN**  \L1_0/abs_reg[13][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3662 ), .force_10(\L1_0/n3663 ), 
        .force_11(1'b0), .QN(n8211) );
  \**FFGEN**  \L1_0/abs_reg[13][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3666 ), .force_10(\L1_0/n3667 ), 
        .force_11(1'b0), .QN(n8212) );
  \**FFGEN**  \L1_0/abs_reg[13][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3670 ), .force_10(\L1_0/n3671 ), 
        .force_11(1'b0), .QN(n8213) );
  \**FFGEN**  \L1_0/abs_reg[13][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3674 ), .force_10(\L1_0/n3675 ), 
        .force_11(1'b0), .QN(n8214) );
  \**FFGEN**  \L1_0/abs_reg[13][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3678 ), .force_10(\L1_0/n3679 ), 
        .force_11(1'b0), .QN(n8215) );
  \**FFGEN**  \L1_0/abs_reg[13][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3682 ), .force_10(\L1_0/n3683 ), 
        .force_11(1'b0), .QN(n8216) );
  \**FFGEN**  \L1_0/abs_reg[13][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3686 ), .force_10(\L1_0/n3687 ), 
        .force_11(1'b0), .QN(n8217) );
  \**FFGEN**  \L1_0/abs_reg[13][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3690 ), .force_10(\L1_0/n3691 ), 
        .force_11(1'b0), .QN(n8218) );
  \**FFGEN**  \L1_0/abs_reg[13][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3694 ), .force_10(\L1_0/n3695 ), 
        .force_11(1'b0), .QN(n8219) );
  \**FFGEN**  \L1_0/abs_reg[13][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3698 ), .force_10(\L1_0/n3699 ), 
        .force_11(1'b0), .QN(n8220) );
  \**FFGEN**  \L1_0/abs_reg[13][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3702 ), .force_10(\L1_0/n3703 ), 
        .force_11(1'b0), .Q(n40829), .QN(n8221) );
  \**FFGEN**  \L1_0/abs_reg[13][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3706 ), .force_10(\L1_0/n3707 ), 
        .force_11(1'b0), .QN(n8222) );
  \**FFGEN**  \L1_0/abs_reg[12][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3710 ), .force_10(\L1_0/n3711 ), 
        .force_11(1'b0), .QN(n8223) );
  \**FFGEN**  \L1_0/abs_reg[12][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3714 ), .force_10(\L1_0/n3715 ), 
        .force_11(1'b0), .QN(n8224) );
  \**FFGEN**  \L1_0/abs_reg[12][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3718 ), .force_10(\L1_0/n3719 ), 
        .force_11(1'b0), .QN(n8225) );
  \**FFGEN**  \L1_0/abs_reg[12][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3722 ), .force_10(\L1_0/n3723 ), 
        .force_11(1'b0), .QN(n8226) );
  \**FFGEN**  \L1_0/abs_reg[12][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3726 ), .force_10(\L1_0/n3727 ), 
        .force_11(1'b0), .QN(n8227) );
  \**FFGEN**  \L1_0/abs_reg[12][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3730 ), .force_10(\L1_0/n3731 ), 
        .force_11(1'b0), .QN(n8228) );
  \**FFGEN**  \L1_0/abs_reg[12][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3734 ), .force_10(\L1_0/n3735 ), 
        .force_11(1'b0), .QN(n8229) );
  \**FFGEN**  \L1_0/abs_reg[12][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3738 ), .force_10(\L1_0/n3739 ), 
        .force_11(1'b0), .QN(n8230) );
  \**FFGEN**  \L1_0/abs_reg[12][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3742 ), .force_10(\L1_0/n3743 ), 
        .force_11(1'b0), .QN(n8231) );
  \**FFGEN**  \L1_0/abs_reg[12][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3746 ), .force_10(\L1_0/n3747 ), 
        .force_11(1'b0), .QN(n8232) );
  \**FFGEN**  \L1_0/abs_reg[12][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3750 ), .force_10(\L1_0/n3751 ), 
        .force_11(1'b0), .QN(n8233) );
  \**FFGEN**  \L1_0/abs_reg[12][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3754 ), .force_10(\L1_0/n3755 ), 
        .force_11(1'b0), .QN(n8234) );
  \**FFGEN**  \L1_0/abs_reg[12][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3758 ), .force_10(\L1_0/n3759 ), 
        .force_11(1'b0), .QN(n8235) );
  \**FFGEN**  \L1_0/abs_reg[12][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3762 ), .force_10(\L1_0/n3763 ), 
        .force_11(1'b0), .QN(n8236) );
  \**FFGEN**  \L1_0/abs_reg[12][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3766 ), .force_10(\L1_0/n3767 ), 
        .force_11(1'b0), .QN(n8237) );
  \**FFGEN**  \L1_0/abs_reg[12][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3770 ), .force_10(\L1_0/n3771 ), 
        .force_11(1'b0), .QN(n8238) );
  \**FFGEN**  \L1_0/abs_reg[12][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3774 ), .force_10(\L1_0/n3775 ), 
        .force_11(1'b0), .QN(n8239) );
  \**FFGEN**  \L1_0/abs_reg[12][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3778 ), .force_10(\L1_0/n3779 ), 
        .force_11(1'b0), .QN(n8240) );
  \**FFGEN**  \L1_0/abs_reg[12][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3782 ), .force_10(\L1_0/n3783 ), 
        .force_11(1'b0), .Q(n40826), .QN(n8241) );
  \**FFGEN**  \L1_0/abs_reg[12][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3786 ), .force_10(\L1_0/n3787 ), 
        .force_11(1'b0), .QN(n8242) );
  \**FFGEN**  \L1_0/abs_reg[11][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3790 ), .force_10(\L1_0/n3791 ), 
        .force_11(1'b0), .QN(n8243) );
  \**FFGEN**  \L1_0/abs_reg[11][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3794 ), .force_10(\L1_0/n3795 ), 
        .force_11(1'b0), .QN(n8244) );
  \**FFGEN**  \L1_0/abs_reg[11][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3798 ), .force_10(\L1_0/n3799 ), 
        .force_11(1'b0), .QN(n8245) );
  \**FFGEN**  \L1_0/abs_reg[11][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3802 ), .force_10(\L1_0/n3803 ), 
        .force_11(1'b0), .QN(n8246) );
  \**FFGEN**  \L1_0/abs_reg[11][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3806 ), .force_10(\L1_0/n3807 ), 
        .force_11(1'b0), .QN(n8247) );
  \**FFGEN**  \L1_0/abs_reg[11][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3810 ), .force_10(\L1_0/n3811 ), 
        .force_11(1'b0), .QN(n8248) );
  \**FFGEN**  \L1_0/abs_reg[11][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3814 ), .force_10(\L1_0/n3815 ), 
        .force_11(1'b0), .QN(n8249) );
  \**FFGEN**  \L1_0/abs_reg[11][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3818 ), .force_10(\L1_0/n3819 ), 
        .force_11(1'b0), .QN(n8250) );
  \**FFGEN**  \L1_0/abs_reg[11][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3822 ), .force_10(\L1_0/n3823 ), 
        .force_11(1'b0), .QN(n8251) );
  \**FFGEN**  \L1_0/abs_reg[11][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3826 ), .force_10(\L1_0/n3827 ), 
        .force_11(1'b0), .QN(n8252) );
  \**FFGEN**  \L1_0/abs_reg[11][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3830 ), .force_10(\L1_0/n3831 ), 
        .force_11(1'b0), .QN(n8253) );
  \**FFGEN**  \L1_0/abs_reg[11][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3834 ), .force_10(\L1_0/n3835 ), 
        .force_11(1'b0), .QN(n8254) );
  \**FFGEN**  \L1_0/abs_reg[11][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3838 ), .force_10(\L1_0/n3839 ), 
        .force_11(1'b0), .QN(n8255) );
  \**FFGEN**  \L1_0/abs_reg[11][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3842 ), .force_10(\L1_0/n3843 ), 
        .force_11(1'b0), .QN(n8256) );
  \**FFGEN**  \L1_0/abs_reg[11][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3846 ), .force_10(\L1_0/n3847 ), 
        .force_11(1'b0), .QN(n8257) );
  \**FFGEN**  \L1_0/abs_reg[11][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3850 ), .force_10(\L1_0/n3851 ), 
        .force_11(1'b0), .QN(n8258) );
  \**FFGEN**  \L1_0/abs_reg[11][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3854 ), .force_10(\L1_0/n3855 ), 
        .force_11(1'b0), .QN(n8259) );
  \**FFGEN**  \L1_0/abs_reg[11][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3858 ), .force_10(\L1_0/n3859 ), 
        .force_11(1'b0), .QN(n8260) );
  \**FFGEN**  \L1_0/abs_reg[11][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3862 ), .force_10(\L1_0/n3863 ), 
        .force_11(1'b0), .Q(n40823), .QN(n8261) );
  \**FFGEN**  \L1_0/abs_reg[11][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3866 ), .force_10(\L1_0/n3867 ), 
        .force_11(1'b0), .QN(n8262) );
  \**FFGEN**  \L1_0/abs_reg[10][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3870 ), .force_10(\L1_0/n3871 ), 
        .force_11(1'b0), .QN(n8263) );
  \**FFGEN**  \L1_0/abs_reg[10][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3874 ), .force_10(\L1_0/n3875 ), 
        .force_11(1'b0), .QN(n8264) );
  \**FFGEN**  \L1_0/abs_reg[10][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3878 ), .force_10(\L1_0/n3879 ), 
        .force_11(1'b0), .QN(n8265) );
  \**FFGEN**  \L1_0/abs_reg[10][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3882 ), .force_10(\L1_0/n3883 ), 
        .force_11(1'b0), .QN(n8266) );
  \**FFGEN**  \L1_0/abs_reg[10][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3886 ), .force_10(\L1_0/n3887 ), 
        .force_11(1'b0), .QN(n8267) );
  \**FFGEN**  \L1_0/abs_reg[10][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3890 ), .force_10(\L1_0/n3891 ), 
        .force_11(1'b0), .QN(n8268) );
  \**FFGEN**  \L1_0/abs_reg[10][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3894 ), .force_10(\L1_0/n3895 ), 
        .force_11(1'b0), .QN(n8269) );
  \**FFGEN**  \L1_0/abs_reg[10][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3898 ), .force_10(\L1_0/n3899 ), 
        .force_11(1'b0), .QN(n8270) );
  \**FFGEN**  \L1_0/abs_reg[10][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3902 ), .force_10(\L1_0/n3903 ), 
        .force_11(1'b0), .QN(n8271) );
  \**FFGEN**  \L1_0/abs_reg[10][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3906 ), .force_10(\L1_0/n3907 ), 
        .force_11(1'b0), .QN(n8272) );
  \**FFGEN**  \L1_0/abs_reg[10][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3910 ), .force_10(\L1_0/n3911 ), 
        .force_11(1'b0), .QN(n8273) );
  \**FFGEN**  \L1_0/abs_reg[10][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3914 ), .force_10(\L1_0/n3915 ), 
        .force_11(1'b0), .QN(n8274) );
  \**FFGEN**  \L1_0/abs_reg[10][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3918 ), .force_10(\L1_0/n3919 ), 
        .force_11(1'b0), .QN(n8275) );
  \**FFGEN**  \L1_0/abs_reg[10][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3922 ), .force_10(\L1_0/n3923 ), 
        .force_11(1'b0), .QN(n8276) );
  \**FFGEN**  \L1_0/abs_reg[10][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3926 ), .force_10(\L1_0/n3927 ), 
        .force_11(1'b0), .QN(n8277) );
  \**FFGEN**  \L1_0/abs_reg[10][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3930 ), .force_10(\L1_0/n3931 ), 
        .force_11(1'b0), .QN(n8278) );
  \**FFGEN**  \L1_0/abs_reg[10][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3934 ), .force_10(\L1_0/n3935 ), 
        .force_11(1'b0), .QN(n8279) );
  \**FFGEN**  \L1_0/abs_reg[10][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3938 ), .force_10(\L1_0/n3939 ), 
        .force_11(1'b0), .QN(n8280) );
  \**FFGEN**  \L1_0/abs_reg[10][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3942 ), .force_10(\L1_0/n3943 ), 
        .force_11(1'b0), .Q(n40820), .QN(n8281) );
  \**FFGEN**  \L1_0/abs_reg[10][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3946 ), .force_10(\L1_0/n3947 ), 
        .force_11(1'b0), .QN(n8282) );
  \**FFGEN**  \L1_0/abs_reg[9][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3950 ), .force_10(\L1_0/n3951 ), 
        .force_11(1'b0), .QN(n8283) );
  \**FFGEN**  \L1_0/abs_reg[9][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3954 ), .force_10(\L1_0/n3955 ), 
        .force_11(1'b0), .QN(n8284) );
  \**FFGEN**  \L1_0/abs_reg[9][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3958 ), .force_10(\L1_0/n3959 ), 
        .force_11(1'b0), .QN(n8285) );
  \**FFGEN**  \L1_0/abs_reg[9][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3962 ), .force_10(\L1_0/n3963 ), 
        .force_11(1'b0), .QN(n8286) );
  \**FFGEN**  \L1_0/abs_reg[9][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3966 ), .force_10(\L1_0/n3967 ), 
        .force_11(1'b0), .QN(n8287) );
  \**FFGEN**  \L1_0/abs_reg[9][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3970 ), .force_10(\L1_0/n3971 ), 
        .force_11(1'b0), .QN(n8288) );
  \**FFGEN**  \L1_0/abs_reg[9][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3974 ), .force_10(\L1_0/n3975 ), 
        .force_11(1'b0), .QN(n8289) );
  \**FFGEN**  \L1_0/abs_reg[9][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3978 ), .force_10(\L1_0/n3979 ), 
        .force_11(1'b0), .QN(n8290) );
  \**FFGEN**  \L1_0/abs_reg[9][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3982 ), .force_10(\L1_0/n3983 ), 
        .force_11(1'b0), .QN(n8291) );
  \**FFGEN**  \L1_0/abs_reg[9][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3986 ), .force_10(\L1_0/n3987 ), 
        .force_11(1'b0), .QN(n8292) );
  \**FFGEN**  \L1_0/abs_reg[9][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3990 ), .force_10(\L1_0/n3991 ), 
        .force_11(1'b0), .QN(n8293) );
  \**FFGEN**  \L1_0/abs_reg[9][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3994 ), .force_10(\L1_0/n3995 ), 
        .force_11(1'b0), .QN(n8294) );
  \**FFGEN**  \L1_0/abs_reg[9][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3998 ), .force_10(\L1_0/n3999 ), 
        .force_11(1'b0), .QN(n8295) );
  \**FFGEN**  \L1_0/abs_reg[9][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4002 ), .force_10(\L1_0/n4003 ), 
        .force_11(1'b0), .QN(n8296) );
  \**FFGEN**  \L1_0/abs_reg[9][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4006 ), .force_10(\L1_0/n4007 ), 
        .force_11(1'b0), .QN(n8297) );
  \**FFGEN**  \L1_0/abs_reg[9][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4010 ), .force_10(\L1_0/n4011 ), 
        .force_11(1'b0), .QN(n8298) );
  \**FFGEN**  \L1_0/abs_reg[9][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4014 ), .force_10(\L1_0/n4015 ), 
        .force_11(1'b0), .QN(n8299) );
  \**FFGEN**  \L1_0/abs_reg[9][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4018 ), .force_10(\L1_0/n4019 ), 
        .force_11(1'b0), .QN(n8300) );
  \**FFGEN**  \L1_0/abs_reg[9][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4022 ), .force_10(\L1_0/n4023 ), 
        .force_11(1'b0), .Q(n40819), .QN(n8301) );
  \**FFGEN**  \L1_0/abs_reg[9][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4026 ), .force_10(\L1_0/n4027 ), 
        .force_11(1'b0), .QN(n8302) );
  \**FFGEN**  \L1_0/abs_reg[8][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4030 ), .force_10(\L1_0/n4031 ), 
        .force_11(1'b0), .QN(n8303) );
  \**FFGEN**  \L1_0/abs_reg[8][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4034 ), .force_10(\L1_0/n4035 ), 
        .force_11(1'b0), .QN(n8304) );
  \**FFGEN**  \L1_0/abs_reg[8][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4038 ), .force_10(\L1_0/n4039 ), 
        .force_11(1'b0), .QN(n8305) );
  \**FFGEN**  \L1_0/abs_reg[8][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4042 ), .force_10(\L1_0/n4043 ), 
        .force_11(1'b0), .QN(n8306) );
  \**FFGEN**  \L1_0/abs_reg[8][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4046 ), .force_10(\L1_0/n4047 ), 
        .force_11(1'b0), .QN(n8307) );
  \**FFGEN**  \L1_0/abs_reg[8][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4050 ), .force_10(\L1_0/n4051 ), 
        .force_11(1'b0), .QN(n8308) );
  \**FFGEN**  \L1_0/abs_reg[8][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4054 ), .force_10(\L1_0/n4055 ), 
        .force_11(1'b0), .QN(n8309) );
  \**FFGEN**  \L1_0/abs_reg[8][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4058 ), .force_10(\L1_0/n4059 ), 
        .force_11(1'b0), .QN(n8310) );
  \**FFGEN**  \L1_0/abs_reg[8][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4062 ), .force_10(\L1_0/n4063 ), 
        .force_11(1'b0), .QN(n8311) );
  \**FFGEN**  \L1_0/abs_reg[8][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4066 ), .force_10(\L1_0/n4067 ), 
        .force_11(1'b0), .QN(n8312) );
  \**FFGEN**  \L1_0/abs_reg[8][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4070 ), .force_10(\L1_0/n4071 ), 
        .force_11(1'b0), .QN(n8313) );
  \**FFGEN**  \L1_0/abs_reg[8][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4074 ), .force_10(\L1_0/n4075 ), 
        .force_11(1'b0), .QN(n8314) );
  \**FFGEN**  \L1_0/abs_reg[8][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4078 ), .force_10(\L1_0/n4079 ), 
        .force_11(1'b0), .QN(n8315) );
  \**FFGEN**  \L1_0/abs_reg[8][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4082 ), .force_10(\L1_0/n4083 ), 
        .force_11(1'b0), .QN(n8316) );
  \**FFGEN**  \L1_0/abs_reg[8][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4086 ), .force_10(\L1_0/n4087 ), 
        .force_11(1'b0), .QN(n8317) );
  \**FFGEN**  \L1_0/abs_reg[8][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4090 ), .force_10(\L1_0/n4091 ), 
        .force_11(1'b0), .QN(n8318) );
  \**FFGEN**  \L1_0/abs_reg[8][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4094 ), .force_10(\L1_0/n4095 ), 
        .force_11(1'b0), .QN(n8319) );
  \**FFGEN**  \L1_0/abs_reg[8][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4098 ), .force_10(\L1_0/n4099 ), 
        .force_11(1'b0), .QN(n8320) );
  \**FFGEN**  \L1_0/abs_reg[8][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4102 ), .force_10(\L1_0/n4103 ), 
        .force_11(1'b0), .Q(n40816), .QN(n8321) );
  \**FFGEN**  \L1_0/abs_reg[8][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4106 ), .force_10(\L1_0/n4107 ), 
        .force_11(1'b0), .QN(n8322) );
  \**FFGEN**  \L1_0/abs_reg[7][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4110 ), .force_10(\L1_0/n4111 ), 
        .force_11(1'b0), .QN(n8323) );
  \**FFGEN**  \L1_0/abs_reg[7][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4114 ), .force_10(\L1_0/n4115 ), 
        .force_11(1'b0), .QN(n8324) );
  \**FFGEN**  \L1_0/abs_reg[7][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4118 ), .force_10(\L1_0/n4119 ), 
        .force_11(1'b0), .QN(n8325) );
  \**FFGEN**  \L1_0/abs_reg[7][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4122 ), .force_10(\L1_0/n4123 ), 
        .force_11(1'b0), .QN(n8326) );
  \**FFGEN**  \L1_0/abs_reg[7][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4126 ), .force_10(\L1_0/n4127 ), 
        .force_11(1'b0), .QN(n8327) );
  \**FFGEN**  \L1_0/abs_reg[7][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4130 ), .force_10(\L1_0/n4131 ), 
        .force_11(1'b0), .QN(n8328) );
  \**FFGEN**  \L1_0/abs_reg[7][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4134 ), .force_10(\L1_0/n4135 ), 
        .force_11(1'b0), .QN(n8329) );
  \**FFGEN**  \L1_0/abs_reg[7][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4138 ), .force_10(\L1_0/n4139 ), 
        .force_11(1'b0), .QN(n8330) );
  \**FFGEN**  \L1_0/abs_reg[7][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4142 ), .force_10(\L1_0/n4143 ), 
        .force_11(1'b0), .QN(n8331) );
  \**FFGEN**  \L1_0/abs_reg[7][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4146 ), .force_10(\L1_0/n4147 ), 
        .force_11(1'b0), .QN(n8332) );
  \**FFGEN**  \L1_0/abs_reg[7][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4150 ), .force_10(\L1_0/n4151 ), 
        .force_11(1'b0), .QN(n8333) );
  \**FFGEN**  \L1_0/abs_reg[7][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4154 ), .force_10(\L1_0/n4155 ), 
        .force_11(1'b0), .QN(n8334) );
  \**FFGEN**  \L1_0/abs_reg[7][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4158 ), .force_10(\L1_0/n4159 ), 
        .force_11(1'b0), .QN(n8335) );
  \**FFGEN**  \L1_0/abs_reg[7][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4162 ), .force_10(\L1_0/n4163 ), 
        .force_11(1'b0), .QN(n8336) );
  \**FFGEN**  \L1_0/abs_reg[7][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4166 ), .force_10(\L1_0/n4167 ), 
        .force_11(1'b0), .QN(n8337) );
  \**FFGEN**  \L1_0/abs_reg[7][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4170 ), .force_10(\L1_0/n4171 ), 
        .force_11(1'b0), .QN(n8338) );
  \**FFGEN**  \L1_0/abs_reg[7][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4174 ), .force_10(\L1_0/n4175 ), 
        .force_11(1'b0), .QN(n8339) );
  \**FFGEN**  \L1_0/abs_reg[7][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4178 ), .force_10(\L1_0/n4179 ), 
        .force_11(1'b0), .QN(n8340) );
  \**FFGEN**  \L1_0/abs_reg[7][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4182 ), .force_10(\L1_0/n4183 ), 
        .force_11(1'b0), .Q(n40814), .QN(n8341) );
  \**FFGEN**  \L1_0/abs_reg[7][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4186 ), .force_10(\L1_0/n4187 ), 
        .force_11(1'b0), .QN(n8342) );
  \**FFGEN**  \L1_0/abs_reg[6][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4190 ), .force_10(\L1_0/n4191 ), 
        .force_11(1'b0), .QN(n8343) );
  \**FFGEN**  \L1_0/abs_reg[6][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4194 ), .force_10(\L1_0/n4195 ), 
        .force_11(1'b0), .Q(n40774), .QN(n8344) );
  \**FFGEN**  \L1_0/abs_reg[6][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4198 ), .force_10(\L1_0/n4199 ), 
        .force_11(1'b0), .Q(n40762), .QN(n8345) );
  \**FFGEN**  \L1_0/abs_reg[6][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4202 ), .force_10(\L1_0/n4203 ), 
        .force_11(1'b0), .Q(n40811), .QN(n8346) );
  \**FFGEN**  \L1_0/abs_reg[6][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4206 ), .force_10(\L1_0/n4207 ), 
        .force_11(1'b0), .Q(n40761), .QN(n8347) );
  \**FFGEN**  \L1_0/abs_reg[6][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4210 ), .force_10(\L1_0/n4211 ), 
        .force_11(1'b0), .Q(n40809), .QN(n8348) );
  \**FFGEN**  \L1_0/abs_reg[6][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4214 ), .force_10(\L1_0/n4215 ), 
        .force_11(1'b0), .Q(n40753), .QN(n8349) );
  \**FFGEN**  \L1_0/abs_reg[6][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4218 ), .force_10(\L1_0/n4219 ), 
        .force_11(1'b0), .Q(n40755), .QN(n8350) );
  \**FFGEN**  \L1_0/abs_reg[6][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4222 ), .force_10(\L1_0/n4223 ), 
        .force_11(1'b0), .Q(n40767), .QN(n8351) );
  \**FFGEN**  \L1_0/abs_reg[6][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4226 ), .force_10(\L1_0/n4227 ), 
        .force_11(1'b0), .Q(n40758), .QN(n8352) );
  \**FFGEN**  \L1_0/abs_reg[6][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4230 ), .force_10(\L1_0/n4231 ), 
        .force_11(1'b0), .Q(n40854), .QN(n8353) );
  \**FFGEN**  \L1_0/abs_reg[6][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4234 ), .force_10(\L1_0/n4235 ), 
        .force_11(1'b0), .Q(n40766), .QN(n8354) );
  \**FFGEN**  \L1_0/abs_reg[6][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4238 ), .force_10(\L1_0/n4239 ), 
        .force_11(1'b0), .Q(n40757), .QN(n8355) );
  \**FFGEN**  \L1_0/abs_reg[6][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4242 ), .force_10(\L1_0/n4243 ), 
        .force_11(1'b0), .Q(n40855), .QN(n8356) );
  \**FFGEN**  \L1_0/abs_reg[6][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4246 ), .force_10(\L1_0/n4247 ), 
        .force_11(1'b0), .Q(n40765), .QN(n8357) );
  \**FFGEN**  \L1_0/abs_reg[6][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4250 ), .force_10(\L1_0/n4251 ), 
        .force_11(1'b0), .Q(n40857), .QN(n8358) );
  \**FFGEN**  \L1_0/abs_reg[6][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4254 ), .force_10(\L1_0/n4255 ), 
        .force_11(1'b0), .Q(n40783), .QN(n8359) );
  \**FFGEN**  \L1_0/abs_reg[6][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4258 ), .force_10(\L1_0/n4259 ), 
        .force_11(1'b0), .QN(n8360) );
  \**FFGEN**  \L1_0/abs_reg[6][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4262 ), .force_10(\L1_0/n4263 ), 
        .force_11(1'b0), .Q(n40834), .QN(n8361) );
  \**FFGEN**  \L1_0/abs_reg[6][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4266 ), .force_10(\L1_0/n4267 ), 
        .force_11(1'b0), .QN(n8362) );
  \**FFGEN**  \L1_0/abs_reg[5][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4270 ), .force_10(\L1_0/n4271 ), 
        .force_11(1'b0), .QN(n8363) );
  \**FFGEN**  \L1_0/abs_reg[5][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4274 ), .force_10(\L1_0/n4275 ), 
        .force_11(1'b0), .QN(n8364) );
  \**FFGEN**  \L1_0/abs_reg[5][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4278 ), .force_10(\L1_0/n4279 ), 
        .force_11(1'b0), .QN(n8365) );
  \**FFGEN**  \L1_0/abs_reg[5][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4282 ), .force_10(\L1_0/n4283 ), 
        .force_11(1'b0), .QN(n8366) );
  \**FFGEN**  \L1_0/abs_reg[5][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4286 ), .force_10(\L1_0/n4287 ), 
        .force_11(1'b0), .QN(n8367) );
  \**FFGEN**  \L1_0/abs_reg[5][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4290 ), .force_10(\L1_0/n4291 ), 
        .force_11(1'b0), .QN(n8368) );
  \**FFGEN**  \L1_0/abs_reg[5][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4294 ), .force_10(\L1_0/n4295 ), 
        .force_11(1'b0), .QN(n8369) );
  \**FFGEN**  \L1_0/abs_reg[5][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4298 ), .force_10(\L1_0/n4299 ), 
        .force_11(1'b0), .QN(n8370) );
  \**FFGEN**  \L1_0/abs_reg[5][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4302 ), .force_10(\L1_0/n4303 ), 
        .force_11(1'b0), .QN(n8371) );
  \**FFGEN**  \L1_0/abs_reg[5][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4306 ), .force_10(\L1_0/n4307 ), 
        .force_11(1'b0), .QN(n8372) );
  \**FFGEN**  \L1_0/abs_reg[5][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4310 ), .force_10(\L1_0/n4311 ), 
        .force_11(1'b0), .QN(n8373) );
  \**FFGEN**  \L1_0/abs_reg[5][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4314 ), .force_10(\L1_0/n4315 ), 
        .force_11(1'b0), .QN(n8374) );
  \**FFGEN**  \L1_0/abs_reg[5][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4318 ), .force_10(\L1_0/n4319 ), 
        .force_11(1'b0), .QN(n8375) );
  \**FFGEN**  \L1_0/abs_reg[5][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4322 ), .force_10(\L1_0/n4323 ), 
        .force_11(1'b0), .QN(n8376) );
  \**FFGEN**  \L1_0/abs_reg[5][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4326 ), .force_10(\L1_0/n4327 ), 
        .force_11(1'b0), .QN(n8377) );
  \**FFGEN**  \L1_0/abs_reg[5][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4330 ), .force_10(\L1_0/n4331 ), 
        .force_11(1'b0), .QN(n8378) );
  \**FFGEN**  \L1_0/abs_reg[5][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4334 ), .force_10(\L1_0/n4335 ), 
        .force_11(1'b0), .QN(n8379) );
  \**FFGEN**  \L1_0/abs_reg[5][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4338 ), .force_10(\L1_0/n4339 ), 
        .force_11(1'b0), .QN(n8380) );
  \**FFGEN**  \L1_0/abs_reg[5][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4342 ), .force_10(\L1_0/n4343 ), 
        .force_11(1'b0), .Q(n40824), .QN(n8381) );
  \**FFGEN**  \L1_0/abs_reg[5][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4346 ), .force_10(\L1_0/n4347 ), 
        .force_11(1'b0), .QN(n8382) );
  \**FFGEN**  \L1_0/abs_reg[4][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4350 ), .force_10(\L1_0/n4351 ), 
        .force_11(1'b0), .QN(n8383) );
  \**FFGEN**  \L1_0/abs_reg[4][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4354 ), .force_10(\L1_0/n4355 ), 
        .force_11(1'b0), .QN(n8384) );
  \**FFGEN**  \L1_0/abs_reg[4][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4358 ), .force_10(\L1_0/n4359 ), 
        .force_11(1'b0), .QN(n8385) );
  \**FFGEN**  \L1_0/abs_reg[4][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4362 ), .force_10(\L1_0/n4363 ), 
        .force_11(1'b0), .QN(n8386) );
  \**FFGEN**  \L1_0/abs_reg[4][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4366 ), .force_10(\L1_0/n4367 ), 
        .force_11(1'b0), .QN(n8387) );
  \**FFGEN**  \L1_0/abs_reg[4][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4370 ), .force_10(\L1_0/n4371 ), 
        .force_11(1'b0), .QN(n8388) );
  \**FFGEN**  \L1_0/abs_reg[4][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4374 ), .force_10(\L1_0/n4375 ), 
        .force_11(1'b0), .QN(n8389) );
  \**FFGEN**  \L1_0/abs_reg[4][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4378 ), .force_10(\L1_0/n4379 ), 
        .force_11(1'b0), .QN(n8390) );
  \**FFGEN**  \L1_0/abs_reg[4][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4382 ), .force_10(\L1_0/n4383 ), 
        .force_11(1'b0), .QN(n8391) );
  \**FFGEN**  \L1_0/abs_reg[4][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4386 ), .force_10(\L1_0/n4387 ), 
        .force_11(1'b0), .QN(n8392) );
  \**FFGEN**  \L1_0/abs_reg[4][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4390 ), .force_10(\L1_0/n4391 ), 
        .force_11(1'b0), .QN(n8393) );
  \**FFGEN**  \L1_0/abs_reg[4][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4394 ), .force_10(\L1_0/n4395 ), 
        .force_11(1'b0), .QN(n8394) );
  \**FFGEN**  \L1_0/abs_reg[4][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4398 ), .force_10(\L1_0/n4399 ), 
        .force_11(1'b0), .QN(n8395) );
  \**FFGEN**  \L1_0/abs_reg[4][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4402 ), .force_10(\L1_0/n4403 ), 
        .force_11(1'b0), .QN(n8396) );
  \**FFGEN**  \L1_0/abs_reg[4][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4406 ), .force_10(\L1_0/n4407 ), 
        .force_11(1'b0), .QN(n8397) );
  \**FFGEN**  \L1_0/abs_reg[4][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4410 ), .force_10(\L1_0/n4411 ), 
        .force_11(1'b0), .QN(n8398) );
  \**FFGEN**  \L1_0/abs_reg[4][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4414 ), .force_10(\L1_0/n4415 ), 
        .force_11(1'b0), .QN(n8399) );
  \**FFGEN**  \L1_0/abs_reg[4][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4418 ), .force_10(\L1_0/n4419 ), 
        .force_11(1'b0), .QN(n8400) );
  \**FFGEN**  \L1_0/abs_reg[4][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4422 ), .force_10(\L1_0/n4423 ), 
        .force_11(1'b0), .Q(n40832), .QN(n8401) );
  \**FFGEN**  \L1_0/abs_reg[4][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4426 ), .force_10(\L1_0/n4427 ), 
        .force_11(1'b0), .QN(n8402) );
  \**FFGEN**  \L1_0/abs_reg[3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4430 ), .force_10(\L1_0/n4431 ), 
        .force_11(1'b0), .QN(n8403) );
  \**FFGEN**  \L1_0/abs_reg[3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4434 ), .force_10(\L1_0/n4435 ), 
        .force_11(1'b0), .QN(n8404) );
  \**FFGEN**  \L1_0/abs_reg[3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4438 ), .force_10(\L1_0/n4439 ), 
        .force_11(1'b0), .QN(n8405) );
  \**FFGEN**  \L1_0/abs_reg[3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4442 ), .force_10(\L1_0/n4443 ), 
        .force_11(1'b0), .QN(n8406) );
  \**FFGEN**  \L1_0/abs_reg[3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4446 ), .force_10(\L1_0/n4447 ), 
        .force_11(1'b0), .QN(n8407) );
  \**FFGEN**  \L1_0/abs_reg[3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4450 ), .force_10(\L1_0/n4451 ), 
        .force_11(1'b0), .QN(n8408) );
  \**FFGEN**  \L1_0/abs_reg[3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4454 ), .force_10(\L1_0/n4455 ), 
        .force_11(1'b0), .QN(n8409) );
  \**FFGEN**  \L1_0/abs_reg[3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4458 ), .force_10(\L1_0/n4459 ), 
        .force_11(1'b0), .QN(n8410) );
  \**FFGEN**  \L1_0/abs_reg[3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4462 ), .force_10(\L1_0/n4463 ), 
        .force_11(1'b0), .QN(n8411) );
  \**FFGEN**  \L1_0/abs_reg[3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4466 ), .force_10(\L1_0/n4467 ), 
        .force_11(1'b0), .QN(n8412) );
  \**FFGEN**  \L1_0/abs_reg[3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4470 ), .force_10(\L1_0/n4471 ), 
        .force_11(1'b0), .QN(n8413) );
  \**FFGEN**  \L1_0/abs_reg[3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4474 ), .force_10(\L1_0/n4475 ), 
        .force_11(1'b0), .QN(n8414) );
  \**FFGEN**  \L1_0/abs_reg[3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4478 ), .force_10(\L1_0/n4479 ), 
        .force_11(1'b0), .QN(n8415) );
  \**FFGEN**  \L1_0/abs_reg[3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4482 ), .force_10(\L1_0/n4483 ), 
        .force_11(1'b0), .QN(n8416) );
  \**FFGEN**  \L1_0/abs_reg[3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4486 ), .force_10(\L1_0/n4487 ), 
        .force_11(1'b0), .QN(n8417) );
  \**FFGEN**  \L1_0/abs_reg[3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4490 ), .force_10(\L1_0/n4491 ), 
        .force_11(1'b0), .QN(n8418) );
  \**FFGEN**  \L1_0/abs_reg[3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4494 ), .force_10(\L1_0/n4495 ), 
        .force_11(1'b0), .QN(n8419) );
  \**FFGEN**  \L1_0/abs_reg[3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4498 ), .force_10(\L1_0/n4499 ), 
        .force_11(1'b0), .QN(n8420) );
  \**FFGEN**  \L1_0/abs_reg[3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4502 ), .force_10(\L1_0/n4503 ), 
        .force_11(1'b0), .Q(n40837), .QN(n8421) );
  \**FFGEN**  \L1_0/abs_reg[3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4506 ), .force_10(\L1_0/n4507 ), 
        .force_11(1'b0), .QN(n8422) );
  \**FFGEN**  \L1_0/abs_reg[2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4510 ), .force_10(\L1_0/n4511 ), 
        .force_11(1'b0), .QN(n8423) );
  \**FFGEN**  \L1_0/abs_reg[2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4514 ), .force_10(\L1_0/n4515 ), 
        .force_11(1'b0), .QN(n8424) );
  \**FFGEN**  \L1_0/abs_reg[2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4518 ), .force_10(\L1_0/n4519 ), 
        .force_11(1'b0), .QN(n8425) );
  \**FFGEN**  \L1_0/abs_reg[2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4522 ), .force_10(\L1_0/n4523 ), 
        .force_11(1'b0), .QN(n8426) );
  \**FFGEN**  \L1_0/abs_reg[2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4526 ), .force_10(\L1_0/n4527 ), 
        .force_11(1'b0), .QN(n8427) );
  \**FFGEN**  \L1_0/abs_reg[2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4530 ), .force_10(\L1_0/n4531 ), 
        .force_11(1'b0), .QN(n8428) );
  \**FFGEN**  \L1_0/abs_reg[2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4534 ), .force_10(\L1_0/n4535 ), 
        .force_11(1'b0), .QN(n8429) );
  \**FFGEN**  \L1_0/abs_reg[2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4538 ), .force_10(\L1_0/n4539 ), 
        .force_11(1'b0), .QN(n8430) );
  \**FFGEN**  \L1_0/abs_reg[2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4542 ), .force_10(\L1_0/n4543 ), 
        .force_11(1'b0), .QN(n8431) );
  \**FFGEN**  \L1_0/abs_reg[2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4546 ), .force_10(\L1_0/n4547 ), 
        .force_11(1'b0), .QN(n8432) );
  \**FFGEN**  \L1_0/abs_reg[2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4550 ), .force_10(\L1_0/n4551 ), 
        .force_11(1'b0), .QN(n8433) );
  \**FFGEN**  \L1_0/abs_reg[2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4554 ), .force_10(\L1_0/n4555 ), 
        .force_11(1'b0), .QN(n8434) );
  \**FFGEN**  \L1_0/abs_reg[2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4558 ), .force_10(\L1_0/n4559 ), 
        .force_11(1'b0), .QN(n8435) );
  \**FFGEN**  \L1_0/abs_reg[2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4562 ), .force_10(\L1_0/n4563 ), 
        .force_11(1'b0), .QN(n8436) );
  \**FFGEN**  \L1_0/abs_reg[2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4566 ), .force_10(\L1_0/n4567 ), 
        .force_11(1'b0), .QN(n8437) );
  \**FFGEN**  \L1_0/abs_reg[2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4570 ), .force_10(\L1_0/n4571 ), 
        .force_11(1'b0), .QN(n8438) );
  \**FFGEN**  \L1_0/abs_reg[2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4574 ), .force_10(\L1_0/n4575 ), 
        .force_11(1'b0), .QN(n8439) );
  \**FFGEN**  \L1_0/abs_reg[2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4578 ), .force_10(\L1_0/n4579 ), 
        .force_11(1'b0), .QN(n8440) );
  \**FFGEN**  \L1_0/abs_reg[2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4582 ), .force_10(\L1_0/n4583 ), 
        .force_11(1'b0), .Q(n40830), .QN(n8441) );
  \**FFGEN**  \L1_0/abs_reg[2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4586 ), .force_10(\L1_0/n4587 ), 
        .force_11(1'b0), .QN(n8442) );
  \**FFGEN**  \L1_0/abs_reg[1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4590 ), .force_10(\L1_0/n4591 ), 
        .force_11(1'b0), .QN(n8443) );
  \**FFGEN**  \L1_0/abs_reg[1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4594 ), .force_10(\L1_0/n4595 ), 
        .force_11(1'b0), .QN(n8444) );
  \**FFGEN**  \L1_0/abs_reg[1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4598 ), .force_10(\L1_0/n4599 ), 
        .force_11(1'b0), .Q(n40777), .QN(n8445) );
  \**FFGEN**  \L1_0/abs_reg[1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4602 ), .force_10(\L1_0/n4603 ), 
        .force_11(1'b0), .Q(n40772), .QN(n8446) );
  \**FFGEN**  \L1_0/abs_reg[1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4606 ), .force_10(\L1_0/n4607 ), 
        .force_11(1'b0), .Q(n40866), .QN(n8447) );
  \**FFGEN**  \L1_0/abs_reg[1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4610 ), .force_10(\L1_0/n4611 ), 
        .force_11(1'b0), .Q(n40776), .QN(n8448) );
  \**FFGEN**  \L1_0/abs_reg[1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4614 ), .force_10(\L1_0/n4615 ), 
        .force_11(1'b0), .Q(n40867), .QN(n8449) );
  \**FFGEN**  \L1_0/abs_reg[1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4618 ), .force_10(\L1_0/n4619 ), 
        .force_11(1'b0), .Q(n40775), .QN(n8450) );
  \**FFGEN**  \L1_0/abs_reg[1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4622 ), .force_10(\L1_0/n4623 ), 
        .force_11(1'b0), .Q(n40868), .QN(n8451) );
  \**FFGEN**  \L1_0/abs_reg[1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4626 ), .force_10(\L1_0/n4627 ), 
        .force_11(1'b0), .Q(n40778), .QN(n8452) );
  \**FFGEN**  \L1_0/abs_reg[1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4630 ), .force_10(\L1_0/n4631 ), 
        .force_11(1'b0), .Q(n40860), .QN(n8453) );
  \**FFGEN**  \L1_0/abs_reg[1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4634 ), .force_10(\L1_0/n4635 ), 
        .force_11(1'b0), .Q(n40865), .QN(n8454) );
  \**FFGEN**  \L1_0/abs_reg[1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4638 ), .force_10(\L1_0/n4639 ), 
        .force_11(1'b0), .QN(n8455) );
  \**FFGEN**  \L1_0/abs_reg[1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4642 ), .force_10(\L1_0/n4643 ), 
        .force_11(1'b0), .QN(n8456) );
  \**FFGEN**  \L1_0/abs_reg[1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4646 ), .force_10(\L1_0/n4647 ), 
        .force_11(1'b0), .QN(n8457) );
  \**FFGEN**  \L1_0/abs_reg[1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4650 ), .force_10(\L1_0/n4651 ), 
        .force_11(1'b0), .QN(n8458) );
  \**FFGEN**  \L1_0/abs_reg[1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4654 ), .force_10(\L1_0/n4655 ), 
        .force_11(1'b0), .QN(n8459) );
  \**FFGEN**  \L1_0/abs_reg[1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4658 ), .force_10(\L1_0/n4659 ), 
        .force_11(1'b0), .QN(n8460) );
  \**FFGEN**  \L1_0/abs_reg[1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4662 ), .force_10(\L1_0/n4663 ), 
        .force_11(1'b0), .Q(n40836), .QN(n8461) );
  \**FFGEN**  \L1_0/abs_reg[1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4666 ), .force_10(\L1_0/n4667 ), 
        .force_11(1'b0), .QN(n8462) );
  \**FFGEN**  \L1_0/abs_reg[0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4670 ), .force_10(\L1_0/n4671 ), 
        .force_11(1'b0), .Q(n40807), .QN(n8463) );
  \**FFGEN**  \L1_0/abs_reg[0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4674 ), .force_10(\L1_0/n4675 ), 
        .force_11(1'b0), .Q(n40742), .QN(n8464) );
  \**FFGEN**  \L1_0/abs_reg[0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4678 ), .force_10(\L1_0/n4679 ), 
        .force_11(1'b0), .QN(n8465) );
  \**FFGEN**  \L1_0/abs_reg[0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4682 ), .force_10(\L1_0/n4683 ), 
        .force_11(1'b0), .Q(n40749), .QN(n8466) );
  \**FFGEN**  \L1_0/abs_reg[0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4686 ), .force_10(\L1_0/n4687 ), 
        .force_11(1'b0), .QN(n8467) );
  \**FFGEN**  \L1_0/abs_reg[0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4690 ), .force_10(\L1_0/n4691 ), 
        .force_11(1'b0), .Q(n40750), .QN(n8468) );
  \**FFGEN**  \L1_0/abs_reg[0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4694 ), .force_10(\L1_0/n4695 ), 
        .force_11(1'b0), .QN(n8469) );
  \**FFGEN**  \L1_0/abs_reg[0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4698 ), .force_10(\L1_0/n4699 ), 
        .force_11(1'b0), .Q(n40751), .QN(n8470) );
  \**FFGEN**  \L1_0/abs_reg[0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4702 ), .force_10(\L1_0/n4703 ), 
        .force_11(1'b0), .QN(n8471) );
  \**FFGEN**  \L1_0/abs_reg[0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4706 ), .force_10(\L1_0/n4707 ), 
        .force_11(1'b0), .Q(n40747), .QN(n8472) );
  \**FFGEN**  \L1_0/abs_reg[0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4710 ), .force_10(\L1_0/n4711 ), 
        .force_11(1'b0), .QN(n8473) );
  \**FFGEN**  \L1_0/abs_reg[0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4714 ), .force_10(\L1_0/n4715 ), 
        .force_11(1'b0), .Q(n40802), .QN(n8474) );
  \**FFGEN**  \L1_0/abs_reg[0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4718 ), .force_10(\L1_0/n4719 ), 
        .force_11(1'b0), .Q(n40798), .QN(n8475) );
  \**FFGEN**  \L1_0/abs_reg[0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4722 ), .force_10(\L1_0/n4723 ), 
        .force_11(1'b0), .Q(n40852), .QN(n8476) );
  \**FFGEN**  \L1_0/abs_reg[0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4726 ), .force_10(\L1_0/n4727 ), 
        .force_11(1'b0), .Q(n40796), .QN(n8477) );
  \**FFGEN**  \L1_0/abs_reg[0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4730 ), .force_10(\L1_0/n4731 ), 
        .force_11(1'b0), .Q(n40738), .QN(n8478) );
  \**FFGEN**  \L1_0/abs_reg[0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4734 ), .force_10(\L1_0/n4735 ), 
        .force_11(1'b0), .Q(n40722), .QN(n8479) );
  \**FFGEN**  \L1_0/abs_reg[0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4738 ), .force_10(\L1_0/n4739 ), 
        .force_11(1'b0), .Q(n40724), .QN(n8480) );
  \**FFGEN**  \L1_0/abs_reg[0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4742 ), .force_10(\L1_0/n4743 ), 
        .force_11(1'b0), .Q(n40752), .QN(n8481) );
  \**FFGEN**  \L1_0/abs_reg[0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4746 ), .force_10(\L1_0/n4747 ), 
        .force_11(1'b0), .QN(n8482) );
  \**FFGEN**  \L1_0/sum_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4750 ), .force_10(\L1_0/n4751 ), 
        .force_11(1'b0), .Q(out_L1[0]), .QN(n40725) );
  \**FFGEN**  \L1_0/sum_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4754 ), .force_10(\L1_0/n4755 ), 
        .force_11(1'b0), .Q(out_L1[1]), .QN(n40736) );
  \**FFGEN**  \L1_0/sum_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4758 ), .force_10(\L1_0/n4759 ), 
        .force_11(1'b0), .Q(out_L1[2]) );
  \**FFGEN**  \L1_0/sum_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4762 ), .force_10(\L1_0/n4763 ), 
        .force_11(1'b0), .Q(out_L1[3]), .QN(n40785) );
  \**FFGEN**  \L1_0/sum_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4766 ), .force_10(\L1_0/n4767 ), 
        .force_11(1'b0), .Q(out_L1[4]), .QN(n40786) );
  \**FFGEN**  \L1_0/sum_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4770 ), .force_10(\L1_0/n4771 ), 
        .force_11(1'b0), .Q(out_L1[5]), .QN(n40794) );
  \**FFGEN**  \L1_0/sum_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4774 ), .force_10(\L1_0/n4775 ), 
        .force_11(1'b0), .Q(out_L1[6]), .QN(n40808) );
  \**FFGEN**  \L1_0/sum_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4778 ), .force_10(\L1_0/n4779 ), 
        .force_11(1'b0), .Q(out_L1[7]), .QN(n40792) );
  \**FFGEN**  \L1_0/sum_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4782 ), .force_10(\L1_0/n4783 ), 
        .force_11(1'b0), .Q(out_L1[8]), .QN(n40801) );
  \**FFGEN**  \L1_0/sum_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4786 ), .force_10(\L1_0/n4787 ), 
        .force_11(1'b0), .Q(out_L1[9]), .QN(n40846) );
  \**FFGEN**  \L1_0/sum_reg[10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4790 ), .force_10(\L1_0/n4791 ), 
        .force_11(1'b0), .Q(out_L1[10]), .QN(n40731) );
  \**FFGEN**  \L1_0/sum_reg[11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4794 ), .force_10(\L1_0/n4795 ), 
        .force_11(1'b0), .Q(out_L1[11]), .QN(n40850) );
  \**FFGEN**  \L1_0/sum_reg[12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4798 ), .force_10(\L1_0/n4799 ), 
        .force_11(1'b0), .Q(out_L1[12]), .QN(n40735) );
  \**FFGEN**  \L1_0/sum_reg[13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4802 ), .force_10(\L1_0/n4803 ), 
        .force_11(1'b0), .Q(out_L1[13]), .QN(n40849) );
  \**FFGEN**  \L1_0/sum_reg[14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4806 ), .force_10(\L1_0/n4807 ), 
        .force_11(1'b0), .Q(out_L1[14]), .QN(n40734) );
  \**FFGEN**  \L1_0/sum_reg[15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4810 ), .force_10(\L1_0/n4811 ), 
        .force_11(1'b0), .Q(out_L1[15]), .QN(n40848) );
  \**FFGEN**  \L1_0/sum_reg[16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4814 ), .force_10(\L1_0/n4815 ), 
        .force_11(1'b0), .Q(out_L1[16]), .QN(n40733) );
  \**FFGEN**  \L1_0/sum_reg[17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4818 ), .force_10(\L1_0/n4819 ), 
        .force_11(1'b0), .Q(out_L1[17]), .QN(n40847) );
  \**FFGEN**  \L1_0/sum_reg[18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4822 ), .force_10(\L1_0/n4823 ), 
        .force_11(1'b0), .Q(out_L1[18]), .QN(n40741) );
  \**FFGEN**  \L1_0/sum_reg[19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3506 ), .force_10(\L1_0/n3507 ), 
        .force_11(1'b0), .Q(out_L1[19]), .QN(n40806) );
  \**FFGEN**  \L2_0/square_reg[14][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8021), .force_10(\L2_0/n2948 ), .force_11(
        1'b0), .QN(n8483) );
  \**FFGEN**  \L2_0/square_reg[14][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8026), .force_10(\L2_0/n2952 ), .force_11(
        1'b0), .QN(n8484) );
  \**FFGEN**  \L2_0/square_reg[14][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8013), .force_10(\L2_0/n2956 ), .force_11(
        1'b0), .QN(n8485) );
  \**FFGEN**  \L2_0/square_reg[14][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8008), .force_10(\L2_0/n2960 ), .force_11(
        1'b0), .QN(n8486) );
  \**FFGEN**  \L2_0/square_reg[14][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8016), .force_10(\L2_0/n2964 ), .force_11(
        1'b0), .QN(n8487) );
  \**FFGEN**  \L2_0/square_reg[14][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8018), .force_10(\L2_0/n2968 ), .force_11(
        1'b0), .QN(n8488) );
  \**FFGEN**  \L2_0/square_reg[14][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8014), .force_10(\L2_0/n2972 ), .force_11(
        1'b0), .QN(n8489) );
  \**FFGEN**  \L2_0/square_reg[14][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8015), .force_10(\L2_0/n2976 ), .force_11(
        1'b0), .QN(n8490) );
  \**FFGEN**  \L2_0/square_reg[14][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8012), .force_10(\L2_0/n2980 ), .force_11(
        1'b0), .QN(n8491) );
  \**FFGEN**  \L2_0/square_reg[14][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8010), .force_10(\L2_0/n2984 ), .force_11(
        1'b0), .QN(n8492) );
  \**FFGEN**  \L2_0/square_reg[14][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8023), .force_10(\L2_0/n2988 ), .force_11(
        1'b0), .QN(n8493) );
  \**FFGEN**  \L2_0/square_reg[14][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8017), .force_10(\L2_0/n2992 ), .force_11(
        1'b0), .QN(n8494) );
  \**FFGEN**  \L2_0/square_reg[14][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8009), .force_10(\L2_0/n2996 ), .force_11(
        1'b0), .QN(n8495) );
  \**FFGEN**  \L2_0/square_reg[14][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8022), .force_10(\L2_0/n3000 ), .force_11(
        1'b0), .QN(n8496) );
  \**FFGEN**  \L2_0/square_reg[14][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8011), .force_10(\L2_0/n3004 ), .force_11(
        1'b0), .QN(n8497) );
  \**FFGEN**  \L2_0/square_reg[14][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8020), .force_10(\L2_0/n3008 ), .force_11(
        1'b0), .QN(n8498) );
  \**FFGEN**  \L2_0/square_reg[14][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8025), .force_10(\L2_0/n3012 ), .force_11(
        1'b0), .QN(n8499) );
  \**FFGEN**  \L2_0/square_reg[14][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8019), .force_10(\L2_0/n3016 ), .force_11(
        1'b0), .QN(n8500) );
  \**FFGEN**  \L2_0/square_reg[14][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46263), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40839), .QN(n8501) );
  \**FFGEN**  \L2_0/square_reg[14][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8024), .force_10(\L2_0/n3024 ), .force_11(
        1'b0), .Q(n40789), .QN(n8502) );
  \**FFGEN**  \L2_0/square_reg[13][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7990), .force_10(\L2_0/n3028 ), .force_11(
        1'b0), .QN(n8503) );
  \**FFGEN**  \L2_0/square_reg[13][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7997), .force_10(\L2_0/n3032 ), .force_11(
        1'b0), .QN(n8504) );
  \**FFGEN**  \L2_0/square_reg[13][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8004), .force_10(\L2_0/n3036 ), .force_11(
        1'b0), .QN(n8505) );
  \**FFGEN**  \L2_0/square_reg[13][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8006), .force_10(\L2_0/n3040 ), .force_11(
        1'b0), .QN(n8506) );
  \**FFGEN**  \L2_0/square_reg[13][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7999), .force_10(\L2_0/n3044 ), .force_11(
        1'b0), .QN(n8507) );
  \**FFGEN**  \L2_0/square_reg[13][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7994), .force_10(\L2_0/n3048 ), .force_11(
        1'b0), .QN(n8508) );
  \**FFGEN**  \L2_0/square_reg[13][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8005), .force_10(\L2_0/n3052 ), .force_11(
        1'b0), .QN(n8509) );
  \**FFGEN**  \L2_0/square_reg[13][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7998), .force_10(\L2_0/n3056 ), .force_11(
        1'b0), .QN(n8510) );
  \**FFGEN**  \L2_0/square_reg[13][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8000), .force_10(\L2_0/n3060 ), .force_11(
        1'b0), .QN(n8511) );
  \**FFGEN**  \L2_0/square_reg[13][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7992), .force_10(\L2_0/n3064 ), .force_11(
        1'b0), .QN(n8512) );
  \**FFGEN**  \L2_0/square_reg[13][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8002), .force_10(\L2_0/n3068 ), .force_11(
        1'b0), .QN(n8513) );
  \**FFGEN**  \L2_0/square_reg[13][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8003), .force_10(\L2_0/n3072 ), .force_11(
        1'b0), .QN(n8514) );
  \**FFGEN**  \L2_0/square_reg[13][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7991), .force_10(\L2_0/n3076 ), .force_11(
        1'b0), .QN(n8515) );
  \**FFGEN**  \L2_0/square_reg[13][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8001), .force_10(\L2_0/n3080 ), .force_11(
        1'b0), .QN(n8516) );
  \**FFGEN**  \L2_0/square_reg[13][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8007), .force_10(\L2_0/n3084 ), .force_11(
        1'b0), .QN(n8517) );
  \**FFGEN**  \L2_0/square_reg[13][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7989), .force_10(\L2_0/n3088 ), .force_11(
        1'b0), .QN(n8518) );
  \**FFGEN**  \L2_0/square_reg[13][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7996), .force_10(\L2_0/n3092 ), .force_11(
        1'b0), .QN(n8519) );
  \**FFGEN**  \L2_0/square_reg[13][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7993), .force_10(\L2_0/n3096 ), .force_11(
        1'b0), .QN(n8520) );
  \**FFGEN**  \L2_0/square_reg[13][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46283), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40827), .QN(n8521) );
  \**FFGEN**  \L2_0/square_reg[13][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7995), .force_10(\L2_0/n3104 ), .force_11(
        1'b0), .QN(n8522) );
  \**FFGEN**  \L2_0/square_reg[12][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7980), .force_10(\L2_0/n3108 ), .force_11(
        1'b0), .QN(n8523) );
  \**FFGEN**  \L2_0/square_reg[12][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7987), .force_10(\L2_0/n3112 ), .force_11(
        1'b0), .QN(n8524) );
  \**FFGEN**  \L2_0/square_reg[12][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7984), .force_10(\L2_0/n3116 ), .force_11(
        1'b0), .QN(n8525) );
  \**FFGEN**  \L2_0/square_reg[12][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7976), .force_10(\L2_0/n3120 ), .force_11(
        1'b0), .QN(n8526) );
  \**FFGEN**  \L2_0/square_reg[12][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7969), .force_10(\L2_0/n3124 ), .force_11(
        1'b0), .QN(n8527) );
  \**FFGEN**  \L2_0/square_reg[12][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7974), .force_10(\L2_0/n3128 ), .force_11(
        1'b0), .QN(n8528) );
  \**FFGEN**  \L2_0/square_reg[12][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7975), .force_10(\L2_0/n3132 ), .force_11(
        1'b0), .QN(n8529) );
  \**FFGEN**  \L2_0/square_reg[12][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7968), .force_10(\L2_0/n3136 ), .force_11(
        1'b0), .QN(n8530) );
  \**FFGEN**  \L2_0/square_reg[12][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7977), .force_10(\L2_0/n3140 ), .force_11(
        1'b0), .QN(n8531) );
  \**FFGEN**  \L2_0/square_reg[12][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7982), .force_10(\L2_0/n3144 ), .force_11(
        1'b0), .QN(n8532) );
  \**FFGEN**  \L2_0/square_reg[12][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7972), .force_10(\L2_0/n3148 ), .force_11(
        1'b0), .QN(n8533) );
  \**FFGEN**  \L2_0/square_reg[12][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7983), .force_10(\L2_0/n3152 ), .force_11(
        1'b0), .QN(n8534) );
  \**FFGEN**  \L2_0/square_reg[12][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7981), .force_10(\L2_0/n3156 ), .force_11(
        1'b0), .QN(n8535) );
  \**FFGEN**  \L2_0/square_reg[12][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7971), .force_10(\L2_0/n3160 ), .force_11(
        1'b0), .QN(n8536) );
  \**FFGEN**  \L2_0/square_reg[12][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7970), .force_10(\L2_0/n3164 ), .force_11(
        1'b0), .QN(n8537) );
  \**FFGEN**  \L2_0/square_reg[12][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7979), .force_10(\L2_0/n3168 ), .force_11(
        1'b0), .QN(n8538) );
  \**FFGEN**  \L2_0/square_reg[12][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7986), .force_10(\L2_0/n3172 ), .force_11(
        1'b0), .QN(n8539) );
  \**FFGEN**  \L2_0/square_reg[12][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7973), .force_10(\L2_0/n3176 ), .force_11(
        1'b0), .QN(n8540) );
  \**FFGEN**  \L2_0/square_reg[12][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46308), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40825), .QN(n8541) );
  \**FFGEN**  \L2_0/square_reg[12][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7985), .force_10(\L2_0/n3184 ), .force_11(
        1'b0), .QN(n8542) );
  \**FFGEN**  \L2_0/square_reg[11][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7950), .force_10(\L2_0/n3188 ), .force_11(
        1'b0), .QN(n8543) );
  \**FFGEN**  \L2_0/square_reg[11][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7957), .force_10(\L2_0/n3192 ), .force_11(
        1'b0), .QN(n8544) );
  \**FFGEN**  \L2_0/square_reg[11][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7964), .force_10(\L2_0/n3196 ), .force_11(
        1'b0), .QN(n8545) );
  \**FFGEN**  \L2_0/square_reg[11][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7966), .force_10(\L2_0/n3200 ), .force_11(
        1'b0), .QN(n8546) );
  \**FFGEN**  \L2_0/square_reg[11][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7959), .force_10(\L2_0/n3204 ), .force_11(
        1'b0), .QN(n8547) );
  \**FFGEN**  \L2_0/square_reg[11][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7954), .force_10(\L2_0/n3208 ), .force_11(
        1'b0), .QN(n8548) );
  \**FFGEN**  \L2_0/square_reg[11][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7965), .force_10(\L2_0/n3212 ), .force_11(
        1'b0), .QN(n8549) );
  \**FFGEN**  \L2_0/square_reg[11][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7958), .force_10(\L2_0/n3216 ), .force_11(
        1'b0), .QN(n8550) );
  \**FFGEN**  \L2_0/square_reg[11][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7960), .force_10(\L2_0/n3220 ), .force_11(
        1'b0), .QN(n8551) );
  \**FFGEN**  \L2_0/square_reg[11][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7952), .force_10(\L2_0/n3224 ), .force_11(
        1'b0), .QN(n8552) );
  \**FFGEN**  \L2_0/square_reg[11][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7962), .force_10(\L2_0/n3228 ), .force_11(
        1'b0), .QN(n8553) );
  \**FFGEN**  \L2_0/square_reg[11][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7963), .force_10(\L2_0/n3232 ), .force_11(
        1'b0), .QN(n8554) );
  \**FFGEN**  \L2_0/square_reg[11][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7951), .force_10(\L2_0/n3236 ), .force_11(
        1'b0), .QN(n8555) );
  \**FFGEN**  \L2_0/square_reg[11][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7961), .force_10(\L2_0/n3240 ), .force_11(
        1'b0), .QN(n8556) );
  \**FFGEN**  \L2_0/square_reg[11][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7967), .force_10(\L2_0/n3244 ), .force_11(
        1'b0), .QN(n8557) );
  \**FFGEN**  \L2_0/square_reg[11][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7949), .force_10(\L2_0/n3248 ), .force_11(
        1'b0), .QN(n8558) );
  \**FFGEN**  \L2_0/square_reg[11][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7956), .force_10(\L2_0/n3252 ), .force_11(
        1'b0), .QN(n8559) );
  \**FFGEN**  \L2_0/square_reg[11][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7953), .force_10(\L2_0/n3256 ), .force_11(
        1'b0), .QN(n8560) );
  \**FFGEN**  \L2_0/square_reg[11][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46327), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40821), .QN(n8561) );
  \**FFGEN**  \L2_0/square_reg[11][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7955), .force_10(\L2_0/n3264 ), .force_11(
        1'b0), .QN(n8562) );
  \**FFGEN**  \L2_0/square_reg[10][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8027), .force_10(\L2_0/n3268 ), .force_11(
        1'b0), .QN(n8563) );
  \**FFGEN**  \L2_0/square_reg[10][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8045), .force_10(\L2_0/n3272 ), .force_11(
        1'b0), .QN(n8564) );
  \**FFGEN**  \L2_0/square_reg[10][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8030), .force_10(\L2_0/n3276 ), .force_11(
        1'b0), .QN(n8565) );
  \**FFGEN**  \L2_0/square_reg[10][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8042), .force_10(\L2_0/n3280 ), .force_11(
        1'b0), .QN(n8566) );
  \**FFGEN**  \L2_0/square_reg[10][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8039), .force_10(\L2_0/n3284 ), .force_11(
        1'b0), .QN(n8567) );
  \**FFGEN**  \L2_0/square_reg[10][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8031), .force_10(\L2_0/n3288 ), .force_11(
        1'b0), .QN(n8568) );
  \**FFGEN**  \L2_0/square_reg[10][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8035), .force_10(\L2_0/n3292 ), .force_11(
        1'b0), .QN(n8569) );
  \**FFGEN**  \L2_0/square_reg[10][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8038), .force_10(\L2_0/n3296 ), .force_11(
        1'b0), .QN(n8570) );
  \**FFGEN**  \L2_0/square_reg[10][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8033), .force_10(\L2_0/n3300 ), .force_11(
        1'b0), .QN(n8571) );
  \**FFGEN**  \L2_0/square_reg[10][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8046), .force_10(\L2_0/n3304 ), .force_11(
        1'b0), .QN(n8572) );
  \**FFGEN**  \L2_0/square_reg[10][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8041), .force_10(\L2_0/n3308 ), .force_11(
        1'b0), .QN(n8573) );
  \**FFGEN**  \L2_0/square_reg[10][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8037), .force_10(\L2_0/n3312 ), .force_11(
        1'b0), .QN(n8574) );
  \**FFGEN**  \L2_0/square_reg[10][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8028), .force_10(\L2_0/n3316 ), .force_11(
        1'b0), .QN(n8575) );
  \**FFGEN**  \L2_0/square_reg[10][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8040), .force_10(\L2_0/n3320 ), .force_11(
        1'b0), .QN(n8576) );
  \**FFGEN**  \L2_0/square_reg[10][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8029), .force_10(\L2_0/n3324 ), .force_11(
        1'b0), .QN(n8577) );
  \**FFGEN**  \L2_0/square_reg[10][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8036), .force_10(\L2_0/n3328 ), .force_11(
        1'b0), .QN(n8578) );
  \**FFGEN**  \L2_0/square_reg[10][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8044), .force_10(\L2_0/n3332 ), .force_11(
        1'b0), .QN(n8579) );
  \**FFGEN**  \L2_0/square_reg[10][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8032), .force_10(\L2_0/n3336 ), .force_11(
        1'b0), .QN(n8580) );
  \**FFGEN**  \L2_0/square_reg[10][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46355), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40818), .QN(n8581) );
  \**FFGEN**  \L2_0/square_reg[10][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8043), .force_10(\L2_0/n3344 ), .force_11(
        1'b0), .QN(n8582) );
  \**FFGEN**  \L2_0/square_reg[9][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7931), .force_10(\L2_0/n3348 ), .force_11(
        1'b0), .QN(n8583) );
  \**FFGEN**  \L2_0/square_reg[9][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7938), .force_10(\L2_0/n3352 ), .force_11(
        1'b0), .QN(n8584) );
  \**FFGEN**  \L2_0/square_reg[9][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7945), .force_10(\L2_0/n3356 ), .force_11(
        1'b0), .QN(n8585) );
  \**FFGEN**  \L2_0/square_reg[9][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7947), .force_10(\L2_0/n3360 ), .force_11(
        1'b0), .QN(n8586) );
  \**FFGEN**  \L2_0/square_reg[9][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7940), .force_10(\L2_0/n3364 ), .force_11(
        1'b0), .QN(n8587) );
  \**FFGEN**  \L2_0/square_reg[9][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7935), .force_10(\L2_0/n3368 ), .force_11(
        1'b0), .QN(n8588) );
  \**FFGEN**  \L2_0/square_reg[9][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7946), .force_10(\L2_0/n3372 ), .force_11(
        1'b0), .QN(n8589) );
  \**FFGEN**  \L2_0/square_reg[9][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7939), .force_10(\L2_0/n3376 ), .force_11(
        1'b0), .QN(n8590) );
  \**FFGEN**  \L2_0/square_reg[9][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7941), .force_10(\L2_0/n3380 ), .force_11(
        1'b0), .QN(n8591) );
  \**FFGEN**  \L2_0/square_reg[9][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7933), .force_10(\L2_0/n3384 ), .force_11(
        1'b0), .QN(n8592) );
  \**FFGEN**  \L2_0/square_reg[9][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7943), .force_10(\L2_0/n3388 ), .force_11(
        1'b0), .QN(n8593) );
  \**FFGEN**  \L2_0/square_reg[9][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7944), .force_10(\L2_0/n3392 ), .force_11(
        1'b0), .QN(n8594) );
  \**FFGEN**  \L2_0/square_reg[9][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7932), .force_10(\L2_0/n3396 ), .force_11(
        1'b0), .QN(n8595) );
  \**FFGEN**  \L2_0/square_reg[9][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7942), .force_10(\L2_0/n3400 ), .force_11(
        1'b0), .QN(n8596) );
  \**FFGEN**  \L2_0/square_reg[9][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7948), .force_10(\L2_0/n3404 ), .force_11(
        1'b0), .QN(n8597) );
  \**FFGEN**  \L2_0/square_reg[9][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7930), .force_10(\L2_0/n3408 ), .force_11(
        1'b0), .QN(n8598) );
  \**FFGEN**  \L2_0/square_reg[9][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7937), .force_10(\L2_0/n3412 ), .force_11(
        1'b0), .QN(n8599) );
  \**FFGEN**  \L2_0/square_reg[9][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7934), .force_10(\L2_0/n3416 ), .force_11(
        1'b0), .QN(n8600) );
  \**FFGEN**  \L2_0/square_reg[9][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46375), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40817), .QN(n8601) );
  \**FFGEN**  \L2_0/square_reg[9][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7936), .force_10(\L2_0/n3424 ), .force_11(
        1'b0), .QN(n8602) );
  \**FFGEN**  \L2_0/square_reg[8][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7911), .force_10(\L2_0/n3428 ), .force_11(
        1'b0), .QN(n8603) );
  \**FFGEN**  \L2_0/square_reg[8][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7919), .force_10(\L2_0/n3432 ), .force_11(
        1'b0), .QN(n8604) );
  \**FFGEN**  \L2_0/square_reg[8][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7926), .force_10(\L2_0/n3436 ), .force_11(
        1'b0), .QN(n8605) );
  \**FFGEN**  \L2_0/square_reg[8][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7928), .force_10(\L2_0/n3440 ), .force_11(
        1'b0), .QN(n8606) );
  \**FFGEN**  \L2_0/square_reg[8][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7921), .force_10(\L2_0/n3444 ), .force_11(
        1'b0), .QN(n8607) );
  \**FFGEN**  \L2_0/square_reg[8][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7916), .force_10(\L2_0/n3448 ), .force_11(
        1'b0), .QN(n8608) );
  \**FFGEN**  \L2_0/square_reg[8][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7927), .force_10(\L2_0/n3452 ), .force_11(
        1'b0), .QN(n8609) );
  \**FFGEN**  \L2_0/square_reg[8][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7920), .force_10(\L2_0/n3456 ), .force_11(
        1'b0), .QN(n8610) );
  \**FFGEN**  \L2_0/square_reg[8][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7922), .force_10(\L2_0/n3460 ), .force_11(
        1'b0), .QN(n8611) );
  \**FFGEN**  \L2_0/square_reg[8][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7914), .force_10(\L2_0/n3464 ), .force_11(
        1'b0), .QN(n8612) );
  \**FFGEN**  \L2_0/square_reg[8][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7924), .force_10(\L2_0/n3468 ), .force_11(
        1'b0), .QN(n8613) );
  \**FFGEN**  \L2_0/square_reg[8][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7925), .force_10(\L2_0/n3472 ), .force_11(
        1'b0), .QN(n8614) );
  \**FFGEN**  \L2_0/square_reg[8][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7913), .force_10(\L2_0/n3476 ), .force_11(
        1'b0), .QN(n8615) );
  \**FFGEN**  \L2_0/square_reg[8][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7923), .force_10(\L2_0/n3480 ), .force_11(
        1'b0), .QN(n8616) );
  \**FFGEN**  \L2_0/square_reg[8][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7929), .force_10(\L2_0/n3484 ), .force_11(
        1'b0), .QN(n8617) );
  \**FFGEN**  \L2_0/square_reg[8][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7912), .force_10(\L2_0/n3488 ), .force_11(
        1'b0), .QN(n8618) );
  \**FFGEN**  \L2_0/square_reg[8][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7918), .force_10(\L2_0/n3492 ), .force_11(
        1'b0), .QN(n8619) );
  \**FFGEN**  \L2_0/square_reg[8][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7915), .force_10(\L2_0/n3496 ), .force_11(
        1'b0), .QN(n8620) );
  \**FFGEN**  \L2_0/square_reg[8][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46398), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40815), .QN(n8621) );
  \**FFGEN**  \L2_0/square_reg[8][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7917), .force_10(\L2_0/n3504 ), .force_11(
        1'b0), .QN(n8622) );
  \**FFGEN**  \L2_0/square_reg[7][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7907), .force_10(\L2_0/n3508 ), .force_11(
        1'b0), .QN(n8623) );
  \**FFGEN**  \L2_0/square_reg[7][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7901), .force_10(\L2_0/n3512 ), .force_11(
        1'b0), .QN(n8624) );
  \**FFGEN**  \L2_0/square_reg[7][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7894), .force_10(\L2_0/n3516 ), .force_11(
        1'b0), .QN(n8625) );
  \**FFGEN**  \L2_0/square_reg[7][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7910), .force_10(\L2_0/n3520 ), .force_11(
        1'b0), .QN(n8626) );
  \**FFGEN**  \L2_0/square_reg[7][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7905), .force_10(\L2_0/n3524 ), .force_11(
        1'b0), .QN(n8627) );
  \**FFGEN**  \L2_0/square_reg[7][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7896), .force_10(\L2_0/n3528 ), .force_11(
        1'b0), .QN(n8628) );
  \**FFGEN**  \L2_0/square_reg[7][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7904), .force_10(\L2_0/n3532 ), .force_11(
        1'b0), .QN(n8629) );
  \**FFGEN**  \L2_0/square_reg[7][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7898), .force_10(\L2_0/n3536 ), .force_11(
        1'b0), .QN(n8630) );
  \**FFGEN**  \L2_0/square_reg[7][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7893), .force_10(\L2_0/n3540 ), .force_11(
        1'b0), .QN(n8631) );
  \**FFGEN**  \L2_0/square_reg[7][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7909), .force_10(\L2_0/n3544 ), .force_11(
        1'b0), .QN(n8632) );
  \**FFGEN**  \L2_0/square_reg[7][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7903), .force_10(\L2_0/n3548 ), .force_11(
        1'b0), .QN(n8633) );
  \**FFGEN**  \L2_0/square_reg[7][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7895), .force_10(\L2_0/n3552 ), .force_11(
        1'b0), .QN(n8634) );
  \**FFGEN**  \L2_0/square_reg[7][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7908), .force_10(\L2_0/n3556 ), .force_11(
        1'b0), .QN(n8635) );
  \**FFGEN**  \L2_0/square_reg[7][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7902), .force_10(\L2_0/n3560 ), .force_11(
        1'b0), .QN(n8636) );
  \**FFGEN**  \L2_0/square_reg[7][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7892), .force_10(\L2_0/n3564 ), .force_11(
        1'b0), .QN(n8637) );
  \**FFGEN**  \L2_0/square_reg[7][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7906), .force_10(\L2_0/n3568 ), .force_11(
        1'b0), .QN(n8638) );
  \**FFGEN**  \L2_0/square_reg[7][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7900), .force_10(\L2_0/n3572 ), .force_11(
        1'b0), .QN(n8639) );
  \**FFGEN**  \L2_0/square_reg[7][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7897), .force_10(\L2_0/n3576 ), .force_11(
        1'b0), .QN(n8640) );
  \**FFGEN**  \L2_0/square_reg[7][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46419), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40813), .QN(n8641) );
  \**FFGEN**  \L2_0/square_reg[7][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n7899), .force_10(\L2_0/n3584 ), .force_11(
        1'b0), .QN(n8642) );
  \**FFGEN**  \L2_0/square_reg[6][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8075), .force_10(\L2_0/n3588 ), .force_11(
        1'b0), .QN(n8643) );
  \**FFGEN**  \L2_0/square_reg[6][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8078), .force_10(\L2_0/n3592 ), .force_11(
        1'b0), .Q(n40773), .QN(n8644) );
  \**FFGEN**  \L2_0/square_reg[6][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8090), .force_10(\L2_0/n3596 ), .force_11(
        1'b0), .Q(n40764), .QN(n8645) );
  \**FFGEN**  \L2_0/square_reg[6][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8092), .force_10(\L2_0/n3600 ), .force_11(
        1'b0), .Q(n40812), .QN(n8646) );
  \**FFGEN**  \L2_0/square_reg[6][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8085), .force_10(\L2_0/n3604 ), .force_11(
        1'b0), .Q(n40763), .QN(n8647) );
  \**FFGEN**  \L2_0/square_reg[6][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8077), .force_10(\L2_0/n3608 ), .force_11(
        1'b0), .Q(n40810), .QN(n8648) );
  \**FFGEN**  \L2_0/square_reg[6][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8091), .force_10(\L2_0/n3612 ), .force_11(
        1'b0), .Q(n40754), .QN(n8649) );
  \**FFGEN**  \L2_0/square_reg[6][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8084), .force_10(\L2_0/n3616 ), .force_11(
        1'b0), .Q(n40756), .QN(n8650) );
  \**FFGEN**  \L2_0/square_reg[6][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8086), .force_10(\L2_0/n3620 ), .force_11(
        1'b0), .Q(n40770), .QN(n8651) );
  \**FFGEN**  \L2_0/square_reg[6][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8082), .force_10(\L2_0/n3624 ), .force_11(
        1'b0), .Q(n40760), .QN(n8652) );
  \**FFGEN**  \L2_0/square_reg[6][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8088), .force_10(\L2_0/n3628 ), .force_11(
        1'b0), .Q(n40853), .QN(n8653) );
  \**FFGEN**  \L2_0/square_reg[6][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8089), .force_10(\L2_0/n3632 ), .force_11(
        1'b0), .Q(n40769), .QN(n8654) );
  \**FFGEN**  \L2_0/square_reg[6][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8079), .force_10(\L2_0/n3636 ), .force_11(
        1'b0), .Q(n40759), .QN(n8655) );
  \**FFGEN**  \L2_0/square_reg[6][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8087), .force_10(\L2_0/n3640 ), .force_11(
        1'b0), .Q(n40856), .QN(n8656) );
  \**FFGEN**  \L2_0/square_reg[6][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8093), .force_10(\L2_0/n3644 ), .force_11(
        1'b0), .Q(n40768), .QN(n8657) );
  \**FFGEN**  \L2_0/square_reg[6][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8080), .force_10(\L2_0/n3648 ), .force_11(
        1'b0), .Q(n40858), .QN(n8658) );
  \**FFGEN**  \L2_0/square_reg[6][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8083), .force_10(\L2_0/n3652 ), .force_11(
        1'b0), .Q(n40784), .QN(n8659) );
  \**FFGEN**  \L2_0/square_reg[6][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8076), .force_10(\L2_0/n3656 ), .force_11(
        1'b0), .QN(n8660) );
  \**FFGEN**  \L2_0/square_reg[6][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46442), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40838), .QN(n8661) );
  \**FFGEN**  \L2_0/square_reg[6][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8081), .force_10(\L2_0/n3664 ), .force_11(
        1'b0), .QN(n8662) );
  \**FFGEN**  \L2_0/square_reg[5][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8068), .force_10(\L2_0/n3668 ), .force_11(
        1'b0), .QN(n8663) );
  \**FFGEN**  \L2_0/square_reg[5][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8072), .force_10(\L2_0/n3672 ), .force_11(
        1'b0), .QN(n8664) );
  \**FFGEN**  \L2_0/square_reg[5][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8101), .force_10(\L2_0/n3676 ), .force_11(
        1'b0), .QN(n8665) );
  \**FFGEN**  \L2_0/square_reg[5][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8103), .force_10(\L2_0/n3680 ), .force_11(
        1'b0), .QN(n8666) );
  \**FFGEN**  \L2_0/square_reg[5][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8097), .force_10(\L2_0/n3684 ), .force_11(
        1'b0), .QN(n8667) );
  \**FFGEN**  \L2_0/square_reg[5][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8073), .force_10(\L2_0/n3688 ), .force_11(
        1'b0), .QN(n8668) );
  \**FFGEN**  \L2_0/square_reg[5][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8102), .force_10(\L2_0/n3692 ), .force_11(
        1'b0), .QN(n8669) );
  \**FFGEN**  \L2_0/square_reg[5][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8096), .force_10(\L2_0/n3696 ), .force_11(
        1'b0), .QN(n8670) );
  \**FFGEN**  \L2_0/square_reg[5][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8098), .force_10(\L2_0/n3700 ), .force_11(
        1'b0), .QN(n8671) );
  \**FFGEN**  \L2_0/square_reg[5][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8095), .force_10(\L2_0/n3704 ), .force_11(
        1'b0), .QN(n8672) );
  \**FFGEN**  \L2_0/square_reg[5][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8100), .force_10(\L2_0/n3708 ), .force_11(
        1'b0), .QN(n8673) );
  \**FFGEN**  \L2_0/square_reg[5][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8105), .force_10(\L2_0/n3712 ), .force_11(
        1'b0), .QN(n8674) );
  \**FFGEN**  \L2_0/square_reg[5][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8094), .force_10(\L2_0/n3716 ), .force_11(
        1'b0), .QN(n8675) );
  \**FFGEN**  \L2_0/square_reg[5][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8099), .force_10(\L2_0/n3720 ), .force_11(
        1'b0), .QN(n8676) );
  \**FFGEN**  \L2_0/square_reg[5][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8104), .force_10(\L2_0/n3724 ), .force_11(
        1'b0), .QN(n8677) );
  \**FFGEN**  \L2_0/square_reg[5][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8067), .force_10(\L2_0/n3728 ), .force_11(
        1'b0), .QN(n8678) );
  \**FFGEN**  \L2_0/square_reg[5][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8071), .force_10(\L2_0/n3732 ), .force_11(
        1'b0), .QN(n8679) );
  \**FFGEN**  \L2_0/square_reg[5][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8069), .force_10(\L2_0/n3736 ), .force_11(
        1'b0), .QN(n8680) );
  \**FFGEN**  \L2_0/square_reg[5][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46465), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40831), .QN(n8681) );
  \**FFGEN**  \L2_0/square_reg[5][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8070), .force_10(\L2_0/n3744 ), .force_11(
        1'b0), .QN(n8682) );
  \**FFGEN**  \L2_0/square_reg[4][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8164), .force_10(\L2_0/n3748 ), .force_11(
        1'b0), .QN(n8683) );
  \**FFGEN**  \L2_0/square_reg[4][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8175), .force_10(\L2_0/n3752 ), .force_11(
        1'b0), .QN(n8684) );
  \**FFGEN**  \L2_0/square_reg[4][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8168), .force_10(\L2_0/n3756 ), .force_11(
        1'b0), .QN(n8685) );
  \**FFGEN**  \L2_0/square_reg[4][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8179), .force_10(\L2_0/n3760 ), .force_11(
        1'b0), .QN(n8686) );
  \**FFGEN**  \L2_0/square_reg[4][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8177), .force_10(\L2_0/n3764 ), .force_11(
        1'b0), .QN(n8687) );
  \**FFGEN**  \L2_0/square_reg[4][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8169), .force_10(\L2_0/n3768 ), .force_11(
        1'b0), .QN(n8688) );
  \**FFGEN**  \L2_0/square_reg[4][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8171), .force_10(\L2_0/n3772 ), .force_11(
        1'b0), .QN(n8689) );
  \**FFGEN**  \L2_0/square_reg[4][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8176), .force_10(\L2_0/n3776 ), .force_11(
        1'b0), .QN(n8690) );
  \**FFGEN**  \L2_0/square_reg[4][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8173), .force_10(\L2_0/n3780 ), .force_11(
        1'b0), .QN(n8691) );
  \**FFGEN**  \L2_0/square_reg[4][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8166), .force_10(\L2_0/n3784 ), .force_11(
        1'b0), .QN(n8692) );
  \**FFGEN**  \L2_0/square_reg[4][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8181), .force_10(\L2_0/n3788 ), .force_11(
        1'b0), .QN(n8693) );
  \**FFGEN**  \L2_0/square_reg[4][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8174), .force_10(\L2_0/n3792 ), .force_11(
        1'b0), .QN(n8694) );
  \**FFGEN**  \L2_0/square_reg[4][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8165), .force_10(\L2_0/n3796 ), .force_11(
        1'b0), .QN(n8695) );
  \**FFGEN**  \L2_0/square_reg[4][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8180), .force_10(\L2_0/n3800 ), .force_11(
        1'b0), .QN(n8696) );
  \**FFGEN**  \L2_0/square_reg[4][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8167), .force_10(\L2_0/n3804 ), .force_11(
        1'b0), .QN(n8697) );
  \**FFGEN**  \L2_0/square_reg[4][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8172), .force_10(\L2_0/n3808 ), .force_11(
        1'b0), .QN(n8698) );
  \**FFGEN**  \L2_0/square_reg[4][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8178), .force_10(\L2_0/n3812 ), .force_11(
        1'b0), .QN(n8699) );
  \**FFGEN**  \L2_0/square_reg[4][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8170), .force_10(\L2_0/n3816 ), .force_11(
        1'b0), .QN(n8700) );
  \**FFGEN**  \L2_0/square_reg[4][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46487), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40828), .QN(n8701) );
  \**FFGEN**  \L2_0/square_reg[4][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8182), .force_10(\L2_0/n3824 ), .force_11(
        1'b0), .QN(n8702) );
  \**FFGEN**  \L2_0/square_reg[3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8145), .force_10(\L2_0/n3828 ), .force_11(
        1'b0), .QN(n8703) );
  \**FFGEN**  \L2_0/square_reg[3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8151), .force_10(\L2_0/n3832 ), .force_11(
        1'b0), .QN(n8704) );
  \**FFGEN**  \L2_0/square_reg[3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8160), .force_10(\L2_0/n3836 ), .force_11(
        1'b0), .QN(n8705) );
  \**FFGEN**  \L2_0/square_reg[3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8162), .force_10(\L2_0/n3840 ), .force_11(
        1'b0), .QN(n8706) );
  \**FFGEN**  \L2_0/square_reg[3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8155), .force_10(\L2_0/n3844 ), .force_11(
        1'b0), .QN(n8707) );
  \**FFGEN**  \L2_0/square_reg[3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8149), .force_10(\L2_0/n3848 ), .force_11(
        1'b0), .QN(n8708) );
  \**FFGEN**  \L2_0/square_reg[3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8161), .force_10(\L2_0/n3852 ), .force_11(
        1'b0), .QN(n8709) );
  \**FFGEN**  \L2_0/square_reg[3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8154), .force_10(\L2_0/n3856 ), .force_11(
        1'b0), .QN(n8710) );
  \**FFGEN**  \L2_0/square_reg[3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8156), .force_10(\L2_0/n3860 ), .force_11(
        1'b0), .QN(n8711) );
  \**FFGEN**  \L2_0/square_reg[3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8147), .force_10(\L2_0/n3864 ), .force_11(
        1'b0), .QN(n8712) );
  \**FFGEN**  \L2_0/square_reg[3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8158), .force_10(\L2_0/n3868 ), .force_11(
        1'b0), .QN(n8713) );
  \**FFGEN**  \L2_0/square_reg[3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8159), .force_10(\L2_0/n3872 ), .force_11(
        1'b0), .QN(n8714) );
  \**FFGEN**  \L2_0/square_reg[3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8146), .force_10(\L2_0/n3876 ), .force_11(
        1'b0), .QN(n8715) );
  \**FFGEN**  \L2_0/square_reg[3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8157), .force_10(\L2_0/n3880 ), .force_11(
        1'b0), .QN(n8716) );
  \**FFGEN**  \L2_0/square_reg[3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8163), .force_10(\L2_0/n3884 ), .force_11(
        1'b0), .QN(n8717) );
  \**FFGEN**  \L2_0/square_reg[3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8152), .force_10(\L2_0/n3888 ), .force_11(
        1'b0), .QN(n8718) );
  \**FFGEN**  \L2_0/square_reg[3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8153), .force_10(\L2_0/n3892 ), .force_11(
        1'b0), .QN(n8719) );
  \**FFGEN**  \L2_0/square_reg[3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8148), .force_10(\L2_0/n3896 ), .force_11(
        1'b0), .QN(n8720) );
  \**FFGEN**  \L2_0/square_reg[3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46510), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40835), .QN(n8721) );
  \**FFGEN**  \L2_0/square_reg[3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8150), .force_10(\L2_0/n3904 ), .force_11(
        1'b0), .QN(n8722) );
  \**FFGEN**  \L2_0/square_reg[2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8110), .force_10(\L2_0/n3908 ), .force_11(
        1'b0), .QN(n8723) );
  \**FFGEN**  \L2_0/square_reg[2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8125), .force_10(\L2_0/n3912 ), .force_11(
        1'b0), .QN(n8724) );
  \**FFGEN**  \L2_0/square_reg[2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8119), .force_10(\L2_0/n3916 ), .force_11(
        1'b0), .QN(n8725) );
  \**FFGEN**  \L2_0/square_reg[2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8111), .force_10(\L2_0/n3920 ), .force_11(
        1'b0), .QN(n8726) );
  \**FFGEN**  \L2_0/square_reg[2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8106), .force_10(\L2_0/n3924 ), .force_11(
        1'b0), .QN(n8727) );
  \**FFGEN**  \L2_0/square_reg[2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8114), .force_10(\L2_0/n3928 ), .force_11(
        1'b0), .QN(n8728) );
  \**FFGEN**  \L2_0/square_reg[2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8122), .force_10(\L2_0/n3932 ), .force_11(
        1'b0), .QN(n8729) );
  \**FFGEN**  \L2_0/square_reg[2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8116), .force_10(\L2_0/n3936 ), .force_11(
        1'b0), .QN(n8730) );
  \**FFGEN**  \L2_0/square_reg[2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8118), .force_10(\L2_0/n3940 ), .force_11(
        1'b0), .QN(n8731) );
  \**FFGEN**  \L2_0/square_reg[2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8112), .force_10(\L2_0/n3944 ), .force_11(
        1'b0), .QN(n8732) );
  \**FFGEN**  \L2_0/square_reg[2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8121), .force_10(\L2_0/n3948 ), .force_11(
        1'b0), .QN(n8733) );
  \**FFGEN**  \L2_0/square_reg[2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8113), .force_10(\L2_0/n3952 ), .force_11(
        1'b0), .QN(n8734) );
  \**FFGEN**  \L2_0/square_reg[2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8107), .force_10(\L2_0/n3956 ), .force_11(
        1'b0), .QN(n8735) );
  \**FFGEN**  \L2_0/square_reg[2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8120), .force_10(\L2_0/n3960 ), .force_11(
        1'b0), .QN(n8736) );
  \**FFGEN**  \L2_0/square_reg[2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8117), .force_10(\L2_0/n3964 ), .force_11(
        1'b0), .QN(n8737) );
  \**FFGEN**  \L2_0/square_reg[2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8109), .force_10(\L2_0/n3968 ), .force_11(
        1'b0), .QN(n8738) );
  \**FFGEN**  \L2_0/square_reg[2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8124), .force_10(\L2_0/n3972 ), .force_11(
        1'b0), .QN(n8739) );
  \**FFGEN**  \L2_0/square_reg[2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8115), .force_10(\L2_0/n3976 ), .force_11(
        1'b0), .QN(n8740) );
  \**FFGEN**  \L2_0/square_reg[2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46531), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40822), .QN(n8741) );
  \**FFGEN**  \L2_0/square_reg[2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8123), .force_10(\L2_0/n3984 ), .force_11(
        1'b0), .QN(n8742) );
  \**FFGEN**  \L2_0/square_reg[1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8127), .force_10(\L2_0/n3988 ), .force_11(
        1'b0), .QN(n8743) );
  \**FFGEN**  \L2_0/square_reg[1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8134), .force_10(\L2_0/n3992 ), .force_11(
        1'b0), .QN(n8744) );
  \**FFGEN**  \L2_0/square_reg[1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8141), .force_10(\L2_0/n3996 ), .force_11(
        1'b0), .Q(n40771), .QN(n8745) );
  \**FFGEN**  \L2_0/square_reg[1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8143), .force_10(\L2_0/n4000 ), .force_11(
        1'b0), .Q(n40779), .QN(n8746) );
  \**FFGEN**  \L2_0/square_reg[1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8136), .force_10(\L2_0/n4004 ), .force_11(
        1'b0), .Q(n40861), .QN(n8747) );
  \**FFGEN**  \L2_0/square_reg[1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8133), .force_10(\L2_0/n4008 ), .force_11(
        1'b0), .Q(n40782), .QN(n8748) );
  \**FFGEN**  \L2_0/square_reg[1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8142), .force_10(\L2_0/n4012 ), .force_11(
        1'b0), .Q(n40862), .QN(n8749) );
  \**FFGEN**  \L2_0/square_reg[1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8135), .force_10(\L2_0/n4016 ), .force_11(
        1'b0), .Q(n40781), .QN(n8750) );
  \**FFGEN**  \L2_0/square_reg[1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8137), .force_10(\L2_0/n4020 ), .force_11(
        1'b0), .Q(n40863), .QN(n8751) );
  \**FFGEN**  \L2_0/square_reg[1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8129), .force_10(\L2_0/n4024 ), .force_11(
        1'b0), .Q(n40780), .QN(n8752) );
  \**FFGEN**  \L2_0/square_reg[1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8139), .force_10(\L2_0/n4028 ), .force_11(
        1'b0), .Q(n40859), .QN(n8753) );
  \**FFGEN**  \L2_0/square_reg[1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8140), .force_10(\L2_0/n4032 ), .force_11(
        1'b0), .Q(n40864), .QN(n8754) );
  \**FFGEN**  \L2_0/square_reg[1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8132), .force_10(\L2_0/n4036 ), .force_11(
        1'b0), .QN(n8755) );
  \**FFGEN**  \L2_0/square_reg[1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8138), .force_10(\L2_0/n4040 ), .force_11(
        1'b0), .QN(n8756) );
  \**FFGEN**  \L2_0/square_reg[1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8144), .force_10(\L2_0/n4044 ), .force_11(
        1'b0), .QN(n8757) );
  \**FFGEN**  \L2_0/square_reg[1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8126), .force_10(\L2_0/n4048 ), .force_11(
        1'b0), .QN(n8758) );
  \**FFGEN**  \L2_0/square_reg[1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8130), .force_10(\L2_0/n4052 ), .force_11(
        1'b0), .QN(n8759) );
  \**FFGEN**  \L2_0/square_reg[1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8128), .force_10(\L2_0/n4056 ), .force_11(
        1'b0), .QN(n8760) );
  \**FFGEN**  \L2_0/square_reg[1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46553), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40833), .QN(n8761) );
  \**FFGEN**  \L2_0/square_reg[1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8131), .force_10(\L2_0/n4064 ), .force_11(
        1'b0), .QN(n8762) );
  \**FFGEN**  \L2_0/square_reg[0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8066), .force_10(\L2_0/n4068 ), .force_11(
        1'b0), .Q(n40804), .QN(n8763) );
  \**FFGEN**  \L2_0/square_reg[0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8065), .force_10(\L2_0/n4072 ), .force_11(
        1'b0), .Q(n40740), .QN(n8764) );
  \**FFGEN**  \L2_0/square_reg[0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8064), .force_10(\L2_0/n4076 ), .force_11(
        1'b0), .QN(n8765) );
  \**FFGEN**  \L2_0/square_reg[0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8051), .force_10(\L2_0/n4080 ), .force_11(
        1'b0), .Q(n40743), .QN(n8766) );
  \**FFGEN**  \L2_0/square_reg[0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8063), .force_10(\L2_0/n4084 ), .force_11(
        1'b0), .QN(n8767) );
  \**FFGEN**  \L2_0/square_reg[0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8062), .force_10(\L2_0/n4088 ), .force_11(
        1'b0), .Q(n40744), .QN(n8768) );
  \**FFGEN**  \L2_0/square_reg[0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8061), .force_10(\L2_0/n4092 ), .force_11(
        1'b0), .QN(n8769) );
  \**FFGEN**  \L2_0/square_reg[0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8053), .force_10(\L2_0/n4096 ), .force_11(
        1'b0), .Q(n40745), .QN(n8770) );
  \**FFGEN**  \L2_0/square_reg[0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8052), .force_10(\L2_0/n4100 ), .force_11(
        1'b0), .QN(n8771) );
  \**FFGEN**  \L2_0/square_reg[0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8060), .force_10(\L2_0/n4104 ), .force_11(
        1'b0), .Q(n40746), .QN(n8772) );
  \**FFGEN**  \L2_0/square_reg[0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8059), .force_10(\L2_0/n4108 ), .force_11(
        1'b0), .QN(n8773) );
  \**FFGEN**  \L2_0/square_reg[0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8048), .force_10(\L2_0/n4112 ), .force_11(
        1'b0), .Q(n40800), .QN(n8774) );
  \**FFGEN**  \L2_0/square_reg[0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8058), .force_10(\L2_0/n4116 ), .force_11(
        1'b0), .Q(n40797), .QN(n8775) );
  \**FFGEN**  \L2_0/square_reg[0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8057), .force_10(\L2_0/n4120 ), .force_11(
        1'b0), .Q(n40851), .QN(n8776) );
  \**FFGEN**  \L2_0/square_reg[0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8056), .force_10(\L2_0/n4124 ), .force_11(
        1'b0), .Q(n40795), .QN(n8777) );
  \**FFGEN**  \L2_0/square_reg[0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8049), .force_10(\L2_0/n4128 ), .force_11(
        1'b0), .Q(n40737), .QN(n8778) );
  \**FFGEN**  \L2_0/square_reg[0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8047), .force_10(\L2_0/n4132 ), .force_11(
        1'b0), .Q(n40721), .QN(n8779) );
  \**FFGEN**  \L2_0/square_reg[0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8055), .force_10(\L2_0/n4136 ), .force_11(
        1'b0), .Q(n40723), .QN(n8780) );
  \**FFGEN**  \L2_0/square_reg[0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n46577), .force_10(1'b0), .force_11(1'b0), 
        .Q(n40748), .QN(n8781) );
  \**FFGEN**  \L2_0/square_reg[0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n8054), .force_10(\L2_0/n4144 ), .force_11(
        1'b0), .QN(n8782) );
  \**FFGEN**  \L2_0/sum_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4147 ), .force_10(\L2_0/n4148 ), 
        .force_11(1'b0), .Q(out_L2[0]), .QN(n40726) );
  \**FFGEN**  \L2_0/sum_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4151 ), .force_10(\L2_0/n4152 ), 
        .force_11(1'b0), .Q(out_L2[1]), .QN(n40732) );
  \**FFGEN**  \L2_0/sum_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4155 ), .force_10(\L2_0/n4156 ), 
        .force_11(1'b0), .Q(out_L2[2]) );
  \**FFGEN**  \L2_0/sum_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4159 ), .force_10(\L2_0/n4160 ), 
        .force_11(1'b0), .Q(out_L2[3]), .QN(n40787) );
  \**FFGEN**  \L2_0/sum_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4163 ), .force_10(\L2_0/n4164 ), 
        .force_11(1'b0), .Q(out_L2[4]), .QN(n40788) );
  \**FFGEN**  \L2_0/sum_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4167 ), .force_10(\L2_0/n4168 ), 
        .force_11(1'b0), .Q(out_L2[5]), .QN(n40793) );
  \**FFGEN**  \L2_0/sum_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4171 ), .force_10(\L2_0/n4172 ), 
        .force_11(1'b0), .Q(out_L2[6]), .QN(n40805) );
  \**FFGEN**  \L2_0/sum_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4175 ), .force_10(\L2_0/n4176 ), 
        .force_11(1'b0), .Q(out_L2[7]), .QN(n40791) );
  \**FFGEN**  \L2_0/sum_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4179 ), .force_10(\L2_0/n4180 ), 
        .force_11(1'b0), .Q(out_L2[8]), .QN(n40799) );
  \**FFGEN**  \L2_0/sum_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4183 ), .force_10(\L2_0/n4184 ), 
        .force_11(1'b0), .Q(out_L2[9]), .QN(n40841) );
  \**FFGEN**  \L2_0/sum_reg[10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4187 ), .force_10(\L2_0/n4188 ), 
        .force_11(1'b0), .Q(out_L2[10]), .QN(n40730) );
  \**FFGEN**  \L2_0/sum_reg[11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4191 ), .force_10(\L2_0/n4192 ), 
        .force_11(1'b0), .Q(out_L2[11]), .QN(n40845) );
  \**FFGEN**  \L2_0/sum_reg[12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4195 ), .force_10(\L2_0/n4196 ), 
        .force_11(1'b0), .Q(out_L2[12]), .QN(n40729) );
  \**FFGEN**  \L2_0/sum_reg[13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4199 ), .force_10(\L2_0/n4200 ), 
        .force_11(1'b0), .Q(out_L2[13]), .QN(n40844) );
  \**FFGEN**  \L2_0/sum_reg[14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4203 ), .force_10(\L2_0/n4204 ), 
        .force_11(1'b0), .Q(out_L2[14]), .QN(n40728) );
  \**FFGEN**  \L2_0/sum_reg[15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4207 ), .force_10(\L2_0/n4208 ), 
        .force_11(1'b0), .Q(out_L2[15]), .QN(n40843) );
  \**FFGEN**  \L2_0/sum_reg[16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4211 ), .force_10(\L2_0/n4212 ), 
        .force_11(1'b0), .Q(out_L2[16]), .QN(n40727) );
  \**FFGEN**  \L2_0/sum_reg[17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4215 ), .force_10(\L2_0/n4216 ), 
        .force_11(1'b0), .Q(out_L2[17]), .QN(n40842) );
  \**FFGEN**  \L2_0/sum_reg[18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n4219 ), .force_10(\L2_0/n4220 ), 
        .force_11(1'b0), .Q(out_L2[18]), .QN(n40739) );
  \**FFGEN**  \L2_0/sum_reg[19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2903 ), .force_10(\L2_0/n2904 ), 
        .force_11(1'b0), .Q(out_L2[19]), .QN(n40803) );
  nand_x8_sg U10131 ( .A(n46579), .B(n46578), .X(n9012) );
  nand_x8_sg U36316 ( .A(n32138), .B(n55511), .X(n39300) );
  nand_x8_sg U10130 ( .A(n11831), .B(n24470), .X(n8050) );
  nand_x8_sg U12251 ( .A(n13393), .B(n24471), .X(n11831) );
  nand_x8_sg U24926 ( .A(n46576), .B(n46579), .X(n13393) );
  nand_x8_sg U32365 ( .A(n55459), .B(n46583), .X(n26078) );
  nand_x8_sg U10129 ( .A(n46582), .B(n13393), .X(n24470) );
  nor_x2_sg U4816 ( .A(n22615), .B(n8543), .X(n22613) );
  nand_x8_sg U5044 ( .A(n22774), .B(n50938), .X(n9391) );
  nand_x8_sg U5039 ( .A(n22870), .B(n22871), .X(n22612) );
  nor_x2_sg U5264 ( .A(n23119), .B(n50862), .X(n23034) );
  nor_x2_sg U5263 ( .A(n22867), .B(n8585), .X(n23119) );
  nand_x8_sg U5262 ( .A(n23121), .B(n23122), .X(n22867) );
  nand_x8_sg U5485 ( .A(n23339), .B(n23340), .X(n23118) );
  nor_x2_sg U5710 ( .A(n23538), .B(n50774), .X(n23471) );
  nor_x2_sg U5709 ( .A(n23336), .B(n8627), .X(n23538) );
  nand_x8_sg U5708 ( .A(n23540), .B(n23541), .X(n23336) );
  nand_x8_sg U5940 ( .A(n23662), .B(n50749), .X(n9572) );
  nand_x8_sg U6161 ( .A(n50701), .B(n23836), .X(n9648) );
  nor_x2_sg U6157 ( .A(n23720), .B(n8669), .X(n23886) );
  nand_x8_sg U6156 ( .A(n23888), .B(n23889), .X(n23720) );
  nand_x8_sg U6385 ( .A(n23992), .B(n50653), .X(n9672) );
  nand_x8_sg U6380 ( .A(n24035), .B(n24036), .X(n23885) );
  nor_x2_sg U6605 ( .A(n24031), .B(n8711), .X(n24170) );
  nand_x8_sg U6604 ( .A(n24172), .B(n24173), .X(n24031) );
  nand_x8_sg U6833 ( .A(n24258), .B(n50554), .X(n24135) );
  nand_x8_sg U6828 ( .A(n24282), .B(n24283), .X(n24169) );
  nor_x2_sg U7054 ( .A(n24279), .B(n8753), .X(n24375) );
  nand_x8_sg U7280 ( .A(n24444), .B(n50458), .X(n24358) );
  nand_x8_sg U7273 ( .A(n24447), .B(n24448), .X(n24372) );
  nand_x8_sg U7742 ( .A(n24453), .B(n24454), .X(n24435) );
  nand_x8_sg U8683 ( .A(n24465), .B(n24466), .X(n24411) );
  nor_x2_sg U8445 ( .A(n24411), .B(n8780), .X(n24464) );
  nor_x2_sg U7976 ( .A(n50227), .B(n8778), .X(n24458) );
  nor_x2_sg U7504 ( .A(n24435), .B(n8776), .X(n24452) );
  nor_x2_sg U7513 ( .A(n24442), .B(n24443), .X(n24440) );
  nand_x8_sg U7523 ( .A(n24383), .B(n24384), .X(n24355) );
  nand_x8_sg U7759 ( .A(n24386), .B(n24387), .X(n24348) );
  nand_x8_sg U7994 ( .A(n24389), .B(n24390), .X(n24342) );
  nor_x2_sg U8219 ( .A(n24424), .B(n24425), .X(n24422) );
  nor_x2_sg U8216 ( .A(n40788), .B(n8778), .X(n24425) );
  nand_x8_sg U8229 ( .A(n24392), .B(n24393), .X(n24335) );
  nor_x2_sg U8450 ( .A(n40787), .B(n8779), .X(n24419) );
  nand_x8_sg U8463 ( .A(n24395), .B(n24396), .X(n24329) );
  nand_x8_sg U8696 ( .A(n24398), .B(n24399), .X(n24323) );
  nand_x8_sg U7046 ( .A(n24366), .B(n50504), .X(n24278) );
  nand_x8_sg U7039 ( .A(n24369), .B(n50456), .X(n24269) );
  nor_x2_sg U7035 ( .A(n24372), .B(n8774), .X(n24371) );
  nand_x8_sg U7063 ( .A(n24285), .B(n24286), .X(n24256) );
  nor_x2_sg U7289 ( .A(n24362), .B(n8754), .X(n24360) );
  nand_x8_sg U7298 ( .A(n24288), .B(n24289), .X(n24250) );
  nor_x2_sg U7524 ( .A(n24355), .B(n8755), .X(n24353) );
  nand_x8_sg U7533 ( .A(n24291), .B(n24292), .X(n24244) );
  nor_x2_sg U7761 ( .A(n24346), .B(n50362), .X(n24345) );
  nor_x2_sg U7760 ( .A(n24348), .B(n8756), .X(n24346) );
  nand_x8_sg U7769 ( .A(n24294), .B(n24295), .X(n24238) );
  nor_x2_sg U7995 ( .A(n24342), .B(n8757), .X(n24340) );
  nand_x8_sg U8004 ( .A(n24297), .B(n24298), .X(n24232) );
  nor_x2_sg U8231 ( .A(n24333), .B(n50271), .X(n24332) );
  nor_x2_sg U8230 ( .A(n24335), .B(n8758), .X(n24333) );
  nand_x8_sg U8239 ( .A(n24300), .B(n24301), .X(n24226) );
  nor_x2_sg U8465 ( .A(n24327), .B(n50226), .X(n24326) );
  nor_x2_sg U8464 ( .A(n24329), .B(n8759), .X(n24327) );
  nand_x8_sg U8473 ( .A(n24303), .B(n24304), .X(n24220) );
  nor_x2_sg U8697 ( .A(n24323), .B(n8760), .X(n24321) );
  nand_x8_sg U8705 ( .A(n24306), .B(n24307), .X(n24214) );
  nand_x8_sg U9039 ( .A(n50110), .B(n24309), .X(n10245) );
  nor_x2_sg U6819 ( .A(n24163), .B(n8752), .X(n24273) );
  nand_x8_sg U6818 ( .A(n24275), .B(n24276), .X(n24163) );
  nand_x8_sg U6811 ( .A(n24264), .B(n24265), .X(n24162) );
  nor_x2_sg U6799 ( .A(n24269), .B(n8773), .X(n24268) );
  nand_x8_sg U6840 ( .A(n24175), .B(n24176), .X(n24138) );
  nand_x8_sg U7075 ( .A(n24178), .B(n24179), .X(n24131) );
  nand_x8_sg U7310 ( .A(n24181), .B(n24182), .X(n24124) );
  nand_x8_sg U7545 ( .A(n24184), .B(n24185), .X(n24117) );
  nand_x8_sg U7781 ( .A(n24187), .B(n24188), .X(n24110) );
  nand_x8_sg U8016 ( .A(n24190), .B(n24191), .X(n24103) );
  nand_x8_sg U8251 ( .A(n24193), .B(n24194), .X(n24096) );
  nand_x8_sg U8485 ( .A(n24196), .B(n24197), .X(n24089) );
  nand_x8_sg U8716 ( .A(n24199), .B(n24200), .X(n24082) );
  nand_x8_sg U6597 ( .A(n24142), .B(n50600), .X(n24032) );
  nand_x8_sg U6592 ( .A(n24166), .B(n24167), .X(n24025) );
  nor_x2_sg U6583 ( .A(n24019), .B(n8751), .X(n24157) );
  nand_x8_sg U6575 ( .A(n24148), .B(n50595), .X(n24018) );
  nand_x8_sg U6568 ( .A(n24151), .B(n24152), .X(n24009) );
  nand_x8_sg U6614 ( .A(n24038), .B(n24039), .X(n23990) );
  nor_x2_sg U6841 ( .A(n24138), .B(n8712), .X(n24136) );
  nand_x8_sg U6850 ( .A(n24041), .B(n24042), .X(n23984) );
  nor_x2_sg U7076 ( .A(n24131), .B(n8713), .X(n24129) );
  nand_x8_sg U7085 ( .A(n24044), .B(n24045), .X(n23978) );
  nor_x2_sg U7311 ( .A(n24124), .B(n8714), .X(n24122) );
  nand_x8_sg U7320 ( .A(n24047), .B(n24048), .X(n23972) );
  nor_x2_sg U7546 ( .A(n24117), .B(n8715), .X(n24115) );
  nand_x8_sg U7555 ( .A(n24050), .B(n24051), .X(n23966) );
  nor_x2_sg U7782 ( .A(n24110), .B(n8716), .X(n24108) );
  nand_x8_sg U7791 ( .A(n24053), .B(n24054), .X(n23960) );
  nor_x2_sg U8017 ( .A(n24103), .B(n8717), .X(n24101) );
  nand_x8_sg U8026 ( .A(n24056), .B(n24057), .X(n23954) );
  nor_x2_sg U8252 ( .A(n24096), .B(n8718), .X(n24094) );
  nand_x8_sg U8261 ( .A(n24059), .B(n24060), .X(n23948) );
  nor_x2_sg U8486 ( .A(n24089), .B(n8719), .X(n24087) );
  nand_x8_sg U8495 ( .A(n24062), .B(n24063), .X(n23942) );
  nor_x2_sg U8717 ( .A(n24082), .B(n8720), .X(n24080) );
  nand_x8_sg U8725 ( .A(n24065), .B(n24066), .X(n23936) );
  nand_x8_sg U9045 ( .A(n50113), .B(n24068), .X(n10241) );
  nor_x2_sg U6371 ( .A(n23878), .B(n8710), .X(n24026) );
  nand_x8_sg U6370 ( .A(n24028), .B(n24029), .X(n23878) );
  nand_x8_sg U6363 ( .A(n23998), .B(n50646), .X(n23879) );
  nand_x8_sg U6358 ( .A(n24022), .B(n24023), .X(n23872) );
  nor_x2_sg U6349 ( .A(n23866), .B(n8750), .X(n24013) );
  nand_x8_sg U6348 ( .A(n24015), .B(n24016), .X(n23866) );
  nand_x8_sg U6341 ( .A(n24004), .B(n24005), .X(n23865) );
  nor_x2_sg U6329 ( .A(n24009), .B(n8771), .X(n24008) );
  nand_x8_sg U6392 ( .A(n23891), .B(n23892), .X(n23835) );
  nand_x8_sg U6619 ( .A(n23986), .B(n50605), .X(n9719) );
  nand_x8_sg U6626 ( .A(n23894), .B(n23895), .X(n23829) );
  nand_x8_sg U6855 ( .A(n23980), .B(n50556), .X(n9767) );
  nand_x8_sg U6862 ( .A(n23897), .B(n23898), .X(n23823) );
  nand_x8_sg U7090 ( .A(n23974), .B(n50509), .X(n9815) );
  nand_x8_sg U7097 ( .A(n23900), .B(n23901), .X(n23817) );
  nand_x8_sg U7325 ( .A(n23968), .B(n50462), .X(n9863) );
  nand_x8_sg U7332 ( .A(n23903), .B(n23904), .X(n23811) );
  nand_x8_sg U7560 ( .A(n23962), .B(n50416), .X(n9911) );
  nand_x8_sg U7567 ( .A(n23906), .B(n23907), .X(n23805) );
  nand_x8_sg U7796 ( .A(n23956), .B(n50369), .X(n9959) );
  nand_x8_sg U7803 ( .A(n23909), .B(n23910), .X(n23799) );
  nand_x8_sg U8031 ( .A(n23950), .B(n50322), .X(n10008) );
  nand_x8_sg U8038 ( .A(n23912), .B(n23913), .X(n23793) );
  nand_x8_sg U8266 ( .A(n23944), .B(n50276), .X(n10056) );
  nand_x8_sg U8273 ( .A(n23915), .B(n23916), .X(n23787) );
  nand_x8_sg U8500 ( .A(n23938), .B(n50230), .X(n10105) );
  nand_x8_sg U8507 ( .A(n23918), .B(n23919), .X(n23781) );
  nand_x8_sg U8730 ( .A(n23932), .B(n50186), .X(n10154) );
  nand_x8_sg U8736 ( .A(n23921), .B(n23922), .X(n23775) );
  nand_x8_sg U8922 ( .A(n23925), .B(n23926), .X(n10200) );
  nand_x8_sg U9048 ( .A(n50114), .B(n23924), .X(n10244) );
  nand_x8_sg U6149 ( .A(n23839), .B(n50698), .X(n9624) );
  nand_x8_sg U6144 ( .A(n23882), .B(n23883), .X(n23714) );
  nor_x2_sg U6135 ( .A(n23707), .B(n8709), .X(n23873) );
  nand_x8_sg U6134 ( .A(n23875), .B(n23876), .X(n23707) );
  nand_x8_sg U6127 ( .A(n23845), .B(n50691), .X(n23708) );
  nand_x8_sg U6122 ( .A(n23869), .B(n23870), .X(n23701) );
  nor_x2_sg U6113 ( .A(n23695), .B(n8749), .X(n23860) );
  nand_x8_sg U6105 ( .A(n23851), .B(n50686), .X(n23694) );
  nand_x8_sg U6098 ( .A(n23854), .B(n23855), .X(n23685) );
  nor_x2_sg U6393 ( .A(n23835), .B(n8670), .X(n23833) );
  nand_x8_sg U6631 ( .A(n50606), .B(n23824), .X(n9743) );
  nor_x2_sg U6627 ( .A(n23829), .B(n8671), .X(n23827) );
  nand_x8_sg U6867 ( .A(n50557), .B(n23818), .X(n9791) );
  nor_x2_sg U6863 ( .A(n23823), .B(n8672), .X(n23821) );
  nand_x8_sg U7102 ( .A(n50510), .B(n23812), .X(n9839) );
  nor_x2_sg U7098 ( .A(n23817), .B(n8673), .X(n23815) );
  nand_x8_sg U7337 ( .A(n50463), .B(n23806), .X(n9887) );
  nor_x2_sg U7333 ( .A(n23811), .B(n8674), .X(n23809) );
  nand_x8_sg U7572 ( .A(n50417), .B(n23800), .X(n9935) );
  nor_x2_sg U7568 ( .A(n23805), .B(n8675), .X(n23803) );
  nand_x8_sg U7808 ( .A(n50370), .B(n23794), .X(n9984) );
  nor_x2_sg U7804 ( .A(n23799), .B(n8676), .X(n23797) );
  nand_x8_sg U8043 ( .A(n50323), .B(n23788), .X(n10032) );
  nor_x2_sg U8039 ( .A(n23793), .B(n8677), .X(n23791) );
  nand_x8_sg U8278 ( .A(n50277), .B(n23782), .X(n10081) );
  nor_x2_sg U8274 ( .A(n23787), .B(n8678), .X(n23785) );
  nand_x8_sg U8512 ( .A(n50231), .B(n23776), .X(n10130) );
  nor_x2_sg U8508 ( .A(n23781), .B(n8679), .X(n23779) );
  nor_x2_sg U8737 ( .A(n23775), .B(n8680), .X(n23773) );
  nand_x8_sg U8746 ( .A(n23760), .B(n23761), .X(n23595) );
  nor_x2_sg U5923 ( .A(n23530), .B(n8668), .X(n23715) );
  nand_x8_sg U5922 ( .A(n23717), .B(n23718), .X(n23530) );
  nand_x8_sg U5915 ( .A(n23668), .B(n50744), .X(n9576) );
  nand_x8_sg U5910 ( .A(n23711), .B(n23712), .X(n23524) );
  nor_x2_sg U5901 ( .A(n23517), .B(n8708), .X(n23702) );
  nand_x8_sg U5900 ( .A(n23704), .B(n23705), .X(n23517) );
  nand_x8_sg U5893 ( .A(n23674), .B(n50737), .X(n23518) );
  nand_x8_sg U5888 ( .A(n23698), .B(n23699), .X(n23511) );
  nor_x2_sg U5879 ( .A(n23505), .B(n8748), .X(n23689) );
  nand_x8_sg U5878 ( .A(n23691), .B(n23692), .X(n23505) );
  nand_x8_sg U5871 ( .A(n23680), .B(n23681), .X(n23504) );
  nor_x2_sg U5859 ( .A(n23685), .B(n8769), .X(n23684) );
  nand_x8_sg U5947 ( .A(n23543), .B(n23544), .X(n23468) );
  nand_x8_sg U6173 ( .A(n50702), .B(n23656), .X(n9620) );
  nor_x2_sg U6169 ( .A(n23661), .B(n8649), .X(n23659) );
  nand_x8_sg U6180 ( .A(n23546), .B(n23547), .X(n23462) );
  nand_x8_sg U6410 ( .A(n50656), .B(n23650), .X(n9668) );
  nand_x8_sg U6417 ( .A(n23549), .B(n23550), .X(n23456) );
  nand_x8_sg U6644 ( .A(n50607), .B(n23644), .X(n9715) );
  nor_x2_sg U6640 ( .A(n50585), .B(n8651), .X(n23647) );
  nand_x8_sg U6651 ( .A(n23552), .B(n23553), .X(n23450) );
  nand_x8_sg U6880 ( .A(n50558), .B(n23638), .X(n9763) );
  nor_x2_sg U6876 ( .A(n50539), .B(n8652), .X(n23641) );
  nand_x8_sg U6887 ( .A(n23555), .B(n23556), .X(n23444) );
  nand_x8_sg U7115 ( .A(n50511), .B(n23632), .X(n9811) );
  nor_x2_sg U7111 ( .A(n43025), .B(n8653), .X(n23635) );
  nand_x8_sg U7122 ( .A(n23558), .B(n23559), .X(n23438) );
  nand_x8_sg U7350 ( .A(n50464), .B(n23626), .X(n9859) );
  nor_x2_sg U7346 ( .A(n50445), .B(n8654), .X(n23629) );
  nand_x8_sg U7357 ( .A(n23561), .B(n23562), .X(n23432) );
  nand_x8_sg U7585 ( .A(n50418), .B(n23620), .X(n9907) );
  nor_x2_sg U7581 ( .A(n50399), .B(n8655), .X(n23623) );
  nand_x8_sg U7592 ( .A(n23564), .B(n23565), .X(n23426) );
  nand_x8_sg U7821 ( .A(n50371), .B(n23614), .X(n9955) );
  nor_x2_sg U7817 ( .A(n43020), .B(n8656), .X(n23617) );
  nand_x8_sg U7828 ( .A(n23567), .B(n23568), .X(n23420) );
  nand_x8_sg U8056 ( .A(n50324), .B(n23608), .X(n10004) );
  nor_x2_sg U8052 ( .A(n50305), .B(n8657), .X(n23611) );
  nand_x8_sg U8063 ( .A(n23570), .B(n23571), .X(n23414) );
  nand_x8_sg U8291 ( .A(n50278), .B(n23602), .X(n10052) );
  nor_x2_sg U8287 ( .A(n23607), .B(n8658), .X(n23605) );
  nand_x8_sg U8298 ( .A(n23573), .B(n23574), .X(n23408) );
  nand_x8_sg U8525 ( .A(n50232), .B(n23596), .X(n10101) );
  nor_x2_sg U8521 ( .A(n23601), .B(n8659), .X(n23599) );
  nand_x8_sg U8532 ( .A(n23576), .B(n23577), .X(n23402) );
  nand_x8_sg U8751 ( .A(n23589), .B(n23590), .X(n10150) );
  nor_x2_sg U8748 ( .A(n23593), .B(n50168), .X(n23591) );
  nor_x2_sg U8747 ( .A(n23595), .B(n8660), .X(n23593) );
  nand_x8_sg U8757 ( .A(n23579), .B(n23580), .X(n23396) );
  nand_x8_sg U8936 ( .A(n23583), .B(n23584), .X(n10197) );
  nand_x8_sg U9054 ( .A(n50117), .B(n23582), .X(n10240) );
  nand_x8_sg U5701 ( .A(n50796), .B(n23472), .X(n9523) );
  nor_x2_sg U5697 ( .A(n23533), .B(n8647), .X(n23531) );
  nand_x8_sg U5689 ( .A(n50793), .B(n23475), .X(n9552) );
  nor_x2_sg U5685 ( .A(n23325), .B(n8667), .X(n23525) );
  nand_x8_sg U5684 ( .A(n23527), .B(n23528), .X(n23325) );
  nand_x8_sg U5677 ( .A(n23478), .B(n50790), .X(n9527) );
  nand_x8_sg U5672 ( .A(n23521), .B(n23522), .X(n23319) );
  nor_x2_sg U5663 ( .A(n23312), .B(n8707), .X(n23512) );
  nand_x8_sg U5662 ( .A(n23514), .B(n23515), .X(n23312) );
  nand_x8_sg U5655 ( .A(n23484), .B(n50783), .X(n23313) );
  nand_x8_sg U5650 ( .A(n23508), .B(n23509), .X(n23306) );
  nor_x2_sg U5641 ( .A(n23300), .B(n8747), .X(n23499) );
  nand_x8_sg U5633 ( .A(n23490), .B(n50778), .X(n23299) );
  nand_x8_sg U5626 ( .A(n23493), .B(n23494), .X(n23290) );
  nand_x8_sg U5718 ( .A(n23342), .B(n23343), .X(n23259) );
  nor_x2_sg U5949 ( .A(n23466), .B(n50728), .X(n23465) );
  nor_x2_sg U5948 ( .A(n23468), .B(n8628), .X(n23466) );
  nand_x8_sg U5957 ( .A(n23345), .B(n23346), .X(n23253) );
  nor_x2_sg U6182 ( .A(n23460), .B(n50680), .X(n23459) );
  nor_x2_sg U6181 ( .A(n23462), .B(n8629), .X(n23460) );
  nand_x8_sg U6190 ( .A(n23348), .B(n23349), .X(n23247) );
  nor_x2_sg U6418 ( .A(n23456), .B(n8630), .X(n23454) );
  nand_x8_sg U6427 ( .A(n23351), .B(n23352), .X(n23241) );
  nor_x2_sg U6653 ( .A(n23448), .B(n50584), .X(n23447) );
  nor_x2_sg U6652 ( .A(n23450), .B(n8631), .X(n23448) );
  nand_x8_sg U6661 ( .A(n23354), .B(n23355), .X(n23235) );
  nor_x2_sg U6889 ( .A(n23442), .B(n50537), .X(n23441) );
  nor_x2_sg U6888 ( .A(n23444), .B(n8632), .X(n23442) );
  nand_x8_sg U6897 ( .A(n23357), .B(n23358), .X(n23229) );
  nor_x2_sg U7124 ( .A(n23436), .B(n50490), .X(n23435) );
  nor_x2_sg U7123 ( .A(n23438), .B(n8633), .X(n23436) );
  nand_x8_sg U7132 ( .A(n23360), .B(n23361), .X(n23223) );
  nor_x2_sg U7359 ( .A(n23430), .B(n50444), .X(n23429) );
  nor_x2_sg U7358 ( .A(n23432), .B(n8634), .X(n23430) );
  nand_x8_sg U7367 ( .A(n23363), .B(n23364), .X(n23217) );
  nor_x2_sg U7594 ( .A(n23424), .B(n50397), .X(n23423) );
  nor_x2_sg U7593 ( .A(n23426), .B(n8635), .X(n23424) );
  nand_x8_sg U7602 ( .A(n23366), .B(n23367), .X(n23211) );
  nor_x2_sg U7830 ( .A(n23418), .B(n50350), .X(n23417) );
  nor_x2_sg U7829 ( .A(n23420), .B(n8636), .X(n23418) );
  nand_x8_sg U7838 ( .A(n23369), .B(n23370), .X(n23205) );
  nor_x2_sg U8065 ( .A(n23412), .B(n50304), .X(n23411) );
  nor_x2_sg U8064 ( .A(n23414), .B(n8637), .X(n23412) );
  nand_x8_sg U8073 ( .A(n23372), .B(n23373), .X(n23199) );
  nor_x2_sg U8300 ( .A(n23406), .B(n50258), .X(n23405) );
  nor_x2_sg U8299 ( .A(n23408), .B(n8638), .X(n23406) );
  nand_x8_sg U8308 ( .A(n23375), .B(n23376), .X(n23193) );
  nor_x2_sg U8534 ( .A(n23400), .B(n50214), .X(n23399) );
  nor_x2_sg U8533 ( .A(n23402), .B(n8639), .X(n23400) );
  nand_x8_sg U8542 ( .A(n23378), .B(n23379), .X(n23187) );
  nor_x2_sg U8759 ( .A(n23394), .B(n50166), .X(n23393) );
  nor_x2_sg U8758 ( .A(n23396), .B(n8640), .X(n23394) );
  nand_x8_sg U8766 ( .A(n23381), .B(n23382), .X(n23181) );
  nand_x8_sg U9057 ( .A(n50118), .B(n23384), .X(n10252) );
  nor_x2_sg U5477 ( .A(n23331), .B(n50798), .X(n23266) );
  nor_x2_sg U5476 ( .A(n23112), .B(n8626), .X(n23331) );
  nand_x8_sg U5475 ( .A(n23333), .B(n23334), .X(n23112) );
  nand_x8_sg U5468 ( .A(n23267), .B(n50839), .X(n9474) );
  nor_x2_sg U5451 ( .A(n23099), .B(n8666), .X(n23320) );
  nand_x8_sg U5450 ( .A(n23322), .B(n23323), .X(n23099) );
  nand_x8_sg U5443 ( .A(n23273), .B(n50834), .X(n9478) );
  nand_x8_sg U5438 ( .A(n23316), .B(n23317), .X(n23093) );
  nor_x2_sg U5429 ( .A(n23086), .B(n8706), .X(n23307) );
  nand_x8_sg U5428 ( .A(n23309), .B(n23310), .X(n23086) );
  nand_x8_sg U5421 ( .A(n23279), .B(n50827), .X(n23087) );
  nand_x8_sg U5416 ( .A(n23303), .B(n23304), .X(n23080) );
  nor_x2_sg U5407 ( .A(n23074), .B(n8746), .X(n23294) );
  nand_x8_sg U5406 ( .A(n23296), .B(n23297), .X(n23074) );
  nand_x8_sg U5399 ( .A(n23285), .B(n23286), .X(n23073) );
  nor_x2_sg U5387 ( .A(n23290), .B(n8767), .X(n23289) );
  nand_x8_sg U5499 ( .A(n23124), .B(n23125), .X(n23031) );
  nand_x8_sg U5732 ( .A(n23127), .B(n23128), .X(n23025) );
  nand_x8_sg U5969 ( .A(n23130), .B(n23131), .X(n23019) );
  nand_x8_sg U6202 ( .A(n23133), .B(n23134), .X(n23012) );
  nand_x8_sg U6439 ( .A(n23136), .B(n23137), .X(n23005) );
  nand_x8_sg U6673 ( .A(n23139), .B(n23140), .X(n22998) );
  nand_x8_sg U6909 ( .A(n23142), .B(n23143), .X(n22991) );
  nand_x8_sg U7144 ( .A(n23145), .B(n23146), .X(n22984) );
  nand_x8_sg U7379 ( .A(n23148), .B(n23149), .X(n22977) );
  nand_x8_sg U7614 ( .A(n23151), .B(n23152), .X(n22970) );
  nand_x8_sg U7850 ( .A(n23154), .B(n23155), .X(n22963) );
  nand_x8_sg U8085 ( .A(n23157), .B(n23158), .X(n22956) );
  nand_x8_sg U8320 ( .A(n23160), .B(n23161), .X(n22949) );
  nand_x8_sg U8554 ( .A(n23163), .B(n23164), .X(n22942) );
  nand_x8_sg U8777 ( .A(n23166), .B(n23167), .X(n22935) );
  nand_x8_sg U9060 ( .A(n50119), .B(n23169), .X(n10255) );
  nand_x8_sg U5248 ( .A(n23115), .B(n23116), .X(n22861) );
  nor_x2_sg U5240 ( .A(n23107), .B(n50841), .X(n23040) );
  nor_x2_sg U5239 ( .A(n22855), .B(n8625), .X(n23107) );
  nand_x8_sg U5238 ( .A(n23109), .B(n23110), .X(n22855) );
  nand_x8_sg U5231 ( .A(n50884), .B(n23041), .X(n9425) );
  nor_x2_sg U5227 ( .A(n23102), .B(n8645), .X(n23100) );
  nand_x8_sg U5219 ( .A(n50881), .B(n23044), .X(n9454) );
  nor_x2_sg U5215 ( .A(n22844), .B(n8665), .X(n23094) );
  nand_x8_sg U5214 ( .A(n23096), .B(n23097), .X(n22844) );
  nand_x8_sg U5207 ( .A(n23047), .B(n50878), .X(n9429) );
  nand_x8_sg U5202 ( .A(n23090), .B(n23091), .X(n22838) );
  nor_x2_sg U5193 ( .A(n22831), .B(n8705), .X(n23081) );
  nand_x8_sg U5192 ( .A(n23083), .B(n23084), .X(n22831) );
  nand_x8_sg U5185 ( .A(n23053), .B(n50871), .X(n22832) );
  nand_x8_sg U5180 ( .A(n23077), .B(n23078), .X(n22825) );
  nor_x2_sg U5171 ( .A(n22819), .B(n8745), .X(n23068) );
  nand_x8_sg U5170 ( .A(n23070), .B(n23071), .X(n22819) );
  nand_x8_sg U5163 ( .A(n23059), .B(n50865), .X(n22818) );
  nand_x8_sg U5156 ( .A(n23062), .B(n23063), .X(n22809) );
  nand_x8_sg U5272 ( .A(n22873), .B(n22874), .X(n22772) );
  nor_x2_sg U5501 ( .A(n23029), .B(n50818), .X(n23028) );
  nor_x2_sg U5500 ( .A(n23031), .B(n8586), .X(n23029) );
  nand_x8_sg U5509 ( .A(n22876), .B(n22877), .X(n22766) );
  nor_x2_sg U5734 ( .A(n23023), .B(n50770), .X(n23022) );
  nor_x2_sg U5733 ( .A(n23025), .B(n8587), .X(n23023) );
  nand_x8_sg U5742 ( .A(n22879), .B(n22880), .X(n22760) );
  nor_x2_sg U5970 ( .A(n23019), .B(n8588), .X(n23017) );
  nand_x8_sg U5979 ( .A(n22882), .B(n22883), .X(n22754) );
  nor_x2_sg U6203 ( .A(n23012), .B(n8589), .X(n23010) );
  nand_x8_sg U6212 ( .A(n22885), .B(n22886), .X(n22748) );
  nor_x2_sg U6440 ( .A(n23005), .B(n8590), .X(n23003) );
  nand_x8_sg U6449 ( .A(n22888), .B(n22889), .X(n22742) );
  nor_x2_sg U6674 ( .A(n22998), .B(n8591), .X(n22996) );
  nand_x8_sg U6683 ( .A(n22891), .B(n22892), .X(n22736) );
  nor_x2_sg U6910 ( .A(n22991), .B(n8592), .X(n22989) );
  nand_x8_sg U6919 ( .A(n22894), .B(n22895), .X(n22730) );
  nor_x2_sg U7145 ( .A(n22984), .B(n8593), .X(n22982) );
  nand_x8_sg U7154 ( .A(n22897), .B(n22898), .X(n22724) );
  nor_x2_sg U7380 ( .A(n22977), .B(n8594), .X(n22975) );
  nand_x8_sg U7389 ( .A(n22900), .B(n22901), .X(n22718) );
  nor_x2_sg U7615 ( .A(n22970), .B(n8595), .X(n22968) );
  nand_x8_sg U7624 ( .A(n22903), .B(n22904), .X(n22712) );
  nor_x2_sg U7851 ( .A(n22963), .B(n8596), .X(n22961) );
  nand_x8_sg U7860 ( .A(n22906), .B(n22907), .X(n22706) );
  nor_x2_sg U8086 ( .A(n22956), .B(n8597), .X(n22954) );
  nand_x8_sg U8095 ( .A(n22909), .B(n22910), .X(n22700) );
  nor_x2_sg U8321 ( .A(n22949), .B(n8598), .X(n22947) );
  nand_x8_sg U8330 ( .A(n22912), .B(n22913), .X(n22694) );
  nor_x2_sg U8555 ( .A(n22942), .B(n8599), .X(n22940) );
  nand_x8_sg U8564 ( .A(n22915), .B(n22916), .X(n22688) );
  nor_x2_sg U8778 ( .A(n22935), .B(n8600), .X(n22933) );
  nand_x8_sg U8786 ( .A(n22918), .B(n22919), .X(n22682) );
  nand_x8_sg U9063 ( .A(n50120), .B(n22921), .X(n10260) );
  nor_x2_sg U5030 ( .A(n22605), .B(n8584), .X(n22862) );
  nand_x8_sg U5029 ( .A(n22864), .B(n22865), .X(n22605) );
  nand_x8_sg U5015 ( .A(n22858), .B(n22859), .X(n22598) );
  nor_x2_sg U5007 ( .A(n22850), .B(n50886), .X(n22785) );
  nor_x2_sg U5006 ( .A(n22591), .B(n8624), .X(n22850) );
  nand_x8_sg U5005 ( .A(n22852), .B(n22853), .X(n22591) );
  nand_x8_sg U4998 ( .A(n50926), .B(n22786), .X(n9364) );
  nor_x2_sg U4981 ( .A(n22576), .B(n8664), .X(n22839) );
  nand_x8_sg U4980 ( .A(n22841), .B(n22842), .X(n22576) );
  nand_x8_sg U4973 ( .A(n22792), .B(n50921), .X(n9370) );
  nand_x8_sg U4968 ( .A(n22835), .B(n22836), .X(n22569) );
  nor_x2_sg U4959 ( .A(n22562), .B(n8704), .X(n22826) );
  nand_x8_sg U4958 ( .A(n22828), .B(n22829), .X(n22562) );
  nand_x8_sg U4951 ( .A(n22798), .B(n50915), .X(n22561) );
  nand_x8_sg U4946 ( .A(n22822), .B(n22823), .X(n22554) );
  nor_x2_sg U4937 ( .A(n22547), .B(n8744), .X(n22813) );
  nand_x8_sg U4936 ( .A(n22815), .B(n22816), .X(n22547) );
  nor_x2_sg U4917 ( .A(n22809), .B(n8765), .X(n22808) );
  nand_x8_sg U5051 ( .A(n22619), .B(n22620), .X(n22184) );
  nand_x8_sg U5277 ( .A(n22768), .B(n50893), .X(n9446) );
  nand_x8_sg U5284 ( .A(n22622), .B(n22623), .X(n22350) );
  nand_x8_sg U5514 ( .A(n22762), .B(n50846), .X(n9495) );
  nand_x8_sg U5521 ( .A(n22625), .B(n22626), .X(n22497) );
  nand_x8_sg U5747 ( .A(n22756), .B(n50801), .X(n9544) );
  nand_x8_sg U5754 ( .A(n22628), .B(n22629), .X(n22491) );
  nand_x8_sg U5984 ( .A(n22750), .B(n50753), .X(n9592) );
  nand_x8_sg U5991 ( .A(n22631), .B(n22632), .X(n22485) );
  nand_x8_sg U6217 ( .A(n22744), .B(n50706), .X(n9640) );
  nand_x8_sg U6224 ( .A(n22634), .B(n22635), .X(n22479) );
  nand_x8_sg U6454 ( .A(n22738), .B(n50659), .X(n9688) );
  nand_x8_sg U6461 ( .A(n22637), .B(n22638), .X(n22473) );
  nand_x8_sg U6688 ( .A(n22732), .B(n50611), .X(n9735) );
  nand_x8_sg U6695 ( .A(n22640), .B(n22641), .X(n22467) );
  nand_x8_sg U6924 ( .A(n22726), .B(n50562), .X(n9783) );
  nand_x8_sg U6931 ( .A(n22643), .B(n22644), .X(n22461) );
  nand_x8_sg U7159 ( .A(n22720), .B(n50515), .X(n9831) );
  nand_x8_sg U7166 ( .A(n22646), .B(n22647), .X(n22455) );
  nand_x8_sg U7394 ( .A(n22714), .B(n50468), .X(n9879) );
  nand_x8_sg U7401 ( .A(n22649), .B(n22650), .X(n22449) );
  nand_x8_sg U7629 ( .A(n22708), .B(n50422), .X(n9927) );
  nand_x8_sg U7636 ( .A(n22652), .B(n22653), .X(n22443) );
  nand_x8_sg U7865 ( .A(n22702), .B(n50375), .X(n9975) );
  nand_x8_sg U7872 ( .A(n22655), .B(n22656), .X(n22437) );
  nand_x8_sg U8100 ( .A(n22696), .B(n50328), .X(n10024) );
  nand_x8_sg U8107 ( .A(n22658), .B(n22659), .X(n22431) );
  nand_x8_sg U8335 ( .A(n22690), .B(n50282), .X(n10072) );
  nand_x8_sg U8342 ( .A(n22661), .B(n22662), .X(n22425) );
  nand_x8_sg U8569 ( .A(n22684), .B(n50236), .X(n10121) );
  nand_x8_sg U8576 ( .A(n22664), .B(n22665), .X(n22419) );
  nand_x8_sg U8791 ( .A(n22678), .B(n50192), .X(n10170) );
  nand_x8_sg U8797 ( .A(n22667), .B(n22668), .X(n22413) );
  nand_x8_sg U8964 ( .A(n22671), .B(n22672), .X(n10213) );
  nand_x8_sg U9066 ( .A(n50121), .B(n22670), .X(n10257) );
  nor_x2_sg U4770 ( .A(n22587), .B(n8623), .X(n22585) );
  nor_x2_sg U4758 ( .A(n22579), .B(n8643), .X(n22577) );
  nor_x2_sg U4747 ( .A(n22572), .B(n8663), .X(n22570) );
  nand_x8_sg U29373 ( .A(n29018), .B(n55460), .X(n9415) );
  nand_x8_sg U36037 ( .A(n46195), .B(n46584), .X(n29151) );
  nor_x2_sg U4664 ( .A(n9406), .B(n21971), .X(n21970) );
  nand_x8_sg U36042 ( .A(n30163), .B(n55460), .X(n9406) );
  nor_x2_sg U4878 ( .A(n21995), .B(n8504), .X(n22191) );
  nand_x8_sg U4877 ( .A(n22193), .B(n22194), .X(n21995) );
  nand_x8_sg U5107 ( .A(n22342), .B(n50897), .X(n22169) );
  nand_x8_sg U5102 ( .A(n22353), .B(n22354), .X(n22190) );
  nor_x2_sg U5523 ( .A(n22495), .B(n50814), .X(n22494) );
  nor_x2_sg U5522 ( .A(n22497), .B(n8546), .X(n22495) );
  nand_x8_sg U5335 ( .A(n22356), .B(n22357), .X(n22340) );
  nor_x2_sg U5756 ( .A(n22489), .B(n50766), .X(n22488) );
  nor_x2_sg U5755 ( .A(n22491), .B(n8547), .X(n22489) );
  nand_x8_sg U5572 ( .A(n22359), .B(n22360), .X(n22334) );
  nor_x2_sg U5993 ( .A(n22483), .B(n50719), .X(n22482) );
  nor_x2_sg U5992 ( .A(n22485), .B(n8548), .X(n22483) );
  nand_x8_sg U5805 ( .A(n22362), .B(n22363), .X(n22328) );
  nor_x2_sg U6226 ( .A(n22477), .B(n50671), .X(n22476) );
  nor_x2_sg U6225 ( .A(n22479), .B(n8549), .X(n22477) );
  nand_x8_sg U6042 ( .A(n22365), .B(n22366), .X(n22322) );
  nor_x2_sg U6462 ( .A(n22473), .B(n8550), .X(n22471) );
  nand_x8_sg U6275 ( .A(n22368), .B(n22369), .X(n22316) );
  nor_x2_sg U6697 ( .A(n22465), .B(n50575), .X(n22464) );
  nor_x2_sg U6696 ( .A(n22467), .B(n8551), .X(n22465) );
  nand_x8_sg U6512 ( .A(n22371), .B(n22372), .X(n22310) );
  nor_x2_sg U6933 ( .A(n22459), .B(n50528), .X(n22458) );
  nor_x2_sg U6932 ( .A(n22461), .B(n8552), .X(n22459) );
  nand_x8_sg U6746 ( .A(n22374), .B(n22375), .X(n22304) );
  nor_x2_sg U7168 ( .A(n22453), .B(n50481), .X(n22452) );
  nor_x2_sg U7167 ( .A(n22455), .B(n8553), .X(n22453) );
  nand_x8_sg U6982 ( .A(n22377), .B(n22378), .X(n22298) );
  nor_x2_sg U7403 ( .A(n22447), .B(n50435), .X(n22446) );
  nor_x2_sg U7402 ( .A(n22449), .B(n8554), .X(n22447) );
  nand_x8_sg U7217 ( .A(n22380), .B(n22381), .X(n22292) );
  nor_x2_sg U7638 ( .A(n22441), .B(n50388), .X(n22440) );
  nor_x2_sg U7637 ( .A(n22443), .B(n8555), .X(n22441) );
  nand_x8_sg U7451 ( .A(n22383), .B(n22384), .X(n22286) );
  nor_x2_sg U7874 ( .A(n22435), .B(n50341), .X(n22434) );
  nor_x2_sg U7873 ( .A(n22437), .B(n8556), .X(n22435) );
  nand_x8_sg U7686 ( .A(n22386), .B(n22387), .X(n22280) );
  nor_x2_sg U8109 ( .A(n22429), .B(n50295), .X(n22428) );
  nor_x2_sg U8108 ( .A(n22431), .B(n8557), .X(n22429) );
  nand_x8_sg U7922 ( .A(n22389), .B(n22390), .X(n22274) );
  nor_x2_sg U8344 ( .A(n22423), .B(n50249), .X(n22422) );
  nor_x2_sg U8343 ( .A(n22425), .B(n8558), .X(n22423) );
  nand_x8_sg U8157 ( .A(n22392), .B(n22393), .X(n22268) );
  nor_x2_sg U8578 ( .A(n22417), .B(n50205), .X(n22416) );
  nor_x2_sg U8577 ( .A(n22419), .B(n8559), .X(n22417) );
  nand_x8_sg U8392 ( .A(n22395), .B(n22396), .X(n22262) );
  nor_x2_sg U8799 ( .A(n22411), .B(n50160), .X(n22410) );
  nor_x2_sg U8798 ( .A(n22413), .B(n8560), .X(n22411) );
  nand_x8_sg U8625 ( .A(n22398), .B(n22399), .X(n22256) );
  nand_x8_sg U9069 ( .A(n50122), .B(n22401), .X(n10279) );
  nor_x2_sg U5286 ( .A(n22348), .B(n50858), .X(n22347) );
  nor_x2_sg U5285 ( .A(n22350), .B(n8545), .X(n22348) );
  nand_x8_sg U5114 ( .A(n22196), .B(n22197), .X(n22172) );
  nand_x8_sg U5347 ( .A(n22199), .B(n22200), .X(n22165) );
  nand_x8_sg U5584 ( .A(n22202), .B(n22203), .X(n22158) );
  nand_x8_sg U5817 ( .A(n22205), .B(n22206), .X(n22151) );
  nand_x8_sg U6054 ( .A(n22208), .B(n22209), .X(n22144) );
  nand_x8_sg U6287 ( .A(n22211), .B(n22212), .X(n22137) );
  nand_x8_sg U6524 ( .A(n22214), .B(n22215), .X(n22130) );
  nand_x8_sg U6758 ( .A(n22217), .B(n22218), .X(n22123) );
  nand_x8_sg U6994 ( .A(n22220), .B(n22221), .X(n22116) );
  nand_x8_sg U7229 ( .A(n22223), .B(n22224), .X(n22109) );
  nand_x8_sg U7463 ( .A(n22226), .B(n22227), .X(n22102) );
  nand_x8_sg U7698 ( .A(n22229), .B(n22230), .X(n22095) );
  nand_x8_sg U7934 ( .A(n22232), .B(n22233), .X(n22088) );
  nand_x8_sg U8169 ( .A(n22235), .B(n22236), .X(n22081) );
  nand_x8_sg U8404 ( .A(n22238), .B(n22239), .X(n22074) );
  nand_x8_sg U8636 ( .A(n22241), .B(n22242), .X(n22067) );
  nand_x8_sg U9072 ( .A(n50123), .B(n22244), .X(n10280) );
  nand_x8_sg U4863 ( .A(n22187), .B(n22188), .X(n21988) );
  nor_x2_sg U5053 ( .A(n22182), .B(n50906), .X(n22181) );
  nor_x2_sg U5052 ( .A(n22184), .B(n8544), .X(n22182) );
  nand_x8_sg U4887 ( .A(n22002), .B(n22003), .X(n9412) );
  nor_x2_sg U5115 ( .A(n22172), .B(n8505), .X(n22170) );
  nand_x8_sg U5124 ( .A(n22005), .B(n22006), .X(n9462) );
  nor_x2_sg U5348 ( .A(n22165), .B(n8506), .X(n22163) );
  nand_x8_sg U5357 ( .A(n22008), .B(n22009), .X(n9511) );
  nor_x2_sg U5585 ( .A(n22158), .B(n8507), .X(n22156) );
  nand_x8_sg U5594 ( .A(n22011), .B(n22012), .X(n9560) );
  nor_x2_sg U5818 ( .A(n22151), .B(n8508), .X(n22149) );
  nand_x8_sg U5827 ( .A(n22014), .B(n22015), .X(n9608) );
  nor_x2_sg U6055 ( .A(n22144), .B(n8509), .X(n22142) );
  nand_x8_sg U6064 ( .A(n22017), .B(n22018), .X(n9656) );
  nor_x2_sg U6288 ( .A(n22137), .B(n8510), .X(n22135) );
  nand_x8_sg U6297 ( .A(n22020), .B(n22021), .X(n9703) );
  nor_x2_sg U6525 ( .A(n22130), .B(n8511), .X(n22128) );
  nand_x8_sg U6534 ( .A(n22023), .B(n22024), .X(n9751) );
  nor_x2_sg U6759 ( .A(n22123), .B(n8512), .X(n22121) );
  nand_x8_sg U6768 ( .A(n22026), .B(n22027), .X(n9799) );
  nor_x2_sg U6995 ( .A(n22116), .B(n8513), .X(n22114) );
  nand_x8_sg U7004 ( .A(n22029), .B(n22030), .X(n9847) );
  nor_x2_sg U7230 ( .A(n22109), .B(n8514), .X(n22107) );
  nand_x8_sg U7239 ( .A(n22032), .B(n22033), .X(n9895) );
  nor_x2_sg U7464 ( .A(n22102), .B(n8515), .X(n22100) );
  nand_x8_sg U7473 ( .A(n22035), .B(n22036), .X(n9943) );
  nor_x2_sg U7699 ( .A(n22095), .B(n8516), .X(n22093) );
  nand_x8_sg U7708 ( .A(n22038), .B(n22039), .X(n9992) );
  nor_x2_sg U7935 ( .A(n22088), .B(n8517), .X(n22086) );
  nand_x8_sg U7944 ( .A(n22041), .B(n22042), .X(n10040) );
  nor_x2_sg U8170 ( .A(n22081), .B(n8518), .X(n22079) );
  nand_x8_sg U8179 ( .A(n22044), .B(n22045), .X(n10089) );
  nor_x2_sg U8405 ( .A(n22074), .B(n8519), .X(n22072) );
  nand_x8_sg U8414 ( .A(n22047), .B(n22048), .X(n10138) );
  nor_x2_sg U8637 ( .A(n22067), .B(n8520), .X(n22065) );
  nand_x8_sg U8645 ( .A(n22050), .B(n22051), .X(n10185) );
  nand_x8_sg U9006 ( .A(n50124), .B(n22053), .X(n10264) );
  nand_x8_sg U32366 ( .A(n26078), .B(n29633), .X(n15726) );
  nand_x8_sg U29343 ( .A(n29619), .B(n29617), .X(n9394) );
  nor_x2_sg U4616 ( .A(n9392), .B(n21958), .X(n21957) );
  nand_x8_sg U29338 ( .A(n29616), .B(n46582), .X(n9392) );
  nand_x8_sg U29335 ( .A(n55462), .B(n27900), .X(n10256) );
  nand_x8_sg U29332 ( .A(n55465), .B(n46584), .X(n9385) );
  nand_x8_sg U29429 ( .A(n29603), .B(n55460), .X(n10281) );
  nor_x2_sg U4606 ( .A(n9365), .B(n21941), .X(n21938) );
  nand_x8_sg U29326 ( .A(n29595), .B(n55469), .X(n9365) );
  nor_x2_sg U4605 ( .A(n9371), .B(n21940), .X(n21939) );
  nand_x8_sg U29323 ( .A(n15726), .B(n29589), .X(n9371) );
  nand_x8_sg U29320 ( .A(n55470), .B(n26078), .X(n9367) );
  nand_x8_sg U29318 ( .A(n29587), .B(n55468), .X(n9373) );
  nor_x2_sg U29317 ( .A(n46582), .B(n46608), .X(n29587) );
  nor_x2_sg U4600 ( .A(n21928), .B(n21929), .X(n21927) );
  nand_x8_sg U9194 ( .A(n46580), .B(n46577), .X(n9355) );
  nor_x2_sg U4893 ( .A(n9406), .B(n9407), .X(n9405) );
  nor_x2_sg U4844 ( .A(n9391), .B(n9392), .X(n9390) );
  nor_x2_sg U4833 ( .A(n9370), .B(n9371), .X(n9369) );
  nor_x2_sg U4830 ( .A(n9364), .B(n9365), .X(n9363) );
  nor_x2_sg U4828 ( .A(n9356), .B(n9357), .X(n9354) );
  nor_x2_sg U5130 ( .A(n9406), .B(n9457), .X(n9456) );
  nor_x2_sg U5080 ( .A(n9392), .B(n9446), .X(n9445) );
  nor_x2_sg U5069 ( .A(n9429), .B(n9371), .X(n9428) );
  nor_x2_sg U5066 ( .A(n9365), .B(n9425), .X(n9424) );
  nor_x2_sg U5064 ( .A(n9417), .B(n9418), .X(n9416) );
  nor_x2_sg U5363 ( .A(n9406), .B(n9506), .X(n9505) );
  nor_x2_sg U5313 ( .A(n9392), .B(n9495), .X(n9494) );
  nor_x2_sg U5302 ( .A(n9478), .B(n9371), .X(n9477) );
  nor_x2_sg U5299 ( .A(n9365), .B(n9474), .X(n9473) );
  nor_x2_sg U5297 ( .A(n9466), .B(n9467), .X(n9465) );
  nor_x2_sg U5600 ( .A(n9406), .B(n9555), .X(n9554) );
  nor_x2_sg U5550 ( .A(n9392), .B(n9544), .X(n9543) );
  nor_x2_sg U5539 ( .A(n9527), .B(n9371), .X(n9526) );
  nor_x2_sg U5536 ( .A(n9365), .B(n9523), .X(n9522) );
  nor_x2_sg U5534 ( .A(n9515), .B(n9516), .X(n9514) );
  nor_x2_sg U5833 ( .A(n9406), .B(n9603), .X(n9602) );
  nor_x2_sg U5783 ( .A(n9392), .B(n9592), .X(n9591) );
  nor_x2_sg U5772 ( .A(n9576), .B(n9371), .X(n9575) );
  nor_x2_sg U5769 ( .A(n9365), .B(n9572), .X(n9571) );
  nor_x2_sg U5767 ( .A(n9564), .B(n9565), .X(n9563) );
  nor_x2_sg U6070 ( .A(n9406), .B(n9651), .X(n9650) );
  nor_x2_sg U6020 ( .A(n9392), .B(n9640), .X(n9639) );
  nor_x2_sg U6009 ( .A(n9624), .B(n9371), .X(n9623) );
  nor_x2_sg U6006 ( .A(n9365), .B(n9620), .X(n9619) );
  nor_x2_sg U6004 ( .A(n9612), .B(n9613), .X(n9611) );
  nor_x2_sg U6303 ( .A(n9406), .B(n9698), .X(n9697) );
  nor_x2_sg U6253 ( .A(n9392), .B(n9688), .X(n9687) );
  nor_x2_sg U6242 ( .A(n9672), .B(n9371), .X(n9671) );
  nor_x2_sg U6239 ( .A(n9365), .B(n9668), .X(n9667) );
  nor_x2_sg U6237 ( .A(n9660), .B(n9661), .X(n9659) );
  nor_x2_sg U6540 ( .A(n9406), .B(n9746), .X(n9745) );
  nor_x2_sg U6490 ( .A(n9392), .B(n9735), .X(n9734) );
  nor_x2_sg U6479 ( .A(n9719), .B(n9371), .X(n9718) );
  nor_x2_sg U6476 ( .A(n9365), .B(n9715), .X(n9714) );
  nor_x2_sg U6474 ( .A(n9707), .B(n9708), .X(n9706) );
  nor_x2_sg U6774 ( .A(n9406), .B(n9794), .X(n9793) );
  nor_x2_sg U6724 ( .A(n9392), .B(n9783), .X(n9782) );
  nor_x2_sg U6713 ( .A(n9767), .B(n9371), .X(n9766) );
  nor_x2_sg U6710 ( .A(n9365), .B(n9763), .X(n9762) );
  nor_x2_sg U6708 ( .A(n9755), .B(n9756), .X(n9754) );
  nor_x2_sg U7010 ( .A(n9406), .B(n9842), .X(n9841) );
  nor_x2_sg U6960 ( .A(n9392), .B(n9831), .X(n9830) );
  nor_x2_sg U6949 ( .A(n9815), .B(n9371), .X(n9814) );
  nor_x2_sg U6946 ( .A(n9365), .B(n9811), .X(n9810) );
  nor_x2_sg U6944 ( .A(n9803), .B(n9804), .X(n9802) );
  nor_x2_sg U7245 ( .A(n9406), .B(n9890), .X(n9889) );
  nor_x2_sg U7195 ( .A(n9392), .B(n9879), .X(n9878) );
  nor_x2_sg U7184 ( .A(n9863), .B(n9371), .X(n9862) );
  nor_x2_sg U7181 ( .A(n9365), .B(n9859), .X(n9858) );
  nor_x2_sg U7179 ( .A(n9851), .B(n9852), .X(n9850) );
  nor_x2_sg U7479 ( .A(n9406), .B(n9938), .X(n9937) );
  nor_x2_sg U7430 ( .A(n9392), .B(n9927), .X(n9926) );
  nor_x2_sg U7419 ( .A(n9911), .B(n9371), .X(n9910) );
  nor_x2_sg U7416 ( .A(n9365), .B(n9907), .X(n9906) );
  nor_x2_sg U7414 ( .A(n9899), .B(n9900), .X(n9898) );
  nor_x2_sg U7714 ( .A(n9406), .B(n9987), .X(n9986) );
  nor_x2_sg U7665 ( .A(n9392), .B(n9975), .X(n9974) );
  nor_x2_sg U7654 ( .A(n9959), .B(n9371), .X(n9958) );
  nor_x2_sg U7651 ( .A(n9365), .B(n9955), .X(n9954) );
  nor_x2_sg U7649 ( .A(n9947), .B(n9948), .X(n9946) );
  nor_x2_sg U7950 ( .A(n9406), .B(n10035), .X(n10034) );
  nor_x2_sg U7901 ( .A(n9392), .B(n10024), .X(n10023) );
  nor_x2_sg U7890 ( .A(n10008), .B(n9371), .X(n10007) );
  nor_x2_sg U7887 ( .A(n9365), .B(n10004), .X(n10003) );
  nor_x2_sg U7885 ( .A(n9996), .B(n9997), .X(n9995) );
  nor_x2_sg U8185 ( .A(n9406), .B(n10084), .X(n10083) );
  nor_x2_sg U8136 ( .A(n9392), .B(n10072), .X(n10071) );
  nor_x2_sg U8125 ( .A(n10056), .B(n9371), .X(n10055) );
  nor_x2_sg U8122 ( .A(n9365), .B(n10052), .X(n10051) );
  nor_x2_sg U8120 ( .A(n10044), .B(n10045), .X(n10043) );
  nor_x2_sg U8420 ( .A(n9406), .B(n10133), .X(n10132) );
  nor_x2_sg U8371 ( .A(n9392), .B(n10121), .X(n10120) );
  nor_x2_sg U8360 ( .A(n10105), .B(n9371), .X(n10104) );
  nor_x2_sg U8357 ( .A(n9365), .B(n10101), .X(n10100) );
  nor_x2_sg U8355 ( .A(n10093), .B(n10094), .X(n10092) );
  nor_x2_sg U8651 ( .A(n9406), .B(n10180), .X(n10179) );
  nor_x2_sg U8605 ( .A(n9392), .B(n10170), .X(n10169) );
  nor_x2_sg U8594 ( .A(n10154), .B(n9371), .X(n10153) );
  nor_x2_sg U8591 ( .A(n9365), .B(n10150), .X(n10149) );
  nor_x2_sg U8589 ( .A(n10142), .B(n10143), .X(n10141) );
  nor_x2_sg U8863 ( .A(n9406), .B(n10223), .X(n10222) );
  nor_x2_sg U8826 ( .A(n9392), .B(n10213), .X(n10212) );
  nor_x2_sg U8815 ( .A(n10200), .B(n9371), .X(n10199) );
  nor_x2_sg U8812 ( .A(n9365), .B(n10197), .X(n10196) );
  nor_x2_sg U8810 ( .A(n10189), .B(n10190), .X(n10188) );
  nor_x2_sg U9073 ( .A(n10280), .B(n10281), .X(n10277) );
  nor_x2_sg U9019 ( .A(n10279), .B(n9415), .X(n10278) );
  nor_x2_sg U9008 ( .A(n9406), .B(n10267), .X(n10261) );
  nor_x2_sg U8994 ( .A(n9392), .B(n10257), .X(n10253) );
  nor_x2_sg U8993 ( .A(n10255), .B(n10256), .X(n10254) );
  nor_x2_sg U8987 ( .A(n10245), .B(n9373), .X(n10242) );
  nor_x2_sg U8986 ( .A(n10244), .B(n9371), .X(n10243) );
  nor_x2_sg U8984 ( .A(n9367), .B(n10241), .X(n10238) );
  nor_x2_sg U8983 ( .A(n9365), .B(n10240), .X(n10239) );
  nor_x2_sg U8981 ( .A(n10232), .B(n10233), .X(n10231) );
  nand_x8_sg U29442 ( .A(n46572), .B(n46574), .X(n10283) );
  nor_x2_sg U29708 ( .A(n51260), .B(n25599), .X(n25598) );
  nor_x2_sg U29695 ( .A(n25589), .B(n25590), .X(n25587) );
  nor_x2_sg U9258 ( .A(n46567), .B(n51281), .X(n10419) );
  nor_x2_sg U29687 ( .A(n25583), .B(n25584), .X(n25581) );
  nor_x2_sg U9255 ( .A(n10421), .B(n46568), .X(n10420) );
  nand_x8_sg U9695 ( .A(n51280), .B(n46572), .X(n10442) );
  nand_x8_sg U29681 ( .A(n25573), .B(n51292), .X(n10518) );
  nand_x8_sg U29831 ( .A(n25649), .B(n25650), .X(n25576) );
  nor_x2_sg U9347 ( .A(n46565), .B(n46568), .X(n10492) );
  nor_x2_sg U9344 ( .A(n46573), .B(n46561), .X(n10489) );
  nor_x2_sg U9340 ( .A(n10480), .B(n10481), .X(n10479) );
  nand_x8_sg U9450 ( .A(n51280), .B(n46564), .X(n10493) );
  nor_x2_sg U9351 ( .A(n46567), .B(n10458), .X(n10485) );
  nand_x8_sg U9844 ( .A(n46558), .B(n46572), .X(n10545) );
  nand_x8_sg U9454 ( .A(n10573), .B(n10574), .X(n10521) );
  nand_x8_sg U10098 ( .A(n51334), .B(n46574), .X(n10522) );
  nand_x8_sg U29658 ( .A(n25555), .B(n51333), .X(n10655) );
  nor_x2_sg U9429 ( .A(n41788), .B(n43221), .X(n10531) );
  nand_x8_sg U29847 ( .A(n25560), .B(n25641), .X(n25551) );
  nor_x2_sg U9409 ( .A(n10537), .B(n10493), .X(n10536) );
  nor_x2_sg U9406 ( .A(n10324), .B(n41740), .X(n10330) );
  nor_x2_sg U9438 ( .A(n43205), .B(n10529), .X(n10329) );
  nand_x8_sg U29647 ( .A(n25545), .B(n51376), .X(n10660) );
  nor_x2_sg U9503 ( .A(n10604), .B(n51384), .X(n10603) );
  nor_x2_sg U9584 ( .A(n10661), .B(n51399), .X(n10643) );
  nor_x2_sg U9553 ( .A(n10645), .B(n10646), .X(n10644) );
  nor_x2_sg U9441 ( .A(n10558), .B(n10559), .X(n10557) );
  nor_x2_sg U9638 ( .A(n43317), .B(n10704), .X(n10685) );
  nand_x8_sg U29636 ( .A(n25533), .B(n51417), .X(n10782) );
  nor_x2_sg U9603 ( .A(n10678), .B(n10679), .X(n10677) );
  nand_x8_sg U29631 ( .A(n25527), .B(n51434), .X(n10843) );
  nor_x2_sg U9706 ( .A(n10749), .B(n10750), .X(n10748) );
  nand_x8_sg U10023 ( .A(n51435), .B(n46572), .X(n10856) );
  nor_x2_sg U9831 ( .A(n10846), .B(n10847), .X(n10835) );
  nand_x8_sg U29625 ( .A(n25521), .B(n51457), .X(n10923) );
  nand_x8_sg U10071 ( .A(n51293), .B(n51334), .X(n10849) );
  nor_x2_sg U9828 ( .A(n10848), .B(n10849), .X(n10847) );
  nor_x2_sg U10043 ( .A(n46555), .B(n46565), .X(n11018) );
  nand_x8_sg U29756 ( .A(n25614), .B(n51480), .X(n10919) );
  nor_x2_sg U10072 ( .A(n10849), .B(n51464), .X(n11025) );
  nor_x2_sg U10054 ( .A(n11027), .B(n11028), .X(n11026) );
  nor_x2_sg U9729 ( .A(n10768), .B(n10769), .X(n10767) );
  nand_x8_sg U10031 ( .A(n51458), .B(n46572), .X(n10994) );
  nand_x8_sg U10029 ( .A(n51306), .B(n51334), .X(n10993) );
  nor_x2_sg U10028 ( .A(n10993), .B(n51459), .X(n11013) );
  nor_x2_sg U9881 ( .A(n51490), .B(n10884), .X(n10881) );
  nor_x2_sg U10039 ( .A(n43355), .B(n42056), .X(n10973) );
  nor_x2_sg U9995 ( .A(n10993), .B(n10994), .X(n10989) );
  nor_x2_sg U9994 ( .A(n46555), .B(n10991), .X(n10990) );
  nor_x2_sg U10106 ( .A(n51334), .B(n51503), .X(n11041) );
  nand_x8_sg U29875 ( .A(n25619), .B(n25634), .X(n25610) );
  nor_x2_sg U10101 ( .A(n11043), .B(n10655), .X(n11042) );
  nor_x2_sg U9862 ( .A(n10869), .B(n51431), .X(n10868) );
  nor_x2_sg U9970 ( .A(n10932), .B(n51484), .X(n10929) );
  nor_x2_sg U9965 ( .A(n10957), .B(n46559), .X(n10953) );
  nor_x2_sg U9956 ( .A(n10955), .B(n10956), .X(n10954) );
  nor_x2_sg U9934 ( .A(n10931), .B(n51502), .X(n10930) );
  nor_x2_sg U9927 ( .A(n10913), .B(n51482), .X(n10910) );
  nor_x2_sg U9913 ( .A(n10912), .B(n51475), .X(n10911) );
  nor_x2_sg U9896 ( .A(n46555), .B(n10518), .X(n10900) );
  nand_x8_sg U11194 ( .A(n46553), .B(n46579), .X(n8860) );
  nand_x8_sg U29900 ( .A(n46547), .B(n46551), .X(n11051) );
  nor_x2_sg U10143 ( .A(n11051), .B(n51538), .X(n11052) );
  nand_x8_sg U10273 ( .A(n51537), .B(n46551), .X(n11054) );
  nor_x2_sg U30166 ( .A(n51536), .B(n25880), .X(n25879) );
  nand_x8_sg U30289 ( .A(n25931), .B(n25932), .X(n25862) );
  nor_x2_sg U30140 ( .A(n25861), .B(n25862), .X(n25860) );
  nor_x2_sg U10296 ( .A(n11183), .B(n51563), .X(n11182) );
  nand_x8_sg U30291 ( .A(n25928), .B(n25929), .X(n25857) );
  nor_x2_sg U10354 ( .A(n11219), .B(n51590), .X(n11205) );
  nand_x8_sg U10413 ( .A(n46539), .B(n51537), .X(n11238) );
  nand_x8_sg U10410 ( .A(n11262), .B(n11263), .X(n11231) );
  nand_x8_sg U30293 ( .A(n25925), .B(n25926), .X(n25850) );
  nor_x2_sg U10401 ( .A(n11256), .B(n11257), .X(n11255) );
  nor_x2_sg U10396 ( .A(n11238), .B(n11254), .X(n11253) );
  nor_x2_sg U10411 ( .A(n51543), .B(n11231), .X(n11261) );
  nor_x2_sg U10437 ( .A(n51607), .B(n51560), .X(n11279) );
  nor_x2_sg U10432 ( .A(n46539), .B(n11281), .X(n11280) );
  nand_x8_sg U10510 ( .A(n46536), .B(n51543), .X(n11344) );
  nand_x8_sg U30114 ( .A(n25836), .B(n51614), .X(n11434) );
  nand_x8_sg U30109 ( .A(n25830), .B(n51629), .X(n11394) );
  nand_x8_sg U11133 ( .A(n51598), .B(n11265), .X(n11810) );
  nor_x2_sg U10515 ( .A(n11339), .B(n11350), .X(n11349) );
  nor_x2_sg U10505 ( .A(n11343), .B(n11344), .X(n11342) );
  nand_x8_sg U30103 ( .A(n25824), .B(n51649), .X(n11438) );
  nand_x8_sg U30098 ( .A(n25818), .B(n51670), .X(n11515) );
  nor_x2_sg U10613 ( .A(n11425), .B(n11426), .X(n11424) );
  nor_x2_sg U10502 ( .A(n11331), .B(n11332), .X(n11330) );
  nor_x2_sg U10703 ( .A(n51697), .B(n11478), .X(n11414) );
  nand_x8_sg U30092 ( .A(n25812), .B(n51692), .X(n11638) );
  nor_x2_sg U10805 ( .A(n11559), .B(n11560), .X(n11488) );
  nand_x8_sg U30087 ( .A(n25806), .B(n51716), .X(n11623) );
  nor_x2_sg U10665 ( .A(n11459), .B(n11460), .X(n11458) );
  nor_x2_sg U10850 ( .A(n51709), .B(n51642), .X(n11579) );
  nor_x2_sg U10829 ( .A(n11581), .B(n11582), .X(n11580) );
  nor_x2_sg U10896 ( .A(n51745), .B(n11626), .X(n11615) );
  nand_x8_sg U30081 ( .A(n25800), .B(n51737), .X(n11768) );
  nor_x2_sg U10893 ( .A(n11627), .B(n11628), .X(n11626) );
  nor_x2_sg U10890 ( .A(n11622), .B(n11623), .X(n11616) );
  nor_x2_sg U10875 ( .A(n11618), .B(n11619), .X(n11617) );
  nor_x2_sg U10784 ( .A(n11541), .B(n51773), .X(n11497) );
  nor_x2_sg U11152 ( .A(n11817), .B(n51765), .X(n11808) );
  nand_x8_sg U30214 ( .A(n25895), .B(n51760), .X(n11703) );
  nor_x2_sg U11122 ( .A(n11810), .B(n11811), .X(n11809) );
  nor_x2_sg U10794 ( .A(n11554), .B(n11555), .X(n11553) );
  nand_x8_sg U11095 ( .A(n11636), .B(n51726), .X(n11786) );
  nor_x2_sg U11091 ( .A(n11787), .B(n11786), .X(n11794) );
  nor_x2_sg U11079 ( .A(n11790), .B(n11791), .X(n11789) );
  nand_x8_sg U10948 ( .A(n11129), .B(n51788), .X(n11138) );
  nor_x2_sg U10945 ( .A(n51769), .B(n11664), .X(n11661) );
  nor_x2_sg U11107 ( .A(n43357), .B(n11785), .X(n11757) );
  nor_x2_sg U11078 ( .A(n11786), .B(n51741), .X(n11785) );
  nor_x2_sg U11063 ( .A(n11777), .B(n11778), .X(n11774) );
  nor_x2_sg U11062 ( .A(n11515), .B(n41161), .X(n11775) );
  nor_x2_sg U11060 ( .A(n11776), .B(n46541), .X(n11767) );
  nand_x8_sg U11168 ( .A(n51738), .B(n51537), .X(n11681) );
  nor_x2_sg U11177 ( .A(n46532), .B(n51783), .X(n11825) );
  nand_x8_sg U30333 ( .A(n25900), .B(n25913), .X(n25891) );
  nor_x2_sg U11172 ( .A(n11827), .B(n11434), .X(n11826) );
  nor_x2_sg U10926 ( .A(n11649), .B(n51712), .X(n11648) );
  nor_x2_sg U10788 ( .A(n11547), .B(n11138), .X(n11546) );
  nor_x2_sg U11181 ( .A(n11747), .B(n51771), .X(n11744) );
  nor_x2_sg U11040 ( .A(n11746), .B(n51793), .X(n11745) );
  nor_x2_sg U11031 ( .A(n11739), .B(n46535), .X(n11737) );
  nor_x2_sg U10970 ( .A(n11691), .B(n43091), .X(n11688) );
  nand_x8_sg U30337 ( .A(n25894), .B(n25912), .X(n11693) );
  nor_x2_sg U10959 ( .A(n46537), .B(n11515), .X(n11680) );
  nand_x8_sg U12253 ( .A(n46531), .B(n46579), .X(n8898) );
  nand_x8_sg U30354 ( .A(n46525), .B(n46529), .X(n11834) );
  nor_x2_sg U30627 ( .A(n51818), .B(n26160), .X(n26159) );
  nor_x2_sg U30614 ( .A(n26150), .B(n26151), .X(n26148) );
  nor_x2_sg U30606 ( .A(n26144), .B(n26145), .X(n26142) );
  nor_x2_sg U11355 ( .A(n11961), .B(n51841), .X(n11960) );
  nand_x8_sg U11436 ( .A(n46517), .B(n51819), .X(n11995) );
  nand_x8_sg U30600 ( .A(n26134), .B(n51853), .X(n12030) );
  nand_x8_sg U30750 ( .A(n26208), .B(n26209), .X(n26137) );
  nor_x2_sg U11414 ( .A(n51870), .B(n11996), .X(n11983) );
  nor_x2_sg U11469 ( .A(n46518), .B(n46521), .X(n12045) );
  nor_x2_sg U11466 ( .A(n46528), .B(n46514), .X(n12042) );
  nor_x2_sg U11462 ( .A(n12033), .B(n12034), .X(n12032) );
  nor_x2_sg U11473 ( .A(n51826), .B(n12008), .X(n12038) );
  nor_x2_sg U11499 ( .A(n51888), .B(n46516), .X(n12058) );
  nor_x2_sg U11494 ( .A(n51839), .B(n12060), .X(n12059) );
  nand_x8_sg U11572 ( .A(n51826), .B(n51854), .X(n12124) );
  nand_x8_sg U30577 ( .A(n26116), .B(n51895), .X(n12214) );
  nand_x8_sg U30572 ( .A(n26110), .B(n51910), .X(n12174) );
  nor_x2_sg U11577 ( .A(n12119), .B(n12130), .X(n12129) );
  nor_x2_sg U11567 ( .A(n12123), .B(n12124), .X(n12122) );
  nand_x8_sg U30566 ( .A(n26104), .B(n51930), .X(n12218) );
  nand_x8_sg U30561 ( .A(n26098), .B(n51951), .X(n12295) );
  nor_x2_sg U11675 ( .A(n12205), .B(n12206), .X(n12204) );
  nor_x2_sg U11564 ( .A(n12111), .B(n12112), .X(n12110) );
  nor_x2_sg U11761 ( .A(n43313), .B(n12265), .X(n12246) );
  nand_x8_sg U30555 ( .A(n26092), .B(n51973), .X(n12344) );
  nor_x2_sg U11888 ( .A(n51965), .B(n12345), .X(n12269) );
  nand_x8_sg U30550 ( .A(n26086), .B(n51994), .X(n12404) );
  nor_x2_sg U11727 ( .A(n12239), .B(n12240), .X(n12238) );
  nor_x2_sg U11892 ( .A(n12361), .B(n12362), .X(n12360) );
  nor_x2_sg U11958 ( .A(n12407), .B(n12408), .X(n12396) );
  nor_x2_sg U30540 ( .A(n26082), .B(n26083), .X(n12602) );
  nand_x8_sg U12191 ( .A(n51896), .B(n51854), .X(n12410) );
  nor_x2_sg U11955 ( .A(n12409), .B(n12410), .X(n12408) );
  nor_x2_sg U11952 ( .A(n12403), .B(n12404), .X(n12397) );
  nor_x2_sg U11937 ( .A(n12399), .B(n12400), .X(n12398) );
  nor_x2_sg U11845 ( .A(n12321), .B(n52053), .X(n12277) );
  nor_x2_sg U12205 ( .A(n12592), .B(n52045), .X(n12583) );
  nand_x8_sg U30675 ( .A(n26175), .B(n52041), .X(n12482) );
  nor_x2_sg U12192 ( .A(n12410), .B(n52026), .X(n12584) );
  nor_x2_sg U11855 ( .A(n12334), .B(n12335), .X(n12333) );
  nor_x2_sg U11964 ( .A(n52024), .B(n12411), .X(n12331) );
  nor_x2_sg U12159 ( .A(n12422), .B(n41768), .X(n12419) );
  nor_x2_sg U12133 ( .A(n12560), .B(n12561), .X(n12559) );
  nand_x8_sg U12010 ( .A(n11912), .B(n52067), .X(n11921) );
  nand_x8_sg U30794 ( .A(n26180), .B(n26193), .X(n26171) );
  nor_x2_sg U11989 ( .A(n12429), .B(n51991), .X(n12428) );
  nor_x2_sg U11849 ( .A(n12327), .B(n11921), .X(n12326) );
  nor_x2_sg U12014 ( .A(n42347), .B(n52055), .X(n11899) );
  nor_x2_sg U12238 ( .A(n12527), .B(n52051), .X(n12524) );
  nor_x2_sg U12101 ( .A(n12526), .B(n52065), .X(n12525) );
  nor_x2_sg U12092 ( .A(n12519), .B(n12214), .X(n12517) );
  nor_x2_sg U12032 ( .A(n12470), .B(n43089), .X(n12467) );
  nand_x8_sg U30798 ( .A(n26174), .B(n26192), .X(n12472) );
  nor_x2_sg U12021 ( .A(n12030), .B(n12295), .X(n12459) );
  nand_x8_sg U13312 ( .A(n46510), .B(n46579), .X(n8822) );
  nand_x8_sg U30815 ( .A(n46503), .B(n46507), .X(n12612) );
  nor_x2_sg U12265 ( .A(n12612), .B(n52095), .X(n12613) );
  nand_x8_sg U12395 ( .A(n46500), .B(n46507), .X(n12615) );
  nor_x2_sg U31085 ( .A(n52094), .B(n26439), .X(n26438) );
  nand_x8_sg U31208 ( .A(n26490), .B(n26491), .X(n26421) );
  nor_x2_sg U31059 ( .A(n26420), .B(n26421), .X(n26419) );
  nor_x2_sg U12418 ( .A(n12744), .B(n52120), .X(n12743) );
  nand_x8_sg U31210 ( .A(n26487), .B(n26488), .X(n26416) );
  nor_x2_sg U12476 ( .A(n12780), .B(n52148), .X(n12766) );
  nand_x8_sg U12535 ( .A(n46495), .B(n46500), .X(n12799) );
  nand_x8_sg U12532 ( .A(n12823), .B(n12824), .X(n12792) );
  nand_x8_sg U31212 ( .A(n26484), .B(n26485), .X(n26409) );
  nor_x2_sg U12523 ( .A(n12817), .B(n12818), .X(n12816) );
  nor_x2_sg U12518 ( .A(n12799), .B(n12815), .X(n12814) );
  nor_x2_sg U12533 ( .A(n52100), .B(n12792), .X(n12822) );
  nor_x2_sg U12559 ( .A(n52165), .B(n52117), .X(n12840) );
  nor_x2_sg U12554 ( .A(n46495), .B(n12842), .X(n12841) );
  nand_x8_sg U12632 ( .A(n52133), .B(n52100), .X(n12905) );
  nand_x8_sg U31033 ( .A(n26395), .B(n52172), .X(n12995) );
  nor_x2_sg U12612 ( .A(n12875), .B(n12874), .X(n12869) );
  nand_x8_sg U31028 ( .A(n26389), .B(n52186), .X(n12955) );
  nor_x2_sg U12637 ( .A(n12900), .B(n12911), .X(n12910) );
  nor_x2_sg U12627 ( .A(n12904), .B(n12905), .X(n12903) );
  nand_x8_sg U31022 ( .A(n26383), .B(n52205), .X(n12999) );
  nand_x8_sg U31017 ( .A(n26377), .B(n52226), .X(n13076) );
  nor_x2_sg U12734 ( .A(n12986), .B(n12987), .X(n12985) );
  nor_x2_sg U12624 ( .A(n12892), .B(n12893), .X(n12891) );
  nor_x2_sg U12824 ( .A(n52253), .B(n13039), .X(n12975) );
  nand_x8_sg U31011 ( .A(n26371), .B(n52248), .X(n13200) );
  nor_x2_sg U12926 ( .A(n13120), .B(n13121), .X(n13049) );
  nand_x8_sg U31006 ( .A(n26365), .B(n52270), .X(n13184) );
  nor_x2_sg U12786 ( .A(n13020), .B(n13021), .X(n13019) );
  nor_x2_sg U12973 ( .A(n52265), .B(n52198), .X(n13140) );
  nor_x2_sg U12952 ( .A(n13142), .B(n13143), .X(n13141) );
  nor_x2_sg U13019 ( .A(n52302), .B(n13187), .X(n13176) );
  nor_x2_sg U30996 ( .A(n26361), .B(n26362), .X(n13384) );
  nor_x2_sg U13016 ( .A(n13188), .B(n13189), .X(n13187) );
  nor_x2_sg U13013 ( .A(n13183), .B(n13184), .X(n13177) );
  nor_x2_sg U12998 ( .A(n13179), .B(n13180), .X(n13178) );
  nor_x2_sg U12905 ( .A(n13102), .B(n52330), .X(n13058) );
  nor_x2_sg U13265 ( .A(n13374), .B(n52321), .X(n13365) );
  nand_x8_sg U31133 ( .A(n26454), .B(n52317), .X(n13263) );
  nor_x2_sg U13235 ( .A(n13367), .B(n13368), .X(n13366) );
  nor_x2_sg U12915 ( .A(n13115), .B(n13116), .X(n13114) );
  nor_x2_sg U13025 ( .A(n13194), .B(n52287), .X(n13191) );
  nor_x2_sg U13195 ( .A(n13342), .B(n13343), .X(n13341) );
  nand_x8_sg U13072 ( .A(n12690), .B(n52344), .X(n12699) );
  nand_x8_sg U31252 ( .A(n26459), .B(n26472), .X(n26450) );
  nor_x2_sg U13051 ( .A(n13210), .B(n52268), .X(n13209) );
  nor_x2_sg U12909 ( .A(n13108), .B(n12699), .X(n13107) );
  nor_x2_sg U13298 ( .A(n13308), .B(n52328), .X(n13305) );
  nor_x2_sg U13163 ( .A(n13307), .B(n52342), .X(n13306) );
  nor_x2_sg U13154 ( .A(n13300), .B(n46491), .X(n13298) );
  nor_x2_sg U13094 ( .A(n13251), .B(n43087), .X(n13248) );
  nand_x8_sg U31256 ( .A(n26453), .B(n26471), .X(n13253) );
  nor_x2_sg U13083 ( .A(n46493), .B(n13076), .X(n13240) );
  nand_x8_sg U14370 ( .A(n46487), .B(n46579), .X(n8783) );
  nand_x8_sg U31274 ( .A(n46481), .B(n46484), .X(n13396) );
  nor_x2_sg U31545 ( .A(n52371), .B(n26717), .X(n26716) );
  nor_x2_sg U31532 ( .A(n26707), .B(n26708), .X(n26705) );
  nor_x2_sg U31524 ( .A(n26701), .B(n26702), .X(n26699) );
  nor_x2_sg U13473 ( .A(n13522), .B(n52393), .X(n13521) );
  nand_x8_sg U13554 ( .A(n46474), .B(n46478), .X(n13556) );
  nand_x8_sg U31667 ( .A(n26765), .B(n26766), .X(n26694) );
  nor_x2_sg U13532 ( .A(n52422), .B(n13557), .X(n13544) );
  nor_x2_sg U13587 ( .A(n46477), .B(n46475), .X(n13606) );
  nor_x2_sg U13584 ( .A(n46485), .B(n46469), .X(n13603) );
  nor_x2_sg U13571 ( .A(n13587), .B(n13588), .X(n13586) );
  nor_x2_sg U13591 ( .A(n52378), .B(n13569), .X(n13599) );
  nor_x2_sg U13617 ( .A(n52439), .B(n13623), .X(n13621) );
  nor_x2_sg U13613 ( .A(n52391), .B(n43170), .X(n13620) );
  nand_x8_sg U13690 ( .A(n52406), .B(n52378), .X(n13685) );
  nand_x8_sg U31495 ( .A(n26673), .B(n52446), .X(n13775) );
  nand_x8_sg U31490 ( .A(n26667), .B(n52462), .X(n13735) );
  nor_x2_sg U13662 ( .A(n46473), .B(n52438), .X(n13656) );
  nor_x2_sg U13695 ( .A(n13680), .B(n13691), .X(n13690) );
  nor_x2_sg U13685 ( .A(n13684), .B(n13685), .X(n13683) );
  nand_x8_sg U31484 ( .A(n26661), .B(n52482), .X(n13779) );
  nand_x8_sg U31479 ( .A(n26655), .B(n52503), .X(n13856) );
  nor_x2_sg U13792 ( .A(n13766), .B(n13767), .X(n13765) );
  nor_x2_sg U13682 ( .A(n13672), .B(n13673), .X(n13671) );
  nor_x2_sg U13882 ( .A(n52529), .B(n13819), .X(n13755) );
  nand_x8_sg U31473 ( .A(n26649), .B(n52524), .X(n13980) );
  nor_x2_sg U13983 ( .A(n13900), .B(n13901), .X(n13829) );
  nand_x8_sg U31468 ( .A(n26643), .B(n52545), .X(n13964) );
  nor_x2_sg U13844 ( .A(n13800), .B(n13801), .X(n13799) );
  nor_x2_sg U14030 ( .A(n52541), .B(n52475), .X(n13920) );
  nor_x2_sg U14009 ( .A(n13922), .B(n13923), .X(n13921) );
  nor_x2_sg U14076 ( .A(n52577), .B(n13967), .X(n13956) );
  nor_x2_sg U31458 ( .A(n26639), .B(n26640), .X(n14164) );
  nor_x2_sg U14073 ( .A(n13968), .B(n13969), .X(n13967) );
  nor_x2_sg U14070 ( .A(n13963), .B(n13964), .X(n13957) );
  nor_x2_sg U14055 ( .A(n13959), .B(n13960), .X(n13958) );
  nor_x2_sg U13962 ( .A(n13882), .B(n52605), .X(n13838) );
  nor_x2_sg U14323 ( .A(n14154), .B(n52596), .X(n14145) );
  nand_x8_sg U31592 ( .A(n26732), .B(n52592), .X(n14043) );
  nor_x2_sg U14292 ( .A(n14147), .B(n14148), .X(n14146) );
  nor_x2_sg U13972 ( .A(n13895), .B(n13896), .X(n13894) );
  nor_x2_sg U14082 ( .A(n13974), .B(n52562), .X(n13971) );
  nor_x2_sg U14252 ( .A(n14122), .B(n14123), .X(n14121) );
  nand_x8_sg U14129 ( .A(n13474), .B(n52619), .X(n13483) );
  nand_x8_sg U31711 ( .A(n26737), .B(n26750), .X(n26728) );
  nor_x2_sg U13966 ( .A(n13888), .B(n13483), .X(n13887) );
  nor_x2_sg U14356 ( .A(n14088), .B(n52603), .X(n14085) );
  nor_x2_sg U14220 ( .A(n14087), .B(n52617), .X(n14086) );
  nor_x2_sg U14211 ( .A(n14080), .B(n13775), .X(n14078) );
  nor_x2_sg U14151 ( .A(n14031), .B(n43085), .X(n14028) );
  nand_x8_sg U31715 ( .A(n26731), .B(n26749), .X(n14033) );
  nor_x2_sg U14140 ( .A(n46471), .B(n13856), .X(n14020) );
  nand_x8_sg U15420 ( .A(n46465), .B(n46579), .X(n8936) );
  nand_x8_sg U31732 ( .A(n46458), .B(n46462), .X(n14175) );
  nor_x2_sg U31996 ( .A(n52647), .B(n26996), .X(n26995) );
  nor_x2_sg U31983 ( .A(n26986), .B(n26987), .X(n26984) );
  nand_x8_sg U15277 ( .A(n46450), .B(n46458), .X(n14316) );
  nor_x2_sg U14547 ( .A(n52655), .B(n52671), .X(n14311) );
  nor_x2_sg U31975 ( .A(n26980), .B(n26981), .X(n26978) );
  nor_x2_sg U14544 ( .A(n14313), .B(n46454), .X(n14312) );
  nand_x8_sg U14981 ( .A(n52670), .B(n46458), .X(n14334) );
  nand_x8_sg U32120 ( .A(n27044), .B(n27045), .X(n26973) );
  nor_x2_sg U14635 ( .A(n46454), .B(n46451), .X(n14384) );
  nor_x2_sg U32123 ( .A(n27041), .B(n44323), .X(n26966) );
  nor_x2_sg U14632 ( .A(n46463), .B(n46445), .X(n14381) );
  nand_x8_sg U31954 ( .A(n26958), .B(n26959), .X(n14411) );
  nor_x2_sg U14628 ( .A(n14372), .B(n14373), .X(n14371) );
  nor_x2_sg U14639 ( .A(n52655), .B(n14347), .X(n14377) );
  nand_x8_sg U14745 ( .A(n52695), .B(n52648), .X(n14439) );
  nand_x8_sg U15135 ( .A(n52707), .B(n46458), .X(n14438) );
  nand_x8_sg U31947 ( .A(n26952), .B(n52723), .X(n14547) );
  nor_x2_sg U14716 ( .A(n41802), .B(n42365), .X(n14423) );
  nand_x8_sg U31942 ( .A(n26946), .B(n52741), .X(n14507) );
  nor_x2_sg U14712 ( .A(n14443), .B(n14444), .X(n14442) );
  nor_x2_sg U14697 ( .A(n14429), .B(n14430), .X(n14428) );
  nor_x2_sg U14725 ( .A(n43219), .B(n14421), .X(n14221) );
  nand_x8_sg U14865 ( .A(n14550), .B(n14551), .X(n14496) );
  nand_x8_sg U31936 ( .A(n26940), .B(n52762), .X(n14552) );
  nor_x2_sg U14790 ( .A(n14496), .B(n52771), .X(n14495) );
  nand_x8_sg U31931 ( .A(n26934), .B(n52782), .X(n14627) );
  nor_x2_sg U14841 ( .A(n14537), .B(n14538), .X(n14536) );
  nor_x2_sg U14728 ( .A(n14450), .B(n14451), .X(n14449) );
  nor_x2_sg U14926 ( .A(n43341), .B(n14596), .X(n14577) );
  nand_x8_sg U31925 ( .A(n26928), .B(n52805), .X(n14674) );
  nor_x2_sg U15051 ( .A(n52796), .B(n14675), .X(n14600) );
  nor_x2_sg U14891 ( .A(n14570), .B(n14571), .X(n14569) );
  nand_x8_sg U31920 ( .A(n26922), .B(n52823), .X(n14735) );
  nor_x2_sg U14992 ( .A(n14641), .B(n14642), .X(n14640) );
  nor_x2_sg U15081 ( .A(n52839), .B(n14703), .X(n14689) );
  nor_x2_sg U15077 ( .A(n14704), .B(n14705), .X(n14703) );
  nor_x2_sg U15122 ( .A(n52854), .B(n14738), .X(n14727) );
  nand_x8_sg U31914 ( .A(n26916), .B(n52847), .X(n14881) );
  nor_x2_sg U15119 ( .A(n14739), .B(n14740), .X(n14738) );
  nor_x2_sg U15116 ( .A(n14734), .B(n14735), .X(n14728) );
  nor_x2_sg U15101 ( .A(n14730), .B(n14731), .X(n14729) );
  nor_x2_sg U15008 ( .A(n14651), .B(n52883), .X(n14608) );
  nand_x8_sg U15344 ( .A(n14916), .B(n14917), .X(n14880) );
  nor_x2_sg U15378 ( .A(n14929), .B(n52874), .X(n14920) );
  nand_x8_sg U32044 ( .A(n27011), .B(n52869), .X(n14815) );
  nor_x2_sg U15347 ( .A(n14922), .B(n14923), .X(n14921) );
  nor_x2_sg U15018 ( .A(n14664), .B(n14665), .X(n14663) );
  nor_x2_sg U15304 ( .A(n14901), .B(n14902), .X(n14900) );
  nand_x8_sg U15175 ( .A(n14253), .B(n52898), .X(n14262) );
  nor_x2_sg U15172 ( .A(n52878), .B(n14776), .X(n14773) );
  nor_x2_sg U15333 ( .A(n43365), .B(n14898), .X(n14869) );
  nor_x2_sg U15289 ( .A(n14890), .B(n14891), .X(n14887) );
  nor_x2_sg U15288 ( .A(n14627), .B(n14889), .X(n14888) );
  nand_x8_sg U15394 ( .A(n52848), .B(n52648), .X(n14793) );
  nor_x2_sg U15403 ( .A(n46443), .B(n52893), .X(n14937) );
  nand_x8_sg U32164 ( .A(n27016), .B(n27029), .X(n27007) );
  nor_x2_sg U15398 ( .A(n14939), .B(n14547), .X(n14938) );
  nor_x2_sg U15153 ( .A(n14761), .B(n52821), .X(n14760) );
  nor_x2_sg U15012 ( .A(n14657), .B(n14262), .X(n14656) );
  nor_x2_sg U15407 ( .A(n14859), .B(n52880), .X(n14856) );
  nor_x2_sg U15267 ( .A(n14858), .B(n52903), .X(n14857) );
  nor_x2_sg U15258 ( .A(n14851), .B(n14411), .X(n14849) );
  nor_x2_sg U15197 ( .A(n14803), .B(n43083), .X(n14800) );
  nand_x8_sg U32168 ( .A(n27010), .B(n27028), .X(n14805) );
  nor_x2_sg U15186 ( .A(n46447), .B(n14627), .X(n14792) );
  nand_x8_sg U16481 ( .A(n46442), .B(n46579), .X(n8961) );
  nand_x8_sg U32186 ( .A(n46435), .B(n46439), .X(n14945) );
  nor_x2_sg U15432 ( .A(n14945), .B(n52929), .X(n14946) );
  nand_x8_sg U15562 ( .A(n46432), .B(n46439), .X(n14948) );
  nor_x2_sg U32462 ( .A(n52928), .B(n27276), .X(n27275) );
  nand_x8_sg U32585 ( .A(n27327), .B(n27328), .X(n27258) );
  nor_x2_sg U32436 ( .A(n27257), .B(n27258), .X(n27256) );
  nor_x2_sg U15585 ( .A(n15077), .B(n52954), .X(n15076) );
  nand_x8_sg U32587 ( .A(n27324), .B(n27325), .X(n27253) );
  nor_x2_sg U15643 ( .A(n15113), .B(n52982), .X(n15099) );
  nand_x8_sg U15702 ( .A(n46427), .B(n46432), .X(n15132) );
  nand_x8_sg U15699 ( .A(n15156), .B(n15157), .X(n15125) );
  nand_x8_sg U32589 ( .A(n27321), .B(n27322), .X(n27246) );
  nor_x2_sg U15690 ( .A(n15150), .B(n15151), .X(n15149) );
  nor_x2_sg U15685 ( .A(n15132), .B(n15148), .X(n15147) );
  nor_x2_sg U15700 ( .A(n52934), .B(n15125), .X(n15155) );
  nor_x2_sg U15726 ( .A(n52999), .B(n52951), .X(n15173) );
  nor_x2_sg U15721 ( .A(n46427), .B(n15175), .X(n15174) );
  nand_x8_sg U15799 ( .A(n52967), .B(n52934), .X(n15238) );
  nand_x8_sg U32410 ( .A(n27232), .B(n53006), .X(n15328) );
  nor_x2_sg U15779 ( .A(n15208), .B(n15207), .X(n15202) );
  nand_x8_sg U32405 ( .A(n27226), .B(n53020), .X(n15288) );
  nor_x2_sg U15804 ( .A(n15233), .B(n15244), .X(n15243) );
  nor_x2_sg U15794 ( .A(n15237), .B(n15238), .X(n15236) );
  nand_x8_sg U32399 ( .A(n27220), .B(n53039), .X(n15332) );
  nand_x8_sg U32394 ( .A(n27214), .B(n53060), .X(n15409) );
  nor_x2_sg U15901 ( .A(n15319), .B(n15320), .X(n15318) );
  nor_x2_sg U15791 ( .A(n15225), .B(n15226), .X(n15224) );
  nor_x2_sg U15991 ( .A(n53087), .B(n15372), .X(n15308) );
  nand_x8_sg U32388 ( .A(n27208), .B(n53082), .X(n15533) );
  nor_x2_sg U16093 ( .A(n15453), .B(n15454), .X(n15382) );
  nand_x8_sg U32383 ( .A(n27202), .B(n53104), .X(n15517) );
  nor_x2_sg U15953 ( .A(n15353), .B(n15354), .X(n15352) );
  nor_x2_sg U16140 ( .A(n53099), .B(n53032), .X(n15473) );
  nor_x2_sg U16119 ( .A(n15475), .B(n15476), .X(n15474) );
  nor_x2_sg U16186 ( .A(n53136), .B(n15520), .X(n15509) );
  nor_x2_sg U32373 ( .A(n27198), .B(n27199), .X(n15717) );
  nor_x2_sg U16183 ( .A(n15521), .B(n15522), .X(n15520) );
  nor_x2_sg U16180 ( .A(n15516), .B(n15517), .X(n15510) );
  nor_x2_sg U16165 ( .A(n15512), .B(n15513), .X(n15511) );
  nor_x2_sg U16072 ( .A(n15435), .B(n53164), .X(n15391) );
  nor_x2_sg U16432 ( .A(n15707), .B(n53155), .X(n15698) );
  nand_x8_sg U32510 ( .A(n27291), .B(n53151), .X(n15596) );
  nor_x2_sg U16402 ( .A(n15700), .B(n15701), .X(n15699) );
  nor_x2_sg U16082 ( .A(n15448), .B(n15449), .X(n15447) );
  nor_x2_sg U16192 ( .A(n15527), .B(n53121), .X(n15524) );
  nor_x2_sg U16362 ( .A(n15675), .B(n15676), .X(n15674) );
  nand_x8_sg U16239 ( .A(n15023), .B(n53178), .X(n15032) );
  nand_x8_sg U32629 ( .A(n27296), .B(n27309), .X(n27287) );
  nor_x2_sg U16218 ( .A(n15543), .B(n53102), .X(n15542) );
  nor_x2_sg U16076 ( .A(n15441), .B(n15032), .X(n15440) );
  nor_x2_sg U16465 ( .A(n15641), .B(n53162), .X(n15638) );
  nor_x2_sg U16330 ( .A(n15640), .B(n53176), .X(n15639) );
  nor_x2_sg U16321 ( .A(n15633), .B(n46423), .X(n15631) );
  nor_x2_sg U16261 ( .A(n15584), .B(n43079), .X(n15581) );
  nand_x8_sg U32633 ( .A(n27290), .B(n27308), .X(n15586) );
  nor_x2_sg U16250 ( .A(n46425), .B(n15409), .X(n15573) );
  nand_x8_sg U17546 ( .A(n46419), .B(n46579), .X(n9316) );
  nand_x8_sg U32650 ( .A(n46413), .B(n46417), .X(n15729) );
  nor_x2_sg U32915 ( .A(n53206), .B(n27555), .X(n27554) );
  nor_x2_sg U32902 ( .A(n27545), .B(n27546), .X(n27543) );
  nor_x2_sg U16646 ( .A(n15854), .B(n15855), .X(n15850) );
  nor_x2_sg U32894 ( .A(n27539), .B(n27540), .X(n27537) );
  nand_x8_sg U16664 ( .A(n15865), .B(n15866), .X(n15856) );
  nor_x2_sg U16643 ( .A(n15856), .B(n40581), .X(n15855) );
  nand_x8_sg U16724 ( .A(n46405), .B(n53207), .X(n15890) );
  nand_x8_sg U32888 ( .A(n27529), .B(n53239), .X(n15925) );
  nand_x8_sg U33038 ( .A(n27603), .B(n27604), .X(n27532) );
  nor_x2_sg U16702 ( .A(n53257), .B(n15891), .X(n15878) );
  nor_x2_sg U16757 ( .A(n46409), .B(n46406), .X(n15940) );
  nor_x2_sg U16754 ( .A(n46416), .B(n46402), .X(n15937) );
  nor_x2_sg U16750 ( .A(n15928), .B(n15929), .X(n15927) );
  nor_x2_sg U16761 ( .A(n53214), .B(n15903), .X(n15933) );
  nor_x2_sg U16787 ( .A(n53275), .B(n46404), .X(n15953) );
  nor_x2_sg U16782 ( .A(n53227), .B(n15955), .X(n15954) );
  nand_x8_sg U16860 ( .A(n53240), .B(n53214), .X(n16019) );
  nand_x8_sg U32865 ( .A(n27511), .B(n53281), .X(n16109) );
  nand_x8_sg U32860 ( .A(n27505), .B(n53297), .X(n16069) );
  nor_x2_sg U16865 ( .A(n16014), .B(n16025), .X(n16024) );
  nor_x2_sg U16855 ( .A(n16018), .B(n16019), .X(n16017) );
  nand_x8_sg U32854 ( .A(n27499), .B(n53318), .X(n16113) );
  nand_x8_sg U32849 ( .A(n27493), .B(n53339), .X(n16190) );
  nor_x2_sg U16964 ( .A(n16100), .B(n16101), .X(n16099) );
  nor_x2_sg U16852 ( .A(n16006), .B(n16007), .X(n16005) );
  nor_x2_sg U17050 ( .A(n43307), .B(n16160), .X(n16141) );
  nand_x8_sg U32843 ( .A(n27487), .B(n53362), .X(n16239) );
  nor_x2_sg U17177 ( .A(n53354), .B(n16240), .X(n16164) );
  nand_x8_sg U32838 ( .A(n27481), .B(n53383), .X(n16299) );
  nor_x2_sg U17016 ( .A(n16134), .B(n16135), .X(n16133) );
  nor_x2_sg U17206 ( .A(n53396), .B(n16267), .X(n16254) );
  nand_x8_sg U17438 ( .A(n53384), .B(n46413), .X(n16312) );
  nor_x2_sg U17202 ( .A(n16268), .B(n16269), .X(n16267) );
  nor_x2_sg U17180 ( .A(n16256), .B(n16257), .X(n16255) );
  nor_x2_sg U17244 ( .A(n53414), .B(n16302), .X(n16291) );
  nand_x8_sg U32832 ( .A(n27475), .B(n53407), .X(n16442) );
  nor_x2_sg U17241 ( .A(n16303), .B(n16304), .X(n16302) );
  nor_x2_sg U17238 ( .A(n16298), .B(n16299), .X(n16292) );
  nor_x2_sg U17223 ( .A(n16294), .B(n16295), .X(n16293) );
  nor_x2_sg U17135 ( .A(n16216), .B(n53443), .X(n16172) );
  nor_x2_sg U17467 ( .A(n16475), .B(n16476), .X(n16274) );
  nor_x2_sg U17457 ( .A(n53360), .B(n16451), .X(n16476) );
  nor_x2_sg U17500 ( .A(n16492), .B(n53435), .X(n16483) );
  nand_x8_sg U32963 ( .A(n27570), .B(n53429), .X(n16378) );
  nor_x2_sg U17469 ( .A(n16485), .B(n16486), .X(n16484) );
  nor_x2_sg U17141 ( .A(n16225), .B(n16226), .X(n16224) );
  nand_x8_sg U17441 ( .A(n16313), .B(n53393), .X(n16461) );
  nor_x2_sg U17437 ( .A(n16470), .B(n16461), .X(n16469) );
  nor_x2_sg U17425 ( .A(n16464), .B(n16465), .X(n16463) );
  nor_x2_sg U17293 ( .A(n53439), .B(n16339), .X(n16336) );
  nor_x2_sg U17454 ( .A(n43353), .B(n16460), .X(n16431) );
  nor_x2_sg U17410 ( .A(n16452), .B(n16453), .X(n16448) );
  nor_x2_sg U17409 ( .A(n16190), .B(n16450), .X(n16449) );
  nand_x8_sg U17517 ( .A(n53408), .B(n53207), .X(n16357) );
  nand_x8_sg U33082 ( .A(n27575), .B(n27588), .X(n27566) );
  nor_x2_sg U17519 ( .A(n16499), .B(n43175), .X(n16334) );
  nor_x2_sg U17274 ( .A(n16324), .B(n53380), .X(n16323) );
  nor_x2_sg U17385 ( .A(n16390), .B(n53433), .X(n16387) );
  nor_x2_sg U17380 ( .A(n16413), .B(n46400), .X(n16411) );
  nor_x2_sg U17349 ( .A(n16389), .B(n53450), .X(n16388) );
  nor_x2_sg U17342 ( .A(n16372), .B(n53431), .X(n16369) );
  nor_x2_sg U17328 ( .A(n16371), .B(n53409), .X(n16370) );
  nor_x2_sg U17319 ( .A(n16365), .B(n43039), .X(n16362) );
  nand_x8_sg U33086 ( .A(n27569), .B(n27587), .X(n16367) );
  nor_x2_sg U17308 ( .A(n15925), .B(n16190), .X(n16354) );
  nand_x8_sg U18606 ( .A(n46398), .B(n46579), .X(n9278) );
  nand_x8_sg U33106 ( .A(n46391), .B(n46395), .X(n16511) );
  nor_x2_sg U17558 ( .A(n16511), .B(n53487), .X(n16512) );
  nand_x8_sg U17688 ( .A(n46388), .B(n46395), .X(n16514) );
  nor_x2_sg U33372 ( .A(n53486), .B(n27834), .X(n27833) );
  nand_x8_sg U33495 ( .A(n27885), .B(n27886), .X(n27816) );
  nor_x2_sg U33346 ( .A(n27815), .B(n27816), .X(n27814) );
  nor_x2_sg U17711 ( .A(n16643), .B(n53512), .X(n16642) );
  nand_x8_sg U33497 ( .A(n27882), .B(n27883), .X(n27811) );
  nor_x2_sg U17769 ( .A(n16679), .B(n53540), .X(n16665) );
  nand_x8_sg U17828 ( .A(n46383), .B(n46388), .X(n16698) );
  nand_x8_sg U17825 ( .A(n16722), .B(n16723), .X(n16691) );
  nand_x8_sg U33499 ( .A(n27879), .B(n27880), .X(n27804) );
  nor_x2_sg U17816 ( .A(n16716), .B(n16717), .X(n16715) );
  nor_x2_sg U17811 ( .A(n16698), .B(n16714), .X(n16713) );
  nor_x2_sg U17826 ( .A(n53492), .B(n16691), .X(n16721) );
  nor_x2_sg U17852 ( .A(n53557), .B(n53509), .X(n16739) );
  nor_x2_sg U17847 ( .A(n46383), .B(n16741), .X(n16740) );
  nand_x8_sg U17925 ( .A(n53525), .B(n53492), .X(n16804) );
  nand_x8_sg U33320 ( .A(n27790), .B(n53564), .X(n16894) );
  nor_x2_sg U17905 ( .A(n16774), .B(n16773), .X(n16768) );
  nand_x8_sg U33315 ( .A(n27784), .B(n53578), .X(n16854) );
  nor_x2_sg U17930 ( .A(n16799), .B(n16810), .X(n16809) );
  nor_x2_sg U17920 ( .A(n16803), .B(n16804), .X(n16802) );
  nand_x8_sg U33309 ( .A(n27778), .B(n53597), .X(n16898) );
  nand_x8_sg U33304 ( .A(n27772), .B(n53618), .X(n16975) );
  nor_x2_sg U18027 ( .A(n16885), .B(n16886), .X(n16884) );
  nor_x2_sg U17917 ( .A(n16791), .B(n16792), .X(n16790) );
  nor_x2_sg U18117 ( .A(n53645), .B(n16938), .X(n16874) );
  nand_x8_sg U33298 ( .A(n27766), .B(n53640), .X(n17099) );
  nor_x2_sg U18219 ( .A(n17019), .B(n17020), .X(n16948) );
  nand_x8_sg U33293 ( .A(n27760), .B(n53662), .X(n17083) );
  nor_x2_sg U18079 ( .A(n16919), .B(n16920), .X(n16918) );
  nor_x2_sg U18266 ( .A(n53657), .B(n53590), .X(n17039) );
  nor_x2_sg U18245 ( .A(n17041), .B(n17042), .X(n17040) );
  nor_x2_sg U18312 ( .A(n53694), .B(n17086), .X(n17075) );
  nor_x2_sg U33283 ( .A(n27756), .B(n27757), .X(n17283) );
  nor_x2_sg U18309 ( .A(n17087), .B(n17088), .X(n17086) );
  nor_x2_sg U18306 ( .A(n17082), .B(n17083), .X(n17076) );
  nor_x2_sg U18291 ( .A(n17078), .B(n17079), .X(n17077) );
  nor_x2_sg U18198 ( .A(n17001), .B(n53722), .X(n16957) );
  nor_x2_sg U18558 ( .A(n17273), .B(n53713), .X(n17264) );
  nand_x8_sg U33420 ( .A(n27849), .B(n53709), .X(n17162) );
  nor_x2_sg U18528 ( .A(n17266), .B(n17267), .X(n17265) );
  nor_x2_sg U18208 ( .A(n17014), .B(n17015), .X(n17013) );
  nor_x2_sg U18318 ( .A(n17093), .B(n53679), .X(n17090) );
  nor_x2_sg U18488 ( .A(n17241), .B(n17242), .X(n17240) );
  nand_x8_sg U18365 ( .A(n16589), .B(n53736), .X(n16598) );
  nand_x8_sg U33539 ( .A(n27854), .B(n27867), .X(n27845) );
  nor_x2_sg U18344 ( .A(n17109), .B(n53660), .X(n17108) );
  nor_x2_sg U18202 ( .A(n17007), .B(n16598), .X(n17006) );
  nor_x2_sg U18591 ( .A(n17207), .B(n53720), .X(n17204) );
  nor_x2_sg U18456 ( .A(n17206), .B(n53734), .X(n17205) );
  nor_x2_sg U18447 ( .A(n17199), .B(n46379), .X(n17197) );
  nor_x2_sg U18387 ( .A(n17150), .B(n43077), .X(n17147) );
  nand_x8_sg U33543 ( .A(n27848), .B(n27866), .X(n17152) );
  nor_x2_sg U18376 ( .A(n46381), .B(n16975), .X(n17139) );
  nand_x8_sg U19658 ( .A(n46375), .B(n46579), .X(n9240) );
  nand_x8_sg U33565 ( .A(n46368), .B(n46372), .X(n17294) );
  nor_x2_sg U33831 ( .A(n53764), .B(n28115), .X(n28114) );
  nor_x2_sg U18785 ( .A(n46363), .B(n53790), .X(n17433) );
  nand_x8_sg U33954 ( .A(n28166), .B(n28167), .X(n28097) );
  nor_x2_sg U33805 ( .A(n28096), .B(n28097), .X(n28095) );
  nor_x2_sg U18782 ( .A(n17435), .B(n46364), .X(n17434) );
  nand_x8_sg U19221 ( .A(n46360), .B(n46368), .X(n17457) );
  nand_x8_sg U33803 ( .A(n28089), .B(n53801), .X(n17596) );
  nand_x8_sg U33956 ( .A(n28163), .B(n28164), .X(n28092) );
  nand_x8_sg U18876 ( .A(n17500), .B(n17501), .X(n17473) );
  nand_x8_sg U33958 ( .A(n28160), .B(n28161), .X(n28085) );
  nor_x2_sg U33787 ( .A(n28084), .B(n28085), .X(n28083) );
  nand_x8_sg U33786 ( .A(n28077), .B(n28078), .X(n17524) );
  nand_x8_sg U18912 ( .A(n53802), .B(n53765), .X(n17492) );
  nor_x2_sg U18867 ( .A(n17494), .B(n17495), .X(n17493) );
  nor_x2_sg U18862 ( .A(n17457), .B(n17492), .X(n17491) );
  nand_x8_sg U18977 ( .A(n46360), .B(n46361), .X(n17505) );
  nor_x2_sg U18877 ( .A(n46363), .B(n17473), .X(n17499) );
  nand_x8_sg U18985 ( .A(n46358), .B(n53765), .X(n17558) );
  nand_x8_sg U19373 ( .A(n53827), .B(n46368), .X(n17557) );
  nand_x8_sg U33779 ( .A(n28071), .B(n53843), .X(n17668) );
  nor_x2_sg U18956 ( .A(n41800), .B(n42363), .X(n17543) );
  nand_x8_sg U33774 ( .A(n28065), .B(n53861), .X(n17628) );
  nor_x2_sg U18952 ( .A(n17563), .B(n17564), .X(n17562) );
  nor_x2_sg U18936 ( .A(n17549), .B(n17505), .X(n17548) );
  nor_x2_sg U18965 ( .A(n43217), .B(n17541), .X(n17340) );
  nand_x8_sg U19105 ( .A(n17671), .B(n17672), .X(n17617) );
  nand_x8_sg U33768 ( .A(n28059), .B(n53882), .X(n17673) );
  nor_x2_sg U19030 ( .A(n17617), .B(n53891), .X(n17616) );
  nand_x8_sg U33763 ( .A(n28053), .B(n53902), .X(n17748) );
  nor_x2_sg U19081 ( .A(n17658), .B(n17659), .X(n17657) );
  nor_x2_sg U18968 ( .A(n17570), .B(n17571), .X(n17569) );
  nor_x2_sg U19166 ( .A(n43337), .B(n17717), .X(n17698) );
  nand_x8_sg U33757 ( .A(n28047), .B(n53925), .X(n17795) );
  nor_x2_sg U19289 ( .A(n53917), .B(n17796), .X(n17721) );
  nor_x2_sg U19131 ( .A(n17691), .B(n17692), .X(n17690) );
  nand_x8_sg U33752 ( .A(n28041), .B(n53943), .X(n17856) );
  nor_x2_sg U19232 ( .A(n17762), .B(n17763), .X(n17761) );
  nor_x2_sg U19319 ( .A(n53959), .B(n17824), .X(n17810) );
  nor_x2_sg U19315 ( .A(n17825), .B(n17826), .X(n17824) );
  nor_x2_sg U19292 ( .A(n17812), .B(n17813), .X(n17811) );
  nor_x2_sg U19360 ( .A(n53974), .B(n17859), .X(n17848) );
  nand_x8_sg U33746 ( .A(n28035), .B(n53967), .X(n18002) );
  nor_x2_sg U19357 ( .A(n17860), .B(n17861), .X(n17859) );
  nor_x2_sg U19354 ( .A(n17855), .B(n17856), .X(n17849) );
  nor_x2_sg U19339 ( .A(n17851), .B(n17852), .X(n17850) );
  nor_x2_sg U19248 ( .A(n17772), .B(n54003), .X(n17729) );
  nand_x8_sg U19583 ( .A(n18037), .B(n18038), .X(n18001) );
  nor_x2_sg U19616 ( .A(n18050), .B(n53994), .X(n18041) );
  nand_x8_sg U33879 ( .A(n28130), .B(n53989), .X(n17936) );
  nor_x2_sg U19586 ( .A(n18043), .B(n18044), .X(n18042) );
  nor_x2_sg U19258 ( .A(n17785), .B(n17786), .X(n17784) );
  nand_x8_sg U19413 ( .A(n17372), .B(n54018), .X(n17381) );
  nor_x2_sg U19410 ( .A(n53998), .B(n17897), .X(n17894) );
  nor_x2_sg U19572 ( .A(n43363), .B(n18019), .X(n17990) );
  nor_x2_sg U19528 ( .A(n18011), .B(n18012), .X(n18008) );
  nor_x2_sg U19527 ( .A(n17748), .B(n18010), .X(n18009) );
  nand_x8_sg U19632 ( .A(n53968), .B(n53765), .X(n17914) );
  nor_x2_sg U19641 ( .A(n46356), .B(n54013), .X(n18058) );
  nand_x8_sg U33998 ( .A(n28135), .B(n28148), .X(n28126) );
  nor_x2_sg U19636 ( .A(n18060), .B(n17668), .X(n18059) );
  nor_x2_sg U19391 ( .A(n17882), .B(n53941), .X(n17881) );
  nor_x2_sg U19252 ( .A(n17778), .B(n17381), .X(n17777) );
  nor_x2_sg U19645 ( .A(n17980), .B(n54000), .X(n17977) );
  nor_x2_sg U19505 ( .A(n17979), .B(n54023), .X(n17978) );
  nor_x2_sg U19496 ( .A(n17972), .B(n17524), .X(n17970) );
  nor_x2_sg U19435 ( .A(n17924), .B(n43075), .X(n17921) );
  nand_x8_sg U34002 ( .A(n28129), .B(n28147), .X(n17926) );
  nor_x2_sg U19424 ( .A(n17596), .B(n17748), .X(n17913) );
  nand_x8_sg U20711 ( .A(n46355), .B(n46579), .X(n9050) );
  nand_x8_sg U34019 ( .A(n46348), .B(n46352), .X(n18066) );
  nand_x8_sg U34412 ( .A(n28454), .B(n28455), .X(n28394) );
  nor_x2_sg U34295 ( .A(n28393), .B(n28394), .X(n28392) );
  nor_x2_sg U34284 ( .A(n28380), .B(n54059), .X(n18239) );
  nand_x8_sg U19864 ( .A(n46343), .B(n46345), .X(n18205) );
  nor_x2_sg U19835 ( .A(n46343), .B(n54071), .X(n18199) );
  nor_x2_sg U19832 ( .A(n18201), .B(n46344), .X(n18200) );
  nand_x8_sg U20267 ( .A(n54070), .B(n46348), .X(n18223) );
  nor_x2_sg U34264 ( .A(n28372), .B(n54082), .X(n28370) );
  nor_x2_sg U19923 ( .A(n40586), .B(n46340), .X(n18274) );
  nand_x8_sg U34423 ( .A(n28439), .B(n28440), .X(n28364) );
  nor_x2_sg U34251 ( .A(n28363), .B(n28364), .X(n28362) );
  nor_x2_sg U19920 ( .A(n46353), .B(n54097), .X(n18271) );
  nand_x8_sg U19960 ( .A(n54084), .B(n46345), .X(n18260) );
  nor_x2_sg U19913 ( .A(n18262), .B(n18263), .X(n18261) );
  nor_x2_sg U19927 ( .A(n46343), .B(n18240), .X(n18266) );
  nand_x8_sg U19930 ( .A(n18254), .B(n18247), .X(n18253) );
  nand_x8_sg U20421 ( .A(n54109), .B(n46348), .X(n18327) );
  nand_x8_sg U34243 ( .A(n28350), .B(n54123), .X(n18437) );
  nor_x2_sg U20003 ( .A(n41794), .B(n43223), .X(n18313) );
  nand_x8_sg U34435 ( .A(n28355), .B(n28434), .X(n28346) );
  nor_x2_sg U19983 ( .A(n18319), .B(n18320), .X(n18318) );
  nor_x2_sg U19980 ( .A(n18107), .B(n41748), .X(n18113) );
  nor_x2_sg U20012 ( .A(n43211), .B(n18311), .X(n18112) );
  nand_x8_sg U20151 ( .A(n18440), .B(n18441), .X(n18386) );
  nand_x8_sg U34232 ( .A(n28340), .B(n54164), .X(n18442) );
  nor_x2_sg U20077 ( .A(n18386), .B(n54172), .X(n18385) );
  nor_x2_sg U20158 ( .A(n18443), .B(n54188), .X(n18425) );
  nand_x8_sg U34227 ( .A(n28334), .B(n54183), .X(n18574) );
  nor_x2_sg U20127 ( .A(n18427), .B(n18428), .X(n18426) );
  nor_x2_sg U20015 ( .A(n18340), .B(n18341), .X(n18339) );
  nand_x8_sg U34221 ( .A(n28328), .B(n54208), .X(n18654) );
  nor_x2_sg U20211 ( .A(n46333), .B(n54211), .X(n18486) );
  nor_x2_sg U20316 ( .A(n18558), .B(n18485), .X(n18489) );
  nor_x2_sg U20177 ( .A(n18460), .B(n18461), .X(n18459) );
  nand_x8_sg U34216 ( .A(n28322), .B(n54228), .X(n18623) );
  nor_x2_sg U20278 ( .A(n18530), .B(n18531), .X(n18529) );
  nand_x8_sg U20593 ( .A(n46329), .B(n54070), .X(n18793) );
  nor_x2_sg U20408 ( .A(n18626), .B(n18627), .X(n18615) );
  nand_x8_sg U34210 ( .A(n28316), .B(n54249), .X(n18771) );
  nand_x8_sg U20650 ( .A(n54124), .B(n54084), .X(n18629) );
  nor_x2_sg U20405 ( .A(n18628), .B(n18629), .X(n18627) );
  nor_x2_sg U20402 ( .A(n18622), .B(n18623), .X(n18616) );
  nor_x2_sg U20387 ( .A(n18618), .B(n18619), .X(n18617) );
  nor_x2_sg U20295 ( .A(n18540), .B(n54285), .X(n18498) );
  nand_x8_sg U34345 ( .A(n28409), .B(n54272), .X(n18705) );
  nor_x2_sg U20651 ( .A(n18629), .B(n54257), .X(n18812) );
  nor_x2_sg U20634 ( .A(n18814), .B(n18815), .X(n18813) );
  nor_x2_sg U20305 ( .A(n18553), .B(n18554), .X(n18552) );
  nand_x8_sg U20606 ( .A(n18636), .B(n54240), .X(n18789) );
  nor_x2_sg U20602 ( .A(n18790), .B(n18789), .X(n18797) );
  nand_x8_sg U20460 ( .A(n18143), .B(n54300), .X(n18152) );
  nor_x2_sg U20457 ( .A(n54281), .B(n18666), .X(n18663) );
  nor_x2_sg U20618 ( .A(n42447), .B(n18788), .X(n18759) );
  nor_x2_sg U20590 ( .A(n18789), .B(n54253), .X(n18788) );
  nor_x2_sg U20576 ( .A(n18780), .B(n18781), .X(n18777) );
  nor_x2_sg U20575 ( .A(n18574), .B(n54246), .X(n18778) );
  nand_x8_sg U20683 ( .A(n54250), .B(n46345), .X(n18683) );
  nor_x2_sg U20692 ( .A(n54124), .B(n54295), .X(n18830) );
  nand_x8_sg U34463 ( .A(n28414), .B(n28427), .X(n28405) );
  nor_x2_sg U20687 ( .A(n18832), .B(n18437), .X(n18831) );
  nor_x2_sg U20438 ( .A(n18656), .B(n18657), .X(n18655) );
  nor_x2_sg U20299 ( .A(n18546), .B(n18152), .X(n18545) );
  nor_x2_sg U20464 ( .A(n42345), .B(n54287), .X(n18131) );
  nor_x2_sg U20696 ( .A(n18749), .B(n54283), .X(n18746) );
  nor_x2_sg U20552 ( .A(n18748), .B(n54304), .X(n18747) );
  nor_x2_sg U20543 ( .A(n18743), .B(n18437), .X(n18739) );
  nor_x2_sg U20534 ( .A(n18741), .B(n18742), .X(n18740) );
  nor_x2_sg U20482 ( .A(n18693), .B(n43069), .X(n18690) );
  nand_x8_sg U34467 ( .A(n28408), .B(n28426), .X(n18695) );
  nor_x2_sg U20471 ( .A(n46335), .B(n18574), .X(n18682) );
  nand_x8_sg U21763 ( .A(n46327), .B(n46579), .X(n9202) );
  nand_x8_sg U23869 ( .A(n21153), .B(n13393), .X(n19608) );
  nand_x8_sg U34484 ( .A(n46321), .B(n46325), .X(n18839) );
  nor_x2_sg U34751 ( .A(n54329), .B(n28673), .X(n28672) );
  nor_x2_sg U20890 ( .A(n46316), .B(n54355), .X(n18978) );
  nand_x8_sg U34874 ( .A(n28724), .B(n28725), .X(n28655) );
  nor_x2_sg U34725 ( .A(n28654), .B(n28655), .X(n28653) );
  nor_x2_sg U20887 ( .A(n18980), .B(n46317), .X(n18979) );
  nand_x8_sg U21326 ( .A(n46313), .B(n46321), .X(n19002) );
  nand_x8_sg U34723 ( .A(n28647), .B(n54366), .X(n19141) );
  nand_x8_sg U34876 ( .A(n28721), .B(n28722), .X(n28650) );
  nand_x8_sg U20981 ( .A(n19045), .B(n19046), .X(n19018) );
  nand_x8_sg U34878 ( .A(n28718), .B(n28719), .X(n28643) );
  nor_x2_sg U34707 ( .A(n28642), .B(n28643), .X(n28641) );
  nand_x8_sg U34706 ( .A(n28635), .B(n28636), .X(n19069) );
  nand_x8_sg U21017 ( .A(n54367), .B(n54330), .X(n19037) );
  nor_x2_sg U20972 ( .A(n19039), .B(n19040), .X(n19038) );
  nor_x2_sg U20967 ( .A(n19002), .B(n19037), .X(n19036) );
  nand_x8_sg U21082 ( .A(n46313), .B(n46314), .X(n19050) );
  nor_x2_sg U20982 ( .A(n46316), .B(n19018), .X(n19044) );
  nand_x8_sg U21090 ( .A(n46311), .B(n54330), .X(n19103) );
  nand_x8_sg U21478 ( .A(n54392), .B(n46321), .X(n19102) );
  nand_x8_sg U34699 ( .A(n28629), .B(n54408), .X(n19213) );
  nor_x2_sg U21061 ( .A(n41798), .B(n42361), .X(n19088) );
  nand_x8_sg U34694 ( .A(n28623), .B(n54426), .X(n19173) );
  nor_x2_sg U21057 ( .A(n19108), .B(n19109), .X(n19107) );
  nor_x2_sg U21041 ( .A(n19094), .B(n19050), .X(n19093) );
  nor_x2_sg U21070 ( .A(n43215), .B(n19086), .X(n18885) );
  nand_x8_sg U21210 ( .A(n19216), .B(n19217), .X(n19162) );
  nand_x8_sg U34688 ( .A(n28617), .B(n54447), .X(n19218) );
  nor_x2_sg U21135 ( .A(n19162), .B(n54456), .X(n19161) );
  nand_x8_sg U34683 ( .A(n28611), .B(n54467), .X(n19293) );
  nor_x2_sg U21186 ( .A(n19203), .B(n19204), .X(n19202) );
  nor_x2_sg U21073 ( .A(n19115), .B(n19116), .X(n19114) );
  nor_x2_sg U21271 ( .A(n43333), .B(n19262), .X(n19243) );
  nand_x8_sg U34677 ( .A(n28605), .B(n54490), .X(n19340) );
  nor_x2_sg U21394 ( .A(n54482), .B(n19341), .X(n19266) );
  nor_x2_sg U21236 ( .A(n19236), .B(n19237), .X(n19235) );
  nand_x8_sg U34672 ( .A(n28599), .B(n54508), .X(n19401) );
  nor_x2_sg U21337 ( .A(n19307), .B(n19308), .X(n19306) );
  nor_x2_sg U21424 ( .A(n54524), .B(n19369), .X(n19355) );
  nor_x2_sg U21420 ( .A(n19370), .B(n19371), .X(n19369) );
  nor_x2_sg U21397 ( .A(n19357), .B(n19358), .X(n19356) );
  nor_x2_sg U21465 ( .A(n54539), .B(n19404), .X(n19393) );
  nand_x8_sg U34666 ( .A(n28593), .B(n54532), .X(n19547) );
  nor_x2_sg U21462 ( .A(n19405), .B(n19406), .X(n19404) );
  nor_x2_sg U21459 ( .A(n19400), .B(n19401), .X(n19394) );
  nor_x2_sg U21444 ( .A(n19396), .B(n19397), .X(n19395) );
  nor_x2_sg U21353 ( .A(n19317), .B(n54568), .X(n19274) );
  nand_x8_sg U21688 ( .A(n19582), .B(n19583), .X(n19546) );
  nor_x2_sg U21721 ( .A(n19595), .B(n54559), .X(n19586) );
  nand_x8_sg U34799 ( .A(n28688), .B(n54554), .X(n19481) );
  nor_x2_sg U21691 ( .A(n19588), .B(n19589), .X(n19587) );
  nor_x2_sg U21363 ( .A(n19330), .B(n19331), .X(n19329) );
  nand_x8_sg U21518 ( .A(n18917), .B(n54583), .X(n18926) );
  nor_x2_sg U21515 ( .A(n54563), .B(n19442), .X(n19439) );
  nor_x2_sg U21677 ( .A(n43361), .B(n19564), .X(n19535) );
  nor_x2_sg U21633 ( .A(n19556), .B(n19557), .X(n19553) );
  nor_x2_sg U21632 ( .A(n19293), .B(n19555), .X(n19554) );
  nand_x8_sg U21737 ( .A(n54533), .B(n54330), .X(n19459) );
  nor_x2_sg U21746 ( .A(n46309), .B(n54578), .X(n19603) );
  nand_x8_sg U34918 ( .A(n28693), .B(n28706), .X(n28684) );
  nor_x2_sg U21741 ( .A(n19605), .B(n19213), .X(n19604) );
  nor_x2_sg U21496 ( .A(n19427), .B(n54506), .X(n19426) );
  nor_x2_sg U21357 ( .A(n19323), .B(n18926), .X(n19322) );
  nor_x2_sg U21750 ( .A(n19525), .B(n54565), .X(n19522) );
  nor_x2_sg U21610 ( .A(n19524), .B(n54588), .X(n19523) );
  nor_x2_sg U21601 ( .A(n19517), .B(n19069), .X(n19515) );
  nor_x2_sg U21540 ( .A(n19469), .B(n43067), .X(n19466) );
  nand_x8_sg U34922 ( .A(n28687), .B(n28705), .X(n19471) );
  nor_x2_sg U21529 ( .A(n19141), .B(n19293), .X(n19458) );
  nand_x8_sg U22818 ( .A(n46308), .B(n46579), .X(n9164) );
  nand_x8_sg U34939 ( .A(n46301), .B(n46305), .X(n19611) );
  nor_x2_sg U35204 ( .A(n54613), .B(n28951), .X(n28950) );
  nor_x2_sg U35191 ( .A(n28941), .B(n28942), .X(n28939) );
  nand_x8_sg U21969 ( .A(n46294), .B(n46301), .X(n19751) );
  nor_x2_sg U21940 ( .A(n46296), .B(n54635), .X(n19746) );
  nor_x2_sg U35183 ( .A(n28935), .B(n28936), .X(n28933) );
  nor_x2_sg U21937 ( .A(n19748), .B(n46297), .X(n19747) );
  nand_x8_sg U22376 ( .A(n54634), .B(n46301), .X(n19769) );
  nand_x8_sg U35327 ( .A(n28999), .B(n29000), .X(n28928) );
  nor_x2_sg U22029 ( .A(n46295), .B(n46297), .X(n19819) );
  nor_x2_sg U22026 ( .A(n46306), .B(n46289), .X(n19816) );
  nor_x2_sg U22022 ( .A(n19807), .B(n19808), .X(n19806) );
  nand_x8_sg U22132 ( .A(n46294), .B(n54634), .X(n19820) );
  nor_x2_sg U22033 ( .A(n46296), .B(n19785), .X(n19812) );
  nand_x8_sg U22140 ( .A(n54660), .B(n54614), .X(n19873) );
  nand_x8_sg U35154 ( .A(n28907), .B(n54687), .X(n19982) );
  nor_x2_sg U22111 ( .A(n41792), .B(n42357), .X(n19858) );
  nand_x8_sg U35343 ( .A(n28912), .B(n28991), .X(n28903) );
  nor_x2_sg U22091 ( .A(n19864), .B(n19820), .X(n19863) );
  nor_x2_sg U22120 ( .A(n43209), .B(n19856), .X(n19657) );
  nand_x8_sg U35143 ( .A(n28897), .B(n54730), .X(n19987) );
  nor_x2_sg U22185 ( .A(n19931), .B(n54738), .X(n19930) );
  nor_x2_sg U22266 ( .A(n19988), .B(n54755), .X(n19970) );
  nand_x8_sg U35138 ( .A(n28891), .B(n54750), .X(n20229) );
  nor_x2_sg U22235 ( .A(n19972), .B(n19973), .X(n19971) );
  nor_x2_sg U22123 ( .A(n19885), .B(n19886), .X(n19884) );
  nor_x2_sg U22320 ( .A(n43325), .B(n20031), .X(n20012) );
  nand_x8_sg U35132 ( .A(n28885), .B(n54775), .X(n20108) );
  nor_x2_sg U22445 ( .A(n54768), .B(n20109), .X(n20035) );
  nor_x2_sg U22285 ( .A(n20005), .B(n20006), .X(n20004) );
  nand_x8_sg U35127 ( .A(n28879), .B(n54793), .X(n20169) );
  nor_x2_sg U22387 ( .A(n20075), .B(n20076), .X(n20074) );
  nor_x2_sg U22475 ( .A(n54809), .B(n44417), .X(n20123) );
  nand_x8_sg U22700 ( .A(n46285), .B(n54634), .X(n20337) );
  nor_x2_sg U22516 ( .A(n20172), .B(n20173), .X(n20161) );
  nand_x8_sg U35121 ( .A(n28873), .B(n54817), .X(n20317) );
  nand_x8_sg U22758 ( .A(n54688), .B(n54647), .X(n20175) );
  nor_x2_sg U22513 ( .A(n20174), .B(n20175), .X(n20173) );
  nor_x2_sg U22510 ( .A(n20168), .B(n20169), .X(n20162) );
  nor_x2_sg U22495 ( .A(n20164), .B(n20165), .X(n20163) );
  nor_x2_sg U22404 ( .A(n20085), .B(n54853), .X(n20043) );
  nand_x8_sg U22737 ( .A(n20352), .B(n20353), .X(n20316) );
  nand_x8_sg U35252 ( .A(n28966), .B(n54839), .X(n20251) );
  nor_x2_sg U22759 ( .A(n20175), .B(n54824), .X(n20357) );
  nor_x2_sg U22741 ( .A(n20359), .B(n20360), .X(n20358) );
  nor_x2_sg U22414 ( .A(n20098), .B(n20099), .X(n20097) );
  nand_x8_sg U22569 ( .A(n19688), .B(n54868), .X(n19697) );
  nor_x2_sg U22566 ( .A(n54848), .B(n20211), .X(n20208) );
  nor_x2_sg U22726 ( .A(n42445), .B(n20334), .X(n20305) );
  nor_x2_sg U22684 ( .A(n20326), .B(n20327), .X(n20323) );
  nor_x2_sg U22683 ( .A(n20229), .B(n20325), .X(n20324) );
  nand_x8_sg U22791 ( .A(n54818), .B(n54614), .X(n20228) );
  nor_x2_sg U22800 ( .A(n54688), .B(n54863), .X(n20375) );
  nand_x8_sg U35371 ( .A(n28971), .B(n28984), .X(n28962) );
  nor_x2_sg U22795 ( .A(n20377), .B(n19982), .X(n20376) );
  nor_x2_sg U22546 ( .A(n20196), .B(n54790), .X(n20195) );
  nor_x2_sg U22408 ( .A(n20091), .B(n19697), .X(n20090) );
  nor_x2_sg U22573 ( .A(n42343), .B(n54855), .X(n19676) );
  nor_x2_sg U22804 ( .A(n20295), .B(n54850), .X(n20292) );
  nor_x2_sg U22661 ( .A(n20294), .B(n54872), .X(n20293) );
  nor_x2_sg U22652 ( .A(n20289), .B(n19982), .X(n20285) );
  nor_x2_sg U22643 ( .A(n20287), .B(n20288), .X(n20286) );
  nor_x2_sg U22591 ( .A(n20239), .B(n43061), .X(n20236) );
  nand_x8_sg U35375 ( .A(n28965), .B(n28983), .X(n20241) );
  nor_x2_sg U22580 ( .A(n46291), .B(n20229), .X(n20227) );
  nand_x8_sg U23871 ( .A(n46283), .B(n46579), .X(n9126) );
  nand_x8_sg U35398 ( .A(n46276), .B(n46280), .X(n20383) );
  nor_x2_sg U35669 ( .A(n54897), .B(n29234), .X(n29233) );
  nor_x2_sg U22997 ( .A(n46271), .B(n54923), .X(n20522) );
  nand_x8_sg U35792 ( .A(n29285), .B(n29286), .X(n29216) );
  nor_x2_sg U35643 ( .A(n29215), .B(n29216), .X(n29214) );
  nor_x2_sg U22994 ( .A(n20524), .B(n46272), .X(n20523) );
  nand_x8_sg U23433 ( .A(n46268), .B(n46276), .X(n20546) );
  nand_x8_sg U35641 ( .A(n29208), .B(n54934), .X(n20685) );
  nand_x8_sg U35794 ( .A(n29282), .B(n29283), .X(n29211) );
  nand_x8_sg U23088 ( .A(n20589), .B(n20590), .X(n20562) );
  nand_x8_sg U35796 ( .A(n29279), .B(n29280), .X(n29204) );
  nor_x2_sg U35625 ( .A(n29203), .B(n29204), .X(n29202) );
  nand_x8_sg U35624 ( .A(n29196), .B(n29197), .X(n20613) );
  nand_x8_sg U23124 ( .A(n54935), .B(n54898), .X(n20581) );
  nor_x2_sg U23079 ( .A(n20583), .B(n20584), .X(n20582) );
  nor_x2_sg U23074 ( .A(n20546), .B(n20581), .X(n20580) );
  nand_x8_sg U23189 ( .A(n46268), .B(n46269), .X(n20594) );
  nor_x2_sg U23089 ( .A(n46271), .B(n20562), .X(n20588) );
  nand_x8_sg U23197 ( .A(n46266), .B(n54898), .X(n20647) );
  nand_x8_sg U23585 ( .A(n54960), .B(n46276), .X(n20646) );
  nand_x8_sg U35617 ( .A(n29190), .B(n54976), .X(n20757) );
  nor_x2_sg U23168 ( .A(n41796), .B(n42359), .X(n20632) );
  nand_x8_sg U35612 ( .A(n29184), .B(n54994), .X(n20717) );
  nor_x2_sg U23164 ( .A(n20652), .B(n20653), .X(n20651) );
  nor_x2_sg U23148 ( .A(n20638), .B(n20594), .X(n20637) );
  nor_x2_sg U23177 ( .A(n43213), .B(n20630), .X(n20429) );
  nand_x8_sg U23317 ( .A(n20760), .B(n20761), .X(n20706) );
  nand_x8_sg U35606 ( .A(n29178), .B(n55015), .X(n20762) );
  nor_x2_sg U23242 ( .A(n20706), .B(n55024), .X(n20705) );
  nand_x8_sg U35601 ( .A(n29172), .B(n55035), .X(n20837) );
  nor_x2_sg U23293 ( .A(n20747), .B(n20748), .X(n20746) );
  nor_x2_sg U23180 ( .A(n20659), .B(n20660), .X(n20658) );
  nor_x2_sg U23378 ( .A(n43329), .B(n20806), .X(n20787) );
  nand_x8_sg U35595 ( .A(n29166), .B(n55058), .X(n20884) );
  nor_x2_sg U23501 ( .A(n55050), .B(n20885), .X(n20810) );
  nor_x2_sg U23343 ( .A(n20780), .B(n20781), .X(n20779) );
  nand_x8_sg U35590 ( .A(n29160), .B(n55076), .X(n20945) );
  nor_x2_sg U23444 ( .A(n20851), .B(n20852), .X(n20850) );
  nor_x2_sg U23531 ( .A(n55092), .B(n20913), .X(n20899) );
  nor_x2_sg U23527 ( .A(n20914), .B(n20915), .X(n20913) );
  nor_x2_sg U23504 ( .A(n20901), .B(n20902), .X(n20900) );
  nor_x2_sg U23572 ( .A(n55107), .B(n20948), .X(n20937) );
  nand_x8_sg U35584 ( .A(n29154), .B(n55100), .X(n21091) );
  nor_x2_sg U23569 ( .A(n20949), .B(n20950), .X(n20948) );
  nor_x2_sg U23566 ( .A(n20944), .B(n20945), .X(n20938) );
  nor_x2_sg U23551 ( .A(n20940), .B(n20941), .X(n20939) );
  nor_x2_sg U23460 ( .A(n20861), .B(n55136), .X(n20818) );
  nand_x8_sg U23795 ( .A(n21126), .B(n21127), .X(n21090) );
  nor_x2_sg U23828 ( .A(n21139), .B(n55127), .X(n21130) );
  nand_x8_sg U35717 ( .A(n29249), .B(n55122), .X(n21025) );
  nor_x2_sg U23798 ( .A(n21132), .B(n21133), .X(n21131) );
  nor_x2_sg U23470 ( .A(n20874), .B(n20875), .X(n20873) );
  nand_x8_sg U23625 ( .A(n20461), .B(n55151), .X(n20470) );
  nor_x2_sg U23622 ( .A(n55131), .B(n20986), .X(n20983) );
  nor_x2_sg U23784 ( .A(n43359), .B(n21108), .X(n21079) );
  nor_x2_sg U23740 ( .A(n21100), .B(n21101), .X(n21097) );
  nor_x2_sg U23739 ( .A(n20837), .B(n21099), .X(n21098) );
  nand_x8_sg U23844 ( .A(n55101), .B(n54898), .X(n21003) );
  nor_x2_sg U23853 ( .A(n46264), .B(n55146), .X(n21147) );
  nand_x8_sg U35836 ( .A(n29254), .B(n29267), .X(n29245) );
  nor_x2_sg U23848 ( .A(n21149), .B(n20757), .X(n21148) );
  nor_x2_sg U23603 ( .A(n20971), .B(n55074), .X(n20970) );
  nor_x2_sg U23464 ( .A(n20867), .B(n20470), .X(n20866) );
  nor_x2_sg U23857 ( .A(n21069), .B(n55133), .X(n21066) );
  nor_x2_sg U23717 ( .A(n21068), .B(n55156), .X(n21067) );
  nor_x2_sg U23708 ( .A(n21061), .B(n20613), .X(n21059) );
  nor_x2_sg U23647 ( .A(n21013), .B(n43059), .X(n21010) );
  nand_x8_sg U35840 ( .A(n29248), .B(n29266), .X(n21015) );
  nor_x2_sg U23636 ( .A(n20685), .B(n20837), .X(n21002) );
  nand_x8_sg U24929 ( .A(n46263), .B(n46579), .X(n9088) );
  nand_x8_sg U35857 ( .A(n46256), .B(n46260), .X(n21156) );
  nor_x2_sg U36132 ( .A(n55181), .B(n29512), .X(n29511) );
  nor_x2_sg U36119 ( .A(n29502), .B(n29503), .X(n29500) );
  nand_x8_sg U24077 ( .A(n46249), .B(n46256), .X(n21296) );
  nor_x2_sg U24048 ( .A(n46251), .B(n55203), .X(n21291) );
  nor_x2_sg U36111 ( .A(n29496), .B(n29497), .X(n29494) );
  nor_x2_sg U24045 ( .A(n21293), .B(n46252), .X(n21292) );
  nand_x8_sg U24484 ( .A(n55202), .B(n46256), .X(n21314) );
  nand_x8_sg U36255 ( .A(n29560), .B(n29561), .X(n29489) );
  nor_x2_sg U24137 ( .A(n46250), .B(n46252), .X(n21364) );
  nor_x2_sg U24134 ( .A(n46261), .B(n46244), .X(n21361) );
  nor_x2_sg U24130 ( .A(n21352), .B(n21353), .X(n21351) );
  nand_x8_sg U24240 ( .A(n46249), .B(n55202), .X(n21365) );
  nor_x2_sg U24141 ( .A(n46251), .B(n21330), .X(n21357) );
  nand_x8_sg U24248 ( .A(n55228), .B(n55182), .X(n21418) );
  nand_x8_sg U36082 ( .A(n29468), .B(n55255), .X(n21527) );
  nor_x2_sg U24219 ( .A(n41790), .B(n42355), .X(n21403) );
  nand_x8_sg U36271 ( .A(n29473), .B(n29552), .X(n29464) );
  nor_x2_sg U24199 ( .A(n21409), .B(n21365), .X(n21408) );
  nor_x2_sg U24228 ( .A(n43207), .B(n21401), .X(n21202) );
  nand_x8_sg U36071 ( .A(n29458), .B(n55298), .X(n21532) );
  nor_x2_sg U24293 ( .A(n21476), .B(n55306), .X(n21475) );
  nor_x2_sg U24374 ( .A(n21533), .B(n55323), .X(n21515) );
  nand_x8_sg U36066 ( .A(n29452), .B(n55318), .X(n21774) );
  nor_x2_sg U24343 ( .A(n21517), .B(n21518), .X(n21516) );
  nor_x2_sg U24231 ( .A(n21430), .B(n21431), .X(n21429) );
  nor_x2_sg U24428 ( .A(n43321), .B(n21576), .X(n21557) );
  nand_x8_sg U36060 ( .A(n29446), .B(n55343), .X(n21653) );
  nor_x2_sg U24553 ( .A(n55336), .B(n21654), .X(n21580) );
  nor_x2_sg U24393 ( .A(n21550), .B(n21551), .X(n21549) );
  nand_x8_sg U36055 ( .A(n29440), .B(n55361), .X(n21714) );
  nor_x2_sg U24495 ( .A(n21620), .B(n21621), .X(n21619) );
  nor_x2_sg U24583 ( .A(n55377), .B(n44415), .X(n21668) );
  nand_x8_sg U24808 ( .A(n46240), .B(n55202), .X(n21882) );
  nor_x2_sg U24624 ( .A(n21717), .B(n21718), .X(n21706) );
  nand_x8_sg U36049 ( .A(n29434), .B(n55385), .X(n21862) );
  nand_x8_sg U24866 ( .A(n55256), .B(n55215), .X(n21720) );
  nor_x2_sg U24621 ( .A(n21719), .B(n21720), .X(n21718) );
  nor_x2_sg U24618 ( .A(n21713), .B(n21714), .X(n21707) );
  nor_x2_sg U24603 ( .A(n21709), .B(n21710), .X(n21708) );
  nor_x2_sg U24512 ( .A(n21630), .B(n55421), .X(n21588) );
  nand_x8_sg U24845 ( .A(n21897), .B(n21898), .X(n21861) );
  nand_x8_sg U36180 ( .A(n29527), .B(n55407), .X(n21796) );
  nor_x2_sg U24867 ( .A(n21720), .B(n55392), .X(n21902) );
  nor_x2_sg U24849 ( .A(n21904), .B(n21905), .X(n21903) );
  nor_x2_sg U24522 ( .A(n21643), .B(n21644), .X(n21642) );
  nand_x8_sg U24677 ( .A(n21233), .B(n55436), .X(n21242) );
  nor_x2_sg U24674 ( .A(n55416), .B(n21756), .X(n21753) );
  nor_x2_sg U24834 ( .A(n42443), .B(n21879), .X(n21850) );
  nor_x2_sg U24792 ( .A(n21871), .B(n21872), .X(n21868) );
  nor_x2_sg U24791 ( .A(n21774), .B(n21870), .X(n21869) );
  nand_x8_sg U24899 ( .A(n55386), .B(n55182), .X(n21773) );
  nor_x2_sg U24908 ( .A(n55256), .B(n55431), .X(n21920) );
  nand_x8_sg U36299 ( .A(n29532), .B(n29545), .X(n29523) );
  nor_x2_sg U24903 ( .A(n21922), .B(n21527), .X(n21921) );
  nor_x2_sg U24654 ( .A(n21741), .B(n55358), .X(n21740) );
  nor_x2_sg U24516 ( .A(n21636), .B(n21242), .X(n21635) );
  nor_x2_sg U24681 ( .A(n42341), .B(n55423), .X(n21221) );
  nor_x2_sg U24912 ( .A(n21840), .B(n55418), .X(n21837) );
  nor_x2_sg U24769 ( .A(n21839), .B(n55440), .X(n21838) );
  nor_x2_sg U24760 ( .A(n21834), .B(n21527), .X(n21830) );
  nor_x2_sg U24751 ( .A(n21832), .B(n21833), .X(n21831) );
  nor_x2_sg U24699 ( .A(n21784), .B(n43053), .X(n21781) );
  nand_x8_sg U36303 ( .A(n29526), .B(n29544), .X(n21786) );
  nor_x2_sg U24688 ( .A(n46246), .B(n21774), .X(n21772) );
  nand_x8_sg U29893 ( .A(n25388), .B(n46236), .X(n24476) );
  nand_x8_sg U29892 ( .A(n46611), .B(n32136), .X(n25388) );
  nand_x8_sg U36036 ( .A(n46576), .B(n46236), .X(n26358) );
  nor_x2_sg U25147 ( .A(n30281), .B(n8243), .X(n30279) );
  nand_x8_sg U25375 ( .A(n30440), .B(n50079), .X(n24505) );
  nand_x8_sg U25370 ( .A(n30536), .B(n30537), .X(n30278) );
  nor_x2_sg U25595 ( .A(n30785), .B(n50003), .X(n30700) );
  nor_x2_sg U25594 ( .A(n30533), .B(n8285), .X(n30785) );
  nand_x8_sg U25593 ( .A(n30787), .B(n30788), .X(n30533) );
  nand_x8_sg U25816 ( .A(n31005), .B(n31006), .X(n30784) );
  nor_x2_sg U26041 ( .A(n31204), .B(n49915), .X(n31137) );
  nor_x2_sg U26040 ( .A(n31002), .B(n8327), .X(n31204) );
  nand_x8_sg U26039 ( .A(n31206), .B(n31207), .X(n31002) );
  nand_x8_sg U26271 ( .A(n31328), .B(n49890), .X(n24685) );
  nand_x8_sg U26492 ( .A(n49842), .B(n31502), .X(n24756) );
  nor_x2_sg U26488 ( .A(n31386), .B(n8369), .X(n31552) );
  nand_x8_sg U26487 ( .A(n31554), .B(n31555), .X(n31386) );
  nand_x8_sg U26716 ( .A(n31658), .B(n49794), .X(n24780) );
  nand_x8_sg U26711 ( .A(n31701), .B(n31702), .X(n31551) );
  nor_x2_sg U26936 ( .A(n31697), .B(n8411), .X(n31836) );
  nand_x8_sg U26935 ( .A(n31838), .B(n31839), .X(n31697) );
  nand_x8_sg U27164 ( .A(n31924), .B(n49695), .X(n31801) );
  nand_x8_sg U27159 ( .A(n31948), .B(n31949), .X(n31835) );
  nor_x2_sg U27385 ( .A(n31945), .B(n8453), .X(n32041) );
  nand_x8_sg U27611 ( .A(n32110), .B(n49599), .X(n32024) );
  nand_x8_sg U27604 ( .A(n32113), .B(n32114), .X(n32038) );
  nand_x8_sg U28073 ( .A(n32119), .B(n32120), .X(n32101) );
  nand_x8_sg U29014 ( .A(n32131), .B(n32132), .X(n32077) );
  nor_x2_sg U28776 ( .A(n32077), .B(n8480), .X(n32130) );
  nor_x2_sg U28307 ( .A(n49368), .B(n8478), .X(n32124) );
  nor_x2_sg U27835 ( .A(n32101), .B(n8476), .X(n32118) );
  nor_x2_sg U27844 ( .A(n32108), .B(n32109), .X(n32106) );
  nand_x8_sg U27854 ( .A(n32049), .B(n32050), .X(n32021) );
  nand_x8_sg U28090 ( .A(n32052), .B(n32053), .X(n32014) );
  nand_x8_sg U28325 ( .A(n32055), .B(n32056), .X(n32008) );
  nor_x2_sg U28550 ( .A(n32090), .B(n32091), .X(n32088) );
  nor_x2_sg U28547 ( .A(n40786), .B(n8478), .X(n32091) );
  nand_x8_sg U28560 ( .A(n32058), .B(n32059), .X(n32001) );
  nor_x2_sg U28781 ( .A(n40785), .B(n8479), .X(n32085) );
  nand_x8_sg U28794 ( .A(n32061), .B(n32062), .X(n31995) );
  nand_x8_sg U29027 ( .A(n32064), .B(n32065), .X(n31989) );
  nand_x8_sg U27377 ( .A(n32032), .B(n49645), .X(n31944) );
  nand_x8_sg U27370 ( .A(n32035), .B(n49597), .X(n31935) );
  nor_x2_sg U27366 ( .A(n32038), .B(n8474), .X(n32037) );
  nand_x8_sg U27394 ( .A(n31951), .B(n31952), .X(n31922) );
  nor_x2_sg U27620 ( .A(n32028), .B(n8454), .X(n32026) );
  nand_x8_sg U27629 ( .A(n31954), .B(n31955), .X(n31916) );
  nor_x2_sg U27855 ( .A(n32021), .B(n8455), .X(n32019) );
  nand_x8_sg U27864 ( .A(n31957), .B(n31958), .X(n31910) );
  nor_x2_sg U28092 ( .A(n32012), .B(n49503), .X(n32011) );
  nor_x2_sg U28091 ( .A(n32014), .B(n8456), .X(n32012) );
  nand_x8_sg U28100 ( .A(n31960), .B(n31961), .X(n31904) );
  nor_x2_sg U28326 ( .A(n32008), .B(n8457), .X(n32006) );
  nand_x8_sg U28335 ( .A(n31963), .B(n31964), .X(n31898) );
  nor_x2_sg U28562 ( .A(n31999), .B(n49412), .X(n31998) );
  nor_x2_sg U28561 ( .A(n32001), .B(n8458), .X(n31999) );
  nand_x8_sg U28570 ( .A(n31966), .B(n31967), .X(n31892) );
  nor_x2_sg U28796 ( .A(n31993), .B(n49367), .X(n31992) );
  nor_x2_sg U28795 ( .A(n31995), .B(n8459), .X(n31993) );
  nand_x8_sg U28804 ( .A(n31969), .B(n31970), .X(n31886) );
  nor_x2_sg U29028 ( .A(n31989), .B(n8460), .X(n31987) );
  nand_x8_sg U29036 ( .A(n31972), .B(n31973), .X(n31880) );
  nand_x8_sg U29394 ( .A(n49251), .B(n31975), .X(n25348) );
  nor_x2_sg U27150 ( .A(n31829), .B(n8452), .X(n31939) );
  nand_x8_sg U27149 ( .A(n31941), .B(n31942), .X(n31829) );
  nand_x8_sg U27142 ( .A(n31930), .B(n31931), .X(n31828) );
  nor_x2_sg U27130 ( .A(n31935), .B(n8473), .X(n31934) );
  nand_x8_sg U27171 ( .A(n31841), .B(n31842), .X(n31804) );
  nand_x8_sg U27406 ( .A(n31844), .B(n31845), .X(n31797) );
  nand_x8_sg U27641 ( .A(n31847), .B(n31848), .X(n31790) );
  nand_x8_sg U27876 ( .A(n31850), .B(n31851), .X(n31783) );
  nand_x8_sg U28112 ( .A(n31853), .B(n31854), .X(n31776) );
  nand_x8_sg U28347 ( .A(n31856), .B(n31857), .X(n31769) );
  nand_x8_sg U28582 ( .A(n31859), .B(n31860), .X(n31762) );
  nand_x8_sg U28816 ( .A(n31862), .B(n31863), .X(n31755) );
  nand_x8_sg U29047 ( .A(n31865), .B(n31866), .X(n31748) );
  nand_x8_sg U26928 ( .A(n31808), .B(n49741), .X(n31698) );
  nand_x8_sg U26923 ( .A(n31832), .B(n31833), .X(n31691) );
  nor_x2_sg U26914 ( .A(n31685), .B(n8451), .X(n31823) );
  nand_x8_sg U26906 ( .A(n31814), .B(n49736), .X(n31684) );
  nand_x8_sg U26899 ( .A(n31817), .B(n31818), .X(n31675) );
  nand_x8_sg U26945 ( .A(n31704), .B(n31705), .X(n31656) );
  nor_x2_sg U27172 ( .A(n31804), .B(n8412), .X(n31802) );
  nand_x8_sg U27181 ( .A(n31707), .B(n31708), .X(n31650) );
  nor_x2_sg U27407 ( .A(n31797), .B(n8413), .X(n31795) );
  nand_x8_sg U27416 ( .A(n31710), .B(n31711), .X(n31644) );
  nor_x2_sg U27642 ( .A(n31790), .B(n8414), .X(n31788) );
  nand_x8_sg U27651 ( .A(n31713), .B(n31714), .X(n31638) );
  nor_x2_sg U27877 ( .A(n31783), .B(n8415), .X(n31781) );
  nand_x8_sg U27886 ( .A(n31716), .B(n31717), .X(n31632) );
  nor_x2_sg U28113 ( .A(n31776), .B(n8416), .X(n31774) );
  nand_x8_sg U28122 ( .A(n31719), .B(n31720), .X(n31626) );
  nor_x2_sg U28348 ( .A(n31769), .B(n8417), .X(n31767) );
  nand_x8_sg U28357 ( .A(n31722), .B(n31723), .X(n31620) );
  nor_x2_sg U28583 ( .A(n31762), .B(n8418), .X(n31760) );
  nand_x8_sg U28592 ( .A(n31725), .B(n31726), .X(n31614) );
  nor_x2_sg U28817 ( .A(n31755), .B(n8419), .X(n31753) );
  nand_x8_sg U28826 ( .A(n31728), .B(n31729), .X(n31608) );
  nor_x2_sg U29048 ( .A(n31748), .B(n8420), .X(n31746) );
  nand_x8_sg U29056 ( .A(n31731), .B(n31732), .X(n31602) );
  nand_x8_sg U29400 ( .A(n49254), .B(n31734), .X(n25349) );
  nor_x2_sg U26702 ( .A(n31544), .B(n8410), .X(n31692) );
  nand_x8_sg U26701 ( .A(n31694), .B(n31695), .X(n31544) );
  nand_x8_sg U26694 ( .A(n31664), .B(n49787), .X(n31545) );
  nand_x8_sg U26689 ( .A(n31688), .B(n31689), .X(n31538) );
  nor_x2_sg U26680 ( .A(n31532), .B(n8450), .X(n31679) );
  nand_x8_sg U26679 ( .A(n31681), .B(n31682), .X(n31532) );
  nand_x8_sg U26672 ( .A(n31670), .B(n31671), .X(n31531) );
  nor_x2_sg U26660 ( .A(n31675), .B(n8471), .X(n31674) );
  nand_x8_sg U26723 ( .A(n31557), .B(n31558), .X(n31501) );
  nand_x8_sg U26950 ( .A(n31652), .B(n49746), .X(n24827) );
  nand_x8_sg U26957 ( .A(n31560), .B(n31561), .X(n31495) );
  nand_x8_sg U27186 ( .A(n31646), .B(n49697), .X(n24875) );
  nand_x8_sg U27193 ( .A(n31563), .B(n31564), .X(n31489) );
  nand_x8_sg U27421 ( .A(n31640), .B(n49650), .X(n24923) );
  nand_x8_sg U27428 ( .A(n31566), .B(n31567), .X(n31483) );
  nand_x8_sg U27656 ( .A(n31634), .B(n49603), .X(n24971) );
  nand_x8_sg U27663 ( .A(n31569), .B(n31570), .X(n31477) );
  nand_x8_sg U27891 ( .A(n31628), .B(n49557), .X(n25019) );
  nand_x8_sg U27898 ( .A(n31572), .B(n31573), .X(n31471) );
  nand_x8_sg U28127 ( .A(n31622), .B(n49510), .X(n25067) );
  nand_x8_sg U28134 ( .A(n31575), .B(n31576), .X(n31465) );
  nand_x8_sg U28362 ( .A(n31616), .B(n49463), .X(n25116) );
  nand_x8_sg U28369 ( .A(n31578), .B(n31579), .X(n31459) );
  nand_x8_sg U28597 ( .A(n31610), .B(n49417), .X(n25164) );
  nand_x8_sg U28604 ( .A(n31581), .B(n31582), .X(n31453) );
  nand_x8_sg U28831 ( .A(n31604), .B(n49371), .X(n25213) );
  nand_x8_sg U28838 ( .A(n31584), .B(n31585), .X(n31447) );
  nand_x8_sg U29061 ( .A(n31598), .B(n49327), .X(n25262) );
  nand_x8_sg U29067 ( .A(n31587), .B(n31588), .X(n31441) );
  nand_x8_sg U29256 ( .A(n31591), .B(n31592), .X(n25307) );
  nand_x8_sg U29403 ( .A(n49255), .B(n31590), .X(n25352) );
  nand_x8_sg U26480 ( .A(n31505), .B(n49839), .X(n24732) );
  nand_x8_sg U26475 ( .A(n31548), .B(n31549), .X(n31380) );
  nor_x2_sg U26466 ( .A(n31373), .B(n8409), .X(n31539) );
  nand_x8_sg U26465 ( .A(n31541), .B(n31542), .X(n31373) );
  nand_x8_sg U26458 ( .A(n31511), .B(n49832), .X(n31374) );
  nand_x8_sg U26453 ( .A(n31535), .B(n31536), .X(n31367) );
  nor_x2_sg U26444 ( .A(n31361), .B(n8449), .X(n31526) );
  nand_x8_sg U26436 ( .A(n31517), .B(n49827), .X(n31360) );
  nand_x8_sg U26429 ( .A(n31520), .B(n31521), .X(n31351) );
  nor_x2_sg U26724 ( .A(n31501), .B(n8370), .X(n31499) );
  nand_x8_sg U26962 ( .A(n49747), .B(n31490), .X(n24851) );
  nor_x2_sg U26958 ( .A(n31495), .B(n8371), .X(n31493) );
  nand_x8_sg U27198 ( .A(n49698), .B(n31484), .X(n24899) );
  nor_x2_sg U27194 ( .A(n31489), .B(n8372), .X(n31487) );
  nand_x8_sg U27433 ( .A(n49651), .B(n31478), .X(n24947) );
  nor_x2_sg U27429 ( .A(n31483), .B(n8373), .X(n31481) );
  nand_x8_sg U27668 ( .A(n49604), .B(n31472), .X(n24995) );
  nor_x2_sg U27664 ( .A(n31477), .B(n8374), .X(n31475) );
  nand_x8_sg U27903 ( .A(n49558), .B(n31466), .X(n25043) );
  nor_x2_sg U27899 ( .A(n31471), .B(n8375), .X(n31469) );
  nand_x8_sg U28139 ( .A(n49511), .B(n31460), .X(n25092) );
  nor_x2_sg U28135 ( .A(n31465), .B(n8376), .X(n31463) );
  nand_x8_sg U28374 ( .A(n49464), .B(n31454), .X(n25140) );
  nor_x2_sg U28370 ( .A(n31459), .B(n8377), .X(n31457) );
  nand_x8_sg U28609 ( .A(n49418), .B(n31448), .X(n25189) );
  nor_x2_sg U28605 ( .A(n31453), .B(n8378), .X(n31451) );
  nand_x8_sg U28843 ( .A(n49372), .B(n31442), .X(n25238) );
  nor_x2_sg U28839 ( .A(n31447), .B(n8379), .X(n31445) );
  nor_x2_sg U29068 ( .A(n31441), .B(n8380), .X(n31439) );
  nand_x8_sg U29077 ( .A(n31426), .B(n31427), .X(n31261) );
  nor_x2_sg U26254 ( .A(n31196), .B(n8368), .X(n31381) );
  nand_x8_sg U26253 ( .A(n31383), .B(n31384), .X(n31196) );
  nand_x8_sg U26246 ( .A(n31334), .B(n49885), .X(n24684) );
  nand_x8_sg U26241 ( .A(n31377), .B(n31378), .X(n31190) );
  nor_x2_sg U26232 ( .A(n31183), .B(n8408), .X(n31368) );
  nand_x8_sg U26231 ( .A(n31370), .B(n31371), .X(n31183) );
  nand_x8_sg U26224 ( .A(n31340), .B(n49878), .X(n31184) );
  nand_x8_sg U26219 ( .A(n31364), .B(n31365), .X(n31177) );
  nor_x2_sg U26210 ( .A(n31171), .B(n8448), .X(n31355) );
  nand_x8_sg U26209 ( .A(n31357), .B(n31358), .X(n31171) );
  nand_x8_sg U26202 ( .A(n31346), .B(n31347), .X(n31170) );
  nor_x2_sg U26190 ( .A(n31351), .B(n8469), .X(n31350) );
  nand_x8_sg U26278 ( .A(n31209), .B(n31210), .X(n31134) );
  nand_x8_sg U26504 ( .A(n49843), .B(n31322), .X(n24733) );
  nor_x2_sg U26500 ( .A(n31327), .B(n8349), .X(n31325) );
  nand_x8_sg U26511 ( .A(n31212), .B(n31213), .X(n31128) );
  nand_x8_sg U26741 ( .A(n49797), .B(n31316), .X(n24781) );
  nand_x8_sg U26748 ( .A(n31215), .B(n31216), .X(n31122) );
  nand_x8_sg U26975 ( .A(n49748), .B(n31310), .X(n24828) );
  nor_x2_sg U26971 ( .A(n49726), .B(n8351), .X(n31313) );
  nand_x8_sg U26982 ( .A(n31218), .B(n31219), .X(n31116) );
  nand_x8_sg U27211 ( .A(n49699), .B(n31304), .X(n24876) );
  nor_x2_sg U27207 ( .A(n49680), .B(n8352), .X(n31307) );
  nand_x8_sg U27218 ( .A(n31221), .B(n31222), .X(n31110) );
  nand_x8_sg U27446 ( .A(n49652), .B(n31298), .X(n24924) );
  nor_x2_sg U27442 ( .A(n42943), .B(n8353), .X(n31301) );
  nand_x8_sg U27453 ( .A(n31224), .B(n31225), .X(n31104) );
  nand_x8_sg U27681 ( .A(n49605), .B(n31292), .X(n24972) );
  nor_x2_sg U27677 ( .A(n49586), .B(n8354), .X(n31295) );
  nand_x8_sg U27688 ( .A(n31227), .B(n31228), .X(n31098) );
  nand_x8_sg U27916 ( .A(n49559), .B(n31286), .X(n25020) );
  nor_x2_sg U27912 ( .A(n49540), .B(n8355), .X(n31289) );
  nand_x8_sg U27923 ( .A(n31230), .B(n31231), .X(n31092) );
  nand_x8_sg U28152 ( .A(n49512), .B(n31280), .X(n25068) );
  nor_x2_sg U28148 ( .A(n42938), .B(n8356), .X(n31283) );
  nand_x8_sg U28159 ( .A(n31233), .B(n31234), .X(n31086) );
  nand_x8_sg U28387 ( .A(n49465), .B(n31274), .X(n25117) );
  nor_x2_sg U28383 ( .A(n49446), .B(n8357), .X(n31277) );
  nand_x8_sg U28394 ( .A(n31236), .B(n31237), .X(n31080) );
  nand_x8_sg U28622 ( .A(n49419), .B(n31268), .X(n25165) );
  nor_x2_sg U28618 ( .A(n31273), .B(n8358), .X(n31271) );
  nand_x8_sg U28629 ( .A(n31239), .B(n31240), .X(n31074) );
  nand_x8_sg U28856 ( .A(n49373), .B(n31262), .X(n25214) );
  nor_x2_sg U28852 ( .A(n31267), .B(n8359), .X(n31265) );
  nand_x8_sg U28863 ( .A(n31242), .B(n31243), .X(n31068) );
  nand_x8_sg U29082 ( .A(n31255), .B(n31256), .X(n25263) );
  nor_x2_sg U29079 ( .A(n31259), .B(n49309), .X(n31257) );
  nor_x2_sg U29078 ( .A(n31261), .B(n8360), .X(n31259) );
  nand_x8_sg U29088 ( .A(n31245), .B(n31246), .X(n31062) );
  nand_x8_sg U29270 ( .A(n31249), .B(n31250), .X(n25308) );
  nand_x8_sg U29409 ( .A(n49258), .B(n31248), .X(n25353) );
  nand_x8_sg U26032 ( .A(n49937), .B(n31138), .X(n24636) );
  nor_x2_sg U26028 ( .A(n31199), .B(n8347), .X(n31197) );
  nand_x8_sg U26020 ( .A(n49934), .B(n31141), .X(n24660) );
  nor_x2_sg U26016 ( .A(n30991), .B(n8367), .X(n31191) );
  nand_x8_sg U26015 ( .A(n31193), .B(n31194), .X(n30991) );
  nand_x8_sg U26008 ( .A(n31144), .B(n49931), .X(n24635) );
  nand_x8_sg U26003 ( .A(n31187), .B(n31188), .X(n30985) );
  nor_x2_sg U25994 ( .A(n30978), .B(n8407), .X(n31178) );
  nand_x8_sg U25993 ( .A(n31180), .B(n31181), .X(n30978) );
  nand_x8_sg U25986 ( .A(n31150), .B(n49924), .X(n30979) );
  nand_x8_sg U25981 ( .A(n31174), .B(n31175), .X(n30972) );
  nor_x2_sg U25972 ( .A(n30966), .B(n8447), .X(n31165) );
  nand_x8_sg U25964 ( .A(n31156), .B(n49919), .X(n30965) );
  nand_x8_sg U25957 ( .A(n31159), .B(n31160), .X(n30956) );
  nand_x8_sg U26049 ( .A(n31008), .B(n31009), .X(n30925) );
  nor_x2_sg U26280 ( .A(n31132), .B(n49869), .X(n31131) );
  nor_x2_sg U26279 ( .A(n31134), .B(n8328), .X(n31132) );
  nand_x8_sg U26288 ( .A(n31011), .B(n31012), .X(n30919) );
  nor_x2_sg U26513 ( .A(n31126), .B(n49821), .X(n31125) );
  nor_x2_sg U26512 ( .A(n31128), .B(n8329), .X(n31126) );
  nand_x8_sg U26521 ( .A(n31014), .B(n31015), .X(n30913) );
  nor_x2_sg U26749 ( .A(n31122), .B(n8330), .X(n31120) );
  nand_x8_sg U26758 ( .A(n31017), .B(n31018), .X(n30907) );
  nor_x2_sg U26984 ( .A(n31114), .B(n49725), .X(n31113) );
  nor_x2_sg U26983 ( .A(n31116), .B(n8331), .X(n31114) );
  nand_x8_sg U26992 ( .A(n31020), .B(n31021), .X(n30901) );
  nor_x2_sg U27220 ( .A(n31108), .B(n49678), .X(n31107) );
  nor_x2_sg U27219 ( .A(n31110), .B(n8332), .X(n31108) );
  nand_x8_sg U27228 ( .A(n31023), .B(n31024), .X(n30895) );
  nor_x2_sg U27455 ( .A(n31102), .B(n49631), .X(n31101) );
  nor_x2_sg U27454 ( .A(n31104), .B(n8333), .X(n31102) );
  nand_x8_sg U27463 ( .A(n31026), .B(n31027), .X(n30889) );
  nor_x2_sg U27690 ( .A(n31096), .B(n49585), .X(n31095) );
  nor_x2_sg U27689 ( .A(n31098), .B(n8334), .X(n31096) );
  nand_x8_sg U27698 ( .A(n31029), .B(n31030), .X(n30883) );
  nor_x2_sg U27925 ( .A(n31090), .B(n49538), .X(n31089) );
  nor_x2_sg U27924 ( .A(n31092), .B(n8335), .X(n31090) );
  nand_x8_sg U27933 ( .A(n31032), .B(n31033), .X(n30877) );
  nor_x2_sg U28161 ( .A(n31084), .B(n49491), .X(n31083) );
  nor_x2_sg U28160 ( .A(n31086), .B(n8336), .X(n31084) );
  nand_x8_sg U28169 ( .A(n31035), .B(n31036), .X(n30871) );
  nor_x2_sg U28396 ( .A(n31078), .B(n49445), .X(n31077) );
  nor_x2_sg U28395 ( .A(n31080), .B(n8337), .X(n31078) );
  nand_x8_sg U28404 ( .A(n31038), .B(n31039), .X(n30865) );
  nor_x2_sg U28631 ( .A(n31072), .B(n49399), .X(n31071) );
  nor_x2_sg U28630 ( .A(n31074), .B(n8338), .X(n31072) );
  nand_x8_sg U28639 ( .A(n31041), .B(n31042), .X(n30859) );
  nor_x2_sg U28865 ( .A(n31066), .B(n49355), .X(n31065) );
  nor_x2_sg U28864 ( .A(n31068), .B(n8339), .X(n31066) );
  nand_x8_sg U28873 ( .A(n31044), .B(n31045), .X(n30853) );
  nor_x2_sg U29090 ( .A(n31060), .B(n49307), .X(n31059) );
  nor_x2_sg U29089 ( .A(n31062), .B(n8340), .X(n31060) );
  nand_x8_sg U29097 ( .A(n31047), .B(n31048), .X(n30847) );
  nand_x8_sg U29412 ( .A(n49259), .B(n31050), .X(n25360) );
  nor_x2_sg U25808 ( .A(n30997), .B(n49939), .X(n30932) );
  nor_x2_sg U25807 ( .A(n30778), .B(n8326), .X(n30997) );
  nand_x8_sg U25806 ( .A(n30999), .B(n31000), .X(n30778) );
  nand_x8_sg U25799 ( .A(n30933), .B(n49980), .X(n24587) );
  nor_x2_sg U25782 ( .A(n30765), .B(n8366), .X(n30986) );
  nand_x8_sg U25781 ( .A(n30988), .B(n30989), .X(n30765) );
  nand_x8_sg U25774 ( .A(n30939), .B(n49975), .X(n24586) );
  nand_x8_sg U25769 ( .A(n30982), .B(n30983), .X(n30759) );
  nor_x2_sg U25760 ( .A(n30752), .B(n8406), .X(n30973) );
  nand_x8_sg U25759 ( .A(n30975), .B(n30976), .X(n30752) );
  nand_x8_sg U25752 ( .A(n30945), .B(n49968), .X(n30753) );
  nand_x8_sg U25747 ( .A(n30969), .B(n30970), .X(n30746) );
  nor_x2_sg U25738 ( .A(n30740), .B(n8446), .X(n30960) );
  nand_x8_sg U25737 ( .A(n30962), .B(n30963), .X(n30740) );
  nand_x8_sg U25730 ( .A(n30951), .B(n30952), .X(n30739) );
  nor_x2_sg U25718 ( .A(n30956), .B(n8467), .X(n30955) );
  nand_x8_sg U25830 ( .A(n30790), .B(n30791), .X(n30697) );
  nand_x8_sg U26063 ( .A(n30793), .B(n30794), .X(n30691) );
  nand_x8_sg U26300 ( .A(n30796), .B(n30797), .X(n30685) );
  nand_x8_sg U26533 ( .A(n30799), .B(n30800), .X(n30678) );
  nand_x8_sg U26770 ( .A(n30802), .B(n30803), .X(n30671) );
  nand_x8_sg U27004 ( .A(n30805), .B(n30806), .X(n30664) );
  nand_x8_sg U27240 ( .A(n30808), .B(n30809), .X(n30657) );
  nand_x8_sg U27475 ( .A(n30811), .B(n30812), .X(n30650) );
  nand_x8_sg U27710 ( .A(n30814), .B(n30815), .X(n30643) );
  nand_x8_sg U27945 ( .A(n30817), .B(n30818), .X(n30636) );
  nand_x8_sg U28181 ( .A(n30820), .B(n30821), .X(n30629) );
  nand_x8_sg U28416 ( .A(n30823), .B(n30824), .X(n30622) );
  nand_x8_sg U28651 ( .A(n30826), .B(n30827), .X(n30615) );
  nand_x8_sg U28885 ( .A(n30829), .B(n30830), .X(n30608) );
  nand_x8_sg U29108 ( .A(n30832), .B(n30833), .X(n30601) );
  nand_x8_sg U29415 ( .A(n49260), .B(n30835), .X(n25363) );
  nand_x8_sg U25579 ( .A(n30781), .B(n30782), .X(n30527) );
  nor_x2_sg U25571 ( .A(n30773), .B(n49982), .X(n30706) );
  nor_x2_sg U25570 ( .A(n30521), .B(n8325), .X(n30773) );
  nand_x8_sg U25569 ( .A(n30775), .B(n30776), .X(n30521) );
  nand_x8_sg U25562 ( .A(n50025), .B(n30707), .X(n24538) );
  nor_x2_sg U25558 ( .A(n30768), .B(n8345), .X(n30766) );
  nand_x8_sg U25550 ( .A(n50022), .B(n30710), .X(n24562) );
  nor_x2_sg U25546 ( .A(n30510), .B(n8365), .X(n30760) );
  nand_x8_sg U25545 ( .A(n30762), .B(n30763), .X(n30510) );
  nand_x8_sg U25538 ( .A(n30713), .B(n50019), .X(n24537) );
  nand_x8_sg U25533 ( .A(n30756), .B(n30757), .X(n30504) );
  nor_x2_sg U25524 ( .A(n30497), .B(n8405), .X(n30747) );
  nand_x8_sg U25523 ( .A(n30749), .B(n30750), .X(n30497) );
  nand_x8_sg U25516 ( .A(n30719), .B(n50012), .X(n30498) );
  nand_x8_sg U25511 ( .A(n30743), .B(n30744), .X(n30491) );
  nor_x2_sg U25502 ( .A(n30485), .B(n8445), .X(n30734) );
  nand_x8_sg U25501 ( .A(n30736), .B(n30737), .X(n30485) );
  nand_x8_sg U25494 ( .A(n30725), .B(n50006), .X(n30484) );
  nand_x8_sg U25487 ( .A(n30728), .B(n30729), .X(n30475) );
  nand_x8_sg U25603 ( .A(n30539), .B(n30540), .X(n30438) );
  nor_x2_sg U25832 ( .A(n30695), .B(n49959), .X(n30694) );
  nor_x2_sg U25831 ( .A(n30697), .B(n8286), .X(n30695) );
  nand_x8_sg U25840 ( .A(n30542), .B(n30543), .X(n30432) );
  nor_x2_sg U26065 ( .A(n30689), .B(n49911), .X(n30688) );
  nor_x2_sg U26064 ( .A(n30691), .B(n8287), .X(n30689) );
  nand_x8_sg U26073 ( .A(n30545), .B(n30546), .X(n30426) );
  nor_x2_sg U26301 ( .A(n30685), .B(n8288), .X(n30683) );
  nand_x8_sg U26310 ( .A(n30548), .B(n30549), .X(n30420) );
  nor_x2_sg U26534 ( .A(n30678), .B(n8289), .X(n30676) );
  nand_x8_sg U26543 ( .A(n30551), .B(n30552), .X(n30414) );
  nor_x2_sg U26771 ( .A(n30671), .B(n8290), .X(n30669) );
  nand_x8_sg U26780 ( .A(n30554), .B(n30555), .X(n30408) );
  nor_x2_sg U27005 ( .A(n30664), .B(n8291), .X(n30662) );
  nand_x8_sg U27014 ( .A(n30557), .B(n30558), .X(n30402) );
  nor_x2_sg U27241 ( .A(n30657), .B(n8292), .X(n30655) );
  nand_x8_sg U27250 ( .A(n30560), .B(n30561), .X(n30396) );
  nor_x2_sg U27476 ( .A(n30650), .B(n8293), .X(n30648) );
  nand_x8_sg U27485 ( .A(n30563), .B(n30564), .X(n30390) );
  nor_x2_sg U27711 ( .A(n30643), .B(n8294), .X(n30641) );
  nand_x8_sg U27720 ( .A(n30566), .B(n30567), .X(n30384) );
  nor_x2_sg U27946 ( .A(n30636), .B(n8295), .X(n30634) );
  nand_x8_sg U27955 ( .A(n30569), .B(n30570), .X(n30378) );
  nor_x2_sg U28182 ( .A(n30629), .B(n8296), .X(n30627) );
  nand_x8_sg U28191 ( .A(n30572), .B(n30573), .X(n30372) );
  nor_x2_sg U28417 ( .A(n30622), .B(n8297), .X(n30620) );
  nand_x8_sg U28426 ( .A(n30575), .B(n30576), .X(n30366) );
  nor_x2_sg U28652 ( .A(n30615), .B(n8298), .X(n30613) );
  nand_x8_sg U28661 ( .A(n30578), .B(n30579), .X(n30360) );
  nor_x2_sg U28886 ( .A(n30608), .B(n8299), .X(n30606) );
  nand_x8_sg U28895 ( .A(n30581), .B(n30582), .X(n30354) );
  nor_x2_sg U29109 ( .A(n30601), .B(n8300), .X(n30599) );
  nand_x8_sg U29117 ( .A(n30584), .B(n30585), .X(n30348) );
  nand_x8_sg U29418 ( .A(n49261), .B(n30587), .X(n25367) );
  nor_x2_sg U25361 ( .A(n30271), .B(n8284), .X(n30528) );
  nand_x8_sg U25360 ( .A(n30530), .B(n30531), .X(n30271) );
  nand_x8_sg U25346 ( .A(n30524), .B(n30525), .X(n30264) );
  nor_x2_sg U25338 ( .A(n30516), .B(n50027), .X(n30451) );
  nor_x2_sg U25337 ( .A(n30257), .B(n8324), .X(n30516) );
  nand_x8_sg U25336 ( .A(n30518), .B(n30519), .X(n30257) );
  nand_x8_sg U25329 ( .A(n50067), .B(n30452), .X(n24488) );
  nor_x2_sg U25312 ( .A(n30242), .B(n8364), .X(n30505) );
  nand_x8_sg U25311 ( .A(n30507), .B(n30508), .X(n30242) );
  nand_x8_sg U25304 ( .A(n30458), .B(n50062), .X(n24487) );
  nand_x8_sg U25299 ( .A(n30501), .B(n30502), .X(n30235) );
  nor_x2_sg U25290 ( .A(n30228), .B(n8404), .X(n30492) );
  nand_x8_sg U25289 ( .A(n30494), .B(n30495), .X(n30228) );
  nand_x8_sg U25282 ( .A(n30464), .B(n50056), .X(n30227) );
  nand_x8_sg U25277 ( .A(n30488), .B(n30489), .X(n30220) );
  nor_x2_sg U25268 ( .A(n30213), .B(n8444), .X(n30479) );
  nand_x8_sg U25267 ( .A(n30481), .B(n30482), .X(n30213) );
  nor_x2_sg U25248 ( .A(n30475), .B(n8465), .X(n30474) );
  nand_x8_sg U25382 ( .A(n30285), .B(n30286), .X(n29849) );
  nand_x8_sg U25608 ( .A(n30434), .B(n50034), .X(n24554) );
  nand_x8_sg U25615 ( .A(n30288), .B(n30289), .X(n30015) );
  nand_x8_sg U25845 ( .A(n30428), .B(n49987), .X(n24603) );
  nand_x8_sg U25852 ( .A(n30291), .B(n30292), .X(n30162) );
  nand_x8_sg U26078 ( .A(n30422), .B(n49942), .X(n24652) );
  nand_x8_sg U26085 ( .A(n30294), .B(n30295), .X(n30156) );
  nand_x8_sg U26315 ( .A(n30416), .B(n49894), .X(n24700) );
  nand_x8_sg U26322 ( .A(n30297), .B(n30298), .X(n30150) );
  nand_x8_sg U26548 ( .A(n30410), .B(n49847), .X(n24748) );
  nand_x8_sg U26555 ( .A(n30300), .B(n30301), .X(n30144) );
  nand_x8_sg U26785 ( .A(n30404), .B(n49800), .X(n24796) );
  nand_x8_sg U26792 ( .A(n30303), .B(n30304), .X(n30138) );
  nand_x8_sg U27019 ( .A(n30398), .B(n49752), .X(n24843) );
  nand_x8_sg U27026 ( .A(n30306), .B(n30307), .X(n30132) );
  nand_x8_sg U27255 ( .A(n30392), .B(n49703), .X(n24891) );
  nand_x8_sg U27262 ( .A(n30309), .B(n30310), .X(n30126) );
  nand_x8_sg U27490 ( .A(n30386), .B(n49656), .X(n24939) );
  nand_x8_sg U27497 ( .A(n30312), .B(n30313), .X(n30120) );
  nand_x8_sg U27725 ( .A(n30380), .B(n49609), .X(n24987) );
  nand_x8_sg U27732 ( .A(n30315), .B(n30316), .X(n30114) );
  nand_x8_sg U27960 ( .A(n30374), .B(n49563), .X(n25035) );
  nand_x8_sg U27967 ( .A(n30318), .B(n30319), .X(n30108) );
  nand_x8_sg U28196 ( .A(n30368), .B(n49516), .X(n25083) );
  nand_x8_sg U28203 ( .A(n30321), .B(n30322), .X(n30102) );
  nand_x8_sg U28431 ( .A(n30362), .B(n49469), .X(n25132) );
  nand_x8_sg U28438 ( .A(n30324), .B(n30325), .X(n30096) );
  nand_x8_sg U28666 ( .A(n30356), .B(n49423), .X(n25180) );
  nand_x8_sg U28673 ( .A(n30327), .B(n30328), .X(n30090) );
  nand_x8_sg U28900 ( .A(n30350), .B(n49377), .X(n25229) );
  nand_x8_sg U28907 ( .A(n30330), .B(n30331), .X(n30084) );
  nand_x8_sg U29122 ( .A(n30344), .B(n49333), .X(n25278) );
  nand_x8_sg U29128 ( .A(n30333), .B(n30334), .X(n30078) );
  nand_x8_sg U29298 ( .A(n30337), .B(n30338), .X(n25321) );
  nand_x8_sg U29421 ( .A(n49262), .B(n30336), .X(n25364) );
  nor_x2_sg U25101 ( .A(n30253), .B(n8323), .X(n30251) );
  nor_x2_sg U25089 ( .A(n30245), .B(n8343), .X(n30243) );
  nor_x2_sg U25078 ( .A(n30238), .B(n8363), .X(n30236) );
  nor_x2_sg U24995 ( .A(n9406), .B(n29636), .X(n29635) );
  nor_x2_sg U25209 ( .A(n29660), .B(n8204), .X(n29856) );
  nand_x8_sg U25208 ( .A(n29858), .B(n29859), .X(n29660) );
  nand_x8_sg U25438 ( .A(n30007), .B(n50038), .X(n29834) );
  nand_x8_sg U25433 ( .A(n30018), .B(n30019), .X(n29855) );
  nor_x2_sg U25854 ( .A(n30160), .B(n49955), .X(n30159) );
  nor_x2_sg U25853 ( .A(n30162), .B(n8246), .X(n30160) );
  nand_x8_sg U25666 ( .A(n30021), .B(n30022), .X(n30005) );
  nor_x2_sg U26087 ( .A(n30154), .B(n49907), .X(n30153) );
  nor_x2_sg U26086 ( .A(n30156), .B(n8247), .X(n30154) );
  nand_x8_sg U25903 ( .A(n30024), .B(n30025), .X(n29999) );
  nor_x2_sg U26324 ( .A(n30148), .B(n49860), .X(n30147) );
  nor_x2_sg U26323 ( .A(n30150), .B(n8248), .X(n30148) );
  nand_x8_sg U26136 ( .A(n30027), .B(n30028), .X(n29993) );
  nor_x2_sg U26557 ( .A(n30142), .B(n49812), .X(n30141) );
  nor_x2_sg U26556 ( .A(n30144), .B(n8249), .X(n30142) );
  nand_x8_sg U26373 ( .A(n30030), .B(n30031), .X(n29987) );
  nor_x2_sg U26793 ( .A(n30138), .B(n8250), .X(n30136) );
  nand_x8_sg U26606 ( .A(n30033), .B(n30034), .X(n29981) );
  nor_x2_sg U27028 ( .A(n30130), .B(n49716), .X(n30129) );
  nor_x2_sg U27027 ( .A(n30132), .B(n8251), .X(n30130) );
  nand_x8_sg U26843 ( .A(n30036), .B(n30037), .X(n29975) );
  nor_x2_sg U27264 ( .A(n30124), .B(n49669), .X(n30123) );
  nor_x2_sg U27263 ( .A(n30126), .B(n8252), .X(n30124) );
  nand_x8_sg U27077 ( .A(n30039), .B(n30040), .X(n29969) );
  nor_x2_sg U27499 ( .A(n30118), .B(n49622), .X(n30117) );
  nor_x2_sg U27498 ( .A(n30120), .B(n8253), .X(n30118) );
  nand_x8_sg U27313 ( .A(n30042), .B(n30043), .X(n29963) );
  nor_x2_sg U27734 ( .A(n30112), .B(n49576), .X(n30111) );
  nor_x2_sg U27733 ( .A(n30114), .B(n8254), .X(n30112) );
  nand_x8_sg U27548 ( .A(n30045), .B(n30046), .X(n29957) );
  nor_x2_sg U27969 ( .A(n30106), .B(n49529), .X(n30105) );
  nor_x2_sg U27968 ( .A(n30108), .B(n8255), .X(n30106) );
  nand_x8_sg U27782 ( .A(n30048), .B(n30049), .X(n29951) );
  nor_x2_sg U28205 ( .A(n30100), .B(n49482), .X(n30099) );
  nor_x2_sg U28204 ( .A(n30102), .B(n8256), .X(n30100) );
  nand_x8_sg U28017 ( .A(n30051), .B(n30052), .X(n29945) );
  nor_x2_sg U28440 ( .A(n30094), .B(n49436), .X(n30093) );
  nor_x2_sg U28439 ( .A(n30096), .B(n8257), .X(n30094) );
  nand_x8_sg U28253 ( .A(n30054), .B(n30055), .X(n29939) );
  nor_x2_sg U28675 ( .A(n30088), .B(n49390), .X(n30087) );
  nor_x2_sg U28674 ( .A(n30090), .B(n8258), .X(n30088) );
  nand_x8_sg U28488 ( .A(n30057), .B(n30058), .X(n29933) );
  nor_x2_sg U28909 ( .A(n30082), .B(n49346), .X(n30081) );
  nor_x2_sg U28908 ( .A(n30084), .B(n8259), .X(n30082) );
  nand_x8_sg U28723 ( .A(n30060), .B(n30061), .X(n29927) );
  nor_x2_sg U29130 ( .A(n30076), .B(n49301), .X(n30075) );
  nor_x2_sg U29129 ( .A(n30078), .B(n8260), .X(n30076) );
  nand_x8_sg U28956 ( .A(n30063), .B(n30064), .X(n29921) );
  nand_x8_sg U29424 ( .A(n49263), .B(n30066), .X(n25385) );
  nor_x2_sg U25617 ( .A(n30013), .B(n49999), .X(n30012) );
  nor_x2_sg U25616 ( .A(n30015), .B(n8245), .X(n30013) );
  nand_x8_sg U25445 ( .A(n29861), .B(n29862), .X(n29837) );
  nand_x8_sg U25678 ( .A(n29864), .B(n29865), .X(n29830) );
  nand_x8_sg U25915 ( .A(n29867), .B(n29868), .X(n29823) );
  nand_x8_sg U26148 ( .A(n29870), .B(n29871), .X(n29816) );
  nand_x8_sg U26385 ( .A(n29873), .B(n29874), .X(n29809) );
  nand_x8_sg U26618 ( .A(n29876), .B(n29877), .X(n29802) );
  nand_x8_sg U26855 ( .A(n29879), .B(n29880), .X(n29795) );
  nand_x8_sg U27089 ( .A(n29882), .B(n29883), .X(n29788) );
  nand_x8_sg U27325 ( .A(n29885), .B(n29886), .X(n29781) );
  nand_x8_sg U27560 ( .A(n29888), .B(n29889), .X(n29774) );
  nand_x8_sg U27794 ( .A(n29891), .B(n29892), .X(n29767) );
  nand_x8_sg U28029 ( .A(n29894), .B(n29895), .X(n29760) );
  nand_x8_sg U28265 ( .A(n29897), .B(n29898), .X(n29753) );
  nand_x8_sg U28500 ( .A(n29900), .B(n29901), .X(n29746) );
  nand_x8_sg U28735 ( .A(n29903), .B(n29904), .X(n29739) );
  nand_x8_sg U28967 ( .A(n29906), .B(n29907), .X(n29732) );
  nand_x8_sg U29427 ( .A(n49264), .B(n29909), .X(n25386) );
  nand_x8_sg U25194 ( .A(n29852), .B(n29853), .X(n29653) );
  nor_x2_sg U25384 ( .A(n29847), .B(n50047), .X(n29846) );
  nor_x2_sg U25383 ( .A(n29849), .B(n8244), .X(n29847) );
  nand_x8_sg U25218 ( .A(n29667), .B(n29668), .X(n24521) );
  nor_x2_sg U25446 ( .A(n29837), .B(n8205), .X(n29835) );
  nand_x8_sg U25455 ( .A(n29670), .B(n29671), .X(n24570) );
  nor_x2_sg U25679 ( .A(n29830), .B(n8206), .X(n29828) );
  nand_x8_sg U25688 ( .A(n29673), .B(n29674), .X(n24619) );
  nor_x2_sg U25916 ( .A(n29823), .B(n8207), .X(n29821) );
  nand_x8_sg U25925 ( .A(n29676), .B(n29677), .X(n24668) );
  nor_x2_sg U26149 ( .A(n29816), .B(n8208), .X(n29814) );
  nand_x8_sg U26158 ( .A(n29679), .B(n29680), .X(n24716) );
  nor_x2_sg U26386 ( .A(n29809), .B(n8209), .X(n29807) );
  nand_x8_sg U26395 ( .A(n29682), .B(n29683), .X(n24764) );
  nor_x2_sg U26619 ( .A(n29802), .B(n8210), .X(n29800) );
  nand_x8_sg U26628 ( .A(n29685), .B(n29686), .X(n24811) );
  nor_x2_sg U26856 ( .A(n29795), .B(n8211), .X(n29793) );
  nand_x8_sg U26865 ( .A(n29688), .B(n29689), .X(n24859) );
  nor_x2_sg U27090 ( .A(n29788), .B(n8212), .X(n29786) );
  nand_x8_sg U27099 ( .A(n29691), .B(n29692), .X(n24907) );
  nor_x2_sg U27326 ( .A(n29781), .B(n8213), .X(n29779) );
  nand_x8_sg U27335 ( .A(n29694), .B(n29695), .X(n24955) );
  nor_x2_sg U27561 ( .A(n29774), .B(n8214), .X(n29772) );
  nand_x8_sg U27570 ( .A(n29697), .B(n29698), .X(n25003) );
  nor_x2_sg U27795 ( .A(n29767), .B(n8215), .X(n29765) );
  nand_x8_sg U27804 ( .A(n29700), .B(n29701), .X(n25051) );
  nor_x2_sg U28030 ( .A(n29760), .B(n8216), .X(n29758) );
  nand_x8_sg U28039 ( .A(n29703), .B(n29704), .X(n25100) );
  nor_x2_sg U28266 ( .A(n29753), .B(n8217), .X(n29751) );
  nand_x8_sg U28275 ( .A(n29706), .B(n29707), .X(n25148) );
  nor_x2_sg U28501 ( .A(n29746), .B(n8218), .X(n29744) );
  nand_x8_sg U28510 ( .A(n29709), .B(n29710), .X(n25197) );
  nor_x2_sg U28736 ( .A(n29739), .B(n8219), .X(n29737) );
  nand_x8_sg U28745 ( .A(n29712), .B(n29713), .X(n25246) );
  nor_x2_sg U28968 ( .A(n29732), .B(n8220), .X(n29730) );
  nand_x8_sg U28976 ( .A(n29715), .B(n29716), .X(n25293) );
  nand_x8_sg U29355 ( .A(n49265), .B(n29718), .X(n25371) );
  nor_x2_sg U24947 ( .A(n9392), .B(n29615), .X(n29614) );
  nor_x2_sg U24937 ( .A(n9365), .B(n29594), .X(n29590) );
  nor_x2_sg U24936 ( .A(n9371), .B(n29592), .X(n29591) );
  nor_x2_sg U24931 ( .A(n29578), .B(n29579), .X(n29577) );
  nand_x8_sg U29617 ( .A(n46235), .B(n25388), .X(n24473) );
  nor_x2_sg U25224 ( .A(n9406), .B(n24516), .X(n24515) );
  nor_x2_sg U25175 ( .A(n9392), .B(n24505), .X(n24504) );
  nor_x2_sg U25165 ( .A(n9365), .B(n24488), .X(n24485) );
  nor_x2_sg U25164 ( .A(n9371), .B(n24487), .X(n24486) );
  nor_x2_sg U25159 ( .A(n24474), .B(n24475), .X(n24472) );
  nor_x2_sg U25461 ( .A(n9406), .B(n24565), .X(n24564) );
  nor_x2_sg U25411 ( .A(n9392), .B(n24554), .X(n24553) );
  nor_x2_sg U25401 ( .A(n9365), .B(n24538), .X(n24535) );
  nor_x2_sg U25400 ( .A(n9371), .B(n24537), .X(n24536) );
  nor_x2_sg U25395 ( .A(n24525), .B(n24526), .X(n24524) );
  nor_x2_sg U25694 ( .A(n9406), .B(n24614), .X(n24613) );
  nor_x2_sg U25644 ( .A(n9392), .B(n24603), .X(n24602) );
  nor_x2_sg U25634 ( .A(n9365), .B(n24587), .X(n24584) );
  nor_x2_sg U25633 ( .A(n9371), .B(n24586), .X(n24585) );
  nor_x2_sg U25628 ( .A(n24574), .B(n24575), .X(n24573) );
  nor_x2_sg U25931 ( .A(n9406), .B(n24663), .X(n24662) );
  nor_x2_sg U25881 ( .A(n9392), .B(n24652), .X(n24651) );
  nor_x2_sg U25871 ( .A(n9365), .B(n24636), .X(n24633) );
  nor_x2_sg U25870 ( .A(n9371), .B(n24635), .X(n24634) );
  nor_x2_sg U25865 ( .A(n24623), .B(n24624), .X(n24622) );
  nor_x2_sg U26164 ( .A(n9406), .B(n24711), .X(n24710) );
  nor_x2_sg U26114 ( .A(n9392), .B(n24700), .X(n24699) );
  nor_x2_sg U26104 ( .A(n9365), .B(n24685), .X(n24682) );
  nor_x2_sg U26103 ( .A(n9371), .B(n24684), .X(n24683) );
  nor_x2_sg U26098 ( .A(n24672), .B(n24673), .X(n24671) );
  nor_x2_sg U26401 ( .A(n9406), .B(n24759), .X(n24758) );
  nor_x2_sg U26351 ( .A(n9392), .B(n24748), .X(n24747) );
  nor_x2_sg U26341 ( .A(n9365), .B(n24733), .X(n24730) );
  nor_x2_sg U26340 ( .A(n9371), .B(n24732), .X(n24731) );
  nor_x2_sg U26335 ( .A(n24720), .B(n24721), .X(n24719) );
  nor_x2_sg U26634 ( .A(n9406), .B(n24806), .X(n24805) );
  nor_x2_sg U26584 ( .A(n9392), .B(n24796), .X(n24795) );
  nor_x2_sg U26574 ( .A(n9365), .B(n24781), .X(n24778) );
  nor_x2_sg U26573 ( .A(n9371), .B(n24780), .X(n24779) );
  nor_x2_sg U26568 ( .A(n24768), .B(n24769), .X(n24767) );
  nor_x2_sg U26871 ( .A(n9406), .B(n24854), .X(n24853) );
  nor_x2_sg U26821 ( .A(n9392), .B(n24843), .X(n24842) );
  nor_x2_sg U26811 ( .A(n9365), .B(n24828), .X(n24825) );
  nor_x2_sg U26810 ( .A(n9371), .B(n24827), .X(n24826) );
  nor_x2_sg U26805 ( .A(n24815), .B(n24816), .X(n24814) );
  nor_x2_sg U27105 ( .A(n9406), .B(n24902), .X(n24901) );
  nor_x2_sg U27055 ( .A(n9392), .B(n24891), .X(n24890) );
  nor_x2_sg U27045 ( .A(n9365), .B(n24876), .X(n24873) );
  nor_x2_sg U27044 ( .A(n9371), .B(n24875), .X(n24874) );
  nor_x2_sg U27039 ( .A(n24863), .B(n24864), .X(n24862) );
  nor_x2_sg U27341 ( .A(n9406), .B(n24950), .X(n24949) );
  nor_x2_sg U27291 ( .A(n9392), .B(n24939), .X(n24938) );
  nor_x2_sg U27281 ( .A(n9365), .B(n24924), .X(n24921) );
  nor_x2_sg U27280 ( .A(n9371), .B(n24923), .X(n24922) );
  nor_x2_sg U27275 ( .A(n24911), .B(n24912), .X(n24910) );
  nor_x2_sg U27576 ( .A(n9406), .B(n24998), .X(n24997) );
  nor_x2_sg U27526 ( .A(n9392), .B(n24987), .X(n24986) );
  nor_x2_sg U27516 ( .A(n9365), .B(n24972), .X(n24969) );
  nor_x2_sg U27515 ( .A(n9371), .B(n24971), .X(n24970) );
  nor_x2_sg U27510 ( .A(n24959), .B(n24960), .X(n24958) );
  nor_x2_sg U27810 ( .A(n9406), .B(n25046), .X(n25045) );
  nor_x2_sg U27761 ( .A(n9392), .B(n25035), .X(n25034) );
  nor_x2_sg U27751 ( .A(n9365), .B(n25020), .X(n25017) );
  nor_x2_sg U27750 ( .A(n9371), .B(n25019), .X(n25018) );
  nor_x2_sg U27745 ( .A(n25007), .B(n25008), .X(n25006) );
  nor_x2_sg U28045 ( .A(n9406), .B(n25095), .X(n25094) );
  nor_x2_sg U27996 ( .A(n9392), .B(n25083), .X(n25082) );
  nor_x2_sg U27986 ( .A(n9365), .B(n25068), .X(n25065) );
  nor_x2_sg U27985 ( .A(n9371), .B(n25067), .X(n25066) );
  nor_x2_sg U27980 ( .A(n25055), .B(n25056), .X(n25054) );
  nor_x2_sg U28281 ( .A(n9406), .B(n25143), .X(n25142) );
  nor_x2_sg U28232 ( .A(n9392), .B(n25132), .X(n25131) );
  nor_x2_sg U28222 ( .A(n9365), .B(n25117), .X(n25114) );
  nor_x2_sg U28221 ( .A(n9371), .B(n25116), .X(n25115) );
  nor_x2_sg U28216 ( .A(n25104), .B(n25105), .X(n25103) );
  nor_x2_sg U28516 ( .A(n9406), .B(n25192), .X(n25191) );
  nor_x2_sg U28467 ( .A(n9392), .B(n25180), .X(n25179) );
  nor_x2_sg U28457 ( .A(n9365), .B(n25165), .X(n25162) );
  nor_x2_sg U28456 ( .A(n9371), .B(n25164), .X(n25163) );
  nor_x2_sg U28451 ( .A(n25152), .B(n25153), .X(n25151) );
  nor_x2_sg U28751 ( .A(n9406), .B(n25241), .X(n25240) );
  nor_x2_sg U28702 ( .A(n9392), .B(n25229), .X(n25228) );
  nor_x2_sg U28692 ( .A(n9365), .B(n25214), .X(n25211) );
  nor_x2_sg U28691 ( .A(n9371), .B(n25213), .X(n25212) );
  nor_x2_sg U28686 ( .A(n25201), .B(n25202), .X(n25200) );
  nor_x2_sg U28982 ( .A(n9406), .B(n25288), .X(n25287) );
  nor_x2_sg U28936 ( .A(n9392), .B(n25278), .X(n25277) );
  nor_x2_sg U28926 ( .A(n9365), .B(n25263), .X(n25260) );
  nor_x2_sg U28925 ( .A(n9371), .B(n25262), .X(n25261) );
  nor_x2_sg U28920 ( .A(n25250), .B(n25251), .X(n25249) );
  nor_x2_sg U29197 ( .A(n9406), .B(n25331), .X(n25330) );
  nor_x2_sg U29160 ( .A(n9392), .B(n25321), .X(n25320) );
  nor_x2_sg U29147 ( .A(n9365), .B(n25308), .X(n25305) );
  nor_x2_sg U29146 ( .A(n9371), .B(n25307), .X(n25306) );
  nor_x2_sg U29141 ( .A(n25297), .B(n25298), .X(n25296) );
  nor_x2_sg U29430 ( .A(n10281), .B(n25386), .X(n25383) );
  nor_x2_sg U29374 ( .A(n9415), .B(n25385), .X(n25384) );
  nor_x2_sg U29357 ( .A(n9406), .B(n25373), .X(n25368) );
  nor_x2_sg U29339 ( .A(n9392), .B(n25364), .X(n25361) );
  nor_x2_sg U29336 ( .A(n10256), .B(n25363), .X(n25362) );
  nor_x2_sg U29327 ( .A(n9365), .B(n25353), .X(n25350) );
  nor_x2_sg U29324 ( .A(n9371), .B(n25352), .X(n25351) );
  nor_x2_sg U29321 ( .A(n9367), .B(n25349), .X(n25346) );
  nor_x2_sg U29319 ( .A(n9373), .B(n25348), .X(n25347) );
  nor_x2_sg U29315 ( .A(n25340), .B(n25341), .X(n25339) );
  nor_x2_sg U29445 ( .A(n46232), .B(n46572), .X(n25393) );
  nor_x2_sg U29759 ( .A(n25621), .B(n25622), .X(n25620) );
  nor_x2_sg U29443 ( .A(n10283), .B(n46231), .X(n25392) );
  nor_x2_sg U29452 ( .A(n46231), .B(n25400), .X(n25399) );
  nor_x2_sg U29465 ( .A(n46567), .B(n46232), .X(n25409) );
  nor_x2_sg U29462 ( .A(n46231), .B(n25407), .X(n25406) );
  nor_x2_sg U29475 ( .A(n46564), .B(n46232), .X(n25416) );
  nor_x2_sg U29472 ( .A(n46231), .B(n25414), .X(n25413) );
  nor_x2_sg U29486 ( .A(n51280), .B(n46232), .X(n25424) );
  nand_x8_sg U29734 ( .A(n51278), .B(n46563), .X(n25423) );
  nor_x2_sg U29482 ( .A(n46231), .B(n25421), .X(n25420) );
  nor_x2_sg U29495 ( .A(n51293), .B(n46232), .X(n25431) );
  nor_x2_sg U29493 ( .A(n46231), .B(n25430), .X(n25429) );
  nand_x8_sg U29738 ( .A(n51316), .B(n46559), .X(n25442) );
  nor_x2_sg U29523 ( .A(n46232), .B(n51334), .X(n25452) );
  nor_x2_sg U29521 ( .A(n10655), .B(n25451), .X(n25450) );
  nor_x2_sg U29540 ( .A(n10660), .B(n25466), .X(n25465) );
  nor_x2_sg U29559 ( .A(n10782), .B(n25480), .X(n25479) );
  nor_x2_sg U29745 ( .A(n25485), .B(n51458), .X(n25492) );
  nor_x2_sg U29578 ( .A(n10923), .B(n25494), .X(n25493) );
  nor_x2_sg U29589 ( .A(n10919), .B(n25500), .X(n25498) );
  nor_x2_sg U29596 ( .A(n46232), .B(n41260), .X(n25504) );
  nor_x2_sg U29897 ( .A(n46552), .B(n46236), .X(n25668) );
  nor_x2_sg U29903 ( .A(n46230), .B(n46547), .X(n25673) );
  nor_x2_sg U30217 ( .A(n25902), .B(n25903), .X(n25901) );
  nor_x2_sg U29901 ( .A(n11051), .B(n46229), .X(n25672) );
  nor_x2_sg U29913 ( .A(n46230), .B(n51537), .X(n25681) );
  nor_x2_sg U29910 ( .A(n46229), .B(n25679), .X(n25678) );
  nor_x2_sg U29923 ( .A(n51543), .B(n46230), .X(n25688) );
  nor_x2_sg U29920 ( .A(n46229), .B(n25686), .X(n25685) );
  nor_x2_sg U29933 ( .A(n46540), .B(n46230), .X(n25695) );
  nor_x2_sg U29930 ( .A(n46229), .B(n25693), .X(n25692) );
  nor_x2_sg U29943 ( .A(n46539), .B(n46230), .X(n25703) );
  nor_x2_sg U29940 ( .A(n46229), .B(n25700), .X(n25699) );
  nor_x2_sg U29952 ( .A(n46536), .B(n46230), .X(n25710) );
  nor_x2_sg U29950 ( .A(n46229), .B(n25709), .X(n25708) );
  nand_x8_sg U30196 ( .A(n51588), .B(n46535), .X(n25721) );
  nor_x2_sg U29980 ( .A(n46230), .B(n46532), .X(n25731) );
  nor_x2_sg U29978 ( .A(n11434), .B(n25730), .X(n25729) );
  nor_x2_sg U29997 ( .A(n11438), .B(n25744), .X(n25743) );
  nor_x2_sg U30016 ( .A(n11638), .B(n25758), .X(n25757) );
  nor_x2_sg U30031 ( .A(n25761), .B(n25762), .X(n25760) );
  nor_x2_sg U30035 ( .A(n11768), .B(n25772), .X(n25771) );
  nor_x2_sg U30046 ( .A(n11703), .B(n25778), .X(n25776) );
  nor_x2_sg U30053 ( .A(n46230), .B(n41274), .X(n25782) );
  nor_x2_sg U30068 ( .A(n25793), .B(n51807), .X(n25790) );
  nand_x8_sg U30345 ( .A(n25910), .B(n25911), .X(n25793) );
  nor_x2_sg U30347 ( .A(n25798), .B(n25795), .X(n25797) );
  nor_x2_sg U30351 ( .A(n46528), .B(n46236), .X(n25946) );
  nor_x2_sg U30357 ( .A(n46228), .B(n46525), .X(n25951) );
  nor_x2_sg U30678 ( .A(n26182), .B(n26183), .X(n26181) );
  nor_x2_sg U30355 ( .A(n11834), .B(n46227), .X(n25950) );
  nor_x2_sg U30367 ( .A(n46228), .B(n51819), .X(n25959) );
  nor_x2_sg U30364 ( .A(n46227), .B(n25957), .X(n25956) );
  nor_x2_sg U30377 ( .A(n51826), .B(n46228), .X(n25966) );
  nor_x2_sg U30374 ( .A(n46227), .B(n25964), .X(n25963) );
  nor_x2_sg U30387 ( .A(n46517), .B(n46228), .X(n25973) );
  nor_x2_sg U30384 ( .A(n46227), .B(n25971), .X(n25970) );
  nor_x2_sg U30398 ( .A(n51839), .B(n46228), .X(n25981) );
  nand_x8_sg U30653 ( .A(n51837), .B(n46516), .X(n25980) );
  nor_x2_sg U30394 ( .A(n46227), .B(n25978), .X(n25977) );
  nor_x2_sg U30407 ( .A(n51854), .B(n46228), .X(n25988) );
  nor_x2_sg U30405 ( .A(n46227), .B(n25987), .X(n25986) );
  nand_x8_sg U30657 ( .A(n51876), .B(n46512), .X(n25999) );
  nor_x2_sg U30435 ( .A(n46228), .B(n51896), .X(n26009) );
  nor_x2_sg U30433 ( .A(n12214), .B(n26008), .X(n26007) );
  nor_x2_sg U30452 ( .A(n12218), .B(n26022), .X(n26021) );
  nor_x2_sg U30471 ( .A(n12344), .B(n26036), .X(n26035) );
  nor_x2_sg U30486 ( .A(n26039), .B(n26040), .X(n26038) );
  nor_x2_sg U30664 ( .A(n26041), .B(n52038), .X(n26048) );
  nor_x2_sg U30490 ( .A(n26050), .B(n26051), .X(n26049) );
  nor_x2_sg U30501 ( .A(n12482), .B(n26057), .X(n26055) );
  nor_x2_sg U30508 ( .A(n46228), .B(n41272), .X(n26061) );
  nor_x2_sg U30523 ( .A(n26072), .B(n52083), .X(n26069) );
  nand_x8_sg U30806 ( .A(n26190), .B(n26191), .X(n26072) );
  nor_x2_sg U30808 ( .A(n26080), .B(n26074), .X(n26077) );
  nor_x2_sg U30812 ( .A(n46508), .B(n46236), .X(n26227) );
  nor_x2_sg U30818 ( .A(n46226), .B(n46503), .X(n26232) );
  nor_x2_sg U31136 ( .A(n26461), .B(n26462), .X(n26460) );
  nor_x2_sg U30816 ( .A(n12612), .B(n46225), .X(n26231) );
  nor_x2_sg U30828 ( .A(n46226), .B(n46500), .X(n26240) );
  nor_x2_sg U30825 ( .A(n46225), .B(n26238), .X(n26237) );
  nor_x2_sg U30838 ( .A(n52100), .B(n46226), .X(n26247) );
  nor_x2_sg U30835 ( .A(n46225), .B(n26245), .X(n26244) );
  nor_x2_sg U30848 ( .A(n46496), .B(n46226), .X(n26254) );
  nor_x2_sg U30845 ( .A(n46225), .B(n26252), .X(n26251) );
  nor_x2_sg U30858 ( .A(n46495), .B(n46226), .X(n26262) );
  nor_x2_sg U30855 ( .A(n46225), .B(n26259), .X(n26258) );
  nor_x2_sg U30867 ( .A(n52133), .B(n46226), .X(n26269) );
  nor_x2_sg U30865 ( .A(n46225), .B(n26268), .X(n26267) );
  nand_x8_sg U31115 ( .A(n52146), .B(n46491), .X(n26280) );
  nor_x2_sg U30895 ( .A(n46226), .B(n46488), .X(n26290) );
  nor_x2_sg U30893 ( .A(n12995), .B(n26289), .X(n26288) );
  nor_x2_sg U30912 ( .A(n12999), .B(n26303), .X(n26302) );
  nor_x2_sg U30931 ( .A(n13200), .B(n26317), .X(n26316) );
  nor_x2_sg U31122 ( .A(n26322), .B(n52314), .X(n26329) );
  nor_x2_sg U30950 ( .A(n26331), .B(n26332), .X(n26330) );
  nor_x2_sg U30961 ( .A(n13263), .B(n26338), .X(n26336) );
  nor_x2_sg U30968 ( .A(n46226), .B(n41270), .X(n26342) );
  nor_x2_sg U30983 ( .A(n26353), .B(n52361), .X(n26350) );
  nand_x8_sg U31264 ( .A(n26469), .B(n26470), .X(n26353) );
  nor_x2_sg U31266 ( .A(n26359), .B(n26355), .X(n26357) );
  nor_x2_sg U31270 ( .A(n46485), .B(n46236), .X(n26506) );
  nor_x2_sg U31277 ( .A(n46224), .B(n46481), .X(n26511) );
  nor_x2_sg U31595 ( .A(n26739), .B(n26740), .X(n26738) );
  nor_x2_sg U31275 ( .A(n13396), .B(n46223), .X(n26510) );
  nor_x2_sg U31287 ( .A(n46224), .B(n46478), .X(n26519) );
  nor_x2_sg U31284 ( .A(n46223), .B(n26517), .X(n26516) );
  nor_x2_sg U31297 ( .A(n52378), .B(n46224), .X(n26526) );
  nor_x2_sg U31294 ( .A(n46223), .B(n26524), .X(n26523) );
  nor_x2_sg U31307 ( .A(n46474), .B(n46224), .X(n26533) );
  nor_x2_sg U31304 ( .A(n46223), .B(n26531), .X(n26530) );
  nor_x2_sg U31318 ( .A(n52391), .B(n46224), .X(n26541) );
  nand_x8_sg U31570 ( .A(n52389), .B(n46473), .X(n26540) );
  nor_x2_sg U31314 ( .A(n46223), .B(n26538), .X(n26537) );
  nor_x2_sg U31327 ( .A(n52406), .B(n46224), .X(n26548) );
  nor_x2_sg U31325 ( .A(n46223), .B(n26547), .X(n26546) );
  nand_x8_sg U31574 ( .A(n52427), .B(n46467), .X(n26559) );
  nor_x2_sg U31355 ( .A(n46224), .B(n52447), .X(n26569) );
  nor_x2_sg U31353 ( .A(n13775), .B(n26568), .X(n26567) );
  nor_x2_sg U31372 ( .A(n13779), .B(n26582), .X(n26581) );
  nor_x2_sg U31391 ( .A(n13980), .B(n26596), .X(n26595) );
  nor_x2_sg U31581 ( .A(n26601), .B(n52589), .X(n26608) );
  nor_x2_sg U31410 ( .A(n26610), .B(n26611), .X(n26609) );
  nor_x2_sg U31421 ( .A(n14043), .B(n26617), .X(n26615) );
  nor_x2_sg U31428 ( .A(n46224), .B(n41268), .X(n26621) );
  nor_x2_sg U31443 ( .A(n26632), .B(n52636), .X(n26629) );
  nand_x8_sg U31723 ( .A(n26747), .B(n26748), .X(n26632) );
  nor_x2_sg U31725 ( .A(n26637), .B(n26634), .X(n26636) );
  nor_x2_sg U31729 ( .A(n46463), .B(n46236), .X(n26784) );
  nor_x2_sg U31735 ( .A(n46222), .B(n46458), .X(n26789) );
  nor_x2_sg U32047 ( .A(n27018), .B(n27019), .X(n27017) );
  nor_x2_sg U31733 ( .A(n14175), .B(n46221), .X(n26788) );
  nor_x2_sg U31745 ( .A(n46222), .B(n52648), .X(n26797) );
  nor_x2_sg U31742 ( .A(n46221), .B(n26795), .X(n26794) );
  nor_x2_sg U31755 ( .A(n52655), .B(n46222), .X(n26804) );
  nor_x2_sg U31752 ( .A(n46221), .B(n26802), .X(n26801) );
  nor_x2_sg U31765 ( .A(n46450), .B(n46222), .X(n26811) );
  nor_x2_sg U31762 ( .A(n46221), .B(n26809), .X(n26808) );
  nor_x2_sg U31776 ( .A(n52670), .B(n46222), .X(n26819) );
  nand_x8_sg U32022 ( .A(n52667), .B(n46449), .X(n26818) );
  nor_x2_sg U31772 ( .A(n46221), .B(n26816), .X(n26815) );
  nor_x2_sg U31785 ( .A(n52683), .B(n46222), .X(n26826) );
  nor_x2_sg U31783 ( .A(n46221), .B(n26825), .X(n26824) );
  nand_x8_sg U32026 ( .A(n52704), .B(n14411), .X(n26837) );
  nor_x2_sg U31813 ( .A(n46222), .B(n46443), .X(n26847) );
  nor_x2_sg U31811 ( .A(n14547), .B(n26846), .X(n26845) );
  nor_x2_sg U31830 ( .A(n14552), .B(n26860), .X(n26859) );
  nor_x2_sg U31849 ( .A(n14674), .B(n26874), .X(n26873) );
  nor_x2_sg U31868 ( .A(n14881), .B(n26888), .X(n26887) );
  nor_x2_sg U31879 ( .A(n14815), .B(n26894), .X(n26892) );
  nor_x2_sg U31886 ( .A(n46222), .B(n41569), .X(n26898) );
  nor_x2_sg U31901 ( .A(n26909), .B(n52917), .X(n26906) );
  nand_x8_sg U32176 ( .A(n27026), .B(n27027), .X(n26909) );
  nor_x2_sg U32178 ( .A(n26914), .B(n26911), .X(n26913) );
  nor_x2_sg U32183 ( .A(n46440), .B(n46236), .X(n27063) );
  nor_x2_sg U32189 ( .A(n46220), .B(n46435), .X(n27068) );
  nor_x2_sg U32513 ( .A(n27298), .B(n27299), .X(n27297) );
  nor_x2_sg U32187 ( .A(n14945), .B(n46219), .X(n27067) );
  nor_x2_sg U32199 ( .A(n46220), .B(n46432), .X(n27076) );
  nor_x2_sg U32196 ( .A(n46219), .B(n27074), .X(n27073) );
  nor_x2_sg U32209 ( .A(n52934), .B(n46220), .X(n27083) );
  nor_x2_sg U32206 ( .A(n46219), .B(n27081), .X(n27080) );
  nor_x2_sg U32219 ( .A(n46428), .B(n46220), .X(n27090) );
  nor_x2_sg U32216 ( .A(n46219), .B(n27088), .X(n27087) );
  nor_x2_sg U32229 ( .A(n46427), .B(n46220), .X(n27098) );
  nor_x2_sg U32226 ( .A(n46219), .B(n27095), .X(n27094) );
  nor_x2_sg U32238 ( .A(n52967), .B(n46220), .X(n27105) );
  nor_x2_sg U32236 ( .A(n46219), .B(n27104), .X(n27103) );
  nand_x8_sg U32492 ( .A(n52980), .B(n46423), .X(n27116) );
  nor_x2_sg U32266 ( .A(n46220), .B(n46420), .X(n27126) );
  nor_x2_sg U32264 ( .A(n15328), .B(n27125), .X(n27124) );
  nor_x2_sg U32283 ( .A(n15332), .B(n27139), .X(n27138) );
  nor_x2_sg U32302 ( .A(n15533), .B(n27153), .X(n27152) );
  nor_x2_sg U32499 ( .A(n27158), .B(n53148), .X(n27165) );
  nor_x2_sg U32321 ( .A(n27167), .B(n27168), .X(n27166) );
  nor_x2_sg U32332 ( .A(n15596), .B(n27174), .X(n27172) );
  nor_x2_sg U32339 ( .A(n46220), .B(n41266), .X(n27178) );
  nor_x2_sg U32354 ( .A(n27189), .B(n53195), .X(n27186) );
  nand_x8_sg U32641 ( .A(n27306), .B(n27307), .X(n27189) );
  nor_x2_sg U32643 ( .A(n27196), .B(n27191), .X(n27193) );
  nor_x2_sg U32647 ( .A(n46416), .B(n46236), .X(n27343) );
  nor_x2_sg U32653 ( .A(n46218), .B(n46413), .X(n27348) );
  nor_x2_sg U32966 ( .A(n27577), .B(n27578), .X(n27576) );
  nor_x2_sg U32651 ( .A(n15729), .B(n46217), .X(n27347) );
  nor_x2_sg U32663 ( .A(n46218), .B(n53207), .X(n27356) );
  nor_x2_sg U32660 ( .A(n46217), .B(n27354), .X(n27353) );
  nor_x2_sg U32673 ( .A(n53214), .B(n46218), .X(n27363) );
  nor_x2_sg U32670 ( .A(n46217), .B(n27361), .X(n27360) );
  nor_x2_sg U32683 ( .A(n46405), .B(n46218), .X(n27370) );
  nor_x2_sg U32680 ( .A(n46217), .B(n27368), .X(n27367) );
  nor_x2_sg U32694 ( .A(n53227), .B(n46218), .X(n27378) );
  nand_x8_sg U32941 ( .A(n53225), .B(n46404), .X(n27377) );
  nor_x2_sg U32690 ( .A(n46217), .B(n27375), .X(n27374) );
  nor_x2_sg U32703 ( .A(n53240), .B(n46218), .X(n27385) );
  nor_x2_sg U32701 ( .A(n46217), .B(n27384), .X(n27383) );
  nand_x8_sg U32945 ( .A(n53263), .B(n46400), .X(n27396) );
  nor_x2_sg U32731 ( .A(n46218), .B(n53282), .X(n27406) );
  nor_x2_sg U32729 ( .A(n16109), .B(n27405), .X(n27404) );
  nor_x2_sg U32748 ( .A(n16113), .B(n27419), .X(n27418) );
  nor_x2_sg U32767 ( .A(n16239), .B(n27433), .X(n27432) );
  nor_x2_sg U32782 ( .A(n27436), .B(n27437), .X(n27435) );
  nor_x2_sg U32786 ( .A(n16442), .B(n27447), .X(n27446) );
  nor_x2_sg U32797 ( .A(n16378), .B(n27453), .X(n27451) );
  nor_x2_sg U32804 ( .A(n46218), .B(n41264), .X(n27457) );
  nor_x2_sg U32819 ( .A(n27468), .B(n53475), .X(n27465) );
  nand_x8_sg U33094 ( .A(n27585), .B(n27586), .X(n27468) );
  nor_x2_sg U33096 ( .A(n27473), .B(n27470), .X(n27472) );
  nor_x2_sg U33103 ( .A(n46396), .B(n46236), .X(n27623) );
  nor_x2_sg U33109 ( .A(n46216), .B(n46391), .X(n27628) );
  nor_x2_sg U33423 ( .A(n27856), .B(n27857), .X(n27855) );
  nor_x2_sg U33107 ( .A(n16511), .B(n46215), .X(n27627) );
  nor_x2_sg U33119 ( .A(n46216), .B(n46388), .X(n27636) );
  nor_x2_sg U33116 ( .A(n46215), .B(n27634), .X(n27633) );
  nor_x2_sg U33129 ( .A(n53492), .B(n46216), .X(n27643) );
  nor_x2_sg U33126 ( .A(n46215), .B(n27641), .X(n27640) );
  nor_x2_sg U33139 ( .A(n46384), .B(n46216), .X(n27650) );
  nor_x2_sg U33136 ( .A(n46215), .B(n27648), .X(n27647) );
  nor_x2_sg U33149 ( .A(n46383), .B(n46216), .X(n27658) );
  nor_x2_sg U33146 ( .A(n46215), .B(n27655), .X(n27654) );
  nor_x2_sg U33158 ( .A(n53525), .B(n46216), .X(n27665) );
  nor_x2_sg U33156 ( .A(n46215), .B(n27664), .X(n27663) );
  nand_x8_sg U33402 ( .A(n53538), .B(n46379), .X(n27676) );
  nor_x2_sg U33186 ( .A(n46216), .B(n46376), .X(n27686) );
  nor_x2_sg U33184 ( .A(n16894), .B(n27685), .X(n27684) );
  nor_x2_sg U33203 ( .A(n16898), .B(n27699), .X(n27698) );
  nor_x2_sg U33222 ( .A(n17099), .B(n27713), .X(n27712) );
  nor_x2_sg U33409 ( .A(n27718), .B(n53706), .X(n27725) );
  nor_x2_sg U33241 ( .A(n27727), .B(n27728), .X(n27726) );
  nor_x2_sg U33252 ( .A(n17162), .B(n27734), .X(n27732) );
  nor_x2_sg U33259 ( .A(n46216), .B(n41262), .X(n27738) );
  nor_x2_sg U33274 ( .A(n27749), .B(n53753), .X(n27746) );
  nand_x8_sg U33551 ( .A(n27864), .B(n27865), .X(n27749) );
  nor_x2_sg U33553 ( .A(n27754), .B(n27751), .X(n27753) );
  nor_x2_sg U33562 ( .A(n46373), .B(n46236), .X(n27903) );
  nor_x2_sg U33568 ( .A(n46214), .B(n46368), .X(n27908) );
  nor_x2_sg U33882 ( .A(n28137), .B(n28138), .X(n28136) );
  nor_x2_sg U33566 ( .A(n17294), .B(n46213), .X(n27907) );
  nor_x2_sg U33578 ( .A(n46214), .B(n53765), .X(n27916) );
  nor_x2_sg U33575 ( .A(n46213), .B(n27914), .X(n27913) );
  nor_x2_sg U33588 ( .A(n46363), .B(n46214), .X(n27923) );
  nor_x2_sg U33585 ( .A(n46213), .B(n27921), .X(n27920) );
  nor_x2_sg U33598 ( .A(n46361), .B(n46214), .X(n27930) );
  nor_x2_sg U33595 ( .A(n46213), .B(n27928), .X(n27927) );
  nor_x2_sg U33608 ( .A(n46360), .B(n46214), .X(n27938) );
  nor_x2_sg U33605 ( .A(n46213), .B(n27935), .X(n27934) );
  nor_x2_sg U33617 ( .A(n53802), .B(n46214), .X(n27945) );
  nor_x2_sg U33615 ( .A(n46213), .B(n27944), .X(n27943) );
  nand_x8_sg U33861 ( .A(n53816), .B(n17524), .X(n27956) );
  nor_x2_sg U33645 ( .A(n46214), .B(n46356), .X(n27966) );
  nor_x2_sg U33643 ( .A(n17668), .B(n27965), .X(n27964) );
  nor_x2_sg U33662 ( .A(n17673), .B(n27979), .X(n27978) );
  nor_x2_sg U33681 ( .A(n17795), .B(n27993), .X(n27992) );
  nor_x2_sg U33700 ( .A(n18002), .B(n28007), .X(n28006) );
  nor_x2_sg U33711 ( .A(n17936), .B(n28013), .X(n28011) );
  nor_x2_sg U33718 ( .A(n46214), .B(n41567), .X(n28017) );
  nor_x2_sg U33733 ( .A(n28028), .B(n54037), .X(n28025) );
  nand_x8_sg U34010 ( .A(n28145), .B(n28146), .X(n28028) );
  nor_x2_sg U34012 ( .A(n28033), .B(n28030), .X(n28032) );
  nor_x2_sg U34016 ( .A(n46353), .B(n46236), .X(n28182) );
  nor_x2_sg U34022 ( .A(n46212), .B(n46348), .X(n28187) );
  nor_x2_sg U34348 ( .A(n28416), .B(n28417), .X(n28415) );
  nor_x2_sg U34020 ( .A(n18066), .B(n46211), .X(n28186) );
  nor_x2_sg U34032 ( .A(n46212), .B(n46345), .X(n28195) );
  nor_x2_sg U34029 ( .A(n46211), .B(n28193), .X(n28192) );
  nor_x2_sg U34041 ( .A(n46343), .B(n46212), .X(n28202) );
  nor_x2_sg U34039 ( .A(n46211), .B(n28200), .X(n28199) );
  nor_x2_sg U34050 ( .A(n46339), .B(n46212), .X(n28209) );
  nor_x2_sg U34048 ( .A(n46211), .B(n28207), .X(n28206) );
  nor_x2_sg U34061 ( .A(n54070), .B(n46212), .X(n28217) );
  nand_x8_sg U34323 ( .A(n54066), .B(n46337), .X(n28216) );
  nor_x2_sg U34057 ( .A(n46211), .B(n28214), .X(n28213) );
  nor_x2_sg U34070 ( .A(n54084), .B(n46212), .X(n28224) );
  nor_x2_sg U34068 ( .A(n46211), .B(n28223), .X(n28222) );
  nand_x8_sg U34327 ( .A(n54098), .B(n46331), .X(n28235) );
  nor_x2_sg U34098 ( .A(n46212), .B(n54124), .X(n28245) );
  nor_x2_sg U34096 ( .A(n18437), .B(n28244), .X(n28243) );
  nor_x2_sg U34115 ( .A(n18442), .B(n28259), .X(n28258) );
  nor_x2_sg U34134 ( .A(n18654), .B(n28273), .X(n28272) );
  nor_x2_sg U34153 ( .A(n18771), .B(n28287), .X(n28286) );
  nor_x2_sg U34164 ( .A(n18705), .B(n28293), .X(n28291) );
  nor_x2_sg U34171 ( .A(n46212), .B(n41565), .X(n28297) );
  nor_x2_sg U34186 ( .A(n28308), .B(n54318), .X(n28305) );
  nand_x8_sg U34475 ( .A(n28424), .B(n28425), .X(n28308) );
  nor_x2_sg U34477 ( .A(n28314), .B(n28310), .X(n28312) );
  nor_x2_sg U34481 ( .A(n46326), .B(n46236), .X(n28461) );
  nand_x8_sg U35577 ( .A(n21153), .B(n26358), .X(n28459) );
  nor_x2_sg U34487 ( .A(n46210), .B(n46321), .X(n28466) );
  nor_x2_sg U34802 ( .A(n28695), .B(n28696), .X(n28694) );
  nor_x2_sg U34485 ( .A(n18839), .B(n46209), .X(n28465) );
  nor_x2_sg U34497 ( .A(n46210), .B(n54330), .X(n28474) );
  nor_x2_sg U34494 ( .A(n46209), .B(n28472), .X(n28471) );
  nor_x2_sg U34507 ( .A(n46316), .B(n46210), .X(n28481) );
  nor_x2_sg U34504 ( .A(n46209), .B(n28479), .X(n28478) );
  nor_x2_sg U34517 ( .A(n46314), .B(n46210), .X(n28488) );
  nor_x2_sg U34514 ( .A(n46209), .B(n28486), .X(n28485) );
  nor_x2_sg U34527 ( .A(n46313), .B(n46210), .X(n28496) );
  nor_x2_sg U34524 ( .A(n46209), .B(n28493), .X(n28492) );
  nor_x2_sg U34536 ( .A(n54367), .B(n46210), .X(n28503) );
  nor_x2_sg U34534 ( .A(n46209), .B(n28502), .X(n28501) );
  nand_x8_sg U34781 ( .A(n54381), .B(n19069), .X(n28514) );
  nor_x2_sg U34564 ( .A(n46210), .B(n46309), .X(n28524) );
  nor_x2_sg U34562 ( .A(n19213), .B(n28523), .X(n28522) );
  nor_x2_sg U34581 ( .A(n19218), .B(n28537), .X(n28536) );
  nor_x2_sg U34600 ( .A(n19340), .B(n28551), .X(n28550) );
  nor_x2_sg U34619 ( .A(n19547), .B(n28565), .X(n28564) );
  nor_x2_sg U34630 ( .A(n19481), .B(n28571), .X(n28569) );
  nor_x2_sg U34637 ( .A(n46210), .B(n41563), .X(n28575) );
  nor_x2_sg U34652 ( .A(n28586), .B(n54602), .X(n28583) );
  nand_x8_sg U34930 ( .A(n28703), .B(n28704), .X(n28586) );
  nor_x2_sg U34932 ( .A(n28591), .B(n28588), .X(n28590) );
  nor_x2_sg U34936 ( .A(n46306), .B(n46236), .X(n28740) );
  nor_x2_sg U34942 ( .A(n46208), .B(n46301), .X(n28745) );
  nor_x2_sg U35255 ( .A(n28973), .B(n28974), .X(n28972) );
  nor_x2_sg U34940 ( .A(n19611), .B(n46207), .X(n28744) );
  nor_x2_sg U34952 ( .A(n46208), .B(n54614), .X(n28753) );
  nor_x2_sg U34949 ( .A(n46207), .B(n28751), .X(n28750) );
  nor_x2_sg U34962 ( .A(n46296), .B(n46208), .X(n28760) );
  nor_x2_sg U34959 ( .A(n46207), .B(n28758), .X(n28757) );
  nor_x2_sg U34972 ( .A(n46294), .B(n46208), .X(n28767) );
  nor_x2_sg U34969 ( .A(n46207), .B(n28765), .X(n28764) );
  nor_x2_sg U34983 ( .A(n54634), .B(n46208), .X(n28775) );
  nand_x8_sg U35230 ( .A(n54632), .B(n46293), .X(n28774) );
  nor_x2_sg U34979 ( .A(n46207), .B(n28772), .X(n28771) );
  nor_x2_sg U34992 ( .A(n54647), .B(n46208), .X(n28782) );
  nor_x2_sg U34990 ( .A(n46207), .B(n28781), .X(n28780) );
  nand_x8_sg U35234 ( .A(n54670), .B(n46287), .X(n28793) );
  nor_x2_sg U35020 ( .A(n46208), .B(n54688), .X(n28803) );
  nor_x2_sg U35018 ( .A(n19982), .B(n28802), .X(n28801) );
  nor_x2_sg U35037 ( .A(n19987), .B(n28817), .X(n28816) );
  nor_x2_sg U35056 ( .A(n20108), .B(n28831), .X(n28830) );
  nor_x2_sg U35075 ( .A(n20317), .B(n28845), .X(n28844) );
  nor_x2_sg U35086 ( .A(n20251), .B(n28851), .X(n28849) );
  nor_x2_sg U35093 ( .A(n46208), .B(n41561), .X(n28855) );
  nor_x2_sg U35108 ( .A(n28866), .B(n54886), .X(n28863) );
  nand_x8_sg U35383 ( .A(n28981), .B(n28982), .X(n28866) );
  nor_x2_sg U35385 ( .A(n28871), .B(n28868), .X(n28870) );
  nor_x2_sg U35395 ( .A(n46281), .B(n46236), .X(n29020) );
  nor_x2_sg U35401 ( .A(n46206), .B(n46276), .X(n29025) );
  nor_x2_sg U35720 ( .A(n29256), .B(n29257), .X(n29255) );
  nor_x2_sg U35399 ( .A(n20383), .B(n46205), .X(n29024) );
  nor_x2_sg U35411 ( .A(n46206), .B(n54898), .X(n29033) );
  nor_x2_sg U35408 ( .A(n46205), .B(n29031), .X(n29030) );
  nor_x2_sg U35421 ( .A(n46271), .B(n46206), .X(n29040) );
  nor_x2_sg U35418 ( .A(n46205), .B(n29038), .X(n29037) );
  nor_x2_sg U35431 ( .A(n46269), .B(n46206), .X(n29047) );
  nor_x2_sg U35428 ( .A(n46205), .B(n29045), .X(n29044) );
  nor_x2_sg U35441 ( .A(n46268), .B(n46206), .X(n29055) );
  nor_x2_sg U35438 ( .A(n46205), .B(n29052), .X(n29051) );
  nor_x2_sg U35450 ( .A(n54935), .B(n46206), .X(n29062) );
  nor_x2_sg U35448 ( .A(n46205), .B(n29061), .X(n29060) );
  nand_x8_sg U35699 ( .A(n54949), .B(n20613), .X(n29073) );
  nor_x2_sg U35478 ( .A(n46206), .B(n46264), .X(n29083) );
  nor_x2_sg U35476 ( .A(n20757), .B(n29082), .X(n29081) );
  nor_x2_sg U35495 ( .A(n20762), .B(n29096), .X(n29095) );
  nor_x2_sg U35514 ( .A(n20884), .B(n29110), .X(n29109) );
  nor_x2_sg U35533 ( .A(n21091), .B(n29124), .X(n29123) );
  nor_x2_sg U35544 ( .A(n21025), .B(n29130), .X(n29128) );
  nor_x2_sg U35551 ( .A(n46206), .B(n41559), .X(n29134) );
  nor_x2_sg U35566 ( .A(n29145), .B(n55170), .X(n29142) );
  nand_x8_sg U35848 ( .A(n29264), .B(n29265), .X(n29145) );
  nor_x2_sg U35850 ( .A(n29152), .B(n29147), .X(n29150) );
  nor_x2_sg U35854 ( .A(n46261), .B(n46236), .X(n29301) );
  nor_x2_sg U35860 ( .A(n46204), .B(n46256), .X(n29306) );
  nor_x2_sg U36183 ( .A(n29534), .B(n29535), .X(n29533) );
  nor_x2_sg U35858 ( .A(n21156), .B(n46203), .X(n29305) );
  nor_x2_sg U35870 ( .A(n46204), .B(n55182), .X(n29314) );
  nor_x2_sg U35867 ( .A(n46203), .B(n29312), .X(n29311) );
  nor_x2_sg U35880 ( .A(n46251), .B(n46204), .X(n29321) );
  nor_x2_sg U35877 ( .A(n46203), .B(n29319), .X(n29318) );
  nor_x2_sg U35890 ( .A(n46249), .B(n46204), .X(n29328) );
  nor_x2_sg U35887 ( .A(n46203), .B(n29326), .X(n29325) );
  nor_x2_sg U35901 ( .A(n55202), .B(n46204), .X(n29336) );
  nand_x8_sg U36158 ( .A(n55200), .B(n46248), .X(n29335) );
  nor_x2_sg U35897 ( .A(n46203), .B(n29333), .X(n29332) );
  nor_x2_sg U35910 ( .A(n55215), .B(n46204), .X(n29343) );
  nor_x2_sg U35908 ( .A(n46203), .B(n29342), .X(n29341) );
  nand_x8_sg U36162 ( .A(n55238), .B(n46242), .X(n29354) );
  nor_x2_sg U35938 ( .A(n46204), .B(n55256), .X(n29364) );
  nor_x2_sg U35936 ( .A(n21527), .B(n29363), .X(n29362) );
  nor_x2_sg U35955 ( .A(n21532), .B(n29378), .X(n29377) );
  nor_x2_sg U35974 ( .A(n21653), .B(n29392), .X(n29391) );
  nor_x2_sg U35993 ( .A(n21862), .B(n29406), .X(n29405) );
  nor_x2_sg U36004 ( .A(n21796), .B(n29412), .X(n29410) );
  nor_x2_sg U36011 ( .A(n46204), .B(n41557), .X(n29416) );
  nor_x2_sg U36026 ( .A(n29427), .B(n55454), .X(n29424) );
  nand_x8_sg U36311 ( .A(n29542), .B(n29543), .X(n29427) );
  nor_x2_sg U36321 ( .A(n29432), .B(n29429), .X(n29431) );
  nand_x2_sg U38217 ( .A(n41699), .B(n12425), .X(n11910) );
  nand_x2_sg U38218 ( .A(n41695), .B(n13206), .X(n12688) );
  nand_x2_sg U38219 ( .A(n41691), .B(n13986), .X(n13472) );
  nand_x2_sg U38220 ( .A(n41687), .B(n15539), .X(n15021) );
  nand_x2_sg U38221 ( .A(n41683), .B(n17105), .X(n16587) );
  inv_x4_sg U38222 ( .A(n46637), .X(n46630) );
  inv_x4_sg U38223 ( .A(n46637), .X(n46636) );
  inv_x8_sg U38224 ( .A(n46630), .X(n40519) );
  inv_x8_sg U38225 ( .A(n40519), .X(n40520) );
  inv_x8_sg U38226 ( .A(n40519), .X(n40521) );
  inv_x8_sg U38227 ( .A(n46636), .X(n40522) );
  inv_x8_sg U38228 ( .A(n40522), .X(n40523) );
  inv_x8_sg U38229 ( .A(n40522), .X(n40524) );
  inv_x4_sg U38230 ( .A(n40581), .X(n15857) );
  inv_x4_sg U38231 ( .A(n40564), .X(n24428) );
  inv_x4_sg U38232 ( .A(n40576), .X(n32094) );
  nor_x1_sg U38233 ( .A(n43143), .B(n43771), .X(n15835) );
  inv_x2_sg U38234 ( .A(n15835), .X(n41173) );
  nor_x1_sg U38235 ( .A(n43157), .B(n43755), .X(n11940) );
  inv_x2_sg U38236 ( .A(n11940), .X(n41175) );
  nor_x1_sg U38237 ( .A(n43149), .B(n41594), .X(n19717) );
  inv_x2_sg U38238 ( .A(n19717), .X(n54629) );
  nor_x1_sg U38239 ( .A(n44403), .B(n43973), .X(n18172) );
  inv_x2_sg U38240 ( .A(n18172), .X(n54061) );
  nor_x1_sg U38241 ( .A(n43153), .B(n43800), .X(n13502) );
  inv_x2_sg U38242 ( .A(n13502), .X(n41174) );
  inv_x1_sg U38243 ( .A(n18807), .X(n43566) );
  nor_x1_sg U38244 ( .A(n54226), .B(n54245), .X(n18807) );
  nand_x4_sg U38245 ( .A(n40893), .B(n43566), .X(n40525) );
  inv_x8_sg U38246 ( .A(n40525), .X(n18770) );
  nand_x4_sg U38247 ( .A(n42301), .B(n42300), .X(n40526) );
  nand_x4_sg U38248 ( .A(n42298), .B(n42297), .X(n40527) );
  nand_x4_sg U38249 ( .A(n42295), .B(n42294), .X(n40528) );
  nand_x4_sg U38250 ( .A(n42292), .B(n42291), .X(n40529) );
  nand_x4_sg U38251 ( .A(n42289), .B(n42288), .X(n40530) );
  nor_x1_sg U38252 ( .A(n9791), .B(n23643), .X(n23733) );
  nand_x1_sg U38253 ( .A(n8652), .B(n23735), .X(n23734) );
  nor_x1_sg U38254 ( .A(n9935), .B(n23625), .X(n23742) );
  nand_x1_sg U38255 ( .A(n8655), .B(n23744), .X(n23743) );
  nor_x1_sg U38256 ( .A(n10081), .B(n50260), .X(n23751) );
  nand_x1_sg U38257 ( .A(n8658), .B(n23753), .X(n23752) );
  nand_x4_sg U38258 ( .A(n42136), .B(n11801), .X(n40531) );
  nand_x4_sg U38259 ( .A(n42134), .B(n12576), .X(n40532) );
  nand_x4_sg U38260 ( .A(n42132), .B(n13358), .X(n40533) );
  nand_x4_sg U38261 ( .A(n42130), .B(n14138), .X(n40534) );
  nand_x4_sg U38262 ( .A(n42128), .B(n15691), .X(n40535) );
  nand_x4_sg U38263 ( .A(n42126), .B(n17257), .X(n40536) );
  nand_x4_sg U38264 ( .A(n42124), .B(n18804), .X(n40537) );
  nor_x1_sg U38265 ( .A(n24899), .B(n31309), .X(n31399) );
  nand_x1_sg U38266 ( .A(n8352), .B(n31401), .X(n31400) );
  nor_x1_sg U38267 ( .A(n25043), .B(n31291), .X(n31408) );
  nand_x1_sg U38268 ( .A(n8355), .B(n31410), .X(n31409) );
  nor_x1_sg U38269 ( .A(n25189), .B(n49401), .X(n31417) );
  nand_x1_sg U38270 ( .A(n8358), .B(n31419), .X(n31418) );
  nand_x4_sg U38271 ( .A(n43565), .B(n23734), .X(n40538) );
  inv_x8_sg U38272 ( .A(n40538), .X(n23649) );
  inv_x2_sg U38273 ( .A(n23733), .X(n43565) );
  nand_x4_sg U38274 ( .A(n43564), .B(n23743), .X(n40539) );
  inv_x8_sg U38275 ( .A(n40539), .X(n23631) );
  inv_x2_sg U38276 ( .A(n23742), .X(n43564) );
  nand_x4_sg U38277 ( .A(n43563), .B(n23752), .X(n40540) );
  inv_x8_sg U38278 ( .A(n40540), .X(n23613) );
  inv_x2_sg U38279 ( .A(n23751), .X(n43563) );
  nor_x1_sg U38280 ( .A(n24458), .B(out_L2[4]), .X(n24457) );
  inv_x1_sg U38281 ( .A(n24456), .X(n41554) );
  nor_x1_sg U38282 ( .A(n40737), .B(n24423), .X(n24456) );
  nor_x1_sg U38283 ( .A(n40723), .B(n50179), .X(n24462) );
  inv_x1_sg U38284 ( .A(n24463), .X(n41863) );
  nor_x1_sg U38285 ( .A(n24464), .B(out_L2[2]), .X(n24463) );
  nand_x4_sg U38286 ( .A(n43101), .B(n10741), .X(n40541) );
  nand_x4_sg U38287 ( .A(n10776), .B(n43343), .X(n40542) );
  nand_x4_sg U38288 ( .A(n42112), .B(n11610), .X(n40543) );
  nand_x4_sg U38289 ( .A(n42110), .B(n12391), .X(n40544) );
  nand_x4_sg U38290 ( .A(n11910), .B(n43287), .X(n40545) );
  nand_x4_sg U38291 ( .A(n42108), .B(n13171), .X(n40546) );
  nand_x4_sg U38292 ( .A(n12688), .B(n43285), .X(n40547) );
  nand_x4_sg U38293 ( .A(n42106), .B(n13951), .X(n40548) );
  nand_x4_sg U38294 ( .A(n13472), .B(n43283), .X(n40549) );
  nand_x4_sg U38295 ( .A(n42076), .B(n13991), .X(n40550) );
  nand_x4_sg U38296 ( .A(n42122), .B(n14722), .X(n40551) );
  nand_x4_sg U38297 ( .A(n42104), .B(n15504), .X(n40552) );
  nand_x4_sg U38298 ( .A(n15021), .B(n43281), .X(n40553) );
  nand_x4_sg U38299 ( .A(n42072), .B(n16286), .X(n40554) );
  nand_x4_sg U38300 ( .A(n42102), .B(n17070), .X(n40555) );
  nand_x4_sg U38301 ( .A(n16587), .B(n43279), .X(n40556) );
  nand_x4_sg U38302 ( .A(n42118), .B(n17843), .X(n40557) );
  nand_x4_sg U38303 ( .A(n42100), .B(n18651), .X(n40558) );
  nand_x4_sg U38304 ( .A(n42116), .B(n19388), .X(n40559) );
  nand_x4_sg U38305 ( .A(n42114), .B(n20932), .X(n40560) );
  nand_x4_sg U38306 ( .A(n43562), .B(n31400), .X(n40561) );
  inv_x8_sg U38307 ( .A(n40561), .X(n31315) );
  inv_x2_sg U38308 ( .A(n31399), .X(n43562) );
  nand_x4_sg U38309 ( .A(n43561), .B(n31409), .X(n40562) );
  inv_x8_sg U38310 ( .A(n40562), .X(n31297) );
  inv_x2_sg U38311 ( .A(n31408), .X(n43561) );
  nand_x4_sg U38312 ( .A(n43560), .B(n31418), .X(n40563) );
  inv_x8_sg U38313 ( .A(n40563), .X(n31279) );
  inv_x2_sg U38314 ( .A(n31417), .X(n43560) );
  nor_x1_sg U38315 ( .A(n32124), .B(out_L1[4]), .X(n32123) );
  inv_x1_sg U38316 ( .A(n32122), .X(n41556) );
  nor_x1_sg U38317 ( .A(n40738), .B(n32089), .X(n32122) );
  nor_x1_sg U38318 ( .A(n40724), .B(n49320), .X(n32128) );
  inv_x1_sg U38319 ( .A(n32129), .X(n41861) );
  nor_x1_sg U38320 ( .A(n32130), .B(out_L1[2]), .X(n32129) );
  nor_x1_sg U38321 ( .A(n52404), .B(n26763), .X(n26762) );
  nand_x1_sg U38322 ( .A(n26694), .B(n51049), .X(n26764) );
  nand_x4_sg U38323 ( .A(n41554), .B(n41553), .X(n40564) );
  inv_x2_sg U38324 ( .A(n24457), .X(n41553) );
  inv_x1_sg U38325 ( .A(n24460), .X(n42522) );
  nor_x1_sg U38326 ( .A(n50180), .B(out_L2[3]), .X(n24460) );
  nand_x4_sg U38327 ( .A(n41864), .B(n41863), .X(n40565) );
  inv_x8_sg U38328 ( .A(n40565), .X(n24417) );
  inv_x2_sg U38329 ( .A(n24462), .X(n41864) );
  nand_x4_sg U38330 ( .A(n10825), .B(n42383), .X(n40566) );
  nand_x4_sg U38331 ( .A(n11605), .B(n42385), .X(n40567) );
  nand_x4_sg U38332 ( .A(n14717), .B(n42393), .X(n40568) );
  inv_x1_sg U38333 ( .A(n15871), .X(n41869) );
  nor_x1_sg U38334 ( .A(n15872), .B(n46409), .X(n15871) );
  nand_x4_sg U38335 ( .A(n16281), .B(n42381), .X(n40569) );
  nand_x4_sg U38336 ( .A(n17838), .B(n42391), .X(n40570) );
  nand_x4_sg U38337 ( .A(n18605), .B(n43301), .X(n40571) );
  nand_x4_sg U38338 ( .A(n19383), .B(n42389), .X(n40572) );
  nand_x4_sg U38339 ( .A(n20151), .B(n43299), .X(n40573) );
  nand_x4_sg U38340 ( .A(n20927), .B(n42387), .X(n40574) );
  nand_x4_sg U38341 ( .A(n21696), .B(n43297), .X(n40575) );
  nand_x4_sg U38342 ( .A(n41556), .B(n41555), .X(n40576) );
  inv_x2_sg U38343 ( .A(n32123), .X(n41555) );
  inv_x1_sg U38344 ( .A(n32126), .X(n42523) );
  nor_x1_sg U38345 ( .A(n49321), .B(out_L1[3]), .X(n32126) );
  nand_x4_sg U38346 ( .A(n41862), .B(n41861), .X(n40577) );
  inv_x8_sg U38347 ( .A(n40577), .X(n32083) );
  inv_x2_sg U38348 ( .A(n32128), .X(n41862) );
  nor_x1_sg U38349 ( .A(n51291), .B(n25647), .X(n25646) );
  nand_x1_sg U38350 ( .A(n25576), .B(n50972), .X(n25648) );
  nor_x1_sg U38351 ( .A(n51852), .B(n26206), .X(n26205) );
  nand_x1_sg U38352 ( .A(n26137), .B(n51010), .X(n26207) );
  nand_x4_sg U38353 ( .A(n26764), .B(n43555), .X(n40578) );
  inv_x8_sg U38354 ( .A(n40578), .X(n26687) );
  inv_x2_sg U38355 ( .A(n26762), .X(n43555) );
  nor_x1_sg U38356 ( .A(n53238), .B(n27601), .X(n27600) );
  nand_x1_sg U38357 ( .A(n27532), .B(n51106), .X(n27602) );
  nor_x1_sg U38358 ( .A(n54645), .B(n28997), .X(n28996) );
  nand_x1_sg U38359 ( .A(n28928), .B(n51200), .X(n28998) );
  nor_x1_sg U38360 ( .A(n55213), .B(n29558), .X(n29557) );
  nand_x1_sg U38361 ( .A(n29489), .B(n51238), .X(n29559) );
  inv_x1_sg U38362 ( .A(n22801), .X(n43732) );
  nor_x1_sg U38363 ( .A(n44647), .B(n50910), .X(n22801) );
  inv_x1_sg U38364 ( .A(n22173), .X(n43675) );
  nor_x1_sg U38365 ( .A(n44653), .B(n50943), .X(n22173) );
  inv_x1_sg U38366 ( .A(n22777), .X(n43676) );
  nor_x1_sg U38367 ( .A(n44633), .B(n50933), .X(n22777) );
  nor_x1_sg U38368 ( .A(n42226), .B(n22818), .X(n23056) );
  nand_x1_sg U38369 ( .A(n22818), .B(n42226), .X(n23057) );
  nor_x1_sg U38370 ( .A(n41954), .B(n50890), .X(n23032) );
  inv_x1_sg U38371 ( .A(n23033), .X(n43674) );
  nor_x1_sg U38372 ( .A(n9443), .B(n41953), .X(n23033) );
  nor_x1_sg U38373 ( .A(n9440), .B(n23036), .X(n23035) );
  nand_x1_sg U38374 ( .A(n23036), .B(n9440), .X(n23037) );
  nor_x1_sg U38375 ( .A(n42224), .B(n23073), .X(n23282) );
  nand_x1_sg U38376 ( .A(n23073), .B(n42224), .X(n23283) );
  nor_x1_sg U38377 ( .A(n44619), .B(n41328), .X(n22159) );
  inv_x1_sg U38378 ( .A(n22160), .X(n43667) );
  nor_x1_sg U38379 ( .A(n50849), .B(n50810), .X(n22160) );
  nor_x1_sg U38380 ( .A(n41952), .B(n50845), .X(n23026) );
  inv_x1_sg U38381 ( .A(n23027), .X(n43670) );
  nor_x1_sg U38382 ( .A(n9492), .B(n41951), .X(n23027) );
  nor_x1_sg U38383 ( .A(n9489), .B(n23262), .X(n23261) );
  nand_x1_sg U38384 ( .A(n23262), .B(n9489), .X(n23263) );
  nor_x1_sg U38385 ( .A(n42220), .B(n23299), .X(n23487) );
  nand_x1_sg U38386 ( .A(n23299), .B(n42220), .X(n23488) );
  nor_x1_sg U38387 ( .A(n44617), .B(n41327), .X(n22152) );
  inv_x1_sg U38388 ( .A(n22153), .X(n43663) );
  nor_x1_sg U38389 ( .A(n50804), .B(n50762), .X(n22153) );
  nor_x1_sg U38390 ( .A(n41950), .B(n50800), .X(n23020) );
  inv_x1_sg U38391 ( .A(n23021), .X(n43666) );
  nor_x1_sg U38392 ( .A(n9541), .B(n41949), .X(n23021) );
  nor_x1_sg U38393 ( .A(n9538), .B(n23256), .X(n23255) );
  nand_x1_sg U38394 ( .A(n23256), .B(n9538), .X(n23257) );
  nor_x1_sg U38395 ( .A(n42218), .B(n23504), .X(n23677) );
  nand_x1_sg U38396 ( .A(n23504), .B(n42218), .X(n23678) );
  nor_x1_sg U38397 ( .A(n44613), .B(n41325), .X(n22145) );
  inv_x1_sg U38398 ( .A(n22146), .X(n43659) );
  nor_x1_sg U38399 ( .A(n50756), .B(n50715), .X(n22146) );
  nor_x1_sg U38400 ( .A(n44615), .B(n41326), .X(n23013) );
  inv_x1_sg U38401 ( .A(n23014), .X(n43661) );
  nor_x1_sg U38402 ( .A(n50752), .B(n50724), .X(n23014) );
  nor_x1_sg U38403 ( .A(n42214), .B(n23694), .X(n23848) );
  nand_x1_sg U38404 ( .A(n23694), .B(n42214), .X(n23849) );
  nor_x1_sg U38405 ( .A(n44609), .B(n41323), .X(n22138) );
  inv_x1_sg U38406 ( .A(n22139), .X(n43655) );
  nor_x1_sg U38407 ( .A(n50709), .B(n50667), .X(n22139) );
  nor_x1_sg U38408 ( .A(n44611), .B(n41324), .X(n23006) );
  inv_x1_sg U38409 ( .A(n23007), .X(n43657) );
  nor_x1_sg U38410 ( .A(n50705), .B(n50676), .X(n23007) );
  nor_x1_sg U38411 ( .A(n42212), .B(n23865), .X(n24001) );
  nand_x1_sg U38412 ( .A(n23865), .B(n42212), .X(n24002) );
  nor_x1_sg U38413 ( .A(n42196), .B(n9668), .X(n23451) );
  nand_x1_sg U38414 ( .A(n9668), .B(n42196), .X(n23452) );
  nor_x1_sg U38415 ( .A(n44607), .B(n41322), .X(n22131) );
  inv_x1_sg U38416 ( .A(n22132), .X(n42556) );
  nor_x1_sg U38417 ( .A(n50661), .B(n50620), .X(n22132) );
  nor_x1_sg U38418 ( .A(n42230), .B(n9688), .X(n22468) );
  nand_x1_sg U38419 ( .A(n9688), .B(n42230), .X(n22469) );
  nor_x1_sg U38420 ( .A(n44645), .B(n41578), .X(n22999) );
  inv_x1_sg U38421 ( .A(n23000), .X(n42558) );
  nor_x1_sg U38422 ( .A(n50658), .B(n50629), .X(n23000) );
  nor_x1_sg U38423 ( .A(n42208), .B(n24018), .X(n24145) );
  nand_x1_sg U38424 ( .A(n24018), .B(n42208), .X(n24146) );
  nor_x1_sg U38425 ( .A(n44603), .B(n41320), .X(n22124) );
  inv_x1_sg U38426 ( .A(n22125), .X(n43651) );
  nor_x1_sg U38427 ( .A(n50614), .B(n50571), .X(n22125) );
  nor_x1_sg U38428 ( .A(n44605), .B(n41321), .X(n22992) );
  inv_x1_sg U38429 ( .A(n22993), .X(n43653) );
  nor_x1_sg U38430 ( .A(n50610), .B(n50580), .X(n22993) );
  nor_x1_sg U38431 ( .A(n42206), .B(n24162), .X(n24261) );
  nand_x1_sg U38432 ( .A(n24162), .B(n42206), .X(n24262) );
  nor_x1_sg U38433 ( .A(n44599), .B(n41318), .X(n22117) );
  inv_x1_sg U38434 ( .A(n22118), .X(n43647) );
  nor_x1_sg U38435 ( .A(n50565), .B(n50524), .X(n22118) );
  nor_x1_sg U38436 ( .A(n44601), .B(n41319), .X(n22985) );
  inv_x1_sg U38437 ( .A(n22986), .X(n43649) );
  nor_x1_sg U38438 ( .A(n50561), .B(n50533), .X(n22986) );
  nor_x1_sg U38439 ( .A(n44527), .B(n41164), .X(n24125) );
  inv_x1_sg U38440 ( .A(n24126), .X(n42534) );
  nor_x1_sg U38441 ( .A(n50508), .B(n50498), .X(n24126) );
  nor_x1_sg U38442 ( .A(n42202), .B(n24278), .X(n24363) );
  nand_x1_sg U38443 ( .A(n24278), .B(n42202), .X(n24364) );
  nor_x1_sg U38444 ( .A(n44595), .B(n41316), .X(n22110) );
  inv_x1_sg U38445 ( .A(n22111), .X(n43643) );
  nor_x1_sg U38446 ( .A(n50518), .B(n50477), .X(n22111) );
  nor_x1_sg U38447 ( .A(n44597), .B(n41317), .X(n22978) );
  inv_x1_sg U38448 ( .A(n22979), .X(n43645) );
  nor_x1_sg U38449 ( .A(n50514), .B(n50486), .X(n22979) );
  nor_x1_sg U38450 ( .A(n44525), .B(n41163), .X(n24118) );
  inv_x1_sg U38451 ( .A(n24119), .X(n42532) );
  nor_x1_sg U38452 ( .A(n50461), .B(n50452), .X(n24119) );
  nor_x1_sg U38453 ( .A(n42198), .B(n24358), .X(n24356) );
  nand_x1_sg U38454 ( .A(n24358), .B(n42198), .X(n24357) );
  nor_x1_sg U38455 ( .A(n44591), .B(n41314), .X(n22103) );
  inv_x1_sg U38456 ( .A(n22104), .X(n43639) );
  nor_x1_sg U38457 ( .A(n50471), .B(n50431), .X(n22104) );
  nor_x1_sg U38458 ( .A(n44593), .B(n41315), .X(n22971) );
  inv_x1_sg U38459 ( .A(n22972), .X(n43641) );
  nor_x1_sg U38460 ( .A(n50467), .B(n50440), .X(n22972) );
  nor_x1_sg U38461 ( .A(n44523), .B(n41576), .X(n24111) );
  inv_x1_sg U38462 ( .A(n24112), .X(n42530) );
  nor_x1_sg U38463 ( .A(n50415), .B(n50406), .X(n24112) );
  inv_x1_sg U38464 ( .A(n24350), .X(n43682) );
  nor_x1_sg U38465 ( .A(n50413), .B(n50411), .X(n24350) );
  nor_x1_sg U38466 ( .A(n44587), .B(n41312), .X(n22096) );
  inv_x1_sg U38467 ( .A(n22097), .X(n43635) );
  nor_x1_sg U38468 ( .A(n50425), .B(n50384), .X(n22097) );
  nor_x1_sg U38469 ( .A(n44589), .B(n41313), .X(n22964) );
  inv_x1_sg U38470 ( .A(n22965), .X(n43637) );
  nor_x1_sg U38471 ( .A(n50421), .B(n50393), .X(n22965) );
  nor_x1_sg U38472 ( .A(n44629), .B(n41282), .X(n24104) );
  inv_x1_sg U38473 ( .A(n24105), .X(n42528) );
  nor_x1_sg U38474 ( .A(n50368), .B(n50358), .X(n24105) );
  inv_x1_sg U38475 ( .A(n24343), .X(n43681) );
  nor_x1_sg U38476 ( .A(n41610), .B(n50366), .X(n24343) );
  nor_x1_sg U38477 ( .A(n44585), .B(n41311), .X(n22089) );
  inv_x1_sg U38478 ( .A(n22090), .X(n43633) );
  nor_x1_sg U38479 ( .A(n50378), .B(n50337), .X(n22090) );
  nor_x1_sg U38480 ( .A(n50365), .B(n50363), .X(n24432) );
  inv_x1_sg U38481 ( .A(n24433), .X(n42519) );
  nor_x1_sg U38482 ( .A(n24434), .B(n24435), .X(n24433) );
  nor_x1_sg U38483 ( .A(n44643), .B(n41336), .X(n22957) );
  inv_x1_sg U38484 ( .A(n22958), .X(n43700) );
  nor_x1_sg U38485 ( .A(n50374), .B(n50346), .X(n22958) );
  nor_x1_sg U38486 ( .A(n44521), .B(n41575), .X(n24097) );
  inv_x1_sg U38487 ( .A(n24098), .X(n42526) );
  nor_x1_sg U38488 ( .A(n50321), .B(n50312), .X(n24098) );
  nor_x1_sg U38489 ( .A(n45495), .B(n41169), .X(n24336) );
  inv_x1_sg U38490 ( .A(n24337), .X(n43679) );
  nor_x1_sg U38491 ( .A(n50319), .B(n50317), .X(n24337) );
  nor_x1_sg U38492 ( .A(n44581), .B(n41309), .X(n22082) );
  inv_x1_sg U38493 ( .A(n22083), .X(n43629) );
  nor_x1_sg U38494 ( .A(n50331), .B(n50291), .X(n22083) );
  nor_x1_sg U38495 ( .A(n44583), .B(n41310), .X(n22950) );
  inv_x1_sg U38496 ( .A(n22951), .X(n43631) );
  nor_x1_sg U38497 ( .A(n50327), .B(n50300), .X(n22951) );
  nor_x1_sg U38498 ( .A(n44627), .B(n41332), .X(n24090) );
  inv_x1_sg U38499 ( .A(n24091), .X(n42588) );
  nor_x1_sg U38500 ( .A(n50275), .B(n50267), .X(n24091) );
  nand_x1_sg U38501 ( .A(n41141), .B(n10078), .X(n40579) );
  nor_x1_sg U38502 ( .A(n44579), .B(n41308), .X(n22075) );
  inv_x1_sg U38503 ( .A(n22076), .X(n43627) );
  nor_x1_sg U38504 ( .A(n50285), .B(n50245), .X(n22076) );
  nand_x4_sg U38505 ( .A(n40906), .B(n42522), .X(n40580) );
  inv_x8_sg U38506 ( .A(n40580), .X(n24423) );
  nor_x1_sg U38507 ( .A(n44641), .B(n41335), .X(n22943) );
  inv_x1_sg U38508 ( .A(n22944), .X(n43698) );
  nor_x1_sg U38509 ( .A(n50281), .B(n50254), .X(n22944) );
  nor_x1_sg U38510 ( .A(n44625), .B(n41168), .X(n24083) );
  inv_x1_sg U38511 ( .A(n24084), .X(n42586) );
  nor_x1_sg U38512 ( .A(n50229), .B(n50222), .X(n24084) );
  nor_x1_sg U38513 ( .A(n41616), .B(n41960), .X(n24324) );
  inv_x1_sg U38514 ( .A(n24325), .X(n43721) );
  nor_x1_sg U38515 ( .A(n10127), .B(n41615), .X(n24325) );
  nor_x1_sg U38516 ( .A(n44577), .B(n41307), .X(n22068) );
  inv_x1_sg U38517 ( .A(n22069), .X(n43625) );
  nor_x1_sg U38518 ( .A(n50239), .B(n50201), .X(n22069) );
  nor_x1_sg U38519 ( .A(n41243), .B(n24417), .X(n24414) );
  nand_x1_sg U38520 ( .A(n41243), .B(n24417), .X(n24415) );
  nor_x1_sg U38521 ( .A(n44651), .B(n41338), .X(n22936) );
  inv_x1_sg U38522 ( .A(n22937), .X(n43722) );
  nor_x1_sg U38523 ( .A(n50235), .B(n50210), .X(n22937) );
  nor_x1_sg U38524 ( .A(n44519), .B(n41281), .X(n24076) );
  inv_x1_sg U38525 ( .A(n24077), .X(n42524) );
  nor_x1_sg U38526 ( .A(n50185), .B(n50174), .X(n24077) );
  nor_x1_sg U38527 ( .A(n44247), .B(n41872), .X(n24317) );
  inv_x1_sg U38528 ( .A(n24318), .X(n43677) );
  nor_x1_sg U38529 ( .A(n50183), .B(n50178), .X(n24318) );
  nor_x1_sg U38530 ( .A(n44070), .B(n41306), .X(n22061) );
  inv_x1_sg U38531 ( .A(n22062), .X(n43623) );
  nor_x1_sg U38532 ( .A(n50195), .B(n50158), .X(n22062) );
  nor_x1_sg U38533 ( .A(n44072), .B(n41340), .X(n22929) );
  inv_x1_sg U38534 ( .A(n22930), .X(n43728) );
  nor_x1_sg U38535 ( .A(n50191), .B(n50164), .X(n22930) );
  nand_x4_sg U38536 ( .A(n44153), .B(n41869), .X(n40581) );
  inv_x1_sg U38537 ( .A(n29838), .X(n43621) );
  nor_x1_sg U38538 ( .A(n44529), .B(n50084), .X(n29838) );
  inv_x1_sg U38539 ( .A(n30443), .X(n43622) );
  nor_x1_sg U38540 ( .A(n44631), .B(n50074), .X(n30443) );
  nor_x1_sg U38541 ( .A(n41948), .B(n50031), .X(n30698) );
  inv_x1_sg U38542 ( .A(n30699), .X(n43620) );
  nor_x1_sg U38543 ( .A(n24551), .B(n41947), .X(n30699) );
  nor_x1_sg U38544 ( .A(n24548), .B(n30702), .X(n30701) );
  nand_x1_sg U38545 ( .A(n30702), .B(n24548), .X(n30703) );
  nor_x1_sg U38546 ( .A(n44573), .B(n41305), .X(n29824) );
  inv_x1_sg U38547 ( .A(n29825), .X(n43613) );
  nor_x1_sg U38548 ( .A(n49990), .B(n49951), .X(n29825) );
  nor_x1_sg U38549 ( .A(n41946), .B(n49986), .X(n30692) );
  inv_x1_sg U38550 ( .A(n30693), .X(n43616) );
  nor_x1_sg U38551 ( .A(n24600), .B(n41945), .X(n30693) );
  nor_x1_sg U38552 ( .A(n24597), .B(n30928), .X(n30927) );
  nand_x1_sg U38553 ( .A(n30928), .B(n24597), .X(n30929) );
  nor_x1_sg U38554 ( .A(n44571), .B(n41304), .X(n29817) );
  inv_x1_sg U38555 ( .A(n29818), .X(n43609) );
  nor_x1_sg U38556 ( .A(n49945), .B(n49903), .X(n29818) );
  nor_x1_sg U38557 ( .A(n41944), .B(n49941), .X(n30686) );
  inv_x1_sg U38558 ( .A(n30687), .X(n43612) );
  nor_x1_sg U38559 ( .A(n24649), .B(n41943), .X(n30687) );
  nor_x1_sg U38560 ( .A(n24646), .B(n30922), .X(n30921) );
  nand_x1_sg U38561 ( .A(n30922), .B(n24646), .X(n30923) );
  nor_x1_sg U38562 ( .A(n44567), .B(n41302), .X(n29810) );
  inv_x1_sg U38563 ( .A(n29811), .X(n43605) );
  nor_x1_sg U38564 ( .A(n49897), .B(n49856), .X(n29811) );
  nor_x1_sg U38565 ( .A(n44569), .B(n41303), .X(n30679) );
  inv_x1_sg U38566 ( .A(n30680), .X(n43607) );
  nor_x1_sg U38567 ( .A(n49893), .B(n49865), .X(n30680) );
  nor_x1_sg U38568 ( .A(n44563), .B(n41300), .X(n29803) );
  inv_x1_sg U38569 ( .A(n29804), .X(n43601) );
  nor_x1_sg U38570 ( .A(n49850), .B(n49808), .X(n29804) );
  nor_x1_sg U38571 ( .A(n44565), .B(n41301), .X(n30672) );
  inv_x1_sg U38572 ( .A(n30673), .X(n43603) );
  nor_x1_sg U38573 ( .A(n49846), .B(n49817), .X(n30673) );
  nor_x1_sg U38574 ( .A(n42194), .B(n24781), .X(n31117) );
  nand_x1_sg U38575 ( .A(n24781), .B(n42194), .X(n31118) );
  nor_x1_sg U38576 ( .A(n44561), .B(n41299), .X(n29796) );
  inv_x1_sg U38577 ( .A(n29797), .X(n42552) );
  nor_x1_sg U38578 ( .A(n49802), .B(n49761), .X(n29797) );
  nor_x1_sg U38579 ( .A(n42228), .B(n24796), .X(n30133) );
  nand_x1_sg U38580 ( .A(n24796), .B(n42228), .X(n30134) );
  nor_x1_sg U38581 ( .A(n44639), .B(n41577), .X(n30665) );
  inv_x1_sg U38582 ( .A(n30666), .X(n42554) );
  nor_x1_sg U38583 ( .A(n49799), .B(n49770), .X(n30666) );
  nor_x1_sg U38584 ( .A(n44557), .B(n41297), .X(n29789) );
  inv_x1_sg U38585 ( .A(n29790), .X(n43597) );
  nor_x1_sg U38586 ( .A(n49755), .B(n49712), .X(n29790) );
  nor_x1_sg U38587 ( .A(n44559), .B(n41298), .X(n30658) );
  inv_x1_sg U38588 ( .A(n30659), .X(n43599) );
  nor_x1_sg U38589 ( .A(n49751), .B(n49721), .X(n30659) );
  nor_x1_sg U38590 ( .A(n44553), .B(n41295), .X(n29782) );
  inv_x1_sg U38591 ( .A(n29783), .X(n43593) );
  nor_x1_sg U38592 ( .A(n49706), .B(n49665), .X(n29783) );
  nor_x1_sg U38593 ( .A(n44555), .B(n41296), .X(n30651) );
  inv_x1_sg U38594 ( .A(n30652), .X(n43595) );
  nor_x1_sg U38595 ( .A(n49702), .B(n49674), .X(n30652) );
  nor_x1_sg U38596 ( .A(n44517), .B(n41167), .X(n31791) );
  inv_x1_sg U38597 ( .A(n31792), .X(n42574) );
  nor_x1_sg U38598 ( .A(n49649), .B(n49639), .X(n31792) );
  nor_x1_sg U38599 ( .A(n44549), .B(n41293), .X(n29775) );
  inv_x1_sg U38600 ( .A(n29776), .X(n43589) );
  nor_x1_sg U38601 ( .A(n49659), .B(n49618), .X(n29776) );
  nor_x1_sg U38602 ( .A(n44551), .B(n41294), .X(n30644) );
  inv_x1_sg U38603 ( .A(n30645), .X(n43591) );
  nor_x1_sg U38604 ( .A(n49655), .B(n49627), .X(n30645) );
  nor_x1_sg U38605 ( .A(n44515), .B(n41166), .X(n31784) );
  inv_x1_sg U38606 ( .A(n31785), .X(n42572) );
  nor_x1_sg U38607 ( .A(n49602), .B(n49593), .X(n31785) );
  nor_x1_sg U38608 ( .A(n44545), .B(n41291), .X(n29768) );
  inv_x1_sg U38609 ( .A(n29769), .X(n43585) );
  nor_x1_sg U38610 ( .A(n49612), .B(n49572), .X(n29769) );
  nor_x1_sg U38611 ( .A(n44547), .B(n41292), .X(n30637) );
  inv_x1_sg U38612 ( .A(n30638), .X(n43587) );
  nor_x1_sg U38613 ( .A(n49608), .B(n49581), .X(n30638) );
  nor_x1_sg U38614 ( .A(n44513), .B(n41580), .X(n31777) );
  inv_x1_sg U38615 ( .A(n31778), .X(n42570) );
  nor_x1_sg U38616 ( .A(n49556), .B(n49547), .X(n31778) );
  nor_x1_sg U38617 ( .A(n44541), .B(n41289), .X(n29761) );
  inv_x1_sg U38618 ( .A(n29762), .X(n43581) );
  nor_x1_sg U38619 ( .A(n49566), .B(n49525), .X(n29762) );
  nor_x1_sg U38620 ( .A(n44543), .B(n41290), .X(n30630) );
  inv_x1_sg U38621 ( .A(n30631), .X(n43583) );
  nor_x1_sg U38622 ( .A(n49562), .B(n49534), .X(n30631) );
  nor_x1_sg U38623 ( .A(n44511), .B(n41331), .X(n31770) );
  inv_x1_sg U38624 ( .A(n31771), .X(n42568) );
  nor_x1_sg U38625 ( .A(n49509), .B(n49499), .X(n31771) );
  nor_x1_sg U38626 ( .A(n44539), .B(n41288), .X(n29754) );
  inv_x1_sg U38627 ( .A(n29755), .X(n43579) );
  nor_x1_sg U38628 ( .A(n49519), .B(n49478), .X(n29755) );
  nor_x1_sg U38629 ( .A(n49506), .B(n49504), .X(n32098) );
  inv_x1_sg U38630 ( .A(n32099), .X(n42521) );
  nor_x1_sg U38631 ( .A(n32100), .B(n32101), .X(n32099) );
  nor_x1_sg U38632 ( .A(n44637), .B(n41334), .X(n30623) );
  inv_x1_sg U38633 ( .A(n30624), .X(n43695) );
  nor_x1_sg U38634 ( .A(n49515), .B(n49487), .X(n30624) );
  nor_x1_sg U38635 ( .A(n44509), .B(n41579), .X(n31763) );
  inv_x1_sg U38636 ( .A(n31764), .X(n42566) );
  nor_x1_sg U38637 ( .A(n49462), .B(n49453), .X(n31764) );
  nor_x1_sg U38638 ( .A(n44535), .B(n41286), .X(n29747) );
  inv_x1_sg U38639 ( .A(n29748), .X(n43575) );
  nor_x1_sg U38640 ( .A(n49472), .B(n49432), .X(n29748) );
  nor_x1_sg U38641 ( .A(n44537), .B(n41287), .X(n30616) );
  inv_x1_sg U38642 ( .A(n30617), .X(n43577) );
  nor_x1_sg U38643 ( .A(n49468), .B(n49441), .X(n30617) );
  nor_x1_sg U38644 ( .A(n44507), .B(n41330), .X(n31756) );
  inv_x1_sg U38645 ( .A(n31757), .X(n42564) );
  nor_x1_sg U38646 ( .A(n49416), .B(n49408), .X(n31757) );
  nor_x1_sg U38647 ( .A(n44533), .B(n41285), .X(n29740) );
  inv_x1_sg U38648 ( .A(n29741), .X(n43573) );
  nor_x1_sg U38649 ( .A(n49426), .B(n49386), .X(n29741) );
  nand_x4_sg U38650 ( .A(n40907), .B(n42523), .X(n40582) );
  inv_x8_sg U38651 ( .A(n40582), .X(n32089) );
  nor_x1_sg U38652 ( .A(n44635), .B(n41333), .X(n30609) );
  inv_x1_sg U38653 ( .A(n30610), .X(n43693) );
  nor_x1_sg U38654 ( .A(n49422), .B(n49395), .X(n30610) );
  nor_x1_sg U38655 ( .A(n44505), .B(n41165), .X(n31749) );
  inv_x1_sg U38656 ( .A(n31750), .X(n42562) );
  nor_x1_sg U38657 ( .A(n49370), .B(n49363), .X(n31750) );
  nor_x1_sg U38658 ( .A(n44531), .B(n41284), .X(n29733) );
  inv_x1_sg U38659 ( .A(n29734), .X(n43571) );
  nor_x1_sg U38660 ( .A(n49380), .B(n49342), .X(n29734) );
  nor_x1_sg U38661 ( .A(n41241), .B(n32083), .X(n32080) );
  nand_x1_sg U38662 ( .A(n41241), .B(n32083), .X(n32081) );
  nor_x1_sg U38663 ( .A(n44649), .B(n41337), .X(n30602) );
  inv_x1_sg U38664 ( .A(n30603), .X(n43709) );
  nor_x1_sg U38665 ( .A(n49376), .B(n49351), .X(n30603) );
  nor_x1_sg U38666 ( .A(n44621), .B(n41329), .X(n31742) );
  inv_x1_sg U38667 ( .A(n31743), .X(n42560) );
  nor_x1_sg U38668 ( .A(n49326), .B(n49315), .X(n31743) );
  nor_x1_sg U38669 ( .A(n44066), .B(n41283), .X(n29726) );
  inv_x1_sg U38670 ( .A(n29727), .X(n43569) );
  nor_x1_sg U38671 ( .A(n49336), .B(n49299), .X(n29727) );
  nor_x1_sg U38672 ( .A(n44068), .B(n41339), .X(n30595) );
  inv_x1_sg U38673 ( .A(n30596), .X(n43726) );
  nor_x1_sg U38674 ( .A(n49332), .B(n49305), .X(n30596) );
  nand_x4_sg U38675 ( .A(n25648), .B(n43558), .X(n40583) );
  inv_x8_sg U38676 ( .A(n40583), .X(n25569) );
  inv_x2_sg U38677 ( .A(n25646), .X(n43558) );
  nand_x2_sg U38678 ( .A(n45127), .B(n51499), .X(n25612) );
  nand_x4_sg U38679 ( .A(n26207), .B(n43556), .X(n40584) );
  inv_x8_sg U38680 ( .A(n40584), .X(n26130) );
  inv_x2_sg U38681 ( .A(n26205), .X(n43556) );
  nand_x4_sg U38682 ( .A(n27602), .B(n43557), .X(n40585) );
  inv_x8_sg U38683 ( .A(n40585), .X(n27525) );
  inv_x2_sg U38684 ( .A(n27600), .X(n43557) );
  nand_x4_sg U38685 ( .A(n41522), .B(n28387), .X(n40586) );
  nand_x4_sg U38686 ( .A(n28998), .B(n43554), .X(n40587) );
  inv_x8_sg U38687 ( .A(n40587), .X(n28921) );
  inv_x2_sg U38688 ( .A(n28996), .X(n43554) );
  nand_x4_sg U38689 ( .A(n29559), .B(n43553), .X(n40588) );
  inv_x8_sg U38690 ( .A(n40588), .X(n29482) );
  inv_x2_sg U38691 ( .A(n29557), .X(n43553) );
  nand_x4_sg U38692 ( .A(n43732), .B(n40902), .X(n40589) );
  inv_x8_sg U38693 ( .A(n40589), .X(n9372) );
  nand_x4_sg U38694 ( .A(n43675), .B(n40900), .X(n40590) );
  inv_x8_sg U38695 ( .A(n40590), .X(n9383) );
  nand_x4_sg U38696 ( .A(n43676), .B(n40898), .X(n40591) );
  inv_x8_sg U38697 ( .A(n40591), .X(n9393) );
  nand_x4_sg U38698 ( .A(n43692), .B(n23057), .X(n40592) );
  inv_x8_sg U38699 ( .A(n40592), .X(n9430) );
  inv_x2_sg U38700 ( .A(n23056), .X(n43692) );
  nand_x4_sg U38701 ( .A(n43673), .B(n43674), .X(n40593) );
  inv_x8_sg U38702 ( .A(n40593), .X(n9447) );
  inv_x2_sg U38703 ( .A(n23032), .X(n43673) );
  nand_x4_sg U38704 ( .A(n23037), .B(n41860), .X(n40594) );
  inv_x8_sg U38705 ( .A(n40594), .X(n9443) );
  inv_x2_sg U38706 ( .A(n23035), .X(n41860) );
  nand_x4_sg U38707 ( .A(n43691), .B(n23283), .X(n40595) );
  inv_x8_sg U38708 ( .A(n40595), .X(n9479) );
  inv_x2_sg U38709 ( .A(n23282), .X(n43691) );
  nand_x4_sg U38710 ( .A(n43668), .B(n43667), .X(n40596) );
  inv_x8_sg U38711 ( .A(n40596), .X(n9488) );
  inv_x2_sg U38712 ( .A(n22159), .X(n43668) );
  nand_x4_sg U38713 ( .A(n43669), .B(n43670), .X(n40597) );
  inv_x8_sg U38714 ( .A(n40597), .X(n9496) );
  inv_x2_sg U38715 ( .A(n23026), .X(n43669) );
  nand_x4_sg U38716 ( .A(n23263), .B(n41859), .X(n40598) );
  inv_x8_sg U38717 ( .A(n40598), .X(n9492) );
  inv_x2_sg U38718 ( .A(n23261), .X(n41859) );
  nand_x4_sg U38719 ( .A(n43690), .B(n23488), .X(n40599) );
  inv_x8_sg U38720 ( .A(n40599), .X(n9528) );
  inv_x2_sg U38721 ( .A(n23487), .X(n43690) );
  nand_x4_sg U38722 ( .A(n43664), .B(n43663), .X(n40600) );
  inv_x8_sg U38723 ( .A(n40600), .X(n9537) );
  inv_x2_sg U38724 ( .A(n22152), .X(n43664) );
  nand_x4_sg U38725 ( .A(n43665), .B(n43666), .X(n40601) );
  inv_x8_sg U38726 ( .A(n40601), .X(n9545) );
  inv_x2_sg U38727 ( .A(n23020), .X(n43665) );
  nand_x4_sg U38728 ( .A(n23257), .B(n41858), .X(n40602) );
  inv_x8_sg U38729 ( .A(n40602), .X(n9541) );
  inv_x2_sg U38730 ( .A(n23255), .X(n41858) );
  nand_x4_sg U38731 ( .A(n43689), .B(n23678), .X(n40603) );
  inv_x8_sg U38732 ( .A(n40603), .X(n9577) );
  inv_x2_sg U38733 ( .A(n23677), .X(n43689) );
  nand_x4_sg U38734 ( .A(n43660), .B(n43659), .X(n40604) );
  inv_x8_sg U38735 ( .A(n40604), .X(n9586) );
  inv_x2_sg U38736 ( .A(n22145), .X(n43660) );
  nand_x4_sg U38737 ( .A(n43662), .B(n43661), .X(n40605) );
  inv_x8_sg U38738 ( .A(n40605), .X(n9593) );
  inv_x2_sg U38739 ( .A(n23013), .X(n43662) );
  nand_x4_sg U38740 ( .A(n43688), .B(n23849), .X(n40606) );
  inv_x8_sg U38741 ( .A(n40606), .X(n9625) );
  inv_x2_sg U38742 ( .A(n23848), .X(n43688) );
  nand_x4_sg U38743 ( .A(n43656), .B(n43655), .X(n40607) );
  inv_x8_sg U38744 ( .A(n40607), .X(n9634) );
  inv_x2_sg U38745 ( .A(n22138), .X(n43656) );
  nand_x4_sg U38746 ( .A(n43658), .B(n43657), .X(n40608) );
  inv_x8_sg U38747 ( .A(n40608), .X(n9641) );
  inv_x2_sg U38748 ( .A(n23006), .X(n43658) );
  nand_x4_sg U38749 ( .A(n43687), .B(n24002), .X(n40609) );
  inv_x8_sg U38750 ( .A(n40609), .X(n9673) );
  inv_x2_sg U38751 ( .A(n24001), .X(n43687) );
  nand_x4_sg U38752 ( .A(n43568), .B(n23452), .X(n40610) );
  inv_x8_sg U38753 ( .A(n40610), .X(n9683) );
  inv_x2_sg U38754 ( .A(n23451), .X(n43568) );
  nand_x4_sg U38755 ( .A(n42557), .B(n42556), .X(n40611) );
  inv_x8_sg U38756 ( .A(n40611), .X(n9682) );
  inv_x2_sg U38757 ( .A(n22131), .X(n42557) );
  nand_x4_sg U38758 ( .A(n43702), .B(n22469), .X(n40612) );
  inv_x8_sg U38759 ( .A(n40612), .X(n9705) );
  inv_x2_sg U38760 ( .A(n22468), .X(n43702) );
  nand_x4_sg U38761 ( .A(n42559), .B(n42558), .X(n40613) );
  inv_x8_sg U38762 ( .A(n40613), .X(n9689) );
  inv_x2_sg U38763 ( .A(n22999), .X(n42559) );
  nand_x4_sg U38764 ( .A(n43686), .B(n24146), .X(n40614) );
  inv_x8_sg U38765 ( .A(n40614), .X(n9720) );
  inv_x2_sg U38766 ( .A(n24145), .X(n43686) );
  nand_x4_sg U38767 ( .A(n43652), .B(n43651), .X(n40615) );
  inv_x8_sg U38768 ( .A(n40615), .X(n9729) );
  inv_x2_sg U38769 ( .A(n22124), .X(n43652) );
  nand_x4_sg U38770 ( .A(n43654), .B(n43653), .X(n40616) );
  inv_x8_sg U38771 ( .A(n40616), .X(n9736) );
  inv_x2_sg U38772 ( .A(n22992), .X(n43654) );
  nand_x4_sg U38773 ( .A(n43685), .B(n24262), .X(n40617) );
  inv_x8_sg U38774 ( .A(n40617), .X(n9768) );
  inv_x2_sg U38775 ( .A(n24261), .X(n43685) );
  nand_x4_sg U38776 ( .A(n43648), .B(n43647), .X(n40618) );
  inv_x8_sg U38777 ( .A(n40618), .X(n9777) );
  inv_x2_sg U38778 ( .A(n22117), .X(n43648) );
  nand_x4_sg U38779 ( .A(n43650), .B(n43649), .X(n40619) );
  inv_x8_sg U38780 ( .A(n40619), .X(n9784) );
  inv_x2_sg U38781 ( .A(n22985), .X(n43650) );
  nand_x4_sg U38782 ( .A(n42535), .B(n42534), .X(n40620) );
  inv_x8_sg U38783 ( .A(n40620), .X(n9812) );
  inv_x2_sg U38784 ( .A(n24125), .X(n42535) );
  nand_x4_sg U38785 ( .A(n43684), .B(n24364), .X(n40621) );
  inv_x8_sg U38786 ( .A(n40621), .X(n9816) );
  inv_x2_sg U38787 ( .A(n24363), .X(n43684) );
  nand_x4_sg U38788 ( .A(n43644), .B(n43643), .X(n40622) );
  inv_x8_sg U38789 ( .A(n40622), .X(n9825) );
  inv_x2_sg U38790 ( .A(n22110), .X(n43644) );
  nand_x4_sg U38791 ( .A(n43646), .B(n43645), .X(n40623) );
  inv_x8_sg U38792 ( .A(n40623), .X(n9832) );
  inv_x2_sg U38793 ( .A(n22978), .X(n43646) );
  nand_x4_sg U38794 ( .A(n42533), .B(n42532), .X(n40624) );
  inv_x8_sg U38795 ( .A(n40624), .X(n9860) );
  inv_x2_sg U38796 ( .A(n24118), .X(n42533) );
  nand_x4_sg U38797 ( .A(n43683), .B(n24357), .X(n40625) );
  inv_x8_sg U38798 ( .A(n40625), .X(n9864) );
  inv_x2_sg U38799 ( .A(n24356), .X(n43683) );
  nand_x4_sg U38800 ( .A(n43640), .B(n43639), .X(n40626) );
  inv_x8_sg U38801 ( .A(n40626), .X(n9873) );
  inv_x2_sg U38802 ( .A(n22103), .X(n43640) );
  nand_x4_sg U38803 ( .A(n43642), .B(n43641), .X(n40627) );
  inv_x8_sg U38804 ( .A(n40627), .X(n9880) );
  inv_x2_sg U38805 ( .A(n22971), .X(n43642) );
  nand_x4_sg U38806 ( .A(n42531), .B(n42530), .X(n40628) );
  inv_x8_sg U38807 ( .A(n40628), .X(n9908) );
  inv_x2_sg U38808 ( .A(n24111), .X(n42531) );
  nand_x4_sg U38809 ( .A(n40904), .B(n43682), .X(n40629) );
  inv_x8_sg U38810 ( .A(n40629), .X(n9912) );
  nand_x4_sg U38811 ( .A(n43636), .B(n43635), .X(n40630) );
  inv_x8_sg U38812 ( .A(n40630), .X(n9921) );
  inv_x2_sg U38813 ( .A(n22096), .X(n43636) );
  nand_x4_sg U38814 ( .A(n43638), .B(n43637), .X(n40631) );
  inv_x8_sg U38815 ( .A(n40631), .X(n9928) );
  inv_x2_sg U38816 ( .A(n22964), .X(n43638) );
  nand_x4_sg U38817 ( .A(n42529), .B(n42528), .X(n40632) );
  inv_x8_sg U38818 ( .A(n40632), .X(n9956) );
  inv_x2_sg U38819 ( .A(n24104), .X(n42529) );
  nand_x4_sg U38820 ( .A(n43681), .B(n40896), .X(n40633) );
  inv_x8_sg U38821 ( .A(n40633), .X(n9960) );
  nand_x4_sg U38822 ( .A(n43634), .B(n43633), .X(n40634) );
  inv_x8_sg U38823 ( .A(n40634), .X(n9969) );
  inv_x2_sg U38824 ( .A(n22089), .X(n43634) );
  nand_x4_sg U38825 ( .A(n42518), .B(n42519), .X(n40635) );
  inv_x8_sg U38826 ( .A(n40635), .X(n9981) );
  inv_x2_sg U38827 ( .A(n24432), .X(n42518) );
  nand_x4_sg U38828 ( .A(n43701), .B(n43700), .X(n40636) );
  inv_x8_sg U38829 ( .A(n40636), .X(n9976) );
  inv_x2_sg U38830 ( .A(n22957), .X(n43701) );
  nand_x4_sg U38831 ( .A(n42527), .B(n42526), .X(n40637) );
  inv_x8_sg U38832 ( .A(n40637), .X(n10005) );
  inv_x2_sg U38833 ( .A(n24097), .X(n42527) );
  nand_x4_sg U38834 ( .A(n43680), .B(n43679), .X(n40638) );
  inv_x8_sg U38835 ( .A(n40638), .X(n10009) );
  inv_x2_sg U38836 ( .A(n24336), .X(n43680) );
  nand_x4_sg U38837 ( .A(n43630), .B(n43629), .X(n40639) );
  inv_x8_sg U38838 ( .A(n40639), .X(n10018) );
  inv_x2_sg U38839 ( .A(n22082), .X(n43630) );
  nand_x4_sg U38840 ( .A(n43632), .B(n43631), .X(n40640) );
  inv_x8_sg U38841 ( .A(n40640), .X(n10025) );
  inv_x2_sg U38842 ( .A(n22950), .X(n43632) );
  nand_x4_sg U38843 ( .A(n42589), .B(n42588), .X(n40641) );
  inv_x8_sg U38844 ( .A(n40641), .X(n10053) );
  inv_x2_sg U38845 ( .A(n24090), .X(n42589) );
  nand_x4_sg U38846 ( .A(n40579), .B(n40894), .X(n40642) );
  inv_x8_sg U38847 ( .A(n40642), .X(n10057) );
  nand_x4_sg U38848 ( .A(n43628), .B(n43627), .X(n40643) );
  inv_x8_sg U38849 ( .A(n40643), .X(n10066) );
  inv_x2_sg U38850 ( .A(n22075), .X(n43628) );
  nand_x4_sg U38851 ( .A(n43699), .B(n43698), .X(n40644) );
  inv_x8_sg U38852 ( .A(n40644), .X(n10073) );
  inv_x2_sg U38853 ( .A(n22943), .X(n43699) );
  nand_x4_sg U38854 ( .A(n42587), .B(n42586), .X(n40645) );
  inv_x8_sg U38855 ( .A(n40645), .X(n10102) );
  inv_x2_sg U38856 ( .A(n24083), .X(n42587) );
  nand_x4_sg U38857 ( .A(n43720), .B(n43721), .X(n40646) );
  inv_x8_sg U38858 ( .A(n40646), .X(n10106) );
  inv_x2_sg U38859 ( .A(n24324), .X(n43720) );
  nand_x4_sg U38860 ( .A(n43626), .B(n43625), .X(n40647) );
  inv_x8_sg U38861 ( .A(n40647), .X(n10115) );
  inv_x2_sg U38862 ( .A(n22068), .X(n43626) );
  nand_x4_sg U38863 ( .A(n41544), .B(n24415), .X(n40648) );
  inv_x8_sg U38864 ( .A(n40648), .X(n10127) );
  inv_x2_sg U38865 ( .A(n24414), .X(n41544) );
  nand_x4_sg U38866 ( .A(n43723), .B(n43722), .X(n40649) );
  inv_x8_sg U38867 ( .A(n40649), .X(n10122) );
  inv_x2_sg U38868 ( .A(n22936), .X(n43723) );
  nand_x4_sg U38869 ( .A(n42525), .B(n42524), .X(n40650) );
  inv_x8_sg U38870 ( .A(n40650), .X(n10151) );
  inv_x2_sg U38871 ( .A(n24076), .X(n42525) );
  nand_x4_sg U38872 ( .A(n43678), .B(n43677), .X(n40651) );
  inv_x8_sg U38873 ( .A(n40651), .X(n10155) );
  inv_x2_sg U38874 ( .A(n24317), .X(n43678) );
  nand_x4_sg U38875 ( .A(n43624), .B(n43623), .X(n40652) );
  inv_x8_sg U38876 ( .A(n40652), .X(n10164) );
  inv_x2_sg U38877 ( .A(n22061), .X(n43624) );
  nand_x4_sg U38878 ( .A(n43729), .B(n43728), .X(n40653) );
  inv_x8_sg U38879 ( .A(n40653), .X(n10171) );
  inv_x2_sg U38880 ( .A(n22929), .X(n43729) );
  inv_x2_sg U38881 ( .A(n41345), .X(n41346) );
  inv_x1_sg U38882 ( .A(n11939), .X(n41345) );
  inv_x2_sg U38883 ( .A(n41343), .X(n41344) );
  inv_x1_sg U38884 ( .A(n13501), .X(n41343) );
  inv_x2_sg U38885 ( .A(n41341), .X(n41342) );
  inv_x1_sg U38886 ( .A(n15834), .X(n41341) );
  inv_x2_sg U38887 ( .A(n41176), .X(n41177) );
  inv_x1_sg U38888 ( .A(n19716), .X(n41176) );
  inv_x1_sg U38889 ( .A(n30467), .X(n43731) );
  nor_x1_sg U38890 ( .A(n44623), .B(n50051), .X(n30467) );
  nand_x4_sg U38891 ( .A(n43621), .B(n40901), .X(n40654) );
  inv_x8_sg U38892 ( .A(n40654), .X(n24498) );
  nand_x4_sg U38893 ( .A(n43622), .B(n40899), .X(n40655) );
  inv_x8_sg U38894 ( .A(n40655), .X(n24506) );
  nor_x1_sg U38895 ( .A(n42254), .B(n30484), .X(n30722) );
  nand_x1_sg U38896 ( .A(n30484), .B(n42254), .X(n30723) );
  nand_x4_sg U38897 ( .A(n43619), .B(n43620), .X(n40656) );
  inv_x8_sg U38898 ( .A(n40656), .X(n24555) );
  inv_x2_sg U38899 ( .A(n30698), .X(n43619) );
  nand_x4_sg U38900 ( .A(n30703), .B(n41857), .X(n40657) );
  inv_x8_sg U38901 ( .A(n40657), .X(n24551) );
  inv_x2_sg U38902 ( .A(n30701), .X(n41857) );
  nor_x1_sg U38903 ( .A(n42258), .B(n30739), .X(n30948) );
  nand_x1_sg U38904 ( .A(n30739), .B(n42258), .X(n30949) );
  nand_x4_sg U38905 ( .A(n43614), .B(n43613), .X(n40658) );
  inv_x8_sg U38906 ( .A(n40658), .X(n24596) );
  inv_x2_sg U38907 ( .A(n29824), .X(n43614) );
  nand_x4_sg U38908 ( .A(n43615), .B(n43616), .X(n40659) );
  inv_x8_sg U38909 ( .A(n40659), .X(n24604) );
  inv_x2_sg U38910 ( .A(n30692), .X(n43615) );
  nand_x4_sg U38911 ( .A(n30929), .B(n41856), .X(n40660) );
  inv_x8_sg U38912 ( .A(n40660), .X(n24600) );
  inv_x2_sg U38913 ( .A(n30927), .X(n41856) );
  nor_x1_sg U38914 ( .A(n42250), .B(n30965), .X(n31153) );
  nand_x1_sg U38915 ( .A(n30965), .B(n42250), .X(n31154) );
  nand_x4_sg U38916 ( .A(n43610), .B(n43609), .X(n40661) );
  inv_x8_sg U38917 ( .A(n40661), .X(n24645) );
  inv_x2_sg U38918 ( .A(n29817), .X(n43610) );
  nand_x4_sg U38919 ( .A(n43611), .B(n43612), .X(n40662) );
  inv_x8_sg U38920 ( .A(n40662), .X(n24653) );
  inv_x2_sg U38921 ( .A(n30686), .X(n43611) );
  nand_x4_sg U38922 ( .A(n30923), .B(n41855), .X(n40663) );
  inv_x8_sg U38923 ( .A(n40663), .X(n24649) );
  inv_x2_sg U38924 ( .A(n30921), .X(n41855) );
  nor_x1_sg U38925 ( .A(n42256), .B(n31170), .X(n31343) );
  nand_x1_sg U38926 ( .A(n31170), .B(n42256), .X(n31344) );
  nand_x4_sg U38927 ( .A(n43606), .B(n43605), .X(n40664) );
  inv_x8_sg U38928 ( .A(n40664), .X(n24694) );
  inv_x2_sg U38929 ( .A(n29810), .X(n43606) );
  nand_x4_sg U38930 ( .A(n43608), .B(n43607), .X(n40665) );
  inv_x8_sg U38931 ( .A(n40665), .X(n24701) );
  inv_x2_sg U38932 ( .A(n30679), .X(n43608) );
  nor_x1_sg U38933 ( .A(n42246), .B(n31360), .X(n31514) );
  nand_x1_sg U38934 ( .A(n31360), .B(n42246), .X(n31515) );
  nand_x4_sg U38935 ( .A(n43602), .B(n43601), .X(n40666) );
  inv_x8_sg U38936 ( .A(n40666), .X(n24742) );
  inv_x2_sg U38937 ( .A(n29803), .X(n43602) );
  nand_x4_sg U38938 ( .A(n43604), .B(n43603), .X(n40667) );
  inv_x8_sg U38939 ( .A(n40667), .X(n24749) );
  inv_x2_sg U38940 ( .A(n30672), .X(n43604) );
  nor_x1_sg U38941 ( .A(n42280), .B(n31531), .X(n31667) );
  nand_x1_sg U38942 ( .A(n31531), .B(n42280), .X(n31668) );
  nand_x4_sg U38943 ( .A(n43567), .B(n31118), .X(n40668) );
  inv_x8_sg U38944 ( .A(n40668), .X(n24791) );
  inv_x2_sg U38945 ( .A(n31117), .X(n43567) );
  nand_x4_sg U38946 ( .A(n42553), .B(n42552), .X(n40669) );
  inv_x8_sg U38947 ( .A(n40669), .X(n24790) );
  inv_x2_sg U38948 ( .A(n29796), .X(n42553) );
  nand_x4_sg U38949 ( .A(n43697), .B(n30134), .X(n40670) );
  inv_x8_sg U38950 ( .A(n40670), .X(n24813) );
  inv_x2_sg U38951 ( .A(n30133), .X(n43697) );
  nand_x4_sg U38952 ( .A(n42555), .B(n42554), .X(n40671) );
  inv_x8_sg U38953 ( .A(n40671), .X(n24797) );
  inv_x2_sg U38954 ( .A(n30665), .X(n42555) );
  nor_x1_sg U38955 ( .A(n42242), .B(n31684), .X(n31811) );
  nand_x1_sg U38956 ( .A(n31684), .B(n42242), .X(n31812) );
  nand_x4_sg U38957 ( .A(n43598), .B(n43597), .X(n40672) );
  inv_x8_sg U38958 ( .A(n40672), .X(n24837) );
  inv_x2_sg U38959 ( .A(n29789), .X(n43598) );
  nand_x4_sg U38960 ( .A(n43600), .B(n43599), .X(n40673) );
  inv_x8_sg U38961 ( .A(n40673), .X(n24844) );
  inv_x2_sg U38962 ( .A(n30658), .X(n43600) );
  nor_x1_sg U38963 ( .A(n42240), .B(n31828), .X(n31927) );
  nand_x1_sg U38964 ( .A(n31828), .B(n42240), .X(n31928) );
  nand_x4_sg U38965 ( .A(n43594), .B(n43593), .X(n40674) );
  inv_x8_sg U38966 ( .A(n40674), .X(n24885) );
  inv_x2_sg U38967 ( .A(n29782), .X(n43594) );
  nand_x4_sg U38968 ( .A(n43596), .B(n43595), .X(n40675) );
  inv_x8_sg U38969 ( .A(n40675), .X(n24892) );
  inv_x2_sg U38970 ( .A(n30651), .X(n43596) );
  nor_x1_sg U38971 ( .A(n42236), .B(n31944), .X(n32029) );
  nand_x1_sg U38972 ( .A(n31944), .B(n42236), .X(n32030) );
  nand_x4_sg U38973 ( .A(n42575), .B(n42574), .X(n40676) );
  inv_x8_sg U38974 ( .A(n40676), .X(n24920) );
  inv_x2_sg U38975 ( .A(n31791), .X(n42575) );
  nand_x4_sg U38976 ( .A(n43590), .B(n43589), .X(n40677) );
  inv_x8_sg U38977 ( .A(n40677), .X(n24933) );
  inv_x2_sg U38978 ( .A(n29775), .X(n43590) );
  nand_x4_sg U38979 ( .A(n43592), .B(n43591), .X(n40678) );
  inv_x8_sg U38980 ( .A(n40678), .X(n24940) );
  inv_x2_sg U38981 ( .A(n30644), .X(n43592) );
  nor_x1_sg U38982 ( .A(n42232), .B(n32024), .X(n32022) );
  nand_x1_sg U38983 ( .A(n32024), .B(n42232), .X(n32023) );
  nand_x4_sg U38984 ( .A(n42573), .B(n42572), .X(n40679) );
  inv_x8_sg U38985 ( .A(n40679), .X(n24968) );
  inv_x2_sg U38986 ( .A(n31784), .X(n42573) );
  nand_x4_sg U38987 ( .A(n43586), .B(n43585), .X(n40680) );
  inv_x8_sg U38988 ( .A(n40680), .X(n24981) );
  inv_x2_sg U38989 ( .A(n29768), .X(n43586) );
  nand_x4_sg U38990 ( .A(n43588), .B(n43587), .X(n40681) );
  inv_x8_sg U38991 ( .A(n40681), .X(n24988) );
  inv_x2_sg U38992 ( .A(n30637), .X(n43588) );
  inv_x1_sg U38993 ( .A(n32016), .X(n43712) );
  nor_x1_sg U38994 ( .A(n49554), .B(n49552), .X(n32016) );
  nand_x4_sg U38995 ( .A(n42571), .B(n42570), .X(n40682) );
  inv_x8_sg U38996 ( .A(n40682), .X(n25016) );
  inv_x2_sg U38997 ( .A(n31777), .X(n42571) );
  nand_x4_sg U38998 ( .A(n43582), .B(n43581), .X(n40683) );
  inv_x8_sg U38999 ( .A(n40683), .X(n25029) );
  inv_x2_sg U39000 ( .A(n29761), .X(n43582) );
  nand_x4_sg U39001 ( .A(n43584), .B(n43583), .X(n40684) );
  inv_x8_sg U39002 ( .A(n40684), .X(n25036) );
  inv_x2_sg U39003 ( .A(n30630), .X(n43584) );
  inv_x1_sg U39004 ( .A(n32009), .X(n43711) );
  nor_x1_sg U39005 ( .A(n41614), .B(n49507), .X(n32009) );
  nand_x4_sg U39006 ( .A(n42569), .B(n42568), .X(n40685) );
  inv_x8_sg U39007 ( .A(n40685), .X(n25064) );
  inv_x2_sg U39008 ( .A(n31770), .X(n42569) );
  nand_x4_sg U39009 ( .A(n43580), .B(n43579), .X(n40686) );
  inv_x8_sg U39010 ( .A(n40686), .X(n25077) );
  inv_x2_sg U39011 ( .A(n29754), .X(n43580) );
  nand_x4_sg U39012 ( .A(n42520), .B(n42521), .X(n40687) );
  inv_x8_sg U39013 ( .A(n40687), .X(n25089) );
  inv_x2_sg U39014 ( .A(n32098), .X(n42520) );
  nand_x4_sg U39015 ( .A(n43696), .B(n43695), .X(n40688) );
  inv_x8_sg U39016 ( .A(n40688), .X(n25084) );
  inv_x2_sg U39017 ( .A(n30623), .X(n43696) );
  nor_x1_sg U39018 ( .A(n45489), .B(n41170), .X(n32002) );
  inv_x1_sg U39019 ( .A(n32003), .X(n43707) );
  nor_x1_sg U39020 ( .A(n49460), .B(n49458), .X(n32003) );
  nand_x4_sg U39021 ( .A(n42567), .B(n42566), .X(n40689) );
  inv_x8_sg U39022 ( .A(n40689), .X(n25113) );
  inv_x2_sg U39023 ( .A(n31763), .X(n42567) );
  nand_x4_sg U39024 ( .A(n43576), .B(n43575), .X(n40690) );
  inv_x8_sg U39025 ( .A(n40690), .X(n25126) );
  inv_x2_sg U39026 ( .A(n29747), .X(n43576) );
  nand_x4_sg U39027 ( .A(n43578), .B(n43577), .X(n40691) );
  inv_x8_sg U39028 ( .A(n40691), .X(n25133) );
  inv_x2_sg U39029 ( .A(n30616), .X(n43578) );
  nand_x1_sg U39030 ( .A(n41140), .B(n25186), .X(n40692) );
  nand_x4_sg U39031 ( .A(n42565), .B(n42564), .X(n40693) );
  inv_x8_sg U39032 ( .A(n40693), .X(n25161) );
  inv_x2_sg U39033 ( .A(n31756), .X(n42565) );
  nand_x4_sg U39034 ( .A(n43574), .B(n43573), .X(n40694) );
  inv_x8_sg U39035 ( .A(n40694), .X(n25174) );
  inv_x2_sg U39036 ( .A(n29740), .X(n43574) );
  nand_x4_sg U39037 ( .A(n43694), .B(n43693), .X(n40695) );
  inv_x8_sg U39038 ( .A(n40695), .X(n25181) );
  inv_x2_sg U39039 ( .A(n30609), .X(n43694) );
  nor_x1_sg U39040 ( .A(n41612), .B(n41959), .X(n31990) );
  inv_x1_sg U39041 ( .A(n31991), .X(n43706) );
  nor_x1_sg U39042 ( .A(n25235), .B(n41611), .X(n31991) );
  nand_x4_sg U39043 ( .A(n42563), .B(n42562), .X(n40696) );
  inv_x8_sg U39044 ( .A(n40696), .X(n25210) );
  inv_x2_sg U39045 ( .A(n31749), .X(n42563) );
  nand_x4_sg U39046 ( .A(n43572), .B(n43571), .X(n40697) );
  inv_x8_sg U39047 ( .A(n40697), .X(n25223) );
  inv_x2_sg U39048 ( .A(n29733), .X(n43572) );
  nand_x4_sg U39049 ( .A(n41543), .B(n32081), .X(n40698) );
  inv_x8_sg U39050 ( .A(n40698), .X(n25235) );
  inv_x2_sg U39051 ( .A(n32080), .X(n41543) );
  nand_x4_sg U39052 ( .A(n43710), .B(n43709), .X(n40699) );
  inv_x8_sg U39053 ( .A(n40699), .X(n25230) );
  inv_x2_sg U39054 ( .A(n30602), .X(n43710) );
  nor_x1_sg U39055 ( .A(n44245), .B(n41873), .X(n31983) );
  inv_x1_sg U39056 ( .A(n31984), .X(n43703) );
  nor_x1_sg U39057 ( .A(n49324), .B(n49319), .X(n31984) );
  nand_x4_sg U39058 ( .A(n42561), .B(n42560), .X(n40700) );
  inv_x8_sg U39059 ( .A(n40700), .X(n25259) );
  inv_x2_sg U39060 ( .A(n31742), .X(n42561) );
  nand_x4_sg U39061 ( .A(n43570), .B(n43569), .X(n40701) );
  inv_x8_sg U39062 ( .A(n40701), .X(n25272) );
  inv_x2_sg U39063 ( .A(n29726), .X(n43570) );
  nand_x4_sg U39064 ( .A(n43727), .B(n43726), .X(n40702) );
  inv_x8_sg U39065 ( .A(n40702), .X(n25279) );
  inv_x2_sg U39066 ( .A(n30595), .X(n43727) );
  nand_x4_sg U39067 ( .A(n25613), .B(n25633), .X(n25627) );
  nand_x1_sg U39068 ( .A(n25610), .B(n25612), .X(n25633) );
  nand_x4_sg U39069 ( .A(n43731), .B(n40903), .X(n40703) );
  inv_x8_sg U39070 ( .A(n40703), .X(n24483) );
  nand_x4_sg U39071 ( .A(n43719), .B(n30723), .X(n40704) );
  inv_x8_sg U39072 ( .A(n40704), .X(n24533) );
  inv_x2_sg U39073 ( .A(n30722), .X(n43719) );
  nand_x4_sg U39074 ( .A(n43725), .B(n30949), .X(n40705) );
  inv_x8_sg U39075 ( .A(n40705), .X(n24582) );
  inv_x2_sg U39076 ( .A(n30948), .X(n43725) );
  nand_x4_sg U39077 ( .A(n43718), .B(n31154), .X(n40706) );
  inv_x8_sg U39078 ( .A(n40706), .X(n24631) );
  inv_x2_sg U39079 ( .A(n31153), .X(n43718) );
  nand_x4_sg U39080 ( .A(n43724), .B(n31344), .X(n40707) );
  inv_x8_sg U39081 ( .A(n40707), .X(n24680) );
  inv_x2_sg U39082 ( .A(n31343), .X(n43724) );
  nand_x4_sg U39083 ( .A(n43717), .B(n31515), .X(n40708) );
  inv_x8_sg U39084 ( .A(n40708), .X(n24728) );
  inv_x2_sg U39085 ( .A(n31514), .X(n43717) );
  nand_x4_sg U39086 ( .A(n43730), .B(n31668), .X(n40709) );
  inv_x8_sg U39087 ( .A(n40709), .X(n24776) );
  inv_x2_sg U39088 ( .A(n31667), .X(n43730) );
  nand_x4_sg U39089 ( .A(n43716), .B(n31812), .X(n40710) );
  inv_x8_sg U39090 ( .A(n40710), .X(n24823) );
  inv_x2_sg U39091 ( .A(n31811), .X(n43716) );
  nand_x4_sg U39092 ( .A(n43715), .B(n31928), .X(n40711) );
  inv_x8_sg U39093 ( .A(n40711), .X(n24871) );
  inv_x2_sg U39094 ( .A(n31927), .X(n43715) );
  nand_x4_sg U39095 ( .A(n43714), .B(n32030), .X(n40712) );
  inv_x8_sg U39096 ( .A(n40712), .X(n24919) );
  inv_x2_sg U39097 ( .A(n32029), .X(n43714) );
  nand_x4_sg U39098 ( .A(n43713), .B(n32023), .X(n40713) );
  inv_x8_sg U39099 ( .A(n40713), .X(n24967) );
  inv_x2_sg U39100 ( .A(n32022), .X(n43713) );
  nand_x4_sg U39101 ( .A(n40905), .B(n43712), .X(n40714) );
  inv_x8_sg U39102 ( .A(n40714), .X(n25015) );
  nand_x4_sg U39103 ( .A(n43711), .B(n40897), .X(n40715) );
  inv_x8_sg U39104 ( .A(n40715), .X(n25063) );
  nand_x4_sg U39105 ( .A(n43708), .B(n43707), .X(n40716) );
  inv_x8_sg U39106 ( .A(n40716), .X(n25112) );
  inv_x2_sg U39107 ( .A(n32002), .X(n43708) );
  nand_x4_sg U39108 ( .A(n40692), .B(n40895), .X(n40717) );
  inv_x8_sg U39109 ( .A(n40717), .X(n25160) );
  nand_x4_sg U39110 ( .A(n43705), .B(n43706), .X(n40718) );
  inv_x8_sg U39111 ( .A(n40718), .X(n25209) );
  inv_x2_sg U39112 ( .A(n31990), .X(n43705) );
  nand_x4_sg U39113 ( .A(n43704), .B(n43703), .X(n40719) );
  inv_x8_sg U39114 ( .A(n40719), .X(n25258) );
  inv_x2_sg U39115 ( .A(n31983), .X(n43704) );
  nor_x1_sg U39116 ( .A(n44249), .B(n51515), .X(n25630) );
  inv_x1_sg U39117 ( .A(n25631), .X(n43733) );
  nor_x1_sg U39118 ( .A(n51516), .B(n25627), .X(n25631) );
  nand_x4_sg U39119 ( .A(n43734), .B(n43733), .X(n40720) );
  inv_x8_sg U39120 ( .A(n40720), .X(n10907) );
  inv_x2_sg U39121 ( .A(n25630), .X(n43734) );
  nor_x1_sg U39122 ( .A(n39300), .B(n46638), .X(n39306) );
  inv_x1_sg U39123 ( .A(n46672), .X(n46662) );
  inv_x4_sg U39124 ( .A(n46659), .X(n46658) );
  inv_x2_sg U39125 ( .A(n39306), .X(n46660) );
  nor_x1_sg U39126 ( .A(n11821), .B(n11782), .X(n11819) );
  nor_x1_sg U39127 ( .A(n51714), .B(n51731), .X(n11804) );
  nor_x1_sg U39128 ( .A(n12596), .B(n12554), .X(n12594) );
  nor_x1_sg U39129 ( .A(n12580), .B(n12550), .X(n12578) );
  inv_x2_sg U39130 ( .A(n52050), .X(n41587) );
  inv_x1_sg U39131 ( .A(n12532), .X(n52050) );
  nor_x1_sg U39132 ( .A(n13378), .B(n13335), .X(n13376) );
  nor_x1_sg U39133 ( .A(n13362), .B(n13331), .X(n13360) );
  inv_x2_sg U39134 ( .A(n52327), .X(n42770) );
  inv_x1_sg U39135 ( .A(n13313), .X(n52327) );
  nor_x1_sg U39136 ( .A(n14158), .B(n14115), .X(n14156) );
  nor_x1_sg U39137 ( .A(n14142), .B(n14111), .X(n14140) );
  inv_x2_sg U39138 ( .A(n52602), .X(n42768) );
  inv_x1_sg U39139 ( .A(n14093), .X(n52602) );
  nor_x1_sg U39140 ( .A(n14933), .B(n14895), .X(n14931) );
  inv_x2_sg U39141 ( .A(n14908), .X(n41821) );
  nor_x1_sg U39142 ( .A(n14748), .B(n52836), .X(n14908) );
  nor_x1_sg U39143 ( .A(n15711), .B(n15668), .X(n15709) );
  nor_x1_sg U39144 ( .A(n15695), .B(n15664), .X(n15693) );
  inv_x2_sg U39145 ( .A(n53161), .X(n42766) );
  inv_x1_sg U39146 ( .A(n15646), .X(n53161) );
  nor_x1_sg U39147 ( .A(n17277), .B(n17234), .X(n17275) );
  nor_x1_sg U39148 ( .A(n17261), .B(n17230), .X(n17259) );
  inv_x2_sg U39149 ( .A(n53719), .X(n42762) );
  inv_x1_sg U39150 ( .A(n17212), .X(n53719) );
  nor_x1_sg U39151 ( .A(n18054), .B(n18016), .X(n18052) );
  inv_x2_sg U39152 ( .A(n18029), .X(n41819) );
  nor_x1_sg U39153 ( .A(n17869), .B(n53956), .X(n18029) );
  inv_x2_sg U39154 ( .A(n18808), .X(n54245) );
  nor_x1_sg U39155 ( .A(n19599), .B(n19561), .X(n19597) );
  inv_x2_sg U39156 ( .A(n19574), .X(n41817) );
  nor_x1_sg U39157 ( .A(n19414), .B(n54521), .X(n19574) );
  inv_x2_sg U39158 ( .A(n20344), .X(n41813) );
  nor_x1_sg U39159 ( .A(n20182), .B(n54806), .X(n20344) );
  nor_x1_sg U39160 ( .A(n21143), .B(n21105), .X(n21141) );
  inv_x2_sg U39161 ( .A(n21118), .X(n41815) );
  nor_x1_sg U39162 ( .A(n20958), .B(n55089), .X(n21118) );
  inv_x2_sg U39163 ( .A(n21889), .X(n41811) );
  nor_x1_sg U39164 ( .A(n21727), .B(n55374), .X(n21889) );
  inv_x2_sg U39165 ( .A(n10862), .X(n41525) );
  nor_x1_sg U39166 ( .A(n51461), .B(n11010), .X(n10862) );
  inv_x2_sg U39167 ( .A(n10861), .X(n41741) );
  nor_x1_sg U39168 ( .A(n11004), .B(n11005), .X(n10861) );
  inv_x2_sg U39169 ( .A(n11819), .X(n43467) );
  inv_x2_sg U39170 ( .A(n11804), .X(n43549) );
  inv_x2_sg U39171 ( .A(n11733), .X(n43048) );
  nor_x1_sg U39172 ( .A(n11737), .B(n11738), .X(n11733) );
  inv_x2_sg U39173 ( .A(n11641), .X(n41769) );
  nor_x1_sg U39174 ( .A(n11788), .B(n11789), .X(n11641) );
  inv_x2_sg U39175 ( .A(n11642), .X(n41533) );
  nor_x1_sg U39176 ( .A(n51742), .B(n11794), .X(n11642) );
  inv_x2_sg U39177 ( .A(n12594), .X(n43457) );
  inv_x2_sg U39178 ( .A(n12578), .X(n43543) );
  inv_x2_sg U39179 ( .A(n12539), .X(n42275) );
  nor_x1_sg U39180 ( .A(n42278), .B(n52020), .X(n12539) );
  inv_x2_sg U39181 ( .A(n12603), .X(n52017) );
  inv_x2_sg U39182 ( .A(n12513), .X(n43046) );
  nor_x1_sg U39183 ( .A(n12517), .B(n12518), .X(n12513) );
  inv_x2_sg U39184 ( .A(n13376), .X(n43455) );
  inv_x2_sg U39185 ( .A(n13360), .X(n43541) );
  inv_x2_sg U39186 ( .A(n13385), .X(n52293) );
  inv_x2_sg U39187 ( .A(n13294), .X(n43044) );
  nor_x1_sg U39188 ( .A(n13298), .B(n13299), .X(n13294) );
  inv_x2_sg U39189 ( .A(n13320), .X(n42271) );
  nor_x1_sg U39190 ( .A(n42274), .B(n52296), .X(n13320) );
  inv_x2_sg U39191 ( .A(n14156), .X(n43453) );
  inv_x2_sg U39192 ( .A(n14140), .X(n43539) );
  inv_x2_sg U39193 ( .A(n14165), .X(n52568) );
  inv_x2_sg U39194 ( .A(n14074), .X(n43042) );
  nor_x1_sg U39195 ( .A(n14078), .B(n14079), .X(n14074) );
  inv_x2_sg U39196 ( .A(n14100), .X(n42267) );
  nor_x1_sg U39197 ( .A(n42270), .B(n52571), .X(n14100) );
  inv_x2_sg U39198 ( .A(n14931), .X(n43465) );
  inv_x2_sg U39199 ( .A(n14753), .X(n41785) );
  nor_x1_sg U39200 ( .A(n14899), .B(n14900), .X(n14753) );
  inv_x2_sg U39201 ( .A(n14754), .X(n41541) );
  nor_x1_sg U39202 ( .A(n14905), .B(n14906), .X(n14754) );
  inv_x2_sg U39203 ( .A(n15709), .X(n43451) );
  inv_x2_sg U39204 ( .A(n15693), .X(n43537) );
  inv_x2_sg U39205 ( .A(n15718), .X(n53127) );
  inv_x2_sg U39206 ( .A(n15627), .X(n43040) );
  nor_x1_sg U39207 ( .A(n15631), .B(n15632), .X(n15627) );
  inv_x2_sg U39208 ( .A(n15653), .X(n42263) );
  nor_x1_sg U39209 ( .A(n42266), .B(n53130), .X(n15653) );
  nor_x1_sg U39210 ( .A(n16496), .B(n16457), .X(n16494) );
  inv_x2_sg U39211 ( .A(n16316), .X(n41737) );
  nor_x1_sg U39212 ( .A(n16462), .B(n16463), .X(n16316) );
  inv_x2_sg U39213 ( .A(n16317), .X(n41523) );
  nor_x1_sg U39214 ( .A(n16468), .B(n16469), .X(n16317) );
  inv_x2_sg U39215 ( .A(n17275), .X(n43449) );
  inv_x2_sg U39216 ( .A(n17259), .X(n43535) );
  inv_x2_sg U39217 ( .A(n17284), .X(n53685) );
  inv_x2_sg U39218 ( .A(n17193), .X(n43036) );
  nor_x1_sg U39219 ( .A(n17197), .B(n17198), .X(n17193) );
  inv_x2_sg U39220 ( .A(n17219), .X(n42259) );
  nor_x1_sg U39221 ( .A(n42262), .B(n53688), .X(n17219) );
  inv_x2_sg U39222 ( .A(n18052), .X(n43463) );
  inv_x2_sg U39223 ( .A(n17966), .X(n43034) );
  nor_x1_sg U39224 ( .A(n17970), .B(n17971), .X(n17966) );
  inv_x2_sg U39225 ( .A(n17874), .X(n41783) );
  nor_x1_sg U39226 ( .A(n18020), .B(n18021), .X(n17874) );
  inv_x2_sg U39227 ( .A(n17875), .X(n41539) );
  nor_x1_sg U39228 ( .A(n18026), .B(n18027), .X(n17875) );
  inv_x2_sg U39229 ( .A(n18641), .X(n41765) );
  nor_x1_sg U39230 ( .A(n18791), .B(n18792), .X(n18641) );
  inv_x2_sg U39231 ( .A(n18642), .X(n41531) );
  nor_x1_sg U39232 ( .A(n54254), .B(n18797), .X(n18642) );
  inv_x2_sg U39233 ( .A(n19597), .X(n43461) );
  inv_x2_sg U39234 ( .A(n19511), .X(n43032) );
  nor_x1_sg U39235 ( .A(n19515), .B(n19516), .X(n19511) );
  inv_x2_sg U39236 ( .A(n19419), .X(n41781) );
  nor_x1_sg U39237 ( .A(n19565), .B(n19566), .X(n19419) );
  inv_x2_sg U39238 ( .A(n19420), .X(n41537) );
  nor_x1_sg U39239 ( .A(n19571), .B(n19572), .X(n19420) );
  inv_x2_sg U39240 ( .A(n20187), .X(n41763) );
  nor_x1_sg U39241 ( .A(n20335), .B(n20336), .X(n20187) );
  inv_x2_sg U39242 ( .A(n20188), .X(n41529) );
  nor_x1_sg U39243 ( .A(n20341), .B(n20342), .X(n20188) );
  inv_x2_sg U39244 ( .A(n21141), .X(n43459) );
  inv_x2_sg U39245 ( .A(n21055), .X(n43030) );
  nor_x1_sg U39246 ( .A(n21059), .B(n21060), .X(n21055) );
  inv_x2_sg U39247 ( .A(n20963), .X(n41779) );
  nor_x1_sg U39248 ( .A(n21109), .B(n21110), .X(n20963) );
  inv_x2_sg U39249 ( .A(n20964), .X(n41535) );
  nor_x1_sg U39250 ( .A(n21115), .B(n21116), .X(n20964) );
  inv_x2_sg U39251 ( .A(n21732), .X(n41761) );
  nor_x1_sg U39252 ( .A(n21880), .B(n21881), .X(n21732) );
  inv_x2_sg U39253 ( .A(n21733), .X(n41527) );
  nor_x1_sg U39254 ( .A(n21886), .B(n21887), .X(n21733) );
  nor_x1_sg U39255 ( .A(n10614), .B(n10613), .X(n10611) );
  inv_x2_sg U39256 ( .A(n10705), .X(n42322) );
  nor_x1_sg U39257 ( .A(n51420), .B(n10779), .X(n10705) );
  inv_x2_sg U39258 ( .A(n10859), .X(n43354) );
  nor_x1_sg U39259 ( .A(n41526), .B(n41742), .X(n10859) );
  inv_x2_sg U39260 ( .A(n11639), .X(n43356) );
  nor_x1_sg U39261 ( .A(n41534), .B(n41770), .X(n11639) );
  inv_x2_sg U39262 ( .A(n12266), .X(n42312) );
  nor_x1_sg U39263 ( .A(n51975), .B(n12341), .X(n12266) );
  inv_x2_sg U39264 ( .A(n13202), .X(n43108) );
  nor_x1_sg U39265 ( .A(n13340), .B(n13341), .X(n13202) );
  inv_x2_sg U39266 ( .A(n13982), .X(n43106) );
  nor_x1_sg U39267 ( .A(n14120), .B(n14121), .X(n13982) );
  inv_x2_sg U39268 ( .A(n14597), .X(n42334) );
  nor_x1_sg U39269 ( .A(n52810), .B(n14671), .X(n14597) );
  inv_x2_sg U39270 ( .A(n14751), .X(n43364) );
  nor_x1_sg U39271 ( .A(n41542), .B(n41786), .X(n14751) );
  inv_x2_sg U39272 ( .A(n15535), .X(n43104) );
  nor_x1_sg U39273 ( .A(n15673), .B(n15674), .X(n15535) );
  inv_x2_sg U39274 ( .A(n16161), .X(n42310) );
  nor_x1_sg U39275 ( .A(n53364), .B(n16236), .X(n16161) );
  inv_x2_sg U39276 ( .A(n16494), .X(n43447) );
  inv_x2_sg U39277 ( .A(n16407), .X(n43050) );
  nor_x1_sg U39278 ( .A(n16411), .B(n16412), .X(n16407) );
  inv_x2_sg U39279 ( .A(n16314), .X(n43352) );
  nor_x1_sg U39280 ( .A(n41524), .B(n41738), .X(n16314) );
  inv_x2_sg U39281 ( .A(n17101), .X(n43102) );
  nor_x1_sg U39282 ( .A(n17239), .B(n17240), .X(n17101) );
  inv_x2_sg U39283 ( .A(n17718), .X(n42332) );
  nor_x1_sg U39284 ( .A(n53930), .B(n17792), .X(n17718) );
  inv_x2_sg U39285 ( .A(n17872), .X(n43362) );
  nor_x1_sg U39286 ( .A(n41540), .B(n41784), .X(n17872) );
  nor_x1_sg U39287 ( .A(n18396), .B(n18395), .X(n18393) );
  nor_x1_sg U39288 ( .A(n54181), .B(n54161), .X(n18794) );
  inv_x2_sg U39289 ( .A(n18795), .X(n43531) );
  nor_x1_sg U39290 ( .A(n18793), .B(n18796), .X(n18795) );
  inv_x2_sg U39291 ( .A(n18639), .X(n42446) );
  nor_x1_sg U39292 ( .A(n41532), .B(n41766), .X(n18639) );
  inv_x2_sg U39293 ( .A(n19263), .X(n42330) );
  nor_x1_sg U39294 ( .A(n54495), .B(n19337), .X(n19263) );
  inv_x2_sg U39295 ( .A(n19417), .X(n43360) );
  nor_x1_sg U39296 ( .A(n41538), .B(n41782), .X(n19417) );
  inv_x2_sg U39297 ( .A(n20032), .X(n42326) );
  nor_x1_sg U39298 ( .A(n54779), .B(n20105), .X(n20032) );
  nor_x1_sg U39299 ( .A(n54748), .B(n54727), .X(n20338) );
  inv_x2_sg U39300 ( .A(n20339), .X(n43527) );
  nor_x1_sg U39301 ( .A(n20337), .B(n20340), .X(n20339) );
  inv_x2_sg U39302 ( .A(n20185), .X(n42444) );
  nor_x1_sg U39303 ( .A(n41530), .B(n41764), .X(n20185) );
  inv_x2_sg U39304 ( .A(n20807), .X(n42328) );
  nor_x1_sg U39305 ( .A(n55063), .B(n20881), .X(n20807) );
  inv_x2_sg U39306 ( .A(n20961), .X(n43358) );
  nor_x1_sg U39307 ( .A(n41536), .B(n41780), .X(n20961) );
  inv_x2_sg U39308 ( .A(n21577), .X(n42324) );
  nor_x1_sg U39309 ( .A(n55347), .B(n21650), .X(n21577) );
  nor_x1_sg U39310 ( .A(n55316), .B(n55295), .X(n21883) );
  inv_x2_sg U39311 ( .A(n21884), .X(n43523) );
  nor_x1_sg U39312 ( .A(n21882), .B(n21885), .X(n21884) );
  inv_x2_sg U39313 ( .A(n21730), .X(n42442) );
  nor_x1_sg U39314 ( .A(n41528), .B(n41762), .X(n21730) );
  inv_x2_sg U39315 ( .A(n50734), .X(n41200) );
  inv_x1_sg U39316 ( .A(n23300), .X(n50734) );
  inv_x2_sg U39317 ( .A(n50643), .X(n41198) );
  inv_x1_sg U39318 ( .A(n23695), .X(n50643) );
  inv_x2_sg U39319 ( .A(n50551), .X(n41196) );
  inv_x1_sg U39320 ( .A(n24019), .X(n50551) );
  inv_x2_sg U39321 ( .A(n50501), .X(n41194) );
  inv_x1_sg U39322 ( .A(n24279), .X(n50501) );
  inv_x2_sg U39323 ( .A(n50455), .X(n41152) );
  inv_x1_sg U39324 ( .A(n24362), .X(n50455) );
  inv_x2_sg U39325 ( .A(n10507), .X(n41214) );
  nor_x1_sg U39326 ( .A(n46563), .B(n51315), .X(n10507) );
  inv_x2_sg U39327 ( .A(n10508), .X(n41146) );
  inv_x2_sg U39328 ( .A(n10611), .X(n43483) );
  nor_x1_sg U39329 ( .A(n10701), .B(n51370), .X(n10700) );
  inv_x2_sg U39330 ( .A(n10701), .X(n51350) );
  inv_x2_sg U39331 ( .A(n10785), .X(n42281) );
  nor_x1_sg U39332 ( .A(n10743), .B(n51408), .X(n10785) );
  inv_x2_sg U39333 ( .A(n10852), .X(n41238) );
  nor_x1_sg U39334 ( .A(n43355), .B(n51462), .X(n10852) );
  nor_x1_sg U39335 ( .A(n11300), .B(n51620), .X(n11298) );
  nor_x1_sg U39336 ( .A(n51646), .B(n51616), .X(n11480) );
  inv_x2_sg U39337 ( .A(n11481), .X(n43441) );
  nor_x1_sg U39338 ( .A(n11482), .B(n11483), .X(n11481) );
  inv_x2_sg U39339 ( .A(n11712), .X(n41425) );
  nor_x1_sg U39340 ( .A(n11744), .B(n11745), .X(n11712) );
  inv_x2_sg U39341 ( .A(n11632), .X(n41250) );
  nor_x1_sg U39342 ( .A(n43357), .B(n51743), .X(n11632) );
  nor_x1_sg U39343 ( .A(n12080), .B(n51902), .X(n12078) );
  nor_x1_sg U39344 ( .A(n51926), .B(n51908), .X(n12260) );
  inv_x2_sg U39345 ( .A(n12261), .X(n42402) );
  nor_x1_sg U39346 ( .A(n12262), .B(n12263), .X(n12261) );
  inv_x2_sg U39347 ( .A(n12421), .X(n41767) );
  nor_x1_sg U39348 ( .A(n12558), .B(n12559), .X(n12421) );
  inv_x2_sg U39349 ( .A(n12442), .X(n41495) );
  nor_x1_sg U39350 ( .A(n12538), .B(n52044), .X(n12442) );
  inv_x2_sg U39351 ( .A(n12492), .X(n41423) );
  nor_x1_sg U39352 ( .A(n12524), .B(n12525), .X(n12492) );
  nor_x1_sg U39353 ( .A(n12861), .B(n52179), .X(n12859) );
  nor_x1_sg U39354 ( .A(n52202), .B(n52174), .X(n13041) );
  inv_x2_sg U39355 ( .A(n13042), .X(n43437) );
  nor_x1_sg U39356 ( .A(n13043), .B(n13044), .X(n13042) );
  inv_x2_sg U39357 ( .A(n13273), .X(n41421) );
  nor_x1_sg U39358 ( .A(n13305), .B(n13306), .X(n13273) );
  inv_x2_sg U39359 ( .A(n13223), .X(n41493) );
  nor_x1_sg U39360 ( .A(n13319), .B(n52320), .X(n13223) );
  nor_x1_sg U39361 ( .A(n13641), .B(n52454), .X(n13639) );
  nor_x1_sg U39362 ( .A(n52479), .B(n52449), .X(n13821) );
  inv_x2_sg U39363 ( .A(n13822), .X(n43433) );
  nor_x1_sg U39364 ( .A(n13823), .B(n13824), .X(n13822) );
  inv_x2_sg U39365 ( .A(n14053), .X(n41419) );
  nor_x1_sg U39366 ( .A(n14085), .B(n14086), .X(n14053) );
  inv_x2_sg U39367 ( .A(n14003), .X(n41218) );
  nor_x1_sg U39368 ( .A(n14099), .B(n52595), .X(n14003) );
  inv_x2_sg U39369 ( .A(n14398), .X(n42700) );
  nor_x1_sg U39370 ( .A(n46449), .B(n14400), .X(n14398) );
  inv_x2_sg U39371 ( .A(n14399), .X(n41188) );
  nor_x1_sg U39372 ( .A(n52758), .B(n52725), .X(n14591) );
  inv_x2_sg U39373 ( .A(n14592), .X(n42424) );
  nor_x1_sg U39374 ( .A(n14593), .B(n14594), .X(n14592) );
  inv_x2_sg U39375 ( .A(n14824), .X(n41417) );
  nor_x1_sg U39376 ( .A(n14856), .B(n14857), .X(n14824) );
  inv_x2_sg U39377 ( .A(n14744), .X(n41258) );
  nor_x1_sg U39378 ( .A(n43365), .B(n52852), .X(n14744) );
  nor_x1_sg U39379 ( .A(n15194), .B(n53013), .X(n15192) );
  nor_x1_sg U39380 ( .A(n53036), .B(n53008), .X(n15374) );
  inv_x2_sg U39381 ( .A(n15375), .X(n43429) );
  nor_x1_sg U39382 ( .A(n15376), .B(n15377), .X(n15375) );
  inv_x2_sg U39383 ( .A(n15606), .X(n41415) );
  nor_x1_sg U39384 ( .A(n15638), .B(n15639), .X(n15606) );
  inv_x2_sg U39385 ( .A(n15556), .X(n41491) );
  nor_x1_sg U39386 ( .A(n15652), .B(n53154), .X(n15556) );
  nor_x1_sg U39387 ( .A(n15975), .B(n53287), .X(n15973) );
  nor_x1_sg U39388 ( .A(n53314), .B(n53295), .X(n16155) );
  inv_x2_sg U39389 ( .A(n16156), .X(n42396) );
  nor_x1_sg U39390 ( .A(n16157), .B(n16158), .X(n16156) );
  inv_x2_sg U39391 ( .A(n53401), .X(n43176) );
  inv_x1_sg U39392 ( .A(n16451), .X(n53401) );
  inv_x2_sg U39393 ( .A(n16308), .X(n41236) );
  nor_x1_sg U39394 ( .A(n43353), .B(n53412), .X(n16308) );
  nor_x1_sg U39395 ( .A(n16760), .B(n53571), .X(n16758) );
  nor_x1_sg U39396 ( .A(n53594), .B(n53566), .X(n16940) );
  inv_x2_sg U39397 ( .A(n16941), .X(n43425) );
  nor_x1_sg U39398 ( .A(n16942), .B(n16943), .X(n16941) );
  inv_x2_sg U39399 ( .A(n17172), .X(n41413) );
  nor_x1_sg U39400 ( .A(n17204), .B(n17205), .X(n17172) );
  inv_x2_sg U39401 ( .A(n17122), .X(n41489) );
  nor_x1_sg U39402 ( .A(n17218), .B(n53712), .X(n17122) );
  inv_x2_sg U39403 ( .A(n17519), .X(n42698) );
  nor_x1_sg U39404 ( .A(n53788), .B(n53815), .X(n17519) );
  inv_x2_sg U39405 ( .A(n17520), .X(n41186) );
  nor_x1_sg U39406 ( .A(n17533), .B(n17534), .X(n17532) );
  nor_x1_sg U39407 ( .A(n53878), .B(n53845), .X(n17712) );
  inv_x2_sg U39408 ( .A(n17713), .X(n42420) );
  nor_x1_sg U39409 ( .A(n17714), .B(n17715), .X(n17713) );
  inv_x2_sg U39410 ( .A(n17945), .X(n41411) );
  nor_x1_sg U39411 ( .A(n17977), .B(n17978), .X(n17945) );
  inv_x2_sg U39412 ( .A(n17865), .X(n41256) );
  nor_x1_sg U39413 ( .A(n43363), .B(n53972), .X(n17865) );
  inv_x2_sg U39414 ( .A(n18289), .X(n41904) );
  nor_x1_sg U39415 ( .A(n46337), .B(n18291), .X(n18289) );
  inv_x2_sg U39416 ( .A(n18290), .X(n41148) );
  inv_x2_sg U39417 ( .A(n18393), .X(n43485) );
  inv_x2_sg U39418 ( .A(n18483), .X(n54126) );
  inv_x2_sg U39419 ( .A(n18794), .X(n43533) );
  inv_x2_sg U39420 ( .A(n18714), .X(n41409) );
  nor_x1_sg U39421 ( .A(n18746), .B(n18747), .X(n18714) );
  inv_x2_sg U39422 ( .A(n18632), .X(n41248) );
  nor_x1_sg U39423 ( .A(n42447), .B(n54255), .X(n18632) );
  inv_x2_sg U39424 ( .A(n19064), .X(n42696) );
  nor_x1_sg U39425 ( .A(n54353), .B(n54380), .X(n19064) );
  inv_x2_sg U39426 ( .A(n19065), .X(n41184) );
  nor_x1_sg U39427 ( .A(n19078), .B(n19079), .X(n19077) );
  nor_x1_sg U39428 ( .A(n54443), .B(n54410), .X(n19257) );
  inv_x2_sg U39429 ( .A(n19258), .X(n42416) );
  nor_x1_sg U39430 ( .A(n19259), .B(n19260), .X(n19258) );
  inv_x2_sg U39431 ( .A(n19490), .X(n41407) );
  nor_x1_sg U39432 ( .A(n19522), .B(n19523), .X(n19490) );
  inv_x2_sg U39433 ( .A(n19410), .X(n41254) );
  nor_x1_sg U39434 ( .A(n43361), .B(n54537), .X(n19410) );
  inv_x2_sg U39435 ( .A(n19834), .X(n42694) );
  nor_x1_sg U39436 ( .A(n46293), .B(n54669), .X(n19834) );
  inv_x2_sg U39437 ( .A(n19835), .X(n41517) );
  nor_x1_sg U39438 ( .A(n19872), .B(n54661), .X(n19871) );
  nor_x1_sg U39439 ( .A(n20059), .B(n20023), .X(n20060) );
  nor_x1_sg U39440 ( .A(n20028), .B(n54724), .X(n20027) );
  inv_x2_sg U39441 ( .A(n20028), .X(n54704) );
  inv_x2_sg U39442 ( .A(n20338), .X(n43529) );
  inv_x2_sg U39443 ( .A(n20260), .X(n41405) );
  nor_x1_sg U39444 ( .A(n20292), .B(n20293), .X(n20260) );
  inv_x2_sg U39445 ( .A(n20178), .X(n41246) );
  nor_x1_sg U39446 ( .A(n42445), .B(n54822), .X(n20178) );
  inv_x2_sg U39447 ( .A(n20608), .X(n42692) );
  nor_x1_sg U39448 ( .A(n54921), .B(n54948), .X(n20608) );
  inv_x2_sg U39449 ( .A(n20609), .X(n41182) );
  nor_x1_sg U39450 ( .A(n20622), .B(n20623), .X(n20621) );
  nor_x1_sg U39451 ( .A(n55011), .B(n54978), .X(n20801) );
  inv_x2_sg U39452 ( .A(n20802), .X(n42412) );
  nor_x1_sg U39453 ( .A(n20803), .B(n20804), .X(n20802) );
  inv_x2_sg U39454 ( .A(n21034), .X(n41403) );
  nor_x1_sg U39455 ( .A(n21066), .B(n21067), .X(n21034) );
  inv_x2_sg U39456 ( .A(n20954), .X(n41252) );
  nor_x1_sg U39457 ( .A(n43359), .B(n55105), .X(n20954) );
  inv_x2_sg U39458 ( .A(n21379), .X(n42690) );
  nor_x1_sg U39459 ( .A(n46248), .B(n55237), .X(n21379) );
  inv_x2_sg U39460 ( .A(n21380), .X(n41513) );
  nor_x1_sg U39461 ( .A(n21417), .B(n55229), .X(n21416) );
  nor_x1_sg U39462 ( .A(n21604), .B(n21568), .X(n21605) );
  nor_x1_sg U39463 ( .A(n21573), .B(n55292), .X(n21572) );
  inv_x2_sg U39464 ( .A(n21573), .X(n55272) );
  inv_x2_sg U39465 ( .A(n21883), .X(n43525) );
  inv_x2_sg U39466 ( .A(n21805), .X(n41401) );
  nor_x1_sg U39467 ( .A(n21837), .B(n21838), .X(n21805) );
  inv_x2_sg U39468 ( .A(n21723), .X(n41244) );
  nor_x1_sg U39469 ( .A(n42443), .B(n55390), .X(n21723) );
  inv_x2_sg U39470 ( .A(n28382), .X(n43160) );
  nor_x1_sg U39471 ( .A(n28384), .B(n28385), .X(n28382) );
  inv_x2_sg U39472 ( .A(n50883), .X(n41887) );
  inv_x1_sg U39473 ( .A(n22583), .X(n50883) );
  inv_x2_sg U39474 ( .A(n22791), .X(n41930) );
  nor_x1_sg U39475 ( .A(n22839), .B(n50880), .X(n22791) );
  inv_x2_sg U39476 ( .A(n50635), .X(n41202) );
  inv_x1_sg U39477 ( .A(n23655), .X(n50635) );
  inv_x2_sg U39478 ( .A(n23832), .X(n41932) );
  nor_x1_sg U39479 ( .A(n23833), .B(n50637), .X(n23832) );
  inv_x2_sg U39480 ( .A(n23772), .X(n41957) );
  nor_x1_sg U39481 ( .A(n23773), .B(n50170), .X(n23772) );
  inv_x2_sg U39482 ( .A(n10700), .X(n42404) );
  inv_x2_sg U39483 ( .A(n10892), .X(n41583) );
  nor_x1_sg U39484 ( .A(n10910), .B(n10911), .X(n10892) );
  inv_x2_sg U39485 ( .A(n10864), .X(n43094) );
  nor_x1_sg U39486 ( .A(n51504), .B(n10877), .X(n10864) );
  inv_x2_sg U39487 ( .A(n11298), .X(n41809) );
  inv_x2_sg U39488 ( .A(n11310), .X(n41509) );
  nor_x1_sg U39489 ( .A(n41512), .B(n11342), .X(n11310) );
  inv_x2_sg U39490 ( .A(n51627), .X(n42191) );
  inv_x1_sg U39491 ( .A(n11340), .X(n51627) );
  inv_x2_sg U39492 ( .A(n11480), .X(n43439) );
  inv_x2_sg U39493 ( .A(n11644), .X(n43092) );
  nor_x1_sg U39494 ( .A(n51784), .B(n11657), .X(n11644) );
  inv_x2_sg U39495 ( .A(n12078), .X(n41807) );
  inv_x2_sg U39496 ( .A(n12090), .X(n41505) );
  nor_x1_sg U39497 ( .A(n41508), .B(n12122), .X(n12090) );
  inv_x2_sg U39498 ( .A(n51907), .X(n42189) );
  inv_x1_sg U39499 ( .A(n12120), .X(n51907) );
  inv_x2_sg U39500 ( .A(n12260), .X(n42400) );
  inv_x2_sg U39501 ( .A(n12424), .X(n41698) );
  nor_x1_sg U39502 ( .A(n12437), .B(n41701), .X(n12424) );
  inv_x2_sg U39503 ( .A(n12859), .X(n41551) );
  inv_x2_sg U39504 ( .A(n12871), .X(n41228) );
  nor_x1_sg U39505 ( .A(n41231), .B(n12903), .X(n12871) );
  inv_x2_sg U39506 ( .A(n12872), .X(n42812) );
  nor_x1_sg U39507 ( .A(n12909), .B(n12910), .X(n12872) );
  inv_x2_sg U39508 ( .A(n52184), .X(n41708) );
  inv_x1_sg U39509 ( .A(n12901), .X(n52184) );
  inv_x2_sg U39510 ( .A(n13041), .X(n43435) );
  inv_x2_sg U39511 ( .A(n13205), .X(n41694) );
  nor_x1_sg U39512 ( .A(n13218), .B(n41697), .X(n13205) );
  nand_x4_sg U39513 ( .A(n52406), .B(n46474), .X(n13607) );
  inv_x2_sg U39514 ( .A(n13639), .X(n41805) );
  inv_x2_sg U39515 ( .A(n13610), .X(n41733) );
  nor_x1_sg U39516 ( .A(n13619), .B(n13620), .X(n13610) );
  inv_x2_sg U39517 ( .A(n13651), .X(n41501) );
  nor_x1_sg U39518 ( .A(n41504), .B(n13683), .X(n13651) );
  inv_x2_sg U39519 ( .A(n13652), .X(n42810) );
  nor_x1_sg U39520 ( .A(n13689), .B(n13690), .X(n13652) );
  inv_x2_sg U39521 ( .A(n52460), .X(n41706) );
  inv_x1_sg U39522 ( .A(n13681), .X(n52460) );
  inv_x2_sg U39523 ( .A(n13821), .X(n43431) );
  inv_x2_sg U39524 ( .A(n13985), .X(n41690) );
  nor_x1_sg U39525 ( .A(n13998), .B(n41693), .X(n13985) );
  inv_x2_sg U39526 ( .A(n14591), .X(n42422) );
  inv_x2_sg U39527 ( .A(n14756), .X(n43080) );
  nor_x1_sg U39528 ( .A(n14769), .B(n52894), .X(n14756) );
  inv_x2_sg U39529 ( .A(n15192), .X(n41549) );
  inv_x2_sg U39530 ( .A(n15204), .X(n41224) );
  nor_x1_sg U39531 ( .A(n41227), .B(n15236), .X(n15204) );
  inv_x2_sg U39532 ( .A(n15205), .X(n42808) );
  nor_x1_sg U39533 ( .A(n15242), .B(n15243), .X(n15205) );
  inv_x2_sg U39534 ( .A(n53018), .X(n41704) );
  inv_x1_sg U39535 ( .A(n15234), .X(n53018) );
  inv_x2_sg U39536 ( .A(n15374), .X(n43427) );
  inv_x2_sg U39537 ( .A(n15538), .X(n41686) );
  nor_x1_sg U39538 ( .A(n15551), .B(n41689), .X(n15538) );
  inv_x2_sg U39539 ( .A(n15973), .X(n41803) );
  inv_x2_sg U39540 ( .A(n15985), .X(n41497) );
  nor_x1_sg U39541 ( .A(n41500), .B(n16017), .X(n15985) );
  inv_x2_sg U39542 ( .A(n53294), .X(n42187) );
  inv_x1_sg U39543 ( .A(n16015), .X(n53294) );
  inv_x2_sg U39544 ( .A(n16155), .X(n42394) );
  inv_x2_sg U39545 ( .A(n16347), .X(n41581) );
  nor_x1_sg U39546 ( .A(n16369), .B(n16370), .X(n16347) );
  inv_x2_sg U39547 ( .A(n16319), .X(n42063) );
  nor_x1_sg U39548 ( .A(n42066), .B(n16333), .X(n16319) );
  inv_x2_sg U39549 ( .A(n16758), .X(n41547) );
  inv_x2_sg U39550 ( .A(n16770), .X(n41220) );
  nor_x1_sg U39551 ( .A(n41223), .B(n16802), .X(n16770) );
  inv_x2_sg U39552 ( .A(n16771), .X(n42806) );
  nor_x1_sg U39553 ( .A(n16808), .B(n16809), .X(n16771) );
  inv_x2_sg U39554 ( .A(n53576), .X(n41702) );
  inv_x1_sg U39555 ( .A(n16800), .X(n53576) );
  inv_x2_sg U39556 ( .A(n16940), .X(n43423) );
  inv_x2_sg U39557 ( .A(n17104), .X(n41682) );
  nor_x1_sg U39558 ( .A(n17117), .B(n41685), .X(n17104) );
  inv_x2_sg U39559 ( .A(n17532), .X(n43254) );
  inv_x2_sg U39560 ( .A(n17712), .X(n42418) );
  inv_x2_sg U39561 ( .A(n17877), .X(n43072) );
  nor_x1_sg U39562 ( .A(n17890), .B(n54014), .X(n17877) );
  inv_x2_sg U39563 ( .A(n18644), .X(n43070) );
  nor_x1_sg U39564 ( .A(n18659), .B(n54296), .X(n18644) );
  inv_x2_sg U39565 ( .A(n19077), .X(n43252) );
  inv_x2_sg U39566 ( .A(n19257), .X(n42414) );
  inv_x2_sg U39567 ( .A(n19422), .X(n43064) );
  nor_x1_sg U39568 ( .A(n19435), .B(n54579), .X(n19422) );
  inv_x2_sg U39569 ( .A(n19871), .X(n41519) );
  inv_x2_sg U39570 ( .A(n20060), .X(n42462) );
  inv_x2_sg U39571 ( .A(n20027), .X(n42408) );
  inv_x2_sg U39572 ( .A(n20190), .X(n43062) );
  nor_x1_sg U39573 ( .A(n20204), .B(n54864), .X(n20190) );
  inv_x2_sg U39574 ( .A(n20621), .X(n43250) );
  inv_x2_sg U39575 ( .A(n20801), .X(n42410) );
  inv_x2_sg U39576 ( .A(n20966), .X(n43056) );
  nor_x1_sg U39577 ( .A(n20979), .B(n55147), .X(n20966) );
  inv_x2_sg U39578 ( .A(n21416), .X(n41515) );
  inv_x2_sg U39579 ( .A(n21605), .X(n42460) );
  inv_x2_sg U39580 ( .A(n21572), .X(n42406) );
  inv_x2_sg U39581 ( .A(n21735), .X(n43054) );
  nor_x1_sg U39582 ( .A(n21749), .B(n55432), .X(n21735) );
  inv_x2_sg U39583 ( .A(n50024), .X(n41885) );
  inv_x1_sg U39584 ( .A(n30249), .X(n50024) );
  inv_x2_sg U39585 ( .A(n30457), .X(n41928) );
  nor_x1_sg U39586 ( .A(n30505), .B(n50021), .X(n30457) );
  inv_x2_sg U39587 ( .A(n49875), .X(n41210) );
  inv_x1_sg U39588 ( .A(n30966), .X(n49875) );
  inv_x2_sg U39589 ( .A(n49784), .X(n41208) );
  inv_x1_sg U39590 ( .A(n31361), .X(n49784) );
  inv_x2_sg U39591 ( .A(n49776), .X(n41150) );
  inv_x1_sg U39592 ( .A(n31321), .X(n49776) );
  inv_x2_sg U39593 ( .A(n31498), .X(n41922) );
  nor_x1_sg U39594 ( .A(n31499), .B(n49778), .X(n31498) );
  inv_x2_sg U39595 ( .A(n49692), .X(n41206) );
  inv_x1_sg U39596 ( .A(n31685), .X(n49692) );
  inv_x2_sg U39597 ( .A(n49642), .X(n41204) );
  inv_x1_sg U39598 ( .A(n31945), .X(n49642) );
  inv_x2_sg U39599 ( .A(n49596), .X(n41159) );
  inv_x1_sg U39600 ( .A(n32028), .X(n49596) );
  inv_x2_sg U39601 ( .A(n31438), .X(n41955) );
  nor_x1_sg U39602 ( .A(n31439), .B(n49311), .X(n31438) );
  inv_x2_sg U39603 ( .A(n26686), .X(n42147) );
  nor_x1_sg U39604 ( .A(n42150), .B(n52417), .X(n26686) );
  inv_x2_sg U39605 ( .A(n28388), .X(n41232) );
  nor_x1_sg U39606 ( .A(n41235), .B(n28391), .X(n28388) );
  inv_x2_sg U39607 ( .A(n21979), .X(n41485) );
  inv_x2_sg U39608 ( .A(n21941), .X(n41180) );
  inv_x2_sg U39609 ( .A(n22512), .X(n42760) );
  nor_x1_sg U39610 ( .A(n22585), .B(n50928), .X(n22512) );
  inv_x2_sg U39611 ( .A(n21936), .X(n41349) );
  inv_x2_sg U39612 ( .A(n21958), .X(n41144) );
  inv_x2_sg U39613 ( .A(n22500), .X(n42758) );
  nor_x1_sg U39614 ( .A(n22613), .B(n50950), .X(n22500) );
  inv_x2_sg U39615 ( .A(n21952), .X(n41487) );
  inv_x2_sg U39616 ( .A(n23058), .X(n42225) );
  nor_x1_sg U39617 ( .A(n23068), .B(n23069), .X(n23058) );
  inv_x2_sg U39618 ( .A(n23284), .X(n42223) );
  nor_x1_sg U39619 ( .A(n23294), .B(n23295), .X(n23284) );
  inv_x2_sg U39620 ( .A(n23489), .X(n42219) );
  nor_x1_sg U39621 ( .A(n23499), .B(n42222), .X(n23489) );
  inv_x2_sg U39622 ( .A(n23679), .X(n42217) );
  nor_x1_sg U39623 ( .A(n23689), .B(n23690), .X(n23679) );
  inv_x2_sg U39624 ( .A(n23850), .X(n42213) );
  nor_x1_sg U39625 ( .A(n23860), .B(n42216), .X(n23850) );
  inv_x2_sg U39626 ( .A(n24003), .X(n42211) );
  nor_x1_sg U39627 ( .A(n24013), .B(n24014), .X(n24003) );
  inv_x2_sg U39628 ( .A(n23453), .X(n42195) );
  nor_x1_sg U39629 ( .A(n23454), .B(n50633), .X(n23453) );
  inv_x2_sg U39630 ( .A(n22470), .X(n42229) );
  nor_x1_sg U39631 ( .A(n22471), .B(n50624), .X(n22470) );
  inv_x2_sg U39632 ( .A(n24147), .X(n42207) );
  nor_x1_sg U39633 ( .A(n24157), .B(n42210), .X(n24147) );
  inv_x2_sg U39634 ( .A(n24263), .X(n42205) );
  nor_x1_sg U39635 ( .A(n24273), .B(n24274), .X(n24263) );
  inv_x2_sg U39636 ( .A(n24365), .X(n42201) );
  nor_x1_sg U39637 ( .A(n24375), .B(n42204), .X(n24365) );
  inv_x2_sg U39638 ( .A(n24359), .X(n42197) );
  nor_x1_sg U39639 ( .A(n24360), .B(n42200), .X(n24359) );
  inv_x2_sg U39640 ( .A(n24427), .X(n41926) );
  nor_x1_sg U39641 ( .A(n24430), .B(n24431), .X(n24427) );
  inv_x2_sg U39642 ( .A(n24416), .X(n41242) );
  nor_x1_sg U39643 ( .A(n24418), .B(n24419), .X(n24416) );
  inv_x2_sg U39644 ( .A(n10540), .X(n43220) );
  nor_x1_sg U39645 ( .A(n51315), .B(n10542), .X(n10540) );
  inv_x2_sg U39646 ( .A(n10541), .X(n41787) );
  nor_x1_sg U39647 ( .A(n10549), .B(n51361), .X(n10541) );
  inv_x2_sg U39648 ( .A(n11668), .X(n43004) );
  nor_x1_sg U39649 ( .A(n43007), .B(n51794), .X(n11668) );
  inv_x2_sg U39650 ( .A(n11951), .X(n41601) );
  nand_x1_sg U39651 ( .A(n51827), .B(n41346), .X(n11951) );
  nand_x4_sg U39652 ( .A(n46517), .B(n51854), .X(n12046) );
  inv_x2_sg U39653 ( .A(n12382), .X(n43166) );
  nor_x1_sg U39654 ( .A(n52049), .B(n43169), .X(n12382) );
  inv_x2_sg U39655 ( .A(n12448), .X(n43000) );
  nor_x1_sg U39656 ( .A(n43003), .B(n52066), .X(n12448) );
  nand_x4_sg U39657 ( .A(n52133), .B(n46496), .X(n12828) );
  inv_x2_sg U39658 ( .A(n13229), .X(n42996) );
  nor_x1_sg U39659 ( .A(n42999), .B(n52343), .X(n13229) );
  inv_x2_sg U39660 ( .A(n13162), .X(n41724) );
  nor_x1_sg U39661 ( .A(n52326), .B(n41727), .X(n13162) );
  nand_x2_sg U39662 ( .A(n26726), .B(n26727), .X(n26724) );
  inv_x2_sg U39663 ( .A(n13513), .X(n41599) );
  nand_x1_sg U39664 ( .A(n52379), .B(n41344), .X(n13513) );
  inv_x2_sg U39665 ( .A(n14009), .X(n42992) );
  nor_x1_sg U39666 ( .A(n42995), .B(n52618), .X(n14009) );
  inv_x2_sg U39667 ( .A(n13942), .X(n41720) );
  nor_x1_sg U39668 ( .A(n52601), .B(n41723), .X(n13942) );
  inv_x2_sg U39669 ( .A(n52645), .X(n42834) );
  inv_x1_sg U39670 ( .A(n26996), .X(n52645) );
  inv_x2_sg U39671 ( .A(n14455), .X(n42145) );
  nor_x1_sg U39672 ( .A(n14494), .B(n14495), .X(n14455) );
  inv_x2_sg U39673 ( .A(n14433), .X(n42364) );
  nor_x1_sg U39674 ( .A(n14400), .B(n14435), .X(n14433) );
  inv_x2_sg U39675 ( .A(n14434), .X(n41801) );
  nor_x1_sg U39676 ( .A(n14441), .B(n14442), .X(n14434) );
  inv_x2_sg U39677 ( .A(n14780), .X(n42988) );
  nor_x1_sg U39678 ( .A(n42991), .B(n52904), .X(n14780) );
  nand_x4_sg U39679 ( .A(n52967), .B(n46428), .X(n15161) );
  inv_x2_sg U39680 ( .A(n15562), .X(n42984) );
  nor_x1_sg U39681 ( .A(n42987), .B(n53177), .X(n15562) );
  inv_x2_sg U39682 ( .A(n15495), .X(n41716) );
  nor_x1_sg U39683 ( .A(n53160), .B(n41719), .X(n15495) );
  inv_x2_sg U39684 ( .A(n53204), .X(n42826) );
  inv_x1_sg U39685 ( .A(n27555), .X(n53204) );
  inv_x2_sg U39686 ( .A(n15846), .X(n41595) );
  nand_x1_sg U39687 ( .A(n53215), .B(n41342), .X(n15846) );
  inv_x1_sg U39688 ( .A(n15870), .X(n44153) );
  nand_x4_sg U39689 ( .A(n53525), .B(n46384), .X(n16727) );
  inv_x2_sg U39690 ( .A(n17128), .X(n42976) );
  nor_x1_sg U39691 ( .A(n42979), .B(n53735), .X(n17128) );
  inv_x2_sg U39692 ( .A(n17061), .X(n41712) );
  nor_x1_sg U39693 ( .A(n53718), .B(n41715), .X(n17061) );
  inv_x2_sg U39694 ( .A(n17575), .X(n42143) );
  nor_x1_sg U39695 ( .A(n17615), .B(n17616), .X(n17575) );
  inv_x2_sg U39696 ( .A(n17552), .X(n42362) );
  nor_x1_sg U39697 ( .A(n53815), .B(n17554), .X(n17552) );
  inv_x2_sg U39698 ( .A(n17553), .X(n41799) );
  nor_x1_sg U39699 ( .A(n17561), .B(n17562), .X(n17553) );
  inv_x2_sg U39700 ( .A(n17901), .X(n42972) );
  nor_x1_sg U39701 ( .A(n42975), .B(n54024), .X(n17901) );
  inv_x2_sg U39702 ( .A(n18236), .X(n43513) );
  inv_x2_sg U39703 ( .A(n18345), .X(n42137) );
  nor_x1_sg U39704 ( .A(n18384), .B(n18385), .X(n18345) );
  inv_x2_sg U39705 ( .A(n18323), .X(n43222) );
  nor_x1_sg U39706 ( .A(n18291), .B(n18325), .X(n18323) );
  inv_x2_sg U39707 ( .A(n18324), .X(n41793) );
  nor_x1_sg U39708 ( .A(n18331), .B(n54150), .X(n18324) );
  inv_x2_sg U39709 ( .A(n18670), .X(n42968) );
  nor_x1_sg U39710 ( .A(n42971), .B(n54305), .X(n18670) );
  inv_x2_sg U39711 ( .A(n19120), .X(n42141) );
  nor_x1_sg U39712 ( .A(n19160), .B(n19161), .X(n19120) );
  inv_x2_sg U39713 ( .A(n19097), .X(n42360) );
  nor_x1_sg U39714 ( .A(n54380), .B(n19099), .X(n19097) );
  inv_x2_sg U39715 ( .A(n19098), .X(n41797) );
  nor_x1_sg U39716 ( .A(n19106), .B(n19107), .X(n19098) );
  inv_x2_sg U39717 ( .A(n19446), .X(n42964) );
  nor_x1_sg U39718 ( .A(n42967), .B(n54589), .X(n19446) );
  inv_x2_sg U39719 ( .A(n19728), .X(n41597) );
  nand_x1_sg U39720 ( .A(n19729), .B(n41177), .X(n19728) );
  inv_x2_sg U39721 ( .A(n19782), .X(n42285) );
  nor_x1_sg U39722 ( .A(n54631), .B(n19769), .X(n19782) );
  inv_x2_sg U39723 ( .A(n19867), .X(n42356) );
  nor_x1_sg U39724 ( .A(n54669), .B(n19869), .X(n19867) );
  inv_x2_sg U39725 ( .A(n19868), .X(n41791) );
  nor_x1_sg U39726 ( .A(n19876), .B(n54715), .X(n19868) );
  inv_x2_sg U39727 ( .A(n20215), .X(n42960) );
  nor_x1_sg U39728 ( .A(n42963), .B(n54873), .X(n20215) );
  inv_x2_sg U39729 ( .A(n20664), .X(n42139) );
  nor_x1_sg U39730 ( .A(n20704), .B(n20705), .X(n20664) );
  inv_x2_sg U39731 ( .A(n20641), .X(n42358) );
  nor_x1_sg U39732 ( .A(n54948), .B(n20643), .X(n20641) );
  inv_x2_sg U39733 ( .A(n20642), .X(n41795) );
  nor_x1_sg U39734 ( .A(n20650), .B(n20651), .X(n20642) );
  inv_x2_sg U39735 ( .A(n20990), .X(n42956) );
  nor_x1_sg U39736 ( .A(n42959), .B(n55157), .X(n20990) );
  inv_x2_sg U39737 ( .A(n21327), .X(n42283) );
  nor_x1_sg U39738 ( .A(n55199), .B(n21314), .X(n21327) );
  inv_x2_sg U39739 ( .A(n21412), .X(n42354) );
  nor_x1_sg U39740 ( .A(n55237), .B(n21414), .X(n21412) );
  inv_x2_sg U39741 ( .A(n21413), .X(n41789) );
  nor_x1_sg U39742 ( .A(n21421), .B(n55283), .X(n21413) );
  inv_x2_sg U39743 ( .A(n21760), .X(n42952) );
  nor_x1_sg U39744 ( .A(n42955), .B(n55441), .X(n21760) );
  inv_x2_sg U39745 ( .A(n29644), .X(n41481) );
  inv_x2_sg U39746 ( .A(n29594), .X(n41178) );
  inv_x2_sg U39747 ( .A(n30178), .X(n42688) );
  nor_x1_sg U39748 ( .A(n30251), .B(n50069), .X(n30178) );
  inv_x2_sg U39749 ( .A(n29586), .X(n41347) );
  inv_x2_sg U39750 ( .A(n29615), .X(n41142) );
  inv_x2_sg U39751 ( .A(n30166), .X(n42686) );
  nor_x1_sg U39752 ( .A(n30279), .B(n50091), .X(n30166) );
  inv_x2_sg U39753 ( .A(n29608), .X(n41483) );
  inv_x2_sg U39754 ( .A(n31119), .X(n42193) );
  nor_x1_sg U39755 ( .A(n31120), .B(n49774), .X(n31119) );
  inv_x2_sg U39756 ( .A(n30135), .X(n42227) );
  nor_x1_sg U39757 ( .A(n30136), .B(n49765), .X(n30135) );
  inv_x2_sg U39758 ( .A(n32093), .X(n41934) );
  nor_x1_sg U39759 ( .A(n32096), .B(n32097), .X(n32093) );
  inv_x2_sg U39760 ( .A(n32082), .X(n41240) );
  nor_x1_sg U39761 ( .A(n32084), .B(n32085), .X(n32082) );
  inv_x2_sg U39762 ( .A(n26965), .X(n43162) );
  nor_x1_sg U39763 ( .A(n43165), .B(n52693), .X(n26965) );
  inv_x1_sg U39764 ( .A(n46059), .X(n42846) );
  inv_x1_sg U39765 ( .A(n46057), .X(n42844) );
  inv_x1_sg U39766 ( .A(n46061), .X(n42842) );
  nor_x1_sg U39767 ( .A(n21964), .B(n22523), .X(n22522) );
  nor_x1_sg U39768 ( .A(n21948), .B(n21976), .X(n21975) );
  nor_x1_sg U39769 ( .A(n21955), .B(n22505), .X(n22504) );
  inv_x2_sg U39770 ( .A(n22787), .X(n43012) );
  nor_x1_sg U39771 ( .A(n43015), .B(n22846), .X(n22787) );
  nor_x1_sg U39772 ( .A(n50909), .B(n22538), .X(n22804) );
  inv_x2_sg U39773 ( .A(n22584), .X(n43186) );
  nor_x1_sg U39774 ( .A(n43189), .B(n50924), .X(n22584) );
  inv_x2_sg U39775 ( .A(n23042), .X(n43028) );
  nor_x1_sg U39776 ( .A(n23100), .B(n23101), .X(n23042) );
  inv_x2_sg U39777 ( .A(n23473), .X(n43026) );
  nor_x1_sg U39778 ( .A(n23531), .B(n23532), .X(n23473) );
  inv_x2_sg U39779 ( .A(n23657), .X(n41680) );
  nor_x1_sg U39780 ( .A(n23659), .B(n23660), .X(n23657) );
  inv_x2_sg U39781 ( .A(n23651), .X(n41676) );
  nor_x1_sg U39782 ( .A(n41679), .B(n23654), .X(n23651) );
  inv_x2_sg U39783 ( .A(n23729), .X(n43190) );
  nor_x1_sg U39784 ( .A(n43193), .B(n50654), .X(n23729) );
  inv_x2_sg U39785 ( .A(n23645), .X(n41619) );
  nor_x1_sg U39786 ( .A(n23647), .B(n23648), .X(n23645) );
  inv_x2_sg U39787 ( .A(n23639), .X(n41446) );
  nor_x1_sg U39788 ( .A(n23641), .B(n23642), .X(n23639) );
  inv_x2_sg U39789 ( .A(n23633), .X(n43021) );
  nor_x1_sg U39790 ( .A(n23635), .B(n43024), .X(n23633) );
  inv_x2_sg U39791 ( .A(n23627), .X(n41444) );
  nor_x1_sg U39792 ( .A(n23629), .B(n23630), .X(n23627) );
  inv_x2_sg U39793 ( .A(n23621), .X(n41442) );
  nor_x1_sg U39794 ( .A(n23623), .B(n23624), .X(n23621) );
  inv_x2_sg U39795 ( .A(n23615), .X(n43016) );
  nor_x1_sg U39796 ( .A(n23617), .B(n43019), .X(n23615) );
  inv_x2_sg U39797 ( .A(n23609), .X(n41440) );
  nor_x1_sg U39798 ( .A(n23611), .B(n23612), .X(n23609) );
  inv_x2_sg U39799 ( .A(n23603), .X(n41672) );
  nor_x1_sg U39800 ( .A(n23605), .B(n41675), .X(n23603) );
  inv_x2_sg U39801 ( .A(n51258), .X(n42828) );
  inv_x1_sg U39802 ( .A(n25599), .X(n51258) );
  nor_x1_sg U39803 ( .A(n10442), .B(n10443), .X(n10441) );
  inv_x2_sg U39804 ( .A(n10446), .X(n42852) );
  nor_x1_sg U39805 ( .A(n51298), .B(n10453), .X(n10446) );
  inv_x2_sg U39806 ( .A(n10591), .X(n41874) );
  nand_x1_sg U39807 ( .A(n41649), .B(n10600), .X(n10591) );
  inv_x2_sg U39808 ( .A(n10820), .X(n42850) );
  nor_x1_sg U39809 ( .A(n10881), .B(n10882), .X(n10820) );
  inv_x2_sg U39810 ( .A(n10887), .X(n43008) );
  nor_x1_sg U39811 ( .A(n43011), .B(n51519), .X(n10887) );
  inv_x2_sg U39812 ( .A(n51511), .X(n41399) );
  inv_x1_sg U39813 ( .A(n10358), .X(n51511) );
  inv_x2_sg U39814 ( .A(n51534), .X(n42822) );
  inv_x1_sg U39815 ( .A(n25880), .X(n51534) );
  nor_x1_sg U39816 ( .A(n11246), .B(n51605), .X(n11245) );
  inv_x2_sg U39817 ( .A(n11244), .X(n43414) );
  nor_x1_sg U39818 ( .A(n11247), .B(n51623), .X(n11244) );
  inv_x2_sg U39819 ( .A(n51791), .X(n41397) );
  inv_x1_sg U39820 ( .A(n11125), .X(n51791) );
  inv_x2_sg U39821 ( .A(n51816), .X(n42824) );
  inv_x1_sg U39822 ( .A(n26160), .X(n51816) );
  nor_x1_sg U39823 ( .A(n51848), .B(n51834), .X(n11993) );
  nor_x1_sg U39824 ( .A(n12022), .B(n51886), .X(n12021) );
  inv_x2_sg U39825 ( .A(n12020), .X(n43410) );
  nor_x1_sg U39826 ( .A(n12023), .B(n51905), .X(n12020) );
  inv_x2_sg U39827 ( .A(n52069), .X(n41395) );
  inv_x1_sg U39828 ( .A(n11908), .X(n52069) );
  inv_x2_sg U39829 ( .A(n52092), .X(n42820) );
  inv_x1_sg U39830 ( .A(n26439), .X(n52092) );
  nor_x1_sg U39831 ( .A(n12807), .B(n52163), .X(n12806) );
  inv_x2_sg U39832 ( .A(n12805), .X(n43406) );
  nor_x1_sg U39833 ( .A(n12808), .B(n52182), .X(n12805) );
  inv_x2_sg U39834 ( .A(n52347), .X(n41393) );
  inv_x1_sg U39835 ( .A(n12686), .X(n52347) );
  inv_x2_sg U39836 ( .A(n52369), .X(n42804) );
  inv_x1_sg U39837 ( .A(n26717), .X(n52369) );
  nor_x1_sg U39838 ( .A(n52400), .B(n52386), .X(n13554) );
  nor_x1_sg U39839 ( .A(n13583), .B(n52437), .X(n13582) );
  inv_x2_sg U39840 ( .A(n13581), .X(n43402) );
  nor_x1_sg U39841 ( .A(n13584), .B(n52458), .X(n13581) );
  inv_x2_sg U39842 ( .A(n13616), .X(n42448) );
  nor_x1_sg U39843 ( .A(n13614), .B(n13613), .X(n13616) );
  inv_x2_sg U39844 ( .A(n52622), .X(n41389) );
  inv_x1_sg U39845 ( .A(n13470), .X(n52622) );
  nor_x1_sg U39846 ( .A(n52666), .B(n52678), .X(n14332) );
  inv_x2_sg U39847 ( .A(n14333), .X(n43509) );
  nor_x1_sg U39848 ( .A(n14334), .B(n14335), .X(n14333) );
  inv_x2_sg U39849 ( .A(n14338), .X(n42854) );
  nor_x1_sg U39850 ( .A(n52688), .B(n14348), .X(n14338) );
  inv_x2_sg U39851 ( .A(n52901), .X(n41387) );
  inv_x1_sg U39852 ( .A(n14249), .X(n52901) );
  inv_x2_sg U39853 ( .A(n52926), .X(n42818) );
  inv_x1_sg U39854 ( .A(n27276), .X(n52926) );
  nor_x1_sg U39855 ( .A(n15140), .B(n52997), .X(n15139) );
  inv_x2_sg U39856 ( .A(n15138), .X(n43394) );
  nor_x1_sg U39857 ( .A(n15141), .B(n53016), .X(n15138) );
  inv_x2_sg U39858 ( .A(n53181), .X(n41385) );
  inv_x1_sg U39859 ( .A(n15019), .X(n53181) );
  nor_x1_sg U39860 ( .A(n53234), .B(n53222), .X(n15888) );
  nor_x1_sg U39861 ( .A(n15917), .B(n53273), .X(n15916) );
  inv_x2_sg U39862 ( .A(n15915), .X(n43390) );
  nor_x1_sg U39863 ( .A(n15918), .B(n53290), .X(n15915) );
  inv_x2_sg U39864 ( .A(n16276), .X(n42848) );
  nor_x1_sg U39865 ( .A(n16336), .B(n16337), .X(n16276) );
  inv_x2_sg U39866 ( .A(n16342), .X(n42980) );
  nor_x1_sg U39867 ( .A(n42983), .B(n53468), .X(n16342) );
  inv_x2_sg U39868 ( .A(n53461), .X(n41381) );
  inv_x1_sg U39869 ( .A(n15804), .X(n53461) );
  inv_x2_sg U39870 ( .A(n53484), .X(n42816) );
  inv_x1_sg U39871 ( .A(n27834), .X(n53484) );
  nor_x1_sg U39872 ( .A(n16706), .B(n53555), .X(n16705) );
  inv_x2_sg U39873 ( .A(n16704), .X(n43386) );
  nor_x1_sg U39874 ( .A(n16707), .B(n53574), .X(n16704) );
  inv_x2_sg U39875 ( .A(n53739), .X(n41379) );
  inv_x1_sg U39876 ( .A(n16585), .X(n53739) );
  inv_x2_sg U39877 ( .A(n53762), .X(n42840) );
  inv_x1_sg U39878 ( .A(n28115), .X(n53762) );
  nor_x1_sg U39879 ( .A(n53782), .B(n53797), .X(n17455) );
  inv_x2_sg U39880 ( .A(n17456), .X(n43505) );
  nor_x1_sg U39881 ( .A(n17457), .B(n17458), .X(n17456) );
  inv_x2_sg U39882 ( .A(n54021), .X(n41375) );
  inv_x1_sg U39883 ( .A(n17368), .X(n54021) );
  nor_x1_sg U39884 ( .A(n54063), .B(n54078), .X(n18221) );
  inv_x2_sg U39885 ( .A(n18222), .X(n42472) );
  nor_x1_sg U39886 ( .A(n18223), .B(n18224), .X(n18222) );
  inv_x2_sg U39887 ( .A(n18227), .X(n43138) );
  nor_x1_sg U39888 ( .A(n54089), .B(n18234), .X(n18227) );
  inv_x2_sg U39889 ( .A(n54302), .X(n41190) );
  inv_x1_sg U39890 ( .A(n18140), .X(n54302) );
  inv_x2_sg U39891 ( .A(n54327), .X(n42838) );
  inv_x1_sg U39892 ( .A(n28673), .X(n54327) );
  nor_x1_sg U39893 ( .A(n54347), .B(n54362), .X(n19000) );
  inv_x2_sg U39894 ( .A(n19001), .X(n43501) );
  nor_x1_sg U39895 ( .A(n19002), .B(n19003), .X(n19001) );
  inv_x2_sg U39896 ( .A(n54586), .X(n41373) );
  inv_x1_sg U39897 ( .A(n18913), .X(n54586) );
  inv_x2_sg U39898 ( .A(n54611), .X(n42832) );
  inv_x1_sg U39899 ( .A(n28951), .X(n54611) );
  nor_x1_sg U39900 ( .A(n54631), .B(n54642), .X(n19767) );
  inv_x2_sg U39901 ( .A(n19768), .X(n43491) );
  nor_x1_sg U39902 ( .A(n19769), .B(n19770), .X(n19768) );
  inv_x2_sg U39903 ( .A(n19773), .X(n43134) );
  nor_x1_sg U39904 ( .A(n54652), .B(n43137), .X(n19773) );
  inv_x2_sg U39905 ( .A(n19918), .X(n41878) );
  nand_x1_sg U39906 ( .A(n41651), .B(n19927), .X(n19918) );
  inv_x2_sg U39907 ( .A(n54870), .X(n41371) );
  inv_x1_sg U39908 ( .A(n19685), .X(n54870) );
  inv_x2_sg U39909 ( .A(n54895), .X(n42836) );
  inv_x1_sg U39910 ( .A(n29234), .X(n54895) );
  nor_x1_sg U39911 ( .A(n54915), .B(n54930), .X(n20544) );
  inv_x2_sg U39912 ( .A(n20545), .X(n43497) );
  nor_x1_sg U39913 ( .A(n20546), .B(n20547), .X(n20545) );
  inv_x2_sg U39914 ( .A(n55154), .X(n41369) );
  inv_x1_sg U39915 ( .A(n20457), .X(n55154) );
  inv_x2_sg U39916 ( .A(n55179), .X(n42830) );
  inv_x1_sg U39917 ( .A(n29512), .X(n55179) );
  nor_x1_sg U39918 ( .A(n55199), .B(n55210), .X(n21312) );
  inv_x2_sg U39919 ( .A(n21313), .X(n43487) );
  nor_x1_sg U39920 ( .A(n21314), .B(n21315), .X(n21313) );
  inv_x2_sg U39921 ( .A(n21318), .X(n43130) );
  nor_x1_sg U39922 ( .A(n55220), .B(n43133), .X(n21318) );
  inv_x2_sg U39923 ( .A(n21463), .X(n41876) );
  nand_x1_sg U39924 ( .A(n41650), .B(n21472), .X(n21463) );
  inv_x2_sg U39925 ( .A(n55438), .X(n41367) );
  inv_x1_sg U39926 ( .A(n21230), .X(n55438) );
  nor_x1_sg U39927 ( .A(n29625), .B(n30189), .X(n30188) );
  nor_x1_sg U39928 ( .A(n29602), .B(n29641), .X(n29640) );
  nor_x1_sg U39929 ( .A(n29611), .B(n30171), .X(n30170) );
  inv_x2_sg U39930 ( .A(n30453), .X(n42948) );
  nor_x1_sg U39931 ( .A(n42951), .B(n30512), .X(n30453) );
  nor_x1_sg U39932 ( .A(n50050), .B(n30204), .X(n30470) );
  inv_x2_sg U39933 ( .A(n30250), .X(n43182) );
  nor_x1_sg U39934 ( .A(n43185), .B(n50065), .X(n30250) );
  inv_x2_sg U39935 ( .A(n30724), .X(n42253) );
  nor_x1_sg U39936 ( .A(n30734), .B(n30735), .X(n30724) );
  inv_x2_sg U39937 ( .A(n30708), .X(n42946) );
  nor_x1_sg U39938 ( .A(n30766), .B(n30767), .X(n30708) );
  inv_x2_sg U39939 ( .A(n30950), .X(n42257) );
  nor_x1_sg U39940 ( .A(n30960), .B(n30961), .X(n30950) );
  inv_x2_sg U39941 ( .A(n31155), .X(n42249) );
  nor_x1_sg U39942 ( .A(n31165), .B(n42252), .X(n31155) );
  inv_x2_sg U39943 ( .A(n31139), .X(n42944) );
  nor_x1_sg U39944 ( .A(n31197), .B(n31198), .X(n31139) );
  inv_x2_sg U39945 ( .A(n31345), .X(n42255) );
  nor_x1_sg U39946 ( .A(n31355), .B(n31356), .X(n31345) );
  inv_x2_sg U39947 ( .A(n31516), .X(n42245) );
  nor_x1_sg U39948 ( .A(n31526), .B(n42248), .X(n31516) );
  inv_x2_sg U39949 ( .A(n31323), .X(n41670) );
  nor_x1_sg U39950 ( .A(n31325), .B(n31326), .X(n31323) );
  inv_x2_sg U39951 ( .A(n31669), .X(n42279) );
  nor_x1_sg U39952 ( .A(n31679), .B(n31680), .X(n31669) );
  inv_x2_sg U39953 ( .A(n31317), .X(n41666) );
  nor_x1_sg U39954 ( .A(n41669), .B(n31320), .X(n31317) );
  inv_x2_sg U39955 ( .A(n31395), .X(n43178) );
  nor_x1_sg U39956 ( .A(n43181), .B(n49795), .X(n31395) );
  inv_x2_sg U39957 ( .A(n31813), .X(n42241) );
  nor_x1_sg U39958 ( .A(n31823), .B(n42244), .X(n31813) );
  inv_x2_sg U39959 ( .A(n31311), .X(n41617) );
  nor_x1_sg U39960 ( .A(n31313), .B(n31314), .X(n31311) );
  inv_x2_sg U39961 ( .A(n31929), .X(n42239) );
  nor_x1_sg U39962 ( .A(n31939), .B(n31940), .X(n31929) );
  inv_x2_sg U39963 ( .A(n31305), .X(n41438) );
  nor_x1_sg U39964 ( .A(n31307), .B(n31308), .X(n31305) );
  inv_x2_sg U39965 ( .A(n32031), .X(n42235) );
  nor_x1_sg U39966 ( .A(n32041), .B(n42238), .X(n32031) );
  inv_x2_sg U39967 ( .A(n31299), .X(n42939) );
  nor_x1_sg U39968 ( .A(n31301), .B(n42942), .X(n31299) );
  inv_x2_sg U39969 ( .A(n32025), .X(n42231) );
  nor_x1_sg U39970 ( .A(n32026), .B(n42234), .X(n32025) );
  inv_x2_sg U39971 ( .A(n31293), .X(n41436) );
  nor_x1_sg U39972 ( .A(n31295), .B(n31296), .X(n31293) );
  inv_x2_sg U39973 ( .A(n31287), .X(n41434) );
  nor_x1_sg U39974 ( .A(n31289), .B(n31290), .X(n31287) );
  inv_x2_sg U39975 ( .A(n31281), .X(n42934) );
  nor_x1_sg U39976 ( .A(n31283), .B(n42937), .X(n31281) );
  inv_x2_sg U39977 ( .A(n31275), .X(n41432) );
  nor_x1_sg U39978 ( .A(n31277), .B(n31278), .X(n31275) );
  inv_x2_sg U39979 ( .A(n31269), .X(n41662) );
  nor_x1_sg U39980 ( .A(n31271), .B(n41665), .X(n31269) );
  inv_x2_sg U39981 ( .A(n25568), .X(n42171) );
  nor_x1_sg U39982 ( .A(n42174), .B(n51304), .X(n25568) );
  nand_x2_sg U39983 ( .A(n25872), .B(n25873), .X(n11163) );
  inv_x2_sg U39984 ( .A(n26129), .X(n42183) );
  nor_x1_sg U39985 ( .A(n42186), .B(n51865), .X(n26129) );
  nand_x2_sg U39986 ( .A(n26431), .B(n26432), .X(n12724) );
  nand_x2_sg U39987 ( .A(n26413), .B(n52132), .X(n12801) );
  nand_x2_sg U39988 ( .A(n26709), .B(n26710), .X(n13509) );
  nand_x2_sg U39989 ( .A(n26691), .B(n52405), .X(n13595) );
  nand_x2_sg U39990 ( .A(n26970), .B(n52682), .X(n14410) );
  nand_x2_sg U39991 ( .A(n27268), .B(n27269), .X(n15057) );
  nand_x2_sg U39992 ( .A(n27250), .B(n52966), .X(n15134) );
  inv_x2_sg U39993 ( .A(n27524), .X(n42167) );
  nor_x1_sg U39994 ( .A(n42170), .B(n53251), .X(n27524) );
  nand_x2_sg U39995 ( .A(n27826), .B(n27827), .X(n16623) );
  nand_x2_sg U39996 ( .A(n27808), .B(n53524), .X(n16700) );
  nand_x2_sg U39997 ( .A(n28368), .B(n28369), .X(n18267) );
  nand_x2_sg U39998 ( .A(n28925), .B(n54646), .X(n19845) );
  inv_x2_sg U39999 ( .A(n28920), .X(n42179) );
  nor_x1_sg U40000 ( .A(n42182), .B(n54658), .X(n28920) );
  nand_x2_sg U40001 ( .A(n29486), .B(n55214), .X(n21390) );
  inv_x2_sg U40002 ( .A(n29481), .X(n42175) );
  nor_x1_sg U40003 ( .A(n42178), .B(n55226), .X(n29481) );
  inv_x2_sg U40004 ( .A(n22522), .X(n43547) );
  nand_x4_sg U40005 ( .A(n22519), .B(n50956), .X(n21940) );
  inv_x1_sg U40006 ( .A(n22520), .X(n50956) );
  nand_x1_sg U40007 ( .A(n22521), .B(n21937), .X(n22519) );
  inv_x2_sg U40008 ( .A(n21975), .X(n43519) );
  inv_x2_sg U40009 ( .A(n22504), .X(n43521) );
  inv_x2_sg U40010 ( .A(n22804), .X(n42502) );
  inv_x2_sg U40011 ( .A(n10416), .X(n42151) );
  nor_x1_sg U40012 ( .A(n51295), .B(n10426), .X(n10416) );
  inv_x2_sg U40013 ( .A(n10441), .X(n43258) );
  inv_x2_sg U40014 ( .A(n10387), .X(n42604) );
  nand_x1_sg U40015 ( .A(n42152), .B(n10417), .X(n10387) );
  nor_x1_sg U40016 ( .A(n10470), .B(n51330), .X(n10469) );
  inv_x2_sg U40017 ( .A(n10468), .X(n43418) );
  nor_x1_sg U40018 ( .A(n10471), .B(n51344), .X(n10468) );
  inv_x2_sg U40019 ( .A(n10530), .X(n43204) );
  nor_x1_sg U40020 ( .A(n10553), .B(n51387), .X(n10530) );
  inv_x2_sg U40021 ( .A(n11188), .X(n42159) );
  nor_x1_sg U40022 ( .A(n51577), .B(n11200), .X(n11188) );
  inv_x2_sg U40023 ( .A(n11154), .X(n42616) );
  nand_x1_sg U40024 ( .A(n42160), .B(n11190), .X(n11154) );
  inv_x2_sg U40025 ( .A(n11245), .X(n43416) );
  inv_x2_sg U40026 ( .A(n11135), .X(n42051) );
  nor_x1_sg U40027 ( .A(n11665), .B(n51801), .X(n11135) );
  inv_x2_sg U40028 ( .A(n11134), .X(n41660) );
  nor_x1_sg U40029 ( .A(n11116), .B(n11137), .X(n11134) );
  inv_x2_sg U40030 ( .A(n11848), .X(n43156) );
  nor_x1_sg U40031 ( .A(n43159), .B(n51835), .X(n11848) );
  nand_x1_sg U40032 ( .A(n51820), .B(n51827), .X(n11939) );
  inv_x2_sg U40033 ( .A(n11993), .X(n43262) );
  inv_x2_sg U40034 ( .A(n12021), .X(n43412) );
  inv_x2_sg U40035 ( .A(n11918), .X(n42049) );
  nor_x1_sg U40036 ( .A(n12445), .B(n52077), .X(n11918) );
  inv_x2_sg U40037 ( .A(n11917), .X(n41658) );
  nor_x1_sg U40038 ( .A(n43231), .B(n11920), .X(n11917) );
  inv_x2_sg U40039 ( .A(n12749), .X(n42157) );
  nor_x1_sg U40040 ( .A(n52135), .B(n12761), .X(n12749) );
  inv_x2_sg U40041 ( .A(n12715), .X(n42614) );
  nand_x1_sg U40042 ( .A(n42158), .B(n12751), .X(n12715) );
  inv_x2_sg U40043 ( .A(n12806), .X(n43408) );
  inv_x2_sg U40044 ( .A(n12696), .X(n42047) );
  nor_x1_sg U40045 ( .A(n13226), .B(n52355), .X(n12696) );
  inv_x2_sg U40046 ( .A(n12695), .X(n41391) );
  nor_x1_sg U40047 ( .A(n12677), .B(n12698), .X(n12695) );
  inv_x2_sg U40048 ( .A(n13410), .X(n43152) );
  nor_x1_sg U40049 ( .A(n43155), .B(n52387), .X(n13410) );
  nand_x1_sg U40050 ( .A(n52372), .B(n52379), .X(n13501) );
  inv_x2_sg U40051 ( .A(n13554), .X(n43495) );
  inv_x2_sg U40052 ( .A(n13582), .X(n43404) );
  inv_x2_sg U40053 ( .A(n13434), .X(n41216) );
  nor_x1_sg U40054 ( .A(n13494), .B(n52467), .X(n13434) );
  inv_x2_sg U40055 ( .A(n13480), .X(n42045) );
  nor_x1_sg U40056 ( .A(n14006), .B(n52630), .X(n13480) );
  inv_x2_sg U40057 ( .A(n13479), .X(n41192) );
  nor_x1_sg U40058 ( .A(n13461), .B(n13482), .X(n13479) );
  inv_x2_sg U40059 ( .A(n14332), .X(n43511) );
  nor_x1_sg U40060 ( .A(n14362), .B(n52720), .X(n14361) );
  inv_x2_sg U40061 ( .A(n14360), .X(n43398) );
  nor_x1_sg U40062 ( .A(n14363), .B(n52734), .X(n14360) );
  inv_x2_sg U40063 ( .A(n14422), .X(n43218) );
  nor_x1_sg U40064 ( .A(n14445), .B(n52774), .X(n14422) );
  inv_x2_sg U40065 ( .A(n14259), .X(n42043) );
  nor_x1_sg U40066 ( .A(n14777), .B(n52911), .X(n14259) );
  inv_x2_sg U40067 ( .A(n15082), .X(n42155) );
  nor_x1_sg U40068 ( .A(n52969), .B(n15094), .X(n15082) );
  inv_x2_sg U40069 ( .A(n15048), .X(n42612) );
  nand_x1_sg U40070 ( .A(n42156), .B(n15084), .X(n15048) );
  inv_x2_sg U40071 ( .A(n15139), .X(n43396) );
  inv_x2_sg U40072 ( .A(n15029), .X(n42041) );
  nor_x1_sg U40073 ( .A(n15559), .B(n53189), .X(n15029) );
  inv_x2_sg U40074 ( .A(n15028), .X(n41383) );
  nor_x1_sg U40075 ( .A(n15010), .B(n15031), .X(n15028) );
  inv_x2_sg U40076 ( .A(n15743), .X(n43142) );
  nor_x1_sg U40077 ( .A(n43145), .B(n53223), .X(n15743) );
  nand_x1_sg U40078 ( .A(n53208), .B(n53215), .X(n15834) );
  inv_x2_sg U40079 ( .A(n15888), .X(n43256) );
  inv_x2_sg U40080 ( .A(n15916), .X(n43392) );
  inv_x2_sg U40081 ( .A(n16648), .X(n42153) );
  nor_x1_sg U40082 ( .A(n53527), .B(n16660), .X(n16648) );
  inv_x2_sg U40083 ( .A(n16614), .X(n42610) );
  nand_x1_sg U40084 ( .A(n42154), .B(n16650), .X(n16614) );
  inv_x2_sg U40085 ( .A(n16705), .X(n43388) );
  inv_x2_sg U40086 ( .A(n16595), .X(n42039) );
  nor_x1_sg U40087 ( .A(n17125), .B(n53747), .X(n16595) );
  inv_x2_sg U40088 ( .A(n16594), .X(n41377) );
  nor_x1_sg U40089 ( .A(n16576), .B(n16597), .X(n16594) );
  inv_x2_sg U40090 ( .A(n17429), .X(n42165) );
  nor_x1_sg U40091 ( .A(n53804), .B(n17441), .X(n17429) );
  inv_x2_sg U40092 ( .A(n17455), .X(n43507) );
  inv_x2_sg U40093 ( .A(n17398), .X(n42623) );
  nand_x1_sg U40094 ( .A(n42166), .B(n17430), .X(n17398) );
  nor_x1_sg U40095 ( .A(n17484), .B(n53834), .X(n17483) );
  inv_x2_sg U40096 ( .A(n17482), .X(n43382) );
  nor_x1_sg U40097 ( .A(n17485), .B(n53854), .X(n17482) );
  inv_x2_sg U40098 ( .A(n17542), .X(n43216) );
  nor_x1_sg U40099 ( .A(n17565), .B(n53894), .X(n17542) );
  inv_x2_sg U40100 ( .A(n17378), .X(n42037) );
  nor_x1_sg U40101 ( .A(n17898), .B(n54031), .X(n17378) );
  inv_x2_sg U40102 ( .A(n18221), .X(n42470) );
  inv_x2_sg U40103 ( .A(n18312), .X(n43210) );
  nor_x1_sg U40104 ( .A(n18335), .B(n54175), .X(n18312) );
  inv_x2_sg U40105 ( .A(n18149), .X(n42035) );
  nor_x1_sg U40106 ( .A(n18667), .B(n54312), .X(n18149) );
  inv_x2_sg U40107 ( .A(n18148), .X(n41656) );
  nor_x1_sg U40108 ( .A(n43229), .B(n18151), .X(n18148) );
  inv_x2_sg U40109 ( .A(n18974), .X(n42163) );
  nor_x1_sg U40110 ( .A(n54369), .B(n18986), .X(n18974) );
  inv_x2_sg U40111 ( .A(n19000), .X(n43503) );
  inv_x2_sg U40112 ( .A(n18943), .X(n42621) );
  nand_x1_sg U40113 ( .A(n42164), .B(n18975), .X(n18943) );
  nor_x1_sg U40114 ( .A(n19029), .B(n54399), .X(n19028) );
  inv_x2_sg U40115 ( .A(n19027), .X(n43378) );
  nor_x1_sg U40116 ( .A(n19030), .B(n54419), .X(n19027) );
  inv_x2_sg U40117 ( .A(n19087), .X(n43214) );
  nor_x1_sg U40118 ( .A(n19110), .B(n54459), .X(n19087) );
  inv_x2_sg U40119 ( .A(n18923), .X(n42033) );
  nor_x1_sg U40120 ( .A(n19443), .B(n54596), .X(n18923) );
  inv_x2_sg U40121 ( .A(n19624), .X(n41593) );
  nor_x1_sg U40122 ( .A(n54616), .B(n19718), .X(n19624) );
  inv_x2_sg U40123 ( .A(n19625), .X(n43148) );
  nor_x1_sg U40124 ( .A(n43151), .B(n54628), .X(n19625) );
  nand_x1_sg U40125 ( .A(n54615), .B(n19729), .X(n19716) );
  inv_x2_sg U40126 ( .A(n19743), .X(n41963) );
  nor_x1_sg U40127 ( .A(n54649), .B(n19753), .X(n19743) );
  inv_x2_sg U40128 ( .A(n19767), .X(n43493) );
  inv_x2_sg U40129 ( .A(n19714), .X(n42608) );
  nand_x1_sg U40130 ( .A(n41964), .B(n19744), .X(n19714) );
  nor_x1_sg U40131 ( .A(n19797), .B(n54684), .X(n19796) );
  inv_x2_sg U40132 ( .A(n19795), .X(n43374) );
  nor_x1_sg U40133 ( .A(n19798), .B(n54698), .X(n19795) );
  inv_x2_sg U40134 ( .A(n19857), .X(n43208) );
  nor_x1_sg U40135 ( .A(n19880), .B(n54741), .X(n19857) );
  inv_x2_sg U40136 ( .A(n19694), .X(n42031) );
  nor_x1_sg U40137 ( .A(n20212), .B(n54880), .X(n19694) );
  inv_x2_sg U40138 ( .A(n19693), .X(n41654) );
  nor_x1_sg U40139 ( .A(n43227), .B(n19696), .X(n19693) );
  inv_x2_sg U40140 ( .A(n20518), .X(n42161) );
  nor_x1_sg U40141 ( .A(n54937), .B(n20530), .X(n20518) );
  inv_x2_sg U40142 ( .A(n20544), .X(n43499) );
  inv_x2_sg U40143 ( .A(n20487), .X(n42619) );
  nand_x1_sg U40144 ( .A(n42162), .B(n20519), .X(n20487) );
  nor_x1_sg U40145 ( .A(n20573), .B(n54967), .X(n20572) );
  inv_x2_sg U40146 ( .A(n20571), .X(n43370) );
  nor_x1_sg U40147 ( .A(n20574), .B(n54987), .X(n20571) );
  inv_x2_sg U40148 ( .A(n20631), .X(n43212) );
  nor_x1_sg U40149 ( .A(n20654), .B(n55027), .X(n20631) );
  inv_x2_sg U40150 ( .A(n20467), .X(n42029) );
  nor_x1_sg U40151 ( .A(n20987), .B(n55164), .X(n20467) );
  inv_x2_sg U40152 ( .A(n21261), .X(n42626) );
  nand_x1_sg U40153 ( .A(n55183), .B(n21274), .X(n21261) );
  inv_x2_sg U40154 ( .A(n21288), .X(n41961) );
  nor_x1_sg U40155 ( .A(n55217), .B(n21298), .X(n21288) );
  inv_x2_sg U40156 ( .A(n21312), .X(n43489) );
  inv_x2_sg U40157 ( .A(n21259), .X(n42606) );
  nand_x1_sg U40158 ( .A(n41962), .B(n21289), .X(n21259) );
  nor_x1_sg U40159 ( .A(n21342), .B(n55252), .X(n21341) );
  inv_x2_sg U40160 ( .A(n21340), .X(n43366) );
  nor_x1_sg U40161 ( .A(n21343), .B(n55266), .X(n21340) );
  inv_x2_sg U40162 ( .A(n21402), .X(n43206) );
  nor_x1_sg U40163 ( .A(n21425), .B(n55309), .X(n21402) );
  inv_x2_sg U40164 ( .A(n21239), .X(n42027) );
  nor_x1_sg U40165 ( .A(n21757), .B(n55448), .X(n21239) );
  inv_x2_sg U40166 ( .A(n21238), .X(n41652) );
  nor_x1_sg U40167 ( .A(n43225), .B(n21241), .X(n21238) );
  inv_x2_sg U40168 ( .A(n30188), .X(n43545) );
  nand_x4_sg U40169 ( .A(n30185), .B(n50097), .X(n29592) );
  inv_x1_sg U40170 ( .A(n30186), .X(n50097) );
  nand_x1_sg U40171 ( .A(n30187), .B(n29588), .X(n30185) );
  inv_x2_sg U40172 ( .A(n29640), .X(n43515) );
  inv_x2_sg U40173 ( .A(n30170), .X(n43517) );
  inv_x2_sg U40174 ( .A(n30470), .X(n42498) );
  nand_x2_sg U40175 ( .A(n25539), .B(n51395), .X(n10735) );
  inv_x2_sg U40176 ( .A(n43812), .X(n43813) );
  inv_x1_sg U40177 ( .A(n11199), .X(n43812) );
  inv_x2_sg U40178 ( .A(n43869), .X(n43870) );
  inv_x1_sg U40179 ( .A(n12760), .X(n43869) );
  inv_x1_sg U40180 ( .A(n26407), .X(n46198) );
  nand_x2_sg U40181 ( .A(n52694), .B(n26964), .X(n14382) );
  inv_x2_sg U40182 ( .A(n43867), .X(n43868) );
  inv_x1_sg U40183 ( .A(n15093), .X(n43867) );
  inv_x1_sg U40184 ( .A(n27244), .X(n46197) );
  inv_x2_sg U40185 ( .A(n43865), .X(n43866) );
  inv_x1_sg U40186 ( .A(n16659), .X(n43865) );
  inv_x1_sg U40187 ( .A(n27802), .X(n46196) );
  nor_x2_sg U40188 ( .A(n44140), .B(n43773), .X(n10390) );
  inv_x2_sg U40189 ( .A(n10301), .X(n43110) );
  nor_x1_sg U40190 ( .A(n43113), .B(n10405), .X(n10301) );
  inv_x2_sg U40191 ( .A(n10469), .X(n43420) );
  inv_x2_sg U40192 ( .A(n10321), .X(n41450) );
  nor_x1_sg U40193 ( .A(n10382), .B(n51363), .X(n10321) );
  inv_x2_sg U40194 ( .A(n10323), .X(n41739) );
  nor_x1_sg U40195 ( .A(n10382), .B(n51365), .X(n10323) );
  inv_x2_sg U40196 ( .A(n10353), .X(n42930) );
  nor_x1_sg U40197 ( .A(n42933), .B(n51512), .X(n10353) );
  inv_x2_sg U40198 ( .A(n11069), .X(n43128) );
  nor_x1_sg U40199 ( .A(n11176), .B(n11177), .X(n11069) );
  inv_x2_sg U40200 ( .A(n51565), .X(n41882) );
  inv_x1_sg U40201 ( .A(n11156), .X(n51565) );
  inv_x2_sg U40202 ( .A(n11089), .X(n41466) );
  nor_x1_sg U40203 ( .A(n11149), .B(n51634), .X(n11089) );
  inv_x2_sg U40204 ( .A(n11091), .X(n41759) );
  nor_x1_sg U40205 ( .A(n11149), .B(n51636), .X(n11091) );
  inv_x2_sg U40206 ( .A(n11117), .X(n43202) );
  nor_x1_sg U40207 ( .A(n11545), .B(n11546), .X(n11117) );
  inv_x2_sg U40208 ( .A(n11120), .X(n42926) );
  nor_x1_sg U40209 ( .A(n42929), .B(n51792), .X(n11120) );
  inv_x2_sg U40210 ( .A(n11872), .X(n41464) );
  nor_x1_sg U40211 ( .A(n11932), .B(n51915), .X(n11872) );
  inv_x2_sg U40212 ( .A(n11874), .X(n41757) );
  nor_x1_sg U40213 ( .A(n11932), .B(n51917), .X(n11874) );
  inv_x2_sg U40214 ( .A(n11900), .X(n42346) );
  nor_x1_sg U40215 ( .A(n12325), .B(n12326), .X(n11900) );
  inv_x2_sg U40216 ( .A(n11903), .X(n42023) );
  nor_x1_sg U40217 ( .A(n42026), .B(n52070), .X(n11903) );
  inv_x2_sg U40218 ( .A(n12630), .X(n43126) );
  nor_x1_sg U40219 ( .A(n12737), .B(n12738), .X(n12630) );
  inv_x2_sg U40220 ( .A(n52122), .X(n41880) );
  inv_x1_sg U40221 ( .A(n12717), .X(n52122) );
  inv_x2_sg U40222 ( .A(n12650), .X(n41462) );
  nor_x1_sg U40223 ( .A(n12710), .B(n52190), .X(n12650) );
  inv_x2_sg U40224 ( .A(n12652), .X(n41755) );
  nor_x1_sg U40225 ( .A(n12710), .B(n52192), .X(n12652) );
  inv_x2_sg U40226 ( .A(n12678), .X(n43200) );
  nor_x1_sg U40227 ( .A(n13106), .B(n13107), .X(n12678) );
  inv_x2_sg U40228 ( .A(n12681), .X(n42019) );
  nor_x1_sg U40229 ( .A(n42022), .B(n52348), .X(n12681) );
  inv_x2_sg U40230 ( .A(n13436), .X(n41753) );
  nor_x1_sg U40231 ( .A(n13494), .B(n52469), .X(n13436) );
  inv_x2_sg U40232 ( .A(n13462), .X(n43198) );
  nor_x1_sg U40233 ( .A(n13886), .B(n13887), .X(n13462) );
  inv_x2_sg U40234 ( .A(n13465), .X(n42015) );
  nor_x1_sg U40235 ( .A(n42018), .B(n52623), .X(n13465) );
  inv_x2_sg U40236 ( .A(n44025), .X(n44026) );
  inv_x1_sg U40237 ( .A(n14182), .X(n44025) );
  nor_x2_sg U40238 ( .A(n44405), .B(n43802), .X(n14282) );
  inv_x2_sg U40239 ( .A(n14193), .X(n43146) );
  nor_x1_sg U40240 ( .A(n14296), .B(n14297), .X(n14193) );
  inv_x2_sg U40241 ( .A(n14361), .X(n43400) );
  inv_x2_sg U40242 ( .A(n14213), .X(n41474) );
  nor_x1_sg U40243 ( .A(n14274), .B(n52753), .X(n14213) );
  inv_x2_sg U40244 ( .A(n14215), .X(n41777) );
  nor_x1_sg U40245 ( .A(n14274), .B(n52755), .X(n14215) );
  inv_x2_sg U40246 ( .A(n14244), .X(n42922) );
  nor_x1_sg U40247 ( .A(n42925), .B(n52902), .X(n14244) );
  inv_x2_sg U40248 ( .A(n14963), .X(n43124) );
  nor_x1_sg U40249 ( .A(n15070), .B(n15071), .X(n14963) );
  nor_x2_sg U40250 ( .A(n43125), .B(n41826), .X(n15050) );
  inv_x2_sg U40251 ( .A(n14983), .X(n41460) );
  nor_x1_sg U40252 ( .A(n15043), .B(n53024), .X(n14983) );
  inv_x2_sg U40253 ( .A(n14985), .X(n41751) );
  nor_x1_sg U40254 ( .A(n15043), .B(n53026), .X(n14985) );
  inv_x2_sg U40255 ( .A(n15011), .X(n43196) );
  nor_x1_sg U40256 ( .A(n15439), .B(n15440), .X(n15011) );
  inv_x2_sg U40257 ( .A(n15014), .X(n42011) );
  nor_x1_sg U40258 ( .A(n42014), .B(n53182), .X(n15014) );
  inv_x2_sg U40259 ( .A(n44021), .X(n44022) );
  inv_x1_sg U40260 ( .A(n15736), .X(n44021) );
  inv_x2_sg U40261 ( .A(n15767), .X(n41448) );
  nor_x1_sg U40262 ( .A(n15827), .B(n53302), .X(n15767) );
  inv_x2_sg U40263 ( .A(n15769), .X(n41735) );
  nor_x1_sg U40264 ( .A(n15827), .B(n53304), .X(n15769) );
  inv_x2_sg U40265 ( .A(n15799), .X(n42918) );
  nor_x1_sg U40266 ( .A(n42921), .B(n53462), .X(n15799) );
  inv_x2_sg U40267 ( .A(n16529), .X(n43122) );
  nor_x1_sg U40268 ( .A(n16636), .B(n16637), .X(n16529) );
  nor_x2_sg U40269 ( .A(n43123), .B(n41824), .X(n16616) );
  inv_x2_sg U40270 ( .A(n16549), .X(n41458) );
  nor_x1_sg U40271 ( .A(n16609), .B(n53582), .X(n16549) );
  inv_x2_sg U40272 ( .A(n16551), .X(n41749) );
  nor_x1_sg U40273 ( .A(n16609), .B(n53584), .X(n16551) );
  inv_x2_sg U40274 ( .A(n16577), .X(n43194) );
  nor_x1_sg U40275 ( .A(n17005), .B(n17006), .X(n16577) );
  inv_x2_sg U40276 ( .A(n16580), .X(n42007) );
  nor_x1_sg U40277 ( .A(n42010), .B(n53740), .X(n16580) );
  inv_x2_sg U40278 ( .A(n17483), .X(n43384) );
  inv_x2_sg U40279 ( .A(n17332), .X(n41472) );
  nor_x1_sg U40280 ( .A(n17393), .B(n53873), .X(n17332) );
  inv_x2_sg U40281 ( .A(n17334), .X(n41775) );
  nor_x1_sg U40282 ( .A(n17393), .B(n53875), .X(n17334) );
  inv_x2_sg U40283 ( .A(n17363), .X(n42914) );
  nor_x1_sg U40284 ( .A(n42917), .B(n54022), .X(n17363) );
  inv_x2_sg U40285 ( .A(n18104), .X(n41456) );
  nor_x1_sg U40286 ( .A(n18164), .B(n54152), .X(n18104) );
  inv_x2_sg U40287 ( .A(n18106), .X(n41747) );
  nor_x1_sg U40288 ( .A(n18164), .B(n54154), .X(n18106) );
  inv_x2_sg U40289 ( .A(n18132), .X(n42344) );
  nor_x1_sg U40290 ( .A(n18544), .B(n18545), .X(n18132) );
  inv_x2_sg U40291 ( .A(n18135), .X(n42910) );
  nor_x1_sg U40292 ( .A(n42913), .B(n54303), .X(n18135) );
  inv_x2_sg U40293 ( .A(n19028), .X(n43380) );
  inv_x2_sg U40294 ( .A(n18877), .X(n41470) );
  nor_x1_sg U40295 ( .A(n18938), .B(n54438), .X(n18877) );
  inv_x2_sg U40296 ( .A(n18879), .X(n41773) );
  nor_x1_sg U40297 ( .A(n18938), .B(n54440), .X(n18879) );
  inv_x2_sg U40298 ( .A(n18908), .X(n42906) );
  nor_x1_sg U40299 ( .A(n42909), .B(n54587), .X(n18908) );
  inv_x2_sg U40300 ( .A(n19629), .X(n43118) );
  nor_x1_sg U40301 ( .A(n43121), .B(n19732), .X(n19629) );
  inv_x2_sg U40302 ( .A(n19796), .X(n43376) );
  inv_x2_sg U40303 ( .A(n19649), .X(n41454) );
  nor_x1_sg U40304 ( .A(n19709), .B(n54717), .X(n19649) );
  inv_x2_sg U40305 ( .A(n19651), .X(n41745) );
  nor_x1_sg U40306 ( .A(n19709), .B(n54719), .X(n19651) );
  inv_x2_sg U40307 ( .A(n19677), .X(n42342) );
  nor_x1_sg U40308 ( .A(n20089), .B(n20090), .X(n19677) );
  inv_x2_sg U40309 ( .A(n19680), .X(n42902) );
  nor_x1_sg U40310 ( .A(n42905), .B(n54871), .X(n19680) );
  inv_x2_sg U40311 ( .A(n20572), .X(n43372) );
  inv_x2_sg U40312 ( .A(n20421), .X(n41468) );
  nor_x1_sg U40313 ( .A(n20482), .B(n55006), .X(n20421) );
  inv_x2_sg U40314 ( .A(n20423), .X(n41771) );
  nor_x1_sg U40315 ( .A(n20482), .B(n55008), .X(n20423) );
  inv_x2_sg U40316 ( .A(n20452), .X(n42898) );
  nor_x1_sg U40317 ( .A(n42901), .B(n55155), .X(n20452) );
  inv_x2_sg U40318 ( .A(n21169), .X(n42814) );
  nor_x1_sg U40319 ( .A(n55184), .B(n21263), .X(n21169) );
  nor_x2_sg U40320 ( .A(n44138), .B(n42815), .X(n21262) );
  inv_x2_sg U40321 ( .A(n21174), .X(n43114) );
  nor_x1_sg U40322 ( .A(n43117), .B(n21277), .X(n21174) );
  inv_x2_sg U40323 ( .A(n21341), .X(n43368) );
  inv_x2_sg U40324 ( .A(n21194), .X(n41452) );
  nor_x1_sg U40325 ( .A(n21254), .B(n55285), .X(n21194) );
  inv_x2_sg U40326 ( .A(n21196), .X(n41743) );
  nor_x1_sg U40327 ( .A(n21254), .B(n55287), .X(n21196) );
  inv_x2_sg U40328 ( .A(n21222), .X(n42340) );
  nor_x1_sg U40329 ( .A(n21634), .B(n21635), .X(n21222) );
  inv_x2_sg U40330 ( .A(n21225), .X(n42894) );
  nor_x1_sg U40331 ( .A(n42897), .B(n55439), .X(n21225) );
  inv_x2_sg U40332 ( .A(n51797), .X(n41647) );
  inv_x1_sg U40333 ( .A(n11694), .X(n51797) );
  inv_x2_sg U40334 ( .A(n52073), .X(n41645) );
  inv_x1_sg U40335 ( .A(n12473), .X(n52073) );
  nand_x2_sg U40336 ( .A(n55468), .B(n46576), .X(n13392) );
  inv_x2_sg U40337 ( .A(n52351), .X(n41643) );
  inv_x1_sg U40338 ( .A(n13254), .X(n52351) );
  nand_x2_sg U40339 ( .A(n55470), .B(n46576), .X(n14172) );
  inv_x2_sg U40340 ( .A(n52626), .X(n41641) );
  inv_x1_sg U40341 ( .A(n14034), .X(n52626) );
  inv_x2_sg U40342 ( .A(n52907), .X(n41639) );
  inv_x1_sg U40343 ( .A(n14806), .X(n52907) );
  inv_x2_sg U40344 ( .A(n53185), .X(n41637) );
  inv_x1_sg U40345 ( .A(n15587), .X(n53185) );
  inv_x2_sg U40346 ( .A(n53465), .X(n41621) );
  inv_x1_sg U40347 ( .A(n16368), .X(n53465) );
  inv_x2_sg U40348 ( .A(n53743), .X(n41635) );
  inv_x1_sg U40349 ( .A(n17153), .X(n53743) );
  inv_x2_sg U40350 ( .A(n54027), .X(n41633) );
  inv_x1_sg U40351 ( .A(n17927), .X(n54027) );
  inv_x2_sg U40352 ( .A(n54308), .X(n41631) );
  inv_x1_sg U40353 ( .A(n18696), .X(n54308) );
  inv_x2_sg U40354 ( .A(n54592), .X(n41629) );
  inv_x1_sg U40355 ( .A(n19472), .X(n54592) );
  inv_x2_sg U40356 ( .A(n54876), .X(n41627) );
  inv_x1_sg U40357 ( .A(n20242), .X(n54876) );
  inv_x2_sg U40358 ( .A(n55160), .X(n41625) );
  inv_x1_sg U40359 ( .A(n21016), .X(n55160) );
  nand_x2_sg U40360 ( .A(n46576), .B(n9406), .X(n21926) );
  inv_x2_sg U40361 ( .A(n55444), .X(n41623) );
  inv_x1_sg U40362 ( .A(n21787), .X(n55444) );
  inv_x2_sg U40363 ( .A(n9026), .X(n42005) );
  nor_x1_sg U40364 ( .A(n10314), .B(n51345), .X(n9026) );
  inv_x2_sg U40365 ( .A(n9022), .X(n42892) );
  nor_x1_sg U40366 ( .A(n10331), .B(n51429), .X(n9022) );
  inv_x2_sg U40367 ( .A(n8889), .X(n42890) );
  nor_x1_sg U40368 ( .A(n11052), .B(n11053), .X(n8889) );
  inv_x2_sg U40369 ( .A(n8891), .X(n42001) );
  nor_x1_sg U40370 ( .A(n42004), .B(n51624), .X(n8891) );
  inv_x2_sg U40371 ( .A(n8884), .X(n42888) );
  nor_x1_sg U40372 ( .A(n11099), .B(n51702), .X(n8884) );
  nand_x2_sg U40373 ( .A(n46580), .B(n46553), .X(n11049) );
  inv_x2_sg U40374 ( .A(n8915), .X(n41365) );
  nand_x1_sg U40375 ( .A(n41175), .B(n11846), .X(n8915) );
  inv_x2_sg U40376 ( .A(n8925), .X(n41997) );
  nor_x1_sg U40377 ( .A(n42000), .B(n51906), .X(n8925) );
  inv_x2_sg U40378 ( .A(n8921), .X(n42886) );
  nor_x1_sg U40379 ( .A(n11882), .B(n51983), .X(n8921) );
  nand_x2_sg U40380 ( .A(n46580), .B(n46531), .X(n11832) );
  inv_x2_sg U40381 ( .A(n8844), .X(n42884) );
  nor_x1_sg U40382 ( .A(n12613), .B(n12614), .X(n8844) );
  inv_x2_sg U40383 ( .A(n8855), .X(n41993) );
  nor_x1_sg U40384 ( .A(n41996), .B(n52183), .X(n8855) );
  inv_x2_sg U40385 ( .A(n8851), .X(n42882) );
  nor_x1_sg U40386 ( .A(n12660), .B(n52258), .X(n8851) );
  nand_x2_sg U40387 ( .A(n46580), .B(n46510), .X(n12610) );
  inv_x2_sg U40388 ( .A(n8815), .X(n41363) );
  nand_x1_sg U40389 ( .A(n41174), .B(n13408), .X(n8815) );
  inv_x2_sg U40390 ( .A(n8817), .X(n41989) );
  nor_x1_sg U40391 ( .A(n41992), .B(n52459), .X(n8817) );
  inv_x2_sg U40392 ( .A(n8803), .X(n41361) );
  nand_x1_sg U40393 ( .A(n13431), .B(n52468), .X(n8803) );
  inv_x2_sg U40394 ( .A(n8811), .X(n42880) );
  nor_x1_sg U40395 ( .A(n13444), .B(n52534), .X(n8811) );
  nand_x2_sg U40396 ( .A(n46580), .B(n46487), .X(n13394) );
  inv_x2_sg U40397 ( .A(n8958), .X(n41987) );
  nor_x1_sg U40398 ( .A(n14206), .B(n52735), .X(n8958) );
  inv_x2_sg U40399 ( .A(n9000), .X(n42878) );
  nor_x1_sg U40400 ( .A(n14223), .B(n52819), .X(n9000) );
  nand_x2_sg U40401 ( .A(n46580), .B(n46465), .X(n14173) );
  inv_x2_sg U40402 ( .A(n8983), .X(n42876) );
  nor_x1_sg U40403 ( .A(n14946), .B(n14947), .X(n8983) );
  inv_x2_sg U40404 ( .A(n8985), .X(n41983) );
  nor_x1_sg U40405 ( .A(n41986), .B(n53017), .X(n8985) );
  inv_x2_sg U40406 ( .A(n8994), .X(n42874) );
  nor_x1_sg U40407 ( .A(n14993), .B(n53092), .X(n8994) );
  nand_x2_sg U40408 ( .A(n46580), .B(n46442), .X(n14943) );
  inv_x2_sg U40409 ( .A(n9353), .X(n41359) );
  nand_x1_sg U40410 ( .A(n41173), .B(n15741), .X(n9353) );
  inv_x2_sg U40411 ( .A(n9320), .X(n41979) );
  nor_x1_sg U40412 ( .A(n41982), .B(n53291), .X(n9320) );
  inv_x2_sg U40413 ( .A(n9345), .X(n42872) );
  nor_x1_sg U40414 ( .A(n15777), .B(n53372), .X(n9345) );
  nand_x2_sg U40415 ( .A(n46580), .B(n46419), .X(n15727) );
  inv_x2_sg U40416 ( .A(n9302), .X(n42870) );
  nor_x1_sg U40417 ( .A(n16512), .B(n16513), .X(n9302) );
  inv_x2_sg U40418 ( .A(n9309), .X(n41975) );
  nor_x1_sg U40419 ( .A(n41978), .B(n53575), .X(n9309) );
  inv_x2_sg U40420 ( .A(n9305), .X(n42868) );
  nor_x1_sg U40421 ( .A(n16559), .B(n53650), .X(n9305) );
  nand_x2_sg U40422 ( .A(n46580), .B(n46398), .X(n16509) );
  inv_x2_sg U40423 ( .A(n9264), .X(n41357) );
  nor_x1_sg U40424 ( .A(n17295), .B(n17296), .X(n9264) );
  inv_x2_sg U40425 ( .A(n9271), .X(n41973) );
  nor_x1_sg U40426 ( .A(n17325), .B(n53855), .X(n9271) );
  inv_x2_sg U40427 ( .A(n9267), .X(n42866) );
  nor_x1_sg U40428 ( .A(n17342), .B(n53939), .X(n9267) );
  nand_x2_sg U40429 ( .A(n46580), .B(n46375), .X(n17292) );
  inv_x2_sg U40430 ( .A(n9083), .X(n42628) );
  nand_x1_sg U40431 ( .A(n54061), .B(n18078), .X(n9083) );
  inv_x2_sg U40432 ( .A(n9079), .X(n42864) );
  nor_x1_sg U40433 ( .A(n18114), .B(n54219), .X(n9079) );
  nand_x2_sg U40434 ( .A(n46580), .B(n46355), .X(n18064) );
  inv_x2_sg U40435 ( .A(n9226), .X(n41355) );
  nor_x1_sg U40436 ( .A(n18840), .B(n18841), .X(n9226) );
  inv_x2_sg U40437 ( .A(n9233), .X(n41971) );
  nor_x1_sg U40438 ( .A(n18870), .B(n54420), .X(n9233) );
  inv_x2_sg U40439 ( .A(n9229), .X(n42862) );
  nor_x1_sg U40440 ( .A(n18887), .B(n54504), .X(n9229) );
  nand_x2_sg U40441 ( .A(n46580), .B(n46327), .X(n18837) );
  inv_x2_sg U40442 ( .A(n9197), .X(n41353) );
  nand_x1_sg U40443 ( .A(n54629), .B(n19623), .X(n9197) );
  inv_x2_sg U40444 ( .A(n9175), .X(n41969) );
  nor_x1_sg U40445 ( .A(n19642), .B(n54699), .X(n9175) );
  inv_x2_sg U40446 ( .A(n9189), .X(n42860) );
  nor_x1_sg U40447 ( .A(n19659), .B(n54788), .X(n9189) );
  nand_x2_sg U40448 ( .A(n46580), .B(n46308), .X(n19609) );
  inv_x2_sg U40449 ( .A(n9150), .X(n41351) );
  nor_x1_sg U40450 ( .A(n20384), .B(n20385), .X(n9150) );
  inv_x2_sg U40451 ( .A(n9157), .X(n41967) );
  nor_x1_sg U40452 ( .A(n20414), .B(n54988), .X(n9157) );
  inv_x2_sg U40453 ( .A(n9153), .X(n42858) );
  nor_x1_sg U40454 ( .A(n20431), .B(n55072), .X(n9153) );
  nand_x2_sg U40455 ( .A(n46580), .B(n46283), .X(n20381) );
  inv_x2_sg U40456 ( .A(n9121), .X(n41965) );
  nor_x1_sg U40457 ( .A(n21187), .B(n55267), .X(n9121) );
  inv_x2_sg U40458 ( .A(n9105), .X(n42856) );
  nor_x1_sg U40459 ( .A(n21204), .B(n55356), .X(n9105) );
  nand_x2_sg U40460 ( .A(n46580), .B(n46263), .X(n21154) );
  nand_x2_sg U40461 ( .A(n13392), .B(n26358), .X(n26225) );
  nand_x2_sg U40462 ( .A(n14172), .B(n26358), .X(n26504) );
  nand_x2_sg U40463 ( .A(n27194), .B(n26783), .X(n27061) );
  nand_x1_sg U40464 ( .A(n26079), .B(n46583), .X(n27194) );
  nand_x2_sg U40465 ( .A(n46592), .B(n28313), .X(n28180) );
  nand_x1_sg U40466 ( .A(n26079), .B(n55459), .X(n28313) );
  nand_x2_sg U40467 ( .A(n21926), .B(n26358), .X(n29299) );
  inv_x4_sg U40468 ( .A(n46640), .X(n46639) );
  inv_x1_sg U40469 ( .A(n46672), .X(n46671) );
  inv_x1_sg U40470 ( .A(n46672), .X(n46661) );
  inv_x1_sg U40471 ( .A(n28459), .X(n46595) );
  inv_x4_sg U40472 ( .A(n46610), .X(n46609) );
  inv_x4_sg U40473 ( .A(n9403), .X(n46601) );
  inv_x4_sg U40474 ( .A(n9399), .X(n46599) );
  inv_x4_sg U40475 ( .A(n28180), .X(n46594) );
  inv_x4_sg U40476 ( .A(n27061), .X(n46590) );
  inv_x4_sg U40477 ( .A(n26225), .X(n46586) );
  inv_x4_sg U40478 ( .A(n26504), .X(n46588) );
  inv_x4_sg U40479 ( .A(n29299), .X(n46597) );
  inv_x4_sg U40480 ( .A(n13394), .X(n46482) );
  inv_x4_sg U40481 ( .A(n16509), .X(n46392) );
  inv_x4_sg U40482 ( .A(n21154), .X(n46257) );
  inv_x4_sg U40483 ( .A(n55789), .X(n46374) );
  inv_x4_sg U40484 ( .A(n44175), .X(n46530) );
  inv_x4_sg U40485 ( .A(n43856), .X(n46307) );
  inv_x4_sg U40486 ( .A(n12610), .X(n46504) );
  inv_x4_sg U40487 ( .A(n15727), .X(n46414) );
  inv_x4_sg U40488 ( .A(n14173), .X(n46459) );
  inv_x4_sg U40489 ( .A(n11164), .X(n46550) );
  inv_x4_sg U40490 ( .A(n16624), .X(n46394) );
  inv_x4_sg U40491 ( .A(n15058), .X(n46438) );
  inv_x4_sg U40492 ( .A(n12725), .X(n46506) );
  inv_x4_sg U40493 ( .A(n11049), .X(n46548) );
  inv_x4_sg U40494 ( .A(n18837), .X(n46322) );
  inv_x4_sg U40495 ( .A(n17292), .X(n46369) );
  inv_x4_sg U40496 ( .A(n10282), .X(n46571) );
  inv_x4_sg U40497 ( .A(n19730), .X(n46304) );
  inv_x4_sg U40498 ( .A(n21275), .X(n46259) );
  inv_x4_sg U40499 ( .A(n55786), .X(n46624) );
  inv_x4_sg U40500 ( .A(n55785), .X(n46622) );
  inv_x4_sg U40501 ( .A(n55784), .X(n46620) );
  inv_x4_sg U40502 ( .A(n46618), .X(n46617) );
  inv_x4_sg U40503 ( .A(n46614), .X(n46613) );
  inv_x4_sg U40504 ( .A(n46605), .X(n46604) );
  inv_x4_sg U40505 ( .A(n43880), .X(n46253) );
  inv_x4_sg U40506 ( .A(n43876), .X(n46298) );
  inv_x4_sg U40507 ( .A(n55793), .X(n46464) );
  inv_x4_sg U40508 ( .A(n55787), .X(n46509) );
  inv_x4_sg U40509 ( .A(n55788), .X(n46486) );
  inv_x4_sg U40510 ( .A(n55792), .X(n46418) );
  inv_x4_sg U40511 ( .A(n55791), .X(n46397) );
  inv_x4_sg U40512 ( .A(n55790), .X(n46262) );
  inv_x4_sg U40513 ( .A(n15842), .X(n46408) );
  inv_x4_sg U40514 ( .A(n13509), .X(n46476) );
  inv_x4_sg U40515 ( .A(n14289), .X(n46453) );
  inv_x4_sg U40516 ( .A(n11947), .X(n46520) );
  inv_x4_sg U40517 ( .A(n44429), .X(n46354) );
  inv_x4_sg U40518 ( .A(n44173), .X(n46441) );
  inv_x4_sg U40519 ( .A(n44171), .X(n46282) );
  inv_x4_sg U40520 ( .A(n20381), .X(n46277) );
  inv_x4_sg U40521 ( .A(n11832), .X(n46526) );
  inv_x4_sg U40522 ( .A(n19609), .X(n46302) );
  inv_x4_sg U40523 ( .A(n14943), .X(n46436) );
  inv_x4_sg U40524 ( .A(n18064), .X(n46349) );
  inv_x4_sg U40525 ( .A(n18065), .X(n46347) );
  inv_x4_sg U40526 ( .A(n14174), .X(n46457) );
  inv_x4_sg U40527 ( .A(n10735), .X(n46554) );
  inv_x4_sg U40528 ( .A(n18184), .X(n46351) );
  inv_x4_sg U40529 ( .A(n41521), .X(n46342) );
  nand_x4_sg U40530 ( .A(n18836), .B(n26358), .X(n27901) );
  inv_x2_sg U40531 ( .A(n42302), .X(n42303) );
  inv_x2_sg U40532 ( .A(n42304), .X(n42305) );
  inv_x1_sg U40533 ( .A(n42093), .X(n42094) );
  inv_x1_sg U40534 ( .A(n42091), .X(n42092) );
  inv_x1_sg U40535 ( .A(n42089), .X(n42090) );
  inv_x1_sg U40536 ( .A(n42085), .X(n42086) );
  inv_x1_sg U40537 ( .A(n42083), .X(n42084) );
  inv_x1_sg U40538 ( .A(n42081), .X(n42082) );
  inv_x4_sg U40539 ( .A(n44022), .X(n46410) );
  inv_x4_sg U40540 ( .A(n44006), .X(n46273) );
  inv_x4_sg U40541 ( .A(n44010), .X(n46318) );
  inv_x4_sg U40542 ( .A(n44014), .X(n46365) );
  inv_x4_sg U40543 ( .A(n44018), .X(n46544) );
  inv_x4_sg U40544 ( .A(n44026), .X(n46455) );
  inv_x4_sg U40545 ( .A(n11163), .X(n46542) );
  inv_x4_sg U40546 ( .A(n12724), .X(n46498) );
  inv_x4_sg U40547 ( .A(n15057), .X(n46430) );
  inv_x4_sg U40548 ( .A(n16623), .X(n46386) );
  inv_x4_sg U40549 ( .A(n44030), .X(n46522) );
  inv_x4_sg U40550 ( .A(n13622), .X(n46472) );
  inv_x4_sg U40551 ( .A(n15956), .X(n46403) );
  inv_x4_sg U40552 ( .A(n12061), .X(n46515) );
  inv_x4_sg U40553 ( .A(n16700), .X(n46380) );
  inv_x4_sg U40554 ( .A(n15134), .X(n46424) );
  inv_x4_sg U40555 ( .A(n13595), .X(n46470) );
  inv_x4_sg U40556 ( .A(n12801), .X(n46492) );
  inv_x4_sg U40557 ( .A(n14356), .X(n46448) );
  inv_x4_sg U40558 ( .A(n43265), .X(n46581) );
  inv_x4_sg U40559 ( .A(n18246), .X(n46336) );
  inv_x4_sg U40560 ( .A(n10464), .X(n46562) );
  inv_x4_sg U40561 ( .A(n19791), .X(n46292) );
  inv_x4_sg U40562 ( .A(n21336), .X(n46247) );
  inv_x4_sg U40563 ( .A(n18267), .X(n46334) );
  inv_x4_sg U40564 ( .A(n14382), .X(n46444) );
  inv_x4_sg U40565 ( .A(n19845), .X(n46290) );
  inv_x4_sg U40566 ( .A(n21390), .X(n46245) );
  inv_x4_sg U40567 ( .A(n14410), .X(n46446) );
  inv_x4_sg U40568 ( .A(n15938), .X(n46401) );
  inv_x4_sg U40569 ( .A(n18301), .X(n46330) );
  inv_x4_sg U40570 ( .A(n12070), .X(n46511) );
  inv_x4_sg U40571 ( .A(n15965), .X(n46399) );
  inv_x4_sg U40572 ( .A(n11290), .X(n46534) );
  inv_x4_sg U40573 ( .A(n12851), .X(n46490) );
  inv_x4_sg U40574 ( .A(n15184), .X(n46422) );
  inv_x4_sg U40575 ( .A(n16750), .X(n46378) );
  inv_x4_sg U40576 ( .A(n13631), .X(n46466) );
  inv_x4_sg U40577 ( .A(n15728), .X(n46412) );
  inv_x4_sg U40578 ( .A(n11833), .X(n46524) );
  inv_x4_sg U40579 ( .A(n21362), .X(n46243) );
  inv_x4_sg U40580 ( .A(n19817), .X(n46288) );
  inv_x4_sg U40581 ( .A(n10490), .X(n46560) );
  inv_x4_sg U40582 ( .A(n20521), .X(n46279) );
  inv_x4_sg U40583 ( .A(n18977), .X(n46324) );
  inv_x4_sg U40584 ( .A(n17432), .X(n46371) );
  inv_x4_sg U40585 ( .A(n43866), .X(n46382) );
  inv_x4_sg U40586 ( .A(n43868), .X(n46426) );
  inv_x4_sg U40587 ( .A(n43870), .X(n46494) );
  inv_x4_sg U40588 ( .A(n43813), .X(n46538) );
  inv_x4_sg U40589 ( .A(n43811), .X(n46332) );
  inv_x4_sg U40590 ( .A(n14295), .X(n46461) );
  inv_x2_sg U40591 ( .A(n41730), .X(n41731) );
  inv_x2_sg U40592 ( .A(n42320), .X(n42321) );
  inv_x2_sg U40593 ( .A(n42318), .X(n42319) );
  inv_x2_sg U40594 ( .A(n42316), .X(n42317) );
  inv_x2_sg U40595 ( .A(n42314), .X(n42315) );
  inv_x2_sg U40596 ( .A(n41728), .X(n41729) );
  inv_x2_sg U40597 ( .A(n42308), .X(n42309) );
  inv_x2_sg U40598 ( .A(n42306), .X(n42307) );
  inv_x4_sg U40599 ( .A(n43860), .X(n46265) );
  inv_x4_sg U40600 ( .A(n43862), .X(n46310) );
  inv_x4_sg U40601 ( .A(n43864), .X(n46357) );
  inv_x4_sg U40602 ( .A(n44000), .X(n46267) );
  inv_x4_sg U40603 ( .A(n44002), .X(n46312) );
  inv_x4_sg U40604 ( .A(n44004), .X(n46359) );
  inv_x2_sg U40605 ( .A(n43230), .X(n43231) );
  inv_x2_sg U40606 ( .A(n43228), .X(n43229) );
  inv_x2_sg U40607 ( .A(n43226), .X(n43227) );
  inv_x2_sg U40608 ( .A(n43224), .X(n43225) );
  inv_x1_sg U40609 ( .A(n42119), .X(n42120) );
  inv_x1_sg U40610 ( .A(n40541), .X(n43100) );
  inv_x1_sg U40611 ( .A(n40543), .X(n42111) );
  inv_x1_sg U40612 ( .A(n40551), .X(n42121) );
  inv_x1_sg U40613 ( .A(n40554), .X(n42071) );
  inv_x1_sg U40614 ( .A(n40544), .X(n42109) );
  inv_x1_sg U40615 ( .A(n40546), .X(n42107) );
  inv_x1_sg U40616 ( .A(n40552), .X(n42103) );
  inv_x1_sg U40617 ( .A(n40555), .X(n42101) );
  inv_x1_sg U40618 ( .A(n40557), .X(n42117) );
  inv_x1_sg U40619 ( .A(n40559), .X(n42115) );
  inv_x1_sg U40620 ( .A(n40560), .X(n42113) );
  inv_x1_sg U40621 ( .A(n42079), .X(n42080) );
  inv_x1_sg U40622 ( .A(n40537), .X(n42123) );
  inv_x1_sg U40623 ( .A(n42087), .X(n42088) );
  inv_x1_sg U40624 ( .A(n40531), .X(n42135) );
  inv_x1_sg U40625 ( .A(n40548), .X(n42105) );
  inv_x1_sg U40626 ( .A(n42069), .X(n42070) );
  inv_x1_sg U40627 ( .A(n40533), .X(n42131) );
  inv_x1_sg U40628 ( .A(n40534), .X(n42129) );
  inv_x1_sg U40629 ( .A(n40535), .X(n42127) );
  inv_x1_sg U40630 ( .A(n40536), .X(n42125) );
  inv_x1_sg U40631 ( .A(n40532), .X(n42133) );
  inv_x1_sg U40632 ( .A(n40558), .X(n42099) );
  inv_x1_sg U40633 ( .A(n42097), .X(n42098) );
  inv_x1_sg U40634 ( .A(n42095), .X(n42096) );
  inv_x1_sg U40635 ( .A(n42077), .X(n42078) );
  inv_x1_sg U40636 ( .A(n40550), .X(n42075) );
  inv_x1_sg U40637 ( .A(n42073), .X(n42074) );
  inv_x1_sg U40638 ( .A(n42067), .X(n42068) );
  inv_x1_sg U40639 ( .A(n42061), .X(n42062) );
  inv_x1_sg U40640 ( .A(n42059), .X(n42060) );
  inv_x1_sg U40641 ( .A(n42057), .X(n42058) );
  inv_x1_sg U40642 ( .A(n43098), .X(n43099) );
  inv_x1_sg U40643 ( .A(n43096), .X(n43097) );
  inv_x1_sg U40644 ( .A(n41865), .X(n41866) );
  inv_x1_sg U40645 ( .A(n41867), .X(n41868) );
  inv_x1_sg U40646 ( .A(n42600), .X(n42601) );
  inv_x1_sg U40647 ( .A(n43140), .X(n43141) );
  inv_x1_sg U40648 ( .A(n42053), .X(n42054) );
  inv_x4_sg U40649 ( .A(n41711), .X(n46338) );
  inv_x4_sg U40650 ( .A(n21487), .X(n46239) );
  inv_x4_sg U40651 ( .A(n19942), .X(n46284) );
  inv_x4_sg U40652 ( .A(n18397), .X(n46328) );
  inv_x2_sg U40653 ( .A(n41557), .X(n41558) );
  inv_x2_sg U40654 ( .A(n41559), .X(n41560) );
  inv_x2_sg U40655 ( .A(n41561), .X(n41562) );
  inv_x2_sg U40656 ( .A(n41563), .X(n41564) );
  inv_x2_sg U40657 ( .A(n41565), .X(n41566) );
  inv_x2_sg U40658 ( .A(n41567), .X(n41568) );
  inv_x2_sg U40659 ( .A(n41262), .X(n41263) );
  inv_x2_sg U40660 ( .A(n41264), .X(n41265) );
  inv_x2_sg U40661 ( .A(n41266), .X(n41267) );
  inv_x2_sg U40662 ( .A(n41569), .X(n41570) );
  inv_x2_sg U40663 ( .A(n41268), .X(n41269) );
  inv_x2_sg U40664 ( .A(n41270), .X(n41271) );
  inv_x2_sg U40665 ( .A(n41272), .X(n41273) );
  inv_x2_sg U40666 ( .A(n41274), .X(n41275) );
  inv_x2_sg U40667 ( .A(n41260), .X(n41261) );
  inv_x2_sg U40668 ( .A(n43170), .X(n43171) );
  inv_x4_sg U40669 ( .A(n45300), .X(n45301) );
  inv_x4_sg U40670 ( .A(n45292), .X(n45293) );
  inv_x4_sg U40671 ( .A(n45272), .X(n45273) );
  inv_x4_sg U40672 ( .A(n45276), .X(n45277) );
  inv_x4_sg U40673 ( .A(n45278), .X(n45279) );
  inv_x4_sg U40674 ( .A(n45282), .X(n45283) );
  inv_x4_sg U40675 ( .A(n45326), .X(n45327) );
  inv_x2_sg U40676 ( .A(n41611), .X(n41612) );
  inv_x2_sg U40677 ( .A(n41615), .X(n41616) );
  inv_x2_sg U40678 ( .A(n41943), .X(n41944) );
  inv_x2_sg U40679 ( .A(n41945), .X(n41946) );
  inv_x2_sg U40680 ( .A(n41947), .X(n41948) );
  inv_x2_sg U40681 ( .A(n41949), .X(n41950) );
  inv_x2_sg U40682 ( .A(n41951), .X(n41952) );
  inv_x2_sg U40683 ( .A(n41953), .X(n41954) );
  inv_x4_sg U40684 ( .A(n45270), .X(n45271) );
  inv_x4_sg U40685 ( .A(n45284), .X(n45285) );
  inv_x4_sg U40686 ( .A(n45308), .X(n45309) );
  inv_x4_sg U40687 ( .A(n45274), .X(n45275) );
  inv_x4_sg U40688 ( .A(n45280), .X(n45281) );
  inv_x4_sg U40689 ( .A(n45286), .X(n45287) );
  inv_x4_sg U40690 ( .A(n45288), .X(n45289) );
  inv_x4_sg U40691 ( .A(n45290), .X(n45291) );
  inv_x4_sg U40692 ( .A(n45240), .X(n45241) );
  inv_x4_sg U40693 ( .A(n45294), .X(n45295) );
  inv_x4_sg U40694 ( .A(n45296), .X(n45297) );
  inv_x4_sg U40695 ( .A(n45298), .X(n45299) );
  inv_x4_sg U40696 ( .A(n45302), .X(n45303) );
  inv_x4_sg U40697 ( .A(n45304), .X(n45305) );
  inv_x4_sg U40698 ( .A(n45306), .X(n45307) );
  inv_x4_sg U40699 ( .A(n45310), .X(n45311) );
  inv_x4_sg U40700 ( .A(n45312), .X(n45313) );
  inv_x4_sg U40701 ( .A(n45314), .X(n45315) );
  inv_x4_sg U40702 ( .A(n45316), .X(n45317) );
  inv_x4_sg U40703 ( .A(n45318), .X(n45319) );
  inv_x4_sg U40704 ( .A(n45320), .X(n45321) );
  inv_x4_sg U40705 ( .A(n45322), .X(n45323) );
  inv_x4_sg U40706 ( .A(n45324), .X(n45325) );
  inv_x4_sg U40707 ( .A(n10615), .X(n46556) );
  inv_x1_sg U40708 ( .A(n41161), .X(n41162) );
  inv_x2_sg U40709 ( .A(n55461), .X(n46606) );
  inv_x2_sg U40710 ( .A(n43172), .X(n43173) );
  inv_x2_sg U40711 ( .A(n40526), .X(n42299) );
  inv_x2_sg U40712 ( .A(n40527), .X(n42296) );
  inv_x2_sg U40713 ( .A(n40528), .X(n42293) );
  inv_x2_sg U40714 ( .A(n40529), .X(n42290) );
  inv_x2_sg U40715 ( .A(n40530), .X(n42287) );
  inv_x2_sg U40716 ( .A(n42398), .X(n42399) );
  inv_x2_sg U40717 ( .A(n43308), .X(n43309) );
  inv_x2_sg U40718 ( .A(n43344), .X(n43345) );
  inv_x2_sg U40719 ( .A(n42434), .X(n42435) );
  inv_x2_sg U40720 ( .A(n42432), .X(n42433) );
  inv_x2_sg U40721 ( .A(n42430), .X(n42431) );
  inv_x2_sg U40722 ( .A(n43276), .X(n43277) );
  inv_x2_sg U40723 ( .A(n42378), .X(n42379) );
  inv_x2_sg U40724 ( .A(n43274), .X(n43275) );
  inv_x2_sg U40725 ( .A(n43272), .X(n43273) );
  inv_x2_sg U40726 ( .A(n43294), .X(n43295) );
  inv_x2_sg U40727 ( .A(n43270), .X(n43271) );
  inv_x2_sg U40728 ( .A(n43266), .X(n43267) );
  inv_x2_sg U40729 ( .A(n43268), .X(n43269) );
  inv_x2_sg U40730 ( .A(n42428), .X(n42429) );
  inv_x2_sg U40731 ( .A(n42426), .X(n42427) );
  inv_x2_sg U40732 ( .A(n43292), .X(n43293) );
  inv_x2_sg U40733 ( .A(n42376), .X(n42377) );
  inv_x2_sg U40734 ( .A(n43290), .X(n43291) );
  inv_x2_sg U40735 ( .A(n42374), .X(n42375) );
  inv_x2_sg U40736 ( .A(n43288), .X(n43289) );
  inv_x2_sg U40737 ( .A(n42372), .X(n42373) );
  inv_x2_sg U40738 ( .A(n43302), .X(n43303) );
  inv_x2_sg U40739 ( .A(n40542), .X(n43342) );
  inv_x2_sg U40740 ( .A(n40566), .X(n42382) );
  inv_x2_sg U40741 ( .A(n40567), .X(n42384) );
  inv_x2_sg U40742 ( .A(n40568), .X(n42392) );
  inv_x2_sg U40743 ( .A(n40569), .X(n42380) );
  inv_x2_sg U40744 ( .A(n40570), .X(n42390) );
  inv_x2_sg U40745 ( .A(n40571), .X(n43300) );
  inv_x2_sg U40746 ( .A(n40572), .X(n42388) );
  inv_x2_sg U40747 ( .A(n40573), .X(n43298) );
  inv_x2_sg U40748 ( .A(n40574), .X(n42386) );
  inv_x2_sg U40749 ( .A(n40575), .X(n43296) );
  inv_x2_sg U40750 ( .A(n40545), .X(n43286) );
  inv_x2_sg U40751 ( .A(n40547), .X(n43284) );
  inv_x2_sg U40752 ( .A(n40549), .X(n43282) );
  inv_x2_sg U40753 ( .A(n40553), .X(n43280) );
  inv_x2_sg U40754 ( .A(n40556), .X(n43278) );
  inv_x2_sg U40755 ( .A(n43310), .X(n43311) );
  inv_x2_sg U40756 ( .A(n43334), .X(n43335) );
  inv_x2_sg U40757 ( .A(n43330), .X(n43331) );
  inv_x2_sg U40758 ( .A(n43326), .X(n43327) );
  inv_x2_sg U40759 ( .A(n43304), .X(n43305) );
  inv_x2_sg U40760 ( .A(n43338), .X(n43339) );
  inv_x2_sg U40761 ( .A(n43314), .X(n43315) );
  inv_x2_sg U40762 ( .A(n43322), .X(n43323) );
  inv_x2_sg U40763 ( .A(n43318), .X(n43319) );
  inv_x4_sg U40764 ( .A(n44320), .X(n44321) );
  inv_x2_sg U40765 ( .A(n41609), .X(n41610) );
  inv_x2_sg U40766 ( .A(n41613), .X(n41614) );
  inv_x2_sg U40767 ( .A(n41605), .X(n41606) );
  inv_x2_sg U40768 ( .A(n41607), .X(n41608) );
  inv_x2_sg U40769 ( .A(n41603), .X(n41604) );
  nor_x2_sg U40770 ( .A(n40890), .B(n10264), .X(n10262) );
  nor_x2_sg U40771 ( .A(n40892), .B(n25371), .X(n25369) );
  inv_x1_sg U40772 ( .A(n10284), .X(n40869) );
  inv_x2_sg U40773 ( .A(n40869), .X(n40870) );
  inv_x1_sg U40774 ( .A(n13242), .X(n40871) );
  inv_x2_sg U40775 ( .A(n40871), .X(n40872) );
  inv_x1_sg U40776 ( .A(n14022), .X(n40873) );
  inv_x2_sg U40777 ( .A(n40873), .X(n40874) );
  inv_x1_sg U40778 ( .A(n15575), .X(n40875) );
  inv_x2_sg U40779 ( .A(n40875), .X(n40876) );
  inv_x1_sg U40780 ( .A(n17141), .X(n40877) );
  inv_x2_sg U40781 ( .A(n40877), .X(n40878) );
  inv_x1_sg U40782 ( .A(n12585), .X(n40879) );
  inv_x2_sg U40783 ( .A(n40879), .X(n40880) );
  inv_x1_sg U40784 ( .A(n21934), .X(n40881) );
  inv_x2_sg U40785 ( .A(n40881), .X(n40882) );
  inv_x1_sg U40786 ( .A(n29584), .X(n40883) );
  inv_x2_sg U40787 ( .A(n40883), .X(n40884) );
  inv_x1_sg U40788 ( .A(n16356), .X(n40885) );
  inv_x2_sg U40789 ( .A(n40885), .X(n40886) );
  inv_x1_sg U40790 ( .A(n12461), .X(n40887) );
  inv_x2_sg U40791 ( .A(n40887), .X(n40888) );
  inv_x1_sg U40792 ( .A(n10263), .X(n40889) );
  inv_x2_sg U40793 ( .A(n40889), .X(n40890) );
  inv_x1_sg U40794 ( .A(n25370), .X(n40891) );
  inv_x2_sg U40795 ( .A(n40891), .X(n40892) );
  inv_x1_sg U40796 ( .A(n18806), .X(n40893) );
  inv_x1_sg U40797 ( .A(n24331), .X(n40894) );
  inv_x1_sg U40798 ( .A(n31997), .X(n40895) );
  inv_x1_sg U40799 ( .A(n24344), .X(n40896) );
  inv_x1_sg U40800 ( .A(n32010), .X(n40897) );
  inv_x1_sg U40801 ( .A(n22778), .X(n40898) );
  inv_x1_sg U40802 ( .A(n30444), .X(n40899) );
  inv_x1_sg U40803 ( .A(n22174), .X(n40900) );
  inv_x1_sg U40804 ( .A(n29839), .X(n40901) );
  inv_x1_sg U40805 ( .A(n22802), .X(n40902) );
  inv_x1_sg U40806 ( .A(n30468), .X(n40903) );
  inv_x1_sg U40807 ( .A(n24349), .X(n40904) );
  inv_x1_sg U40808 ( .A(n32015), .X(n40905) );
  inv_x1_sg U40809 ( .A(n24459), .X(n40906) );
  inv_x1_sg U40810 ( .A(n32125), .X(n40907) );
  inv_x1_sg U40811 ( .A(reg_model), .X(n40908) );
  inv_x2_sg U40812 ( .A(n40908), .X(n40909) );
  inv_x1_sg U40813 ( .A(\reg_yHat[0][0] ), .X(n40910) );
  inv_x2_sg U40814 ( .A(n40910), .X(n40911) );
  inv_x1_sg U40815 ( .A(\reg_yHat[0][2] ), .X(n40912) );
  inv_x2_sg U40816 ( .A(n40912), .X(n40913) );
  inv_x1_sg U40817 ( .A(\reg_yHat[0][4] ), .X(n40914) );
  inv_x2_sg U40818 ( .A(n40914), .X(n40915) );
  inv_x1_sg U40819 ( .A(\reg_yHat[0][5] ), .X(n40916) );
  inv_x2_sg U40820 ( .A(n40916), .X(n40917) );
  inv_x1_sg U40821 ( .A(\reg_yHat[0][7] ), .X(n40918) );
  inv_x2_sg U40822 ( .A(n40918), .X(n40919) );
  inv_x1_sg U40823 ( .A(\reg_yHat[0][18] ), .X(n40920) );
  inv_x2_sg U40824 ( .A(n40920), .X(n40921) );
  inv_x1_sg U40825 ( .A(\reg_yHat[1][0] ), .X(n40922) );
  inv_x2_sg U40826 ( .A(n40922), .X(n40923) );
  inv_x1_sg U40827 ( .A(\reg_yHat[1][2] ), .X(n40924) );
  inv_x2_sg U40828 ( .A(n40924), .X(n40925) );
  inv_x1_sg U40829 ( .A(\reg_yHat[1][18] ), .X(n40926) );
  inv_x2_sg U40830 ( .A(n40926), .X(n40927) );
  inv_x1_sg U40831 ( .A(\reg_yHat[2][0] ), .X(n40928) );
  inv_x2_sg U40832 ( .A(n40928), .X(n40929) );
  inv_x1_sg U40833 ( .A(\reg_yHat[2][2] ), .X(n40930) );
  inv_x2_sg U40834 ( .A(n40930), .X(n40931) );
  inv_x1_sg U40835 ( .A(\reg_yHat[2][4] ), .X(n40932) );
  inv_x2_sg U40836 ( .A(n40932), .X(n40933) );
  inv_x1_sg U40837 ( .A(\reg_yHat[2][5] ), .X(n40934) );
  inv_x2_sg U40838 ( .A(n40934), .X(n40935) );
  inv_x1_sg U40839 ( .A(\reg_yHat[2][7] ), .X(n40936) );
  inv_x2_sg U40840 ( .A(n40936), .X(n40937) );
  inv_x1_sg U40841 ( .A(\reg_yHat[2][18] ), .X(n40938) );
  inv_x2_sg U40842 ( .A(n40938), .X(n40939) );
  inv_x1_sg U40843 ( .A(\reg_yHat[3][0] ), .X(n40940) );
  inv_x2_sg U40844 ( .A(n40940), .X(n40941) );
  inv_x1_sg U40845 ( .A(\reg_yHat[3][2] ), .X(n40942) );
  inv_x2_sg U40846 ( .A(n40942), .X(n40943) );
  inv_x1_sg U40847 ( .A(\reg_yHat[3][18] ), .X(n40944) );
  inv_x2_sg U40848 ( .A(n40944), .X(n40945) );
  inv_x1_sg U40849 ( .A(\reg_yHat[4][2] ), .X(n40946) );
  inv_x2_sg U40850 ( .A(n40946), .X(n40947) );
  inv_x1_sg U40851 ( .A(\reg_yHat[4][4] ), .X(n40948) );
  inv_x2_sg U40852 ( .A(n40948), .X(n40949) );
  inv_x1_sg U40853 ( .A(\reg_yHat[4][5] ), .X(n40950) );
  inv_x2_sg U40854 ( .A(n40950), .X(n40951) );
  inv_x1_sg U40855 ( .A(\reg_yHat[4][7] ), .X(n40952) );
  inv_x2_sg U40856 ( .A(n40952), .X(n40953) );
  inv_x1_sg U40857 ( .A(\reg_yHat[4][18] ), .X(n40954) );
  inv_x2_sg U40858 ( .A(n40954), .X(n40955) );
  inv_x1_sg U40859 ( .A(\reg_yHat[5][0] ), .X(n40956) );
  inv_x2_sg U40860 ( .A(n40956), .X(n40957) );
  inv_x1_sg U40861 ( .A(\reg_yHat[5][2] ), .X(n40958) );
  inv_x2_sg U40862 ( .A(n40958), .X(n40959) );
  inv_x1_sg U40863 ( .A(\reg_yHat[5][4] ), .X(n40960) );
  inv_x2_sg U40864 ( .A(n40960), .X(n40961) );
  inv_x1_sg U40865 ( .A(\reg_yHat[5][5] ), .X(n40962) );
  inv_x2_sg U40866 ( .A(n40962), .X(n40963) );
  inv_x1_sg U40867 ( .A(\reg_yHat[5][6] ), .X(n40964) );
  inv_x2_sg U40868 ( .A(n40964), .X(n40965) );
  inv_x1_sg U40869 ( .A(\reg_yHat[5][18] ), .X(n40966) );
  inv_x2_sg U40870 ( .A(n40966), .X(n40967) );
  inv_x1_sg U40871 ( .A(\reg_yHat[6][0] ), .X(n40968) );
  inv_x2_sg U40872 ( .A(n40968), .X(n40969) );
  inv_x1_sg U40873 ( .A(\reg_yHat[6][2] ), .X(n40970) );
  inv_x2_sg U40874 ( .A(n40970), .X(n40971) );
  inv_x1_sg U40875 ( .A(\reg_yHat[6][18] ), .X(n40972) );
  inv_x2_sg U40876 ( .A(n40972), .X(n40973) );
  inv_x1_sg U40877 ( .A(\reg_yHat[7][0] ), .X(n40974) );
  inv_x2_sg U40878 ( .A(n40974), .X(n40975) );
  inv_x1_sg U40879 ( .A(\reg_yHat[7][2] ), .X(n40976) );
  inv_x2_sg U40880 ( .A(n40976), .X(n40977) );
  inv_x1_sg U40881 ( .A(\reg_yHat[7][4] ), .X(n40978) );
  inv_x2_sg U40882 ( .A(n40978), .X(n40979) );
  inv_x1_sg U40883 ( .A(\reg_yHat[7][5] ), .X(n40980) );
  inv_x2_sg U40884 ( .A(n40980), .X(n40981) );
  inv_x1_sg U40885 ( .A(\reg_yHat[7][7] ), .X(n40982) );
  inv_x2_sg U40886 ( .A(n40982), .X(n40983) );
  inv_x1_sg U40887 ( .A(\reg_yHat[7][18] ), .X(n40984) );
  inv_x2_sg U40888 ( .A(n40984), .X(n40985) );
  inv_x1_sg U40889 ( .A(\reg_yHat[8][0] ), .X(n40986) );
  inv_x2_sg U40890 ( .A(n40986), .X(n40987) );
  inv_x1_sg U40891 ( .A(\reg_yHat[8][2] ), .X(n40988) );
  inv_x2_sg U40892 ( .A(n40988), .X(n40989) );
  inv_x1_sg U40893 ( .A(\reg_yHat[8][18] ), .X(n40990) );
  inv_x2_sg U40894 ( .A(n40990), .X(n40991) );
  inv_x1_sg U40895 ( .A(\reg_yHat[9][0] ), .X(n40992) );
  inv_x2_sg U40896 ( .A(n40992), .X(n40993) );
  inv_x1_sg U40897 ( .A(\reg_yHat[9][2] ), .X(n40994) );
  inv_x2_sg U40898 ( .A(n40994), .X(n40995) );
  inv_x1_sg U40899 ( .A(\reg_yHat[9][18] ), .X(n40996) );
  inv_x2_sg U40900 ( .A(n40996), .X(n40997) );
  inv_x1_sg U40901 ( .A(\reg_yHat[10][0] ), .X(n40998) );
  inv_x2_sg U40902 ( .A(n40998), .X(n40999) );
  inv_x1_sg U40903 ( .A(\reg_yHat[10][2] ), .X(n41000) );
  inv_x2_sg U40904 ( .A(n41000), .X(n41001) );
  inv_x1_sg U40905 ( .A(\reg_yHat[10][3] ), .X(n41002) );
  inv_x2_sg U40906 ( .A(n41002), .X(n41003) );
  inv_x1_sg U40907 ( .A(\reg_yHat[10][4] ), .X(n41004) );
  inv_x2_sg U40908 ( .A(n41004), .X(n41005) );
  inv_x1_sg U40909 ( .A(\reg_yHat[10][18] ), .X(n41006) );
  inv_x2_sg U40910 ( .A(n41006), .X(n41007) );
  inv_x1_sg U40911 ( .A(\reg_yHat[11][0] ), .X(n41008) );
  inv_x2_sg U40912 ( .A(n41008), .X(n41009) );
  inv_x1_sg U40913 ( .A(\reg_yHat[11][2] ), .X(n41010) );
  inv_x2_sg U40914 ( .A(n41010), .X(n41011) );
  inv_x1_sg U40915 ( .A(\reg_yHat[11][18] ), .X(n41012) );
  inv_x2_sg U40916 ( .A(n41012), .X(n41013) );
  inv_x1_sg U40917 ( .A(\reg_yHat[12][0] ), .X(n41014) );
  inv_x2_sg U40918 ( .A(n41014), .X(n41015) );
  inv_x1_sg U40919 ( .A(\reg_yHat[12][2] ), .X(n41016) );
  inv_x2_sg U40920 ( .A(n41016), .X(n41017) );
  inv_x1_sg U40921 ( .A(\reg_yHat[12][4] ), .X(n41018) );
  inv_x2_sg U40922 ( .A(n41018), .X(n41019) );
  inv_x1_sg U40923 ( .A(\reg_yHat[12][5] ), .X(n41020) );
  inv_x2_sg U40924 ( .A(n41020), .X(n41021) );
  inv_x1_sg U40925 ( .A(\reg_yHat[12][7] ), .X(n41022) );
  inv_x2_sg U40926 ( .A(n41022), .X(n41023) );
  inv_x1_sg U40927 ( .A(\reg_yHat[12][18] ), .X(n41024) );
  inv_x2_sg U40928 ( .A(n41024), .X(n41025) );
  inv_x1_sg U40929 ( .A(\reg_yHat[13][0] ), .X(n41026) );
  inv_x2_sg U40930 ( .A(n41026), .X(n41027) );
  inv_x1_sg U40931 ( .A(\reg_yHat[13][2] ), .X(n41028) );
  inv_x2_sg U40932 ( .A(n41028), .X(n41029) );
  inv_x1_sg U40933 ( .A(\reg_yHat[13][18] ), .X(n41030) );
  inv_x2_sg U40934 ( .A(n41030), .X(n41031) );
  inv_x1_sg U40935 ( .A(\reg_yHat[14][0] ), .X(n41032) );
  inv_x2_sg U40936 ( .A(n41032), .X(n41033) );
  inv_x1_sg U40937 ( .A(\reg_yHat[14][2] ), .X(n41034) );
  inv_x2_sg U40938 ( .A(n41034), .X(n41035) );
  inv_x1_sg U40939 ( .A(\reg_yHat[14][4] ), .X(n41036) );
  inv_x2_sg U40940 ( .A(n41036), .X(n41037) );
  inv_x1_sg U40941 ( .A(\reg_yHat[14][5] ), .X(n41038) );
  inv_x2_sg U40942 ( .A(n41038), .X(n41039) );
  inv_x1_sg U40943 ( .A(\reg_yHat[14][7] ), .X(n41040) );
  inv_x2_sg U40944 ( .A(n41040), .X(n41041) );
  inv_x1_sg U40945 ( .A(\reg_yHat[14][18] ), .X(n41042) );
  inv_x2_sg U40946 ( .A(n41042), .X(n41043) );
  inv_x1_sg U40947 ( .A(\reg_y[0][2] ), .X(n41044) );
  inv_x2_sg U40948 ( .A(n41044), .X(n41045) );
  inv_x1_sg U40949 ( .A(\reg_y[0][4] ), .X(n41046) );
  inv_x2_sg U40950 ( .A(n41046), .X(n41047) );
  inv_x1_sg U40951 ( .A(\reg_y[0][5] ), .X(n41048) );
  inv_x2_sg U40952 ( .A(n41048), .X(n41049) );
  inv_x1_sg U40953 ( .A(\reg_y[0][18] ), .X(n41050) );
  inv_x2_sg U40954 ( .A(n41050), .X(n41051) );
  inv_x1_sg U40955 ( .A(\reg_y[1][2] ), .X(n41052) );
  inv_x2_sg U40956 ( .A(n41052), .X(n41053) );
  inv_x1_sg U40957 ( .A(\reg_y[1][18] ), .X(n41054) );
  inv_x2_sg U40958 ( .A(n41054), .X(n41055) );
  inv_x1_sg U40959 ( .A(\reg_y[2][2] ), .X(n41056) );
  inv_x2_sg U40960 ( .A(n41056), .X(n41057) );
  inv_x1_sg U40961 ( .A(\reg_y[2][4] ), .X(n41058) );
  inv_x2_sg U40962 ( .A(n41058), .X(n41059) );
  inv_x1_sg U40963 ( .A(\reg_y[2][5] ), .X(n41060) );
  inv_x2_sg U40964 ( .A(n41060), .X(n41061) );
  inv_x1_sg U40965 ( .A(\reg_y[2][18] ), .X(n41062) );
  inv_x2_sg U40966 ( .A(n41062), .X(n41063) );
  inv_x1_sg U40967 ( .A(\reg_y[3][2] ), .X(n41064) );
  inv_x2_sg U40968 ( .A(n41064), .X(n41065) );
  inv_x1_sg U40969 ( .A(\reg_y[3][18] ), .X(n41066) );
  inv_x2_sg U40970 ( .A(n41066), .X(n41067) );
  inv_x1_sg U40971 ( .A(\reg_y[4][2] ), .X(n41068) );
  inv_x2_sg U40972 ( .A(n41068), .X(n41069) );
  inv_x1_sg U40973 ( .A(\reg_y[4][4] ), .X(n41070) );
  inv_x2_sg U40974 ( .A(n41070), .X(n41071) );
  inv_x1_sg U40975 ( .A(\reg_y[4][5] ), .X(n41072) );
  inv_x2_sg U40976 ( .A(n41072), .X(n41073) );
  inv_x1_sg U40977 ( .A(\reg_y[4][18] ), .X(n41074) );
  inv_x2_sg U40978 ( .A(n41074), .X(n41075) );
  inv_x1_sg U40979 ( .A(\reg_y[5][2] ), .X(n41076) );
  inv_x2_sg U40980 ( .A(n41076), .X(n41077) );
  inv_x1_sg U40981 ( .A(\reg_y[5][4] ), .X(n41078) );
  inv_x2_sg U40982 ( .A(n41078), .X(n41079) );
  inv_x1_sg U40983 ( .A(\reg_y[5][5] ), .X(n41080) );
  inv_x2_sg U40984 ( .A(n41080), .X(n41081) );
  inv_x1_sg U40985 ( .A(\reg_y[5][18] ), .X(n41082) );
  inv_x2_sg U40986 ( .A(n41082), .X(n41083) );
  inv_x1_sg U40987 ( .A(\reg_y[6][2] ), .X(n41084) );
  inv_x2_sg U40988 ( .A(n41084), .X(n41085) );
  inv_x1_sg U40989 ( .A(\reg_y[6][18] ), .X(n41086) );
  inv_x2_sg U40990 ( .A(n41086), .X(n41087) );
  inv_x1_sg U40991 ( .A(\reg_y[7][2] ), .X(n41088) );
  inv_x2_sg U40992 ( .A(n41088), .X(n41089) );
  inv_x1_sg U40993 ( .A(\reg_y[7][4] ), .X(n41090) );
  inv_x2_sg U40994 ( .A(n41090), .X(n41091) );
  inv_x1_sg U40995 ( .A(\reg_y[7][5] ), .X(n41092) );
  inv_x2_sg U40996 ( .A(n41092), .X(n41093) );
  inv_x1_sg U40997 ( .A(\reg_y[7][18] ), .X(n41094) );
  inv_x2_sg U40998 ( .A(n41094), .X(n41095) );
  inv_x1_sg U40999 ( .A(\reg_y[8][2] ), .X(n41096) );
  inv_x2_sg U41000 ( .A(n41096), .X(n41097) );
  inv_x1_sg U41001 ( .A(\reg_y[8][18] ), .X(n41098) );
  inv_x2_sg U41002 ( .A(n41098), .X(n41099) );
  inv_x1_sg U41003 ( .A(\reg_y[9][2] ), .X(n41100) );
  inv_x2_sg U41004 ( .A(n41100), .X(n41101) );
  inv_x1_sg U41005 ( .A(\reg_y[9][18] ), .X(n41102) );
  inv_x2_sg U41006 ( .A(n41102), .X(n41103) );
  inv_x1_sg U41007 ( .A(\reg_y[10][4] ), .X(n41104) );
  inv_x2_sg U41008 ( .A(n41104), .X(n41105) );
  inv_x1_sg U41009 ( .A(\reg_y[10][18] ), .X(n41106) );
  inv_x2_sg U41010 ( .A(n41106), .X(n41107) );
  inv_x1_sg U41011 ( .A(\reg_y[11][2] ), .X(n41108) );
  inv_x2_sg U41012 ( .A(n41108), .X(n41109) );
  inv_x1_sg U41013 ( .A(\reg_y[11][18] ), .X(n41110) );
  inv_x2_sg U41014 ( .A(n41110), .X(n41111) );
  inv_x1_sg U41015 ( .A(\reg_y[12][2] ), .X(n41112) );
  inv_x2_sg U41016 ( .A(n41112), .X(n41113) );
  inv_x1_sg U41017 ( .A(\reg_y[12][4] ), .X(n41114) );
  inv_x2_sg U41018 ( .A(n41114), .X(n41115) );
  inv_x1_sg U41019 ( .A(\reg_y[12][5] ), .X(n41116) );
  inv_x2_sg U41020 ( .A(n41116), .X(n41117) );
  inv_x1_sg U41021 ( .A(\reg_y[12][18] ), .X(n41118) );
  inv_x2_sg U41022 ( .A(n41118), .X(n41119) );
  inv_x1_sg U41023 ( .A(\reg_y[13][2] ), .X(n41120) );
  inv_x2_sg U41024 ( .A(n41120), .X(n41121) );
  inv_x1_sg U41025 ( .A(\reg_y[13][18] ), .X(n41122) );
  inv_x2_sg U41026 ( .A(n41122), .X(n41123) );
  inv_x1_sg U41027 ( .A(\reg_y[14][2] ), .X(n41124) );
  inv_x2_sg U41028 ( .A(n41124), .X(n41125) );
  inv_x1_sg U41029 ( .A(\reg_y[14][4] ), .X(n41126) );
  inv_x2_sg U41030 ( .A(n41126), .X(n41127) );
  inv_x1_sg U41031 ( .A(\reg_y[14][5] ), .X(n41128) );
  inv_x2_sg U41032 ( .A(n41128), .X(n41129) );
  inv_x1_sg U41033 ( .A(\reg_y[14][18] ), .X(n41130) );
  inv_x2_sg U41034 ( .A(n41130), .X(n41131) );
  inv_x1_sg U41035 ( .A(reg_num[1]), .X(n41132) );
  inv_x2_sg U41036 ( .A(n41132), .X(n41133) );
  inv_x1_sg U41037 ( .A(reg_num[2]), .X(n41134) );
  inv_x2_sg U41038 ( .A(n41134), .X(n41135) );
  inv_x1_sg U41039 ( .A(n55799), .X(n41136) );
  inv_x2_sg U41040 ( .A(n41136), .X(n41137) );
  inv_x1_sg U41041 ( .A(n55798), .X(n41138) );
  inv_x2_sg U41042 ( .A(n41138), .X(n41139) );
  inv_x8_sg U41043 ( .A(n43179), .X(n49796) );
  inv_x2_sg U41044 ( .A(n28450), .X(n54046) );
  nand_x4_sg U41045 ( .A(n41490), .B(n17123), .X(n17124) );
  nand_x4_sg U41046 ( .A(n41492), .B(n15557), .X(n15558) );
  nand_x4_sg U41047 ( .A(n41219), .B(n14004), .X(n14005) );
  nand_x4_sg U41048 ( .A(n41494), .B(n13224), .X(n13225) );
  nand_x4_sg U41049 ( .A(n41496), .B(n12443), .X(n12444) );
  nand_x4_sg U41050 ( .A(n42064), .B(n16320), .X(n15806) );
  nand_x2_sg U41051 ( .A(n49796), .B(n41667), .X(n31316) );
  inv_x8_sg U41052 ( .A(n43191), .X(n50655) );
  inv_x4_sg U41053 ( .A(n31998), .X(n41140) );
  inv_x4_sg U41054 ( .A(n24332), .X(n41141) );
  inv_x1_sg U41055 ( .A(n28386), .X(n41522) );
  nand_x2_sg U41056 ( .A(n44158), .B(n25508), .X(n25515) );
  nor_x2_sg U41057 ( .A(n28577), .B(n46209), .X(n28574) );
  nor_x2_sg U41058 ( .A(n27740), .B(n46215), .X(n27737) );
  nor_x2_sg U41059 ( .A(n27459), .B(n46217), .X(n27456) );
  nor_x2_sg U41060 ( .A(n27180), .B(n46219), .X(n27177) );
  nor_x2_sg U41061 ( .A(n26623), .B(n46223), .X(n26620) );
  nor_x2_sg U41062 ( .A(n26344), .B(n46225), .X(n26341) );
  nor_x2_sg U41063 ( .A(n26063), .B(n46227), .X(n26060) );
  nor_x2_sg U41064 ( .A(n25784), .B(n46229), .X(n25781) );
  nor_x2_sg U41065 ( .A(n25506), .B(n46231), .X(n25503) );
  nand_x4_sg U41066 ( .A(n43071), .B(n18645), .X(n18142) );
  nand_x4_sg U41067 ( .A(n41171), .B(n16615), .X(n16533) );
  nand_x4_sg U41068 ( .A(n41172), .B(n15049), .X(n14967) );
  inv_x4_sg U41069 ( .A(n41142), .X(n41143) );
  inv_x4_sg U41070 ( .A(n41144), .X(n41145) );
  inv_x4_sg U41071 ( .A(n41146), .X(n41147) );
  inv_x4_sg U41072 ( .A(n41148), .X(n41149) );
  nand_x2_sg U41073 ( .A(n50655), .B(n41677), .X(n23650) );
  nand_x4_sg U41074 ( .A(n42304), .B(n18105), .X(n9067) );
  nand_x4_sg U41075 ( .A(n42302), .B(n10322), .X(n9039) );
  inv_x4_sg U41076 ( .A(n41150), .X(n41151) );
  inv_x4_sg U41077 ( .A(n41152), .X(n41153) );
  inv_x2_sg U41078 ( .A(n17142), .X(n41154) );
  nand_x8_sg U41079 ( .A(n17167), .B(n46388), .X(n17142) );
  inv_x1_sg U41080 ( .A(n17142), .X(n53705) );
  inv_x2_sg U41081 ( .A(n15576), .X(n41155) );
  nand_x8_sg U41082 ( .A(n15601), .B(n46432), .X(n15576) );
  inv_x1_sg U41083 ( .A(n15576), .X(n53147) );
  inv_x2_sg U41084 ( .A(n14023), .X(n41156) );
  nand_x8_sg U41085 ( .A(n14048), .B(n46478), .X(n14023) );
  inv_x1_sg U41086 ( .A(n14023), .X(n52588) );
  inv_x2_sg U41087 ( .A(n13243), .X(n41157) );
  nand_x8_sg U41088 ( .A(n13268), .B(n46500), .X(n13243) );
  inv_x1_sg U41089 ( .A(n13243), .X(n52313) );
  inv_x2_sg U41090 ( .A(n12462), .X(n41158) );
  nand_x8_sg U41091 ( .A(n12487), .B(n51819), .X(n12462) );
  inv_x1_sg U41092 ( .A(n12462), .X(n52037) );
  inv_x4_sg U41093 ( .A(n41159), .X(n41160) );
  nand_x4_sg U41094 ( .A(n41217), .B(n13433), .X(n13431) );
  inv_x8_sg U41095 ( .A(n43183), .X(n50066) );
  inv_x8_sg U41096 ( .A(n43187), .X(n50925) );
  inv_x1_sg U41097 ( .A(n17121), .X(n41714) );
  inv_x1_sg U41098 ( .A(n15555), .X(n41718) );
  inv_x1_sg U41099 ( .A(n13222), .X(n41726) );
  inv_x1_sg U41100 ( .A(n12441), .X(n43168) );
  inv_x1_sg U41101 ( .A(n17103), .X(n43279) );
  inv_x1_sg U41102 ( .A(n15537), .X(n43281) );
  inv_x1_sg U41103 ( .A(n13984), .X(n43283) );
  inv_x1_sg U41104 ( .A(n13204), .X(n43285) );
  inv_x1_sg U41105 ( .A(n12423), .X(n43287) );
  inv_x1_sg U41106 ( .A(n16306), .X(n42381) );
  inv_x1_sg U41107 ( .A(n10850), .X(n42383) );
  inv_x1_sg U41108 ( .A(n11001), .X(n42055) );
  inv_x1_sg U41109 ( .A(n21721), .X(n43297) );
  inv_x1_sg U41110 ( .A(n20176), .X(n43299) );
  inv_x1_sg U41111 ( .A(n18630), .X(n43301) );
  inv_x1_sg U41112 ( .A(n11630), .X(n42385) );
  inv_x1_sg U41113 ( .A(n14102), .X(n42269) );
  inv_x1_sg U41114 ( .A(n20952), .X(n42387) );
  inv_x1_sg U41115 ( .A(n19408), .X(n42389) );
  inv_x1_sg U41116 ( .A(n17863), .X(n42391) );
  inv_x1_sg U41117 ( .A(n14742), .X(n42393) );
  inv_x1_sg U41118 ( .A(n16801), .X(n41222) );
  inv_x1_sg U41119 ( .A(n15235), .X(n41226) );
  inv_x1_sg U41120 ( .A(n12902), .X(n41230) );
  inv_x1_sg U41121 ( .A(n28390), .X(n41234) );
  inv_x8_sg U41122 ( .A(n41589), .X(n41590) );
  inv_x8_sg U41123 ( .A(n41591), .X(n41592) );
  nor_x2_sg U41124 ( .A(n29418), .B(n46203), .X(n29415) );
  nor_x2_sg U41125 ( .A(n29136), .B(n46205), .X(n29133) );
  nor_x2_sg U41126 ( .A(n28857), .B(n46207), .X(n28854) );
  nor_x2_sg U41127 ( .A(n28299), .B(n46211), .X(n28296) );
  nor_x2_sg U41128 ( .A(n28019), .B(n46213), .X(n28016) );
  nor_x2_sg U41129 ( .A(n26900), .B(n46221), .X(n26897) );
  nor_x2_sg U41130 ( .A(n27741), .B(n27742), .X(n27740) );
  nor_x2_sg U41131 ( .A(n27743), .B(n41263), .X(n27741) );
  nor_x2_sg U41132 ( .A(n27460), .B(n27461), .X(n27459) );
  nor_x2_sg U41133 ( .A(n27462), .B(n41265), .X(n27460) );
  nor_x2_sg U41134 ( .A(n27181), .B(n27182), .X(n27180) );
  nor_x2_sg U41135 ( .A(n27183), .B(n41267), .X(n27181) );
  nor_x2_sg U41136 ( .A(n26624), .B(n26625), .X(n26623) );
  nor_x2_sg U41137 ( .A(n26626), .B(n41269), .X(n26624) );
  nor_x2_sg U41138 ( .A(n26345), .B(n26346), .X(n26344) );
  nor_x2_sg U41139 ( .A(n26347), .B(n41271), .X(n26345) );
  nor_x2_sg U41140 ( .A(n26064), .B(n26065), .X(n26063) );
  nor_x2_sg U41141 ( .A(n26066), .B(n41273), .X(n26064) );
  nor_x2_sg U41142 ( .A(n25785), .B(n25786), .X(n25784) );
  nor_x2_sg U41143 ( .A(n25787), .B(n41275), .X(n25785) );
  nor_x2_sg U41144 ( .A(n25507), .B(n25508), .X(n25506) );
  nor_x2_sg U41145 ( .A(n25509), .B(n41261), .X(n25507) );
  nor_x2_sg U41146 ( .A(n21305), .B(n21306), .X(n21304) );
  nor_x2_sg U41147 ( .A(n19760), .B(n19761), .X(n19759) );
  nand_x4_sg U41148 ( .A(n53561), .B(n16738), .X(n16732) );
  nand_x4_sg U41149 ( .A(n53003), .B(n15172), .X(n15166) );
  nand_x4_sg U41150 ( .A(n52169), .B(n12839), .X(n12833) );
  nand_x4_sg U41151 ( .A(n43055), .B(n21736), .X(n21232) );
  nand_x4_sg U41152 ( .A(n43057), .B(n20967), .X(n20459) );
  nand_x4_sg U41153 ( .A(n43063), .B(n20191), .X(n19687) );
  nand_x4_sg U41154 ( .A(n43065), .B(n19423), .X(n18915) );
  nand_x4_sg U41155 ( .A(n43073), .B(n17878), .X(n17370) );
  nand_x4_sg U41156 ( .A(n43081), .B(n14757), .X(n14251) );
  nand_x4_sg U41157 ( .A(n43093), .B(n11645), .X(n11127) );
  nand_x4_sg U41158 ( .A(n43095), .B(n10865), .X(n10360) );
  inv_x4_sg U41159 ( .A(n11767), .X(n41161) );
  nor_x1_sg U41160 ( .A(n18485), .B(n18486), .X(n18467) );
  nand_x4_sg U41161 ( .A(n41881), .B(n12716), .X(n12634) );
  nand_x4_sg U41162 ( .A(n41883), .B(n11155), .X(n11073) );
  inv_x2_sg U41163 ( .A(n50461), .X(n41163) );
  inv_x8_sg U41164 ( .A(n24121), .X(n50461) );
  inv_x2_sg U41165 ( .A(n50508), .X(n41164) );
  inv_x8_sg U41166 ( .A(n24128), .X(n50508) );
  inv_x2_sg U41167 ( .A(n49370), .X(n41165) );
  inv_x8_sg U41168 ( .A(n31752), .X(n49370) );
  inv_x2_sg U41169 ( .A(n49602), .X(n41166) );
  inv_x8_sg U41170 ( .A(n31787), .X(n49602) );
  inv_x2_sg U41171 ( .A(n49649), .X(n41167) );
  inv_x8_sg U41172 ( .A(n31794), .X(n49649) );
  inv_x2_sg U41173 ( .A(n50229), .X(n41168) );
  inv_x8_sg U41174 ( .A(n24086), .X(n50229) );
  inv_x2_sg U41175 ( .A(n50319), .X(n41169) );
  inv_x8_sg U41176 ( .A(n24339), .X(n50319) );
  inv_x2_sg U41177 ( .A(n49460), .X(n41170) );
  inv_x8_sg U41178 ( .A(n32005), .X(n49460) );
  nand_x4_sg U41179 ( .A(n18373), .B(n18379), .X(n18369) );
  nand_x4_sg U41180 ( .A(n41476), .B(n18382), .X(n18373) );
  nand_x4_sg U41181 ( .A(n20693), .B(n20699), .X(n20689) );
  nand_x4_sg U41182 ( .A(n41477), .B(n20702), .X(n20693) );
  nand_x4_sg U41183 ( .A(n19149), .B(n19155), .X(n19145) );
  nand_x4_sg U41184 ( .A(n41478), .B(n19158), .X(n19149) );
  nand_x4_sg U41185 ( .A(n17604), .B(n17610), .X(n17600) );
  nand_x4_sg U41186 ( .A(n41479), .B(n17613), .X(n17604) );
  nand_x4_sg U41187 ( .A(n14483), .B(n14489), .X(n14479) );
  nand_x4_sg U41188 ( .A(n41480), .B(n14492), .X(n14483) );
  inv_x1_sg U41189 ( .A(n16616), .X(n41171) );
  inv_x1_sg U41190 ( .A(n16616), .X(n53514) );
  inv_x1_sg U41191 ( .A(n15050), .X(n41172) );
  inv_x1_sg U41192 ( .A(n15050), .X(n52956) );
  inv_x4_sg U41193 ( .A(n41178), .X(n41179) );
  inv_x4_sg U41194 ( .A(n41180), .X(n41181) );
  inv_x4_sg U41195 ( .A(n41182), .X(n41183) );
  inv_x4_sg U41196 ( .A(n41184), .X(n41185) );
  inv_x4_sg U41197 ( .A(n41186), .X(n41187) );
  inv_x4_sg U41198 ( .A(n41188), .X(n41189) );
  nand_x2_sg U41199 ( .A(n50066), .B(n42949), .X(n30452) );
  nand_x2_sg U41200 ( .A(n50925), .B(n43013), .X(n22786) );
  nand_x4_sg U41201 ( .A(n21191), .B(n55286), .X(n9117) );
  nand_x4_sg U41202 ( .A(n41453), .B(n21193), .X(n21191) );
  nand_x4_sg U41203 ( .A(n20418), .B(n55007), .X(n9142) );
  nand_x4_sg U41204 ( .A(n41469), .B(n20420), .X(n20418) );
  nand_x4_sg U41205 ( .A(n19646), .B(n54718), .X(n9183) );
  nand_x4_sg U41206 ( .A(n41455), .B(n19648), .X(n19646) );
  nand_x4_sg U41207 ( .A(n18874), .B(n54439), .X(n9218) );
  nand_x4_sg U41208 ( .A(n41471), .B(n18876), .X(n18874) );
  nand_x4_sg U41209 ( .A(n17329), .B(n53874), .X(n9256) );
  nand_x4_sg U41210 ( .A(n41473), .B(n17331), .X(n17329) );
  nand_x4_sg U41211 ( .A(n14210), .B(n52754), .X(n8952) );
  nand_x4_sg U41212 ( .A(n41475), .B(n14212), .X(n14210) );
  inv_x4_sg U41213 ( .A(n41190), .X(n41191) );
  inv_x4_sg U41214 ( .A(n41192), .X(n41193) );
  inv_x4_sg U41215 ( .A(n41194), .X(n41195) );
  inv_x4_sg U41216 ( .A(n41196), .X(n41197) );
  inv_x4_sg U41217 ( .A(n41198), .X(n41199) );
  inv_x4_sg U41218 ( .A(n41200), .X(n41201) );
  inv_x4_sg U41219 ( .A(n41202), .X(n41203) );
  inv_x4_sg U41220 ( .A(n41204), .X(n41205) );
  inv_x4_sg U41221 ( .A(n41206), .X(n41207) );
  inv_x4_sg U41222 ( .A(n41208), .X(n41209) );
  inv_x4_sg U41223 ( .A(n41210), .X(n41211) );
  nor_x4_sg U41224 ( .A(n13980), .B(n46475), .X(n13992) );
  nor_x4_sg U41225 ( .A(n18654), .B(n46340), .X(n18652) );
  inv_x4_sg U41226 ( .A(n30204), .X(n41212) );
  inv_x4_sg U41227 ( .A(n22538), .X(n41213) );
  nor_x4_sg U41228 ( .A(n11515), .B(n46541), .X(n11802) );
  nand_x4_sg U41229 ( .A(n15764), .B(n53303), .X(n9351) );
  nand_x4_sg U41230 ( .A(n41449), .B(n15766), .X(n15764) );
  nand_x4_sg U41231 ( .A(n10318), .B(n51364), .X(n9041) );
  nand_x4_sg U41232 ( .A(n41451), .B(n10320), .X(n10318) );
  nand_x4_sg U41233 ( .A(n18101), .B(n54153), .X(n9075) );
  nand_x4_sg U41234 ( .A(n41457), .B(n18103), .X(n18101) );
  nand_x4_sg U41235 ( .A(n16546), .B(n53583), .X(n9294) );
  nand_x4_sg U41236 ( .A(n41459), .B(n16548), .X(n16546) );
  nand_x4_sg U41237 ( .A(n14980), .B(n53025), .X(n8977) );
  nand_x4_sg U41238 ( .A(n41461), .B(n14982), .X(n14980) );
  nand_x4_sg U41239 ( .A(n12647), .B(n52191), .X(n8838) );
  nand_x4_sg U41240 ( .A(n41463), .B(n12649), .X(n12647) );
  nand_x4_sg U41241 ( .A(n11869), .B(n51916), .X(n8913) );
  nand_x4_sg U41242 ( .A(n41465), .B(n11871), .X(n11869) );
  nand_x4_sg U41243 ( .A(n11086), .B(n51635), .X(n8876) );
  nand_x4_sg U41244 ( .A(n41467), .B(n11088), .X(n11086) );
  inv_x4_sg U41245 ( .A(n41214), .X(n41215) );
  inv_x4_sg U41246 ( .A(n41216), .X(n41217) );
  inv_x2_sg U41247 ( .A(n30173), .X(n41847) );
  inv_x2_sg U41248 ( .A(n29643), .X(n41849) );
  inv_x2_sg U41249 ( .A(n22507), .X(n41851) );
  inv_x2_sg U41250 ( .A(n21978), .X(n41853) );
  inv_x1_sg U41251 ( .A(n31319), .X(n41668) );
  inv_x2_sg U41252 ( .A(n21377), .X(n41831) );
  inv_x2_sg U41253 ( .A(n19832), .X(n41835) );
  inv_x2_sg U41254 ( .A(n18287), .X(n41545) );
  inv_x1_sg U41255 ( .A(n17118), .X(n41684) );
  inv_x1_sg U41256 ( .A(n15552), .X(n41688) );
  inv_x1_sg U41257 ( .A(n13999), .X(n41692) );
  inv_x1_sg U41258 ( .A(n13219), .X(n41696) );
  inv_x1_sg U41259 ( .A(n12438), .X(n41700) );
  inv_x1_sg U41260 ( .A(n16332), .X(n42065) );
  inv_x1_sg U41261 ( .A(n17221), .X(n42261) );
  inv_x1_sg U41262 ( .A(n15655), .X(n42265) );
  inv_x1_sg U41263 ( .A(n13322), .X(n42273) );
  inv_x1_sg U41264 ( .A(n12541), .X(n42277) );
  inv_x1_sg U41265 ( .A(n16016), .X(n41499) );
  inv_x1_sg U41266 ( .A(n13682), .X(n41503) );
  inv_x1_sg U41267 ( .A(n12121), .X(n41507) );
  inv_x1_sg U41268 ( .A(n11341), .X(n41511) );
  inv_x4_sg U41269 ( .A(n41218), .X(n41219) );
  nor_x2_sg U41270 ( .A(n14101), .B(n42268), .X(n14099) );
  inv_x4_sg U41271 ( .A(n41220), .X(n41221) );
  inv_x2_sg U41272 ( .A(n41222), .X(n41223) );
  inv_x4_sg U41273 ( .A(n41224), .X(n41225) );
  inv_x2_sg U41274 ( .A(n41226), .X(n41227) );
  inv_x4_sg U41275 ( .A(n41228), .X(n41229) );
  inv_x2_sg U41276 ( .A(n41230), .X(n41231) );
  inv_x4_sg U41277 ( .A(n41232), .X(n41233) );
  inv_x2_sg U41278 ( .A(n41234), .X(n41235) );
  inv_x4_sg U41279 ( .A(n41236), .X(n41237) );
  inv_x4_sg U41280 ( .A(n41238), .X(n41239) );
  inv_x4_sg U41281 ( .A(n41240), .X(n41241) );
  inv_x4_sg U41282 ( .A(n41242), .X(n41243) );
  inv_x4_sg U41283 ( .A(n41244), .X(n41245) );
  inv_x4_sg U41284 ( .A(n41246), .X(n41247) );
  inv_x4_sg U41285 ( .A(n41248), .X(n41249) );
  inv_x4_sg U41286 ( .A(n41250), .X(n41251) );
  inv_x4_sg U41287 ( .A(n41252), .X(n41253) );
  inv_x4_sg U41288 ( .A(n41254), .X(n41255) );
  inv_x4_sg U41289 ( .A(n41256), .X(n41257) );
  inv_x4_sg U41290 ( .A(n41258), .X(n41259) );
  nor_x4_sg U41291 ( .A(n21197), .B(n41744), .X(n21203) );
  nor_x4_sg U41292 ( .A(n19652), .B(n41746), .X(n19658) );
  nor_x4_sg U41293 ( .A(n20424), .B(n41772), .X(n20430) );
  nor_x4_sg U41294 ( .A(n18880), .B(n41774), .X(n18886) );
  nor_x4_sg U41295 ( .A(n17335), .B(n41776), .X(n17341) );
  nor_x4_sg U41296 ( .A(n14216), .B(n41778), .X(n14222) );
  inv_x8_sg U41297 ( .A(n32087), .X(n49413) );
  nor_x8_sg U41298 ( .A(n41590), .B(n32089), .X(n32086) );
  nand_x4_sg U41299 ( .A(n41590), .B(n32089), .X(n32087) );
  inv_x8_sg U41300 ( .A(n24421), .X(n50272) );
  nor_x8_sg U41301 ( .A(n41592), .B(n24423), .X(n24420) );
  nand_x4_sg U41302 ( .A(n41592), .B(n24423), .X(n24421) );
  nor_x2_sg U41303 ( .A(n29419), .B(n29420), .X(n29418) );
  nor_x2_sg U41304 ( .A(n29421), .B(n41558), .X(n29419) );
  nor_x2_sg U41305 ( .A(n29137), .B(n29138), .X(n29136) );
  nor_x2_sg U41306 ( .A(n29139), .B(n41560), .X(n29137) );
  nor_x2_sg U41307 ( .A(n28858), .B(n28859), .X(n28857) );
  nor_x2_sg U41308 ( .A(n28860), .B(n41562), .X(n28858) );
  nor_x2_sg U41309 ( .A(n28578), .B(n28579), .X(n28577) );
  nor_x2_sg U41310 ( .A(n28580), .B(n41564), .X(n28578) );
  nor_x2_sg U41311 ( .A(n28300), .B(n28301), .X(n28299) );
  nor_x2_sg U41312 ( .A(n28302), .B(n41566), .X(n28300) );
  nor_x2_sg U41313 ( .A(n28020), .B(n28021), .X(n28019) );
  nor_x2_sg U41314 ( .A(n28022), .B(n41568), .X(n28020) );
  nor_x2_sg U41315 ( .A(n26901), .B(n26902), .X(n26900) );
  nor_x2_sg U41316 ( .A(n26903), .B(n41570), .X(n26901) );
  nand_x4_sg U41317 ( .A(n53279), .B(n15952), .X(n15946) );
  nand_x4_sg U41318 ( .A(n51892), .B(n12057), .X(n12051) );
  nand_x4_sg U41319 ( .A(n51611), .B(n11278), .X(n11272) );
  nand_x4_sg U41320 ( .A(n41875), .B(n10597), .X(n10587) );
  nand_x4_sg U41321 ( .A(n41877), .B(n21469), .X(n21459) );
  nand_x4_sg U41322 ( .A(n41879), .B(n19924), .X(n19914) );
  inv_x4_sg U41323 ( .A(n25505), .X(n41260) );
  inv_x4_sg U41324 ( .A(n27739), .X(n41262) );
  inv_x4_sg U41325 ( .A(n27458), .X(n41264) );
  inv_x4_sg U41326 ( .A(n27179), .X(n41266) );
  inv_x4_sg U41327 ( .A(n26622), .X(n41268) );
  inv_x4_sg U41328 ( .A(n26343), .X(n41270) );
  inv_x4_sg U41329 ( .A(n26062), .X(n41272) );
  inv_x4_sg U41330 ( .A(n25783), .X(n41274) );
  nand_x4_sg U41331 ( .A(n10298), .B(n10388), .X(n10305) );
  nand_x4_sg U41332 ( .A(n21171), .B(n21260), .X(n21178) );
  nand_x4_sg U41333 ( .A(n19626), .B(n19715), .X(n19633) );
  inv_x4_sg U41334 ( .A(n51350), .X(n41276) );
  inv_x8_sg U41335 ( .A(n41276), .X(n41277) );
  inv_x4_sg U41336 ( .A(n20529), .X(n41278) );
  nor_x8_sg U41337 ( .A(n46272), .B(n46274), .X(n20529) );
  inv_x2_sg U41338 ( .A(n20529), .X(n54907) );
  inv_x4_sg U41339 ( .A(n18985), .X(n41279) );
  nor_x8_sg U41340 ( .A(n46317), .B(n46319), .X(n18985) );
  inv_x2_sg U41341 ( .A(n18985), .X(n54339) );
  inv_x4_sg U41342 ( .A(n17440), .X(n41280) );
  nor_x8_sg U41343 ( .A(n46364), .B(n46366), .X(n17440) );
  inv_x2_sg U41344 ( .A(n17440), .X(n53774) );
  inv_x2_sg U41345 ( .A(n50185), .X(n41281) );
  inv_x8_sg U41346 ( .A(n24079), .X(n50185) );
  inv_x2_sg U41347 ( .A(n50368), .X(n41282) );
  inv_x8_sg U41348 ( .A(n24107), .X(n50368) );
  inv_x2_sg U41349 ( .A(n49336), .X(n41283) );
  inv_x8_sg U41350 ( .A(n29729), .X(n49336) );
  inv_x2_sg U41351 ( .A(n49380), .X(n41284) );
  inv_x8_sg U41352 ( .A(n29736), .X(n49380) );
  inv_x2_sg U41353 ( .A(n49426), .X(n41285) );
  inv_x8_sg U41354 ( .A(n29743), .X(n49426) );
  inv_x2_sg U41355 ( .A(n49472), .X(n41286) );
  inv_x8_sg U41356 ( .A(n29750), .X(n49472) );
  inv_x2_sg U41357 ( .A(n49468), .X(n41287) );
  inv_x8_sg U41358 ( .A(n30619), .X(n49468) );
  inv_x2_sg U41359 ( .A(n49519), .X(n41288) );
  inv_x8_sg U41360 ( .A(n29757), .X(n49519) );
  inv_x2_sg U41361 ( .A(n49566), .X(n41289) );
  inv_x8_sg U41362 ( .A(n29764), .X(n49566) );
  inv_x2_sg U41363 ( .A(n49562), .X(n41290) );
  inv_x8_sg U41364 ( .A(n30633), .X(n49562) );
  inv_x2_sg U41365 ( .A(n49612), .X(n41291) );
  inv_x8_sg U41366 ( .A(n29771), .X(n49612) );
  inv_x2_sg U41367 ( .A(n49608), .X(n41292) );
  inv_x8_sg U41368 ( .A(n30640), .X(n49608) );
  inv_x2_sg U41369 ( .A(n49659), .X(n41293) );
  inv_x8_sg U41370 ( .A(n29778), .X(n49659) );
  inv_x2_sg U41371 ( .A(n49655), .X(n41294) );
  inv_x8_sg U41372 ( .A(n30647), .X(n49655) );
  inv_x2_sg U41373 ( .A(n49706), .X(n41295) );
  inv_x8_sg U41374 ( .A(n29785), .X(n49706) );
  inv_x2_sg U41375 ( .A(n49702), .X(n41296) );
  inv_x8_sg U41376 ( .A(n30654), .X(n49702) );
  inv_x2_sg U41377 ( .A(n49755), .X(n41297) );
  inv_x8_sg U41378 ( .A(n29792), .X(n49755) );
  inv_x2_sg U41379 ( .A(n49751), .X(n41298) );
  inv_x8_sg U41380 ( .A(n30661), .X(n49751) );
  inv_x2_sg U41381 ( .A(n49802), .X(n41299) );
  inv_x8_sg U41382 ( .A(n29799), .X(n49802) );
  inv_x2_sg U41383 ( .A(n49850), .X(n41300) );
  inv_x8_sg U41384 ( .A(n29806), .X(n49850) );
  inv_x2_sg U41385 ( .A(n49846), .X(n41301) );
  inv_x8_sg U41386 ( .A(n30675), .X(n49846) );
  inv_x2_sg U41387 ( .A(n49897), .X(n41302) );
  inv_x8_sg U41388 ( .A(n29813), .X(n49897) );
  inv_x2_sg U41389 ( .A(n49893), .X(n41303) );
  inv_x8_sg U41390 ( .A(n30682), .X(n49893) );
  inv_x2_sg U41391 ( .A(n49945), .X(n41304) );
  inv_x8_sg U41392 ( .A(n29820), .X(n49945) );
  inv_x2_sg U41393 ( .A(n49990), .X(n41305) );
  inv_x8_sg U41394 ( .A(n29827), .X(n49990) );
  inv_x2_sg U41395 ( .A(n50195), .X(n41306) );
  inv_x8_sg U41396 ( .A(n22064), .X(n50195) );
  inv_x2_sg U41397 ( .A(n50239), .X(n41307) );
  inv_x8_sg U41398 ( .A(n22071), .X(n50239) );
  inv_x2_sg U41399 ( .A(n50285), .X(n41308) );
  inv_x8_sg U41400 ( .A(n22078), .X(n50285) );
  inv_x2_sg U41401 ( .A(n50331), .X(n41309) );
  inv_x8_sg U41402 ( .A(n22085), .X(n50331) );
  inv_x2_sg U41403 ( .A(n50327), .X(n41310) );
  inv_x8_sg U41404 ( .A(n22953), .X(n50327) );
  inv_x2_sg U41405 ( .A(n50378), .X(n41311) );
  inv_x8_sg U41406 ( .A(n22092), .X(n50378) );
  inv_x2_sg U41407 ( .A(n50425), .X(n41312) );
  inv_x8_sg U41408 ( .A(n22099), .X(n50425) );
  inv_x2_sg U41409 ( .A(n50421), .X(n41313) );
  inv_x8_sg U41410 ( .A(n22967), .X(n50421) );
  inv_x2_sg U41411 ( .A(n50471), .X(n41314) );
  inv_x8_sg U41412 ( .A(n22106), .X(n50471) );
  inv_x2_sg U41413 ( .A(n50467), .X(n41315) );
  inv_x8_sg U41414 ( .A(n22974), .X(n50467) );
  inv_x2_sg U41415 ( .A(n50518), .X(n41316) );
  inv_x8_sg U41416 ( .A(n22113), .X(n50518) );
  inv_x2_sg U41417 ( .A(n50514), .X(n41317) );
  inv_x8_sg U41418 ( .A(n22981), .X(n50514) );
  inv_x2_sg U41419 ( .A(n50565), .X(n41318) );
  inv_x8_sg U41420 ( .A(n22120), .X(n50565) );
  inv_x2_sg U41421 ( .A(n50561), .X(n41319) );
  inv_x8_sg U41422 ( .A(n22988), .X(n50561) );
  inv_x2_sg U41423 ( .A(n50614), .X(n41320) );
  inv_x8_sg U41424 ( .A(n22127), .X(n50614) );
  inv_x2_sg U41425 ( .A(n50610), .X(n41321) );
  inv_x8_sg U41426 ( .A(n22995), .X(n50610) );
  inv_x2_sg U41427 ( .A(n50661), .X(n41322) );
  inv_x8_sg U41428 ( .A(n22134), .X(n50661) );
  inv_x2_sg U41429 ( .A(n50709), .X(n41323) );
  inv_x8_sg U41430 ( .A(n22141), .X(n50709) );
  inv_x2_sg U41431 ( .A(n50705), .X(n41324) );
  inv_x8_sg U41432 ( .A(n23009), .X(n50705) );
  inv_x2_sg U41433 ( .A(n50756), .X(n41325) );
  inv_x8_sg U41434 ( .A(n22148), .X(n50756) );
  inv_x2_sg U41435 ( .A(n50752), .X(n41326) );
  inv_x8_sg U41436 ( .A(n23016), .X(n50752) );
  inv_x2_sg U41437 ( .A(n50804), .X(n41327) );
  inv_x8_sg U41438 ( .A(n22155), .X(n50804) );
  inv_x2_sg U41439 ( .A(n50849), .X(n41328) );
  inv_x8_sg U41440 ( .A(n22162), .X(n50849) );
  inv_x2_sg U41441 ( .A(n49326), .X(n41329) );
  inv_x8_sg U41442 ( .A(n31745), .X(n49326) );
  inv_x2_sg U41443 ( .A(n49416), .X(n41330) );
  inv_x8_sg U41444 ( .A(n31759), .X(n49416) );
  inv_x2_sg U41445 ( .A(n49509), .X(n41331) );
  inv_x8_sg U41446 ( .A(n31773), .X(n49509) );
  inv_x2_sg U41447 ( .A(n50275), .X(n41332) );
  inv_x8_sg U41448 ( .A(n24093), .X(n50275) );
  inv_x2_sg U41449 ( .A(n49422), .X(n41333) );
  inv_x8_sg U41450 ( .A(n30612), .X(n49422) );
  inv_x2_sg U41451 ( .A(n49515), .X(n41334) );
  inv_x8_sg U41452 ( .A(n30626), .X(n49515) );
  inv_x2_sg U41453 ( .A(n50281), .X(n41335) );
  inv_x8_sg U41454 ( .A(n22946), .X(n50281) );
  inv_x2_sg U41455 ( .A(n50374), .X(n41336) );
  inv_x8_sg U41456 ( .A(n22960), .X(n50374) );
  inv_x2_sg U41457 ( .A(n49376), .X(n41337) );
  inv_x8_sg U41458 ( .A(n30605), .X(n49376) );
  inv_x2_sg U41459 ( .A(n50235), .X(n41338) );
  inv_x8_sg U41460 ( .A(n22939), .X(n50235) );
  inv_x2_sg U41461 ( .A(n49332), .X(n41339) );
  inv_x8_sg U41462 ( .A(n30598), .X(n49332) );
  inv_x2_sg U41463 ( .A(n50191), .X(n41340) );
  inv_x8_sg U41464 ( .A(n22932), .X(n50191) );
  nand_x4_sg U41465 ( .A(n21319), .B(n43131), .X(n21316) );
  nand_x4_sg U41466 ( .A(n19774), .B(n43135), .X(n19771) );
  inv_x4_sg U41467 ( .A(n41347), .X(n41348) );
  inv_x4_sg U41468 ( .A(n41349), .X(n41350) );
  nor_x8_sg U41469 ( .A(n46381), .B(n46377), .X(n17019) );
  nor_x8_sg U41470 ( .A(n46425), .B(n46421), .X(n15453) );
  nor_x8_sg U41471 ( .A(n46469), .B(n46471), .X(n13900) );
  nor_x8_sg U41472 ( .A(n46493), .B(n46489), .X(n13120) );
  nor_x8_sg U41473 ( .A(n46537), .B(n46533), .X(n11559) );
  nor_x8_sg U41474 ( .A(n54097), .B(n46335), .X(n18558) );
  nand_x4_sg U41475 ( .A(n21171), .B(n55207), .X(n9097) );
  nand_x4_sg U41476 ( .A(n43115), .B(n21173), .X(n21171) );
  nand_x4_sg U41477 ( .A(n54927), .B(n20399), .X(n9140) );
  inv_x4_sg U41478 ( .A(n41351), .X(n41352) );
  nand_x4_sg U41479 ( .A(n19626), .B(n54639), .X(n9195) );
  nand_x4_sg U41480 ( .A(n43119), .B(n19628), .X(n19626) );
  inv_x4_sg U41481 ( .A(n41353), .X(n41354) );
  inv_x4_sg U41482 ( .A(n41355), .X(n41356) );
  inv_x4_sg U41483 ( .A(n41357), .X(n41358) );
  inv_x4_sg U41484 ( .A(n41359), .X(n41360) );
  inv_x4_sg U41485 ( .A(n41361), .X(n41362) );
  inv_x4_sg U41486 ( .A(n41363), .X(n41364) );
  inv_x4_sg U41487 ( .A(n41365), .X(n41366) );
  nand_x4_sg U41488 ( .A(n10298), .B(n51285), .X(n9032) );
  nand_x4_sg U41489 ( .A(n43111), .B(n10300), .X(n10298) );
  inv_x4_sg U41490 ( .A(n16545), .X(n53554) );
  inv_x4_sg U41491 ( .A(n15763), .X(n53272) );
  inv_x4_sg U41492 ( .A(n14979), .X(n52996) );
  inv_x4_sg U41493 ( .A(n13430), .X(n52436) );
  inv_x4_sg U41494 ( .A(n12646), .X(n52162) );
  inv_x4_sg U41495 ( .A(n11868), .X(n51885) );
  inv_x4_sg U41496 ( .A(n11085), .X(n51604) );
  inv_x4_sg U41497 ( .A(n41367), .X(n41368) );
  inv_x4_sg U41498 ( .A(n41369), .X(n41370) );
  inv_x4_sg U41499 ( .A(n41371), .X(n41372) );
  inv_x4_sg U41500 ( .A(n41373), .X(n41374) );
  inv_x4_sg U41501 ( .A(n41375), .X(n41376) );
  inv_x4_sg U41502 ( .A(n41377), .X(n41378) );
  inv_x4_sg U41503 ( .A(n41379), .X(n41380) );
  inv_x4_sg U41504 ( .A(n41381), .X(n41382) );
  inv_x4_sg U41505 ( .A(n41383), .X(n41384) );
  inv_x4_sg U41506 ( .A(n41385), .X(n41386) );
  inv_x4_sg U41507 ( .A(n41387), .X(n41388) );
  inv_x4_sg U41508 ( .A(n41389), .X(n41390) );
  inv_x4_sg U41509 ( .A(n41391), .X(n41392) );
  inv_x4_sg U41510 ( .A(n41393), .X(n41394) );
  inv_x4_sg U41511 ( .A(n41395), .X(n41396) );
  inv_x4_sg U41512 ( .A(n41397), .X(n41398) );
  inv_x4_sg U41513 ( .A(n41399), .X(n41400) );
  inv_x4_sg U41514 ( .A(n41401), .X(n41402) );
  inv_x4_sg U41515 ( .A(n41403), .X(n41404) );
  inv_x4_sg U41516 ( .A(n41405), .X(n41406) );
  inv_x4_sg U41517 ( .A(n41407), .X(n41408) );
  inv_x4_sg U41518 ( .A(n41409), .X(n41410) );
  inv_x4_sg U41519 ( .A(n41411), .X(n41412) );
  inv_x4_sg U41520 ( .A(n41413), .X(n41414) );
  inv_x4_sg U41521 ( .A(n41415), .X(n41416) );
  inv_x4_sg U41522 ( .A(n41417), .X(n41418) );
  inv_x4_sg U41523 ( .A(n41419), .X(n41420) );
  inv_x4_sg U41524 ( .A(n41421), .X(n41422) );
  inv_x4_sg U41525 ( .A(n41423), .X(n41424) );
  inv_x4_sg U41526 ( .A(n41425), .X(n41426) );
  inv_x1_sg U41527 ( .A(n17163), .X(n41427) );
  nand_x4_sg U41528 ( .A(n17164), .B(n17165), .X(n17163) );
  inv_x1_sg U41529 ( .A(n16358), .X(n41428) );
  nand_x4_sg U41530 ( .A(n16359), .B(n16360), .X(n16358) );
  inv_x1_sg U41531 ( .A(n15597), .X(n41429) );
  nand_x4_sg U41532 ( .A(n15598), .B(n15599), .X(n15597) );
  inv_x1_sg U41533 ( .A(n13264), .X(n41430) );
  nand_x4_sg U41534 ( .A(n13265), .B(n13266), .X(n13264) );
  inv_x1_sg U41535 ( .A(n12483), .X(n41431) );
  nand_x4_sg U41536 ( .A(n12484), .B(n12485), .X(n12483) );
  nor_x4_sg U41537 ( .A(n18574), .B(n46340), .X(n18805) );
  nor_x4_sg U41538 ( .A(n16975), .B(n46385), .X(n17258) );
  nor_x4_sg U41539 ( .A(n15409), .B(n46429), .X(n15692) );
  nor_x4_sg U41540 ( .A(n13856), .B(n46475), .X(n14139) );
  nor_x4_sg U41541 ( .A(n13076), .B(n46497), .X(n13359) );
  nor_x4_sg U41542 ( .A(n12295), .B(n46518), .X(n12577) );
  nand_x4_sg U41543 ( .A(n20877), .B(n20878), .X(n20825) );
  nand_x4_sg U41544 ( .A(n43347), .B(n20886), .X(n20878) );
  nand_x4_sg U41545 ( .A(n19333), .B(n19334), .X(n19281) );
  nand_x4_sg U41546 ( .A(n43349), .B(n19342), .X(n19334) );
  nand_x4_sg U41547 ( .A(n17788), .B(n17789), .X(n17736) );
  nand_x4_sg U41548 ( .A(n43351), .B(n17797), .X(n17789) );
  inv_x4_sg U41549 ( .A(n41432), .X(n41433) );
  inv_x4_sg U41550 ( .A(n41434), .X(n41435) );
  inv_x4_sg U41551 ( .A(n41436), .X(n41437) );
  inv_x4_sg U41552 ( .A(n41438), .X(n41439) );
  inv_x4_sg U41553 ( .A(n41440), .X(n41441) );
  inv_x4_sg U41554 ( .A(n41442), .X(n41443) );
  inv_x4_sg U41555 ( .A(n41444), .X(n41445) );
  inv_x4_sg U41556 ( .A(n41446), .X(n41447) );
  inv_x4_sg U41557 ( .A(n41448), .X(n41449) );
  inv_x4_sg U41558 ( .A(n41450), .X(n41451) );
  inv_x4_sg U41559 ( .A(n41452), .X(n41453) );
  inv_x4_sg U41560 ( .A(n41454), .X(n41455) );
  inv_x4_sg U41561 ( .A(n41456), .X(n41457) );
  inv_x4_sg U41562 ( .A(n41458), .X(n41459) );
  inv_x4_sg U41563 ( .A(n41460), .X(n41461) );
  inv_x4_sg U41564 ( .A(n41462), .X(n41463) );
  inv_x4_sg U41565 ( .A(n41464), .X(n41465) );
  inv_x4_sg U41566 ( .A(n41466), .X(n41467) );
  inv_x4_sg U41567 ( .A(n41468), .X(n41469) );
  inv_x4_sg U41568 ( .A(n41470), .X(n41471) );
  inv_x4_sg U41569 ( .A(n41472), .X(n41473) );
  inv_x4_sg U41570 ( .A(n41474), .X(n41475) );
  inv_x1_sg U41571 ( .A(n18398), .X(n41476) );
  nand_x4_sg U41572 ( .A(n54167), .B(n18399), .X(n18398) );
  inv_x4_sg U41573 ( .A(n10732), .X(n51396) );
  nor_x4_sg U41574 ( .A(n46555), .B(n46573), .X(n10732) );
  inv_x1_sg U41575 ( .A(n20718), .X(n41477) );
  nand_x4_sg U41576 ( .A(n55018), .B(n20719), .X(n20718) );
  inv_x1_sg U41577 ( .A(n19174), .X(n41478) );
  nand_x4_sg U41578 ( .A(n54450), .B(n19175), .X(n19174) );
  inv_x1_sg U41579 ( .A(n17629), .X(n41479) );
  nand_x4_sg U41580 ( .A(n53885), .B(n17630), .X(n17629) );
  inv_x1_sg U41581 ( .A(n14508), .X(n41480) );
  nand_x4_sg U41582 ( .A(n52765), .B(n14509), .X(n14508) );
  inv_x1_sg U41583 ( .A(n31272), .X(n41664) );
  inv_x1_sg U41584 ( .A(n31284), .X(n42936) );
  inv_x1_sg U41585 ( .A(n31302), .X(n42941) );
  inv_x4_sg U41586 ( .A(n41481), .X(n41482) );
  inv_x2_sg U41587 ( .A(n30164), .X(n42490) );
  inv_x4_sg U41588 ( .A(n41483), .X(n41484) );
  inv_x2_sg U41589 ( .A(n30176), .X(n42492) );
  inv_x2_sg U41590 ( .A(n20606), .X(n41833) );
  inv_x2_sg U41591 ( .A(n19062), .X(n41837) );
  inv_x2_sg U41592 ( .A(n17517), .X(n41839) );
  inv_x2_sg U41593 ( .A(n14396), .X(n41841) );
  inv_x2_sg U41594 ( .A(n10505), .X(n41843) );
  inv_x1_sg U41595 ( .A(n23606), .X(n41674) );
  inv_x4_sg U41596 ( .A(n41485), .X(n41486) );
  inv_x2_sg U41597 ( .A(n22498), .X(n42494) );
  inv_x4_sg U41598 ( .A(n41487), .X(n41488) );
  inv_x2_sg U41599 ( .A(n22510), .X(n42496) );
  inv_x1_sg U41600 ( .A(n14002), .X(n41722) );
  inv_x1_sg U41601 ( .A(n23618), .X(n43018) );
  inv_x1_sg U41602 ( .A(n23636), .X(n43023) );
  inv_x1_sg U41603 ( .A(n23653), .X(n41678) );
  inv_x1_sg U41604 ( .A(n31496), .X(n43180) );
  inv_x1_sg U41605 ( .A(n23830), .X(n43192) );
  inv_x1_sg U41606 ( .A(n16285), .X(n42072) );
  inv_x1_sg U41607 ( .A(n17281), .X(n42288) );
  inv_x1_sg U41608 ( .A(n17280), .X(n42289) );
  inv_x1_sg U41609 ( .A(n15715), .X(n42291) );
  inv_x1_sg U41610 ( .A(n15714), .X(n42292) );
  inv_x1_sg U41611 ( .A(n14162), .X(n42294) );
  inv_x1_sg U41612 ( .A(n14161), .X(n42295) );
  inv_x1_sg U41613 ( .A(n13382), .X(n42297) );
  inv_x1_sg U41614 ( .A(n13381), .X(n42298) );
  inv_x1_sg U41615 ( .A(n12600), .X(n42300) );
  inv_x1_sg U41616 ( .A(n12599), .X(n42301) );
  inv_x1_sg U41617 ( .A(n18650), .X(n42100) );
  inv_x1_sg U41618 ( .A(n16500), .X(n43174) );
  inv_x1_sg U41619 ( .A(n12390), .X(n42110) );
  inv_x1_sg U41620 ( .A(n11609), .X(n42112) );
  inv_x1_sg U41621 ( .A(n20931), .X(n42114) );
  inv_x1_sg U41622 ( .A(n19387), .X(n42116) );
  inv_x1_sg U41623 ( .A(n17842), .X(n42118) );
  inv_x1_sg U41624 ( .A(n14721), .X(n42122) );
  inv_x1_sg U41625 ( .A(n11800), .X(n42136) );
  inv_x2_sg U41626 ( .A(n16528), .X(n41823) );
  inv_x2_sg U41627 ( .A(n14962), .X(n41825) );
  inv_x2_sg U41628 ( .A(n12629), .X(n41827) );
  inv_x2_sg U41629 ( .A(n11068), .X(n41829) );
  inv_x4_sg U41630 ( .A(n41489), .X(n41490) );
  nor_x2_sg U41631 ( .A(n17220), .B(n42260), .X(n17218) );
  inv_x4_sg U41632 ( .A(n41491), .X(n41492) );
  nor_x2_sg U41633 ( .A(n15654), .B(n42264), .X(n15652) );
  inv_x4_sg U41634 ( .A(n41493), .X(n41494) );
  nor_x2_sg U41635 ( .A(n13321), .B(n42272), .X(n13319) );
  inv_x4_sg U41636 ( .A(n41495), .X(n41496) );
  nor_x2_sg U41637 ( .A(n12540), .B(n42276), .X(n12538) );
  inv_x4_sg U41638 ( .A(n41497), .X(n41498) );
  inv_x2_sg U41639 ( .A(n41499), .X(n41500) );
  inv_x4_sg U41640 ( .A(n41501), .X(n41502) );
  inv_x2_sg U41641 ( .A(n41503), .X(n41504) );
  inv_x4_sg U41642 ( .A(n41505), .X(n41506) );
  inv_x2_sg U41643 ( .A(n41507), .X(n41508) );
  inv_x4_sg U41644 ( .A(n41509), .X(n41510) );
  inv_x2_sg U41645 ( .A(n41511), .X(n41512) );
  inv_x4_sg U41646 ( .A(n41513), .X(n41514) );
  inv_x4_sg U41647 ( .A(n41515), .X(n41516) );
  inv_x4_sg U41648 ( .A(n41517), .X(n41518) );
  inv_x4_sg U41649 ( .A(n41519), .X(n41520) );
  inv_x4_sg U41650 ( .A(n40586), .X(n41521) );
  inv_x4_sg U41651 ( .A(n14104), .X(n52570) );
  nand_x2_sg U41652 ( .A(n14105), .B(n14048), .X(n14104) );
  nor_x2_sg U41653 ( .A(n12412), .B(n12413), .X(n12411) );
  nor_x4_sg U41654 ( .A(n42367), .B(n52022), .X(n12413) );
  inv_x4_sg U41655 ( .A(n12420), .X(n52022) );
  nand_x2_sg U41656 ( .A(n41768), .B(n12422), .X(n12420) );
  nor_x4_sg U41657 ( .A(n15770), .B(n41736), .X(n15776) );
  nor_x4_sg U41658 ( .A(n16552), .B(n41750), .X(n16558) );
  nor_x4_sg U41659 ( .A(n14986), .B(n41752), .X(n14992) );
  nor_x4_sg U41660 ( .A(n13437), .B(n41754), .X(n13443) );
  nor_x4_sg U41661 ( .A(n12653), .B(n41756), .X(n12659) );
  nor_x4_sg U41662 ( .A(n11875), .B(n41758), .X(n11881) );
  nor_x4_sg U41663 ( .A(n11092), .B(n41760), .X(n11098) );
  nor_x2_sg U41664 ( .A(n51527), .B(n51481), .X(n25499) );
  nor_x2_sg U41665 ( .A(n51481), .B(n51474), .X(n25509) );
  inv_x4_sg U41666 ( .A(n10919), .X(n51481) );
  inv_x4_sg U41667 ( .A(n41523), .X(n41524) );
  inv_x4_sg U41668 ( .A(n41525), .X(n41526) );
  inv_x4_sg U41669 ( .A(n41527), .X(n41528) );
  nor_x2_sg U41670 ( .A(n55389), .B(n41812), .X(n21886) );
  inv_x4_sg U41671 ( .A(n41529), .X(n41530) );
  nor_x2_sg U41672 ( .A(n54821), .B(n41814), .X(n20341) );
  inv_x4_sg U41673 ( .A(n41531), .X(n41532) );
  inv_x4_sg U41674 ( .A(n41533), .X(n41534) );
  nor_x4_sg U41675 ( .A(n10527), .B(n42369), .X(n10529) );
  nor_x4_sg U41676 ( .A(n21399), .B(n43233), .X(n21401) );
  inv_x4_sg U41677 ( .A(n41535), .X(n41536) );
  nor_x2_sg U41678 ( .A(n55104), .B(n41816), .X(n21115) );
  nor_x4_sg U41679 ( .A(n19854), .B(n43235), .X(n19856) );
  inv_x4_sg U41680 ( .A(n41537), .X(n41538) );
  nor_x2_sg U41681 ( .A(n54536), .B(n41818), .X(n19571) );
  nor_x4_sg U41682 ( .A(n18309), .B(n42371), .X(n18311) );
  inv_x4_sg U41683 ( .A(n41539), .X(n41540) );
  nor_x2_sg U41684 ( .A(n53971), .B(n41820), .X(n18026) );
  inv_x4_sg U41685 ( .A(n41541), .X(n41542) );
  nor_x2_sg U41686 ( .A(n52851), .B(n41822), .X(n14905) );
  nor_x4_sg U41687 ( .A(n20628), .B(n43243), .X(n20630) );
  nor_x4_sg U41688 ( .A(n19084), .B(n43245), .X(n19086) );
  nor_x4_sg U41689 ( .A(n17539), .B(n43247), .X(n17541) );
  nor_x4_sg U41690 ( .A(n14419), .B(n43249), .X(n14421) );
  nor_x4_sg U41691 ( .A(n41734), .B(n52456), .X(n13613) );
  inv_x4_sg U41692 ( .A(n13612), .X(n52456) );
  nand_x4_sg U41693 ( .A(n52443), .B(n13618), .X(n13612) );
  inv_x8_sg U41694 ( .A(n42672), .X(n42673) );
  inv_x8_sg U41695 ( .A(n42676), .X(n42677) );
  inv_x8_sg U41696 ( .A(n42680), .X(n42681) );
  inv_x8_sg U41697 ( .A(n42682), .X(n42683) );
  inv_x8_sg U41698 ( .A(n42684), .X(n42685) );
  inv_x8_sg U41699 ( .A(n42744), .X(n42745) );
  inv_x8_sg U41700 ( .A(n42748), .X(n42749) );
  inv_x8_sg U41701 ( .A(n42752), .X(n42753) );
  inv_x8_sg U41702 ( .A(n42754), .X(n42755) );
  inv_x8_sg U41703 ( .A(n42756), .X(n42757) );
  inv_x4_sg U41704 ( .A(n41545), .X(n41546) );
  nor_x4_sg U41705 ( .A(n41546), .B(n54113), .X(n18277) );
  inv_x4_sg U41706 ( .A(n18288), .X(n54113) );
  nand_x2_sg U41707 ( .A(n41905), .B(n41149), .X(n18288) );
  inv_x4_sg U41708 ( .A(n41547), .X(n41548) );
  nor_x4_sg U41709 ( .A(n41548), .B(n53572), .X(n16738) );
  inv_x4_sg U41710 ( .A(n16759), .X(n53572) );
  nand_x2_sg U41711 ( .A(n16760), .B(n53571), .X(n16759) );
  inv_x4_sg U41712 ( .A(n41549), .X(n41550) );
  nor_x4_sg U41713 ( .A(n41550), .B(n53014), .X(n15172) );
  inv_x4_sg U41714 ( .A(n15193), .X(n53014) );
  nand_x2_sg U41715 ( .A(n15194), .B(n53013), .X(n15193) );
  inv_x4_sg U41716 ( .A(n41551), .X(n41552) );
  nor_x4_sg U41717 ( .A(n41552), .B(n52180), .X(n12839) );
  inv_x4_sg U41718 ( .A(n12860), .X(n52180) );
  nand_x2_sg U41719 ( .A(n12861), .B(n52179), .X(n12860) );
  nor_x2_sg U41720 ( .A(n46218), .B(n53363), .X(n27434) );
  nor_x2_sg U41721 ( .A(n46228), .B(n51974), .X(n26037) );
  nor_x2_sg U41722 ( .A(n46230), .B(n51693), .X(n25759) );
  nor_x2_sg U41723 ( .A(n51476), .B(n51498), .X(n10902) );
  nor_x2_sg U41724 ( .A(n13546), .B(n13547), .X(n13545) );
  nor_x2_sg U41725 ( .A(n20537), .B(n20538), .X(n20536) );
  nor_x2_sg U41726 ( .A(n18993), .B(n18994), .X(n18992) );
  nor_x2_sg U41727 ( .A(n17448), .B(n17449), .X(n17447) );
  nor_x2_sg U41728 ( .A(n14325), .B(n14326), .X(n14324) );
  nand_x4_sg U41729 ( .A(n51508), .B(n10362), .X(n10765) );
  nand_x4_sg U41730 ( .A(n42851), .B(n10821), .X(n10362) );
  inv_x4_sg U41731 ( .A(n29417), .X(n41557) );
  inv_x4_sg U41732 ( .A(n29135), .X(n41559) );
  inv_x4_sg U41733 ( .A(n28856), .X(n41561) );
  inv_x4_sg U41734 ( .A(n28576), .X(n41563) );
  inv_x4_sg U41735 ( .A(n28298), .X(n41565) );
  inv_x4_sg U41736 ( .A(n28018), .X(n41567) );
  inv_x4_sg U41737 ( .A(n26899), .X(n41569) );
  nand_x4_sg U41738 ( .A(n18556), .B(n18557), .X(n18505) );
  inv_x4_sg U41739 ( .A(n55272), .X(n41571) );
  inv_x8_sg U41740 ( .A(n41571), .X(n41572) );
  inv_x4_sg U41741 ( .A(n54704), .X(n41573) );
  inv_x8_sg U41742 ( .A(n41573), .X(n41574) );
  inv_x2_sg U41743 ( .A(n50321), .X(n41575) );
  inv_x8_sg U41744 ( .A(n24100), .X(n50321) );
  inv_x2_sg U41745 ( .A(n50415), .X(n41576) );
  inv_x8_sg U41746 ( .A(n24114), .X(n50415) );
  inv_x2_sg U41747 ( .A(n49799), .X(n41577) );
  inv_x8_sg U41748 ( .A(n30668), .X(n49799) );
  inv_x2_sg U41749 ( .A(n50658), .X(n41578) );
  inv_x8_sg U41750 ( .A(n23002), .X(n50658) );
  inv_x2_sg U41751 ( .A(n49462), .X(n41579) );
  inv_x8_sg U41752 ( .A(n31766), .X(n49462) );
  inv_x2_sg U41753 ( .A(n49556), .X(n41580) );
  inv_x8_sg U41754 ( .A(n31780), .X(n49556) );
  nand_x2_sg U41755 ( .A(n46584), .B(n43265), .X(n29612) );
  inv_x4_sg U41756 ( .A(n41581), .X(n41582) );
  inv_x4_sg U41757 ( .A(n41583), .X(n41584) );
  inv_x1_sg U41758 ( .A(n14044), .X(n41585) );
  nand_x4_sg U41759 ( .A(n14045), .B(n14046), .X(n14044) );
  inv_x1_sg U41760 ( .A(n10903), .X(n41586) );
  nand_x4_sg U41761 ( .A(n10904), .B(n10905), .X(n10903) );
  inv_x4_sg U41762 ( .A(n41587), .X(n41588) );
  inv_x4_sg U41763 ( .A(n32088), .X(n41589) );
  inv_x4_sg U41764 ( .A(n24422), .X(n41591) );
  nor_x2_sg U41765 ( .A(n20974), .B(n20973), .X(n20971) );
  nor_x4_sg U41766 ( .A(n20884), .B(n46270), .X(n20973) );
  nor_x2_sg U41767 ( .A(n19430), .B(n19429), .X(n19427) );
  nor_x4_sg U41768 ( .A(n19340), .B(n46315), .X(n19429) );
  nor_x2_sg U41769 ( .A(n17885), .B(n17884), .X(n17882) );
  nor_x4_sg U41770 ( .A(n17795), .B(n46362), .X(n17884) );
  nor_x2_sg U41771 ( .A(n14764), .B(n14763), .X(n14761) );
  nor_x4_sg U41772 ( .A(n14674), .B(n46451), .X(n14763) );
  nor_x2_sg U41773 ( .A(n11652), .B(n11651), .X(n11649) );
  nor_x4_sg U41774 ( .A(n11638), .B(n46541), .X(n11651) );
  nor_x2_sg U41775 ( .A(n10872), .B(n10871), .X(n10869) );
  nor_x4_sg U41776 ( .A(n46565), .B(n10782), .X(n10871) );
  inv_x4_sg U41777 ( .A(n21442), .X(n55269) );
  inv_x4_sg U41778 ( .A(n19897), .X(n54701) );
  inv_x4_sg U41779 ( .A(n18352), .X(n54137) );
  inv_x4_sg U41780 ( .A(n10407), .X(n51276) );
  inv_x4_sg U41781 ( .A(n21279), .X(n55198) );
  inv_x4_sg U41782 ( .A(n20671), .X(n54990) );
  inv_x4_sg U41783 ( .A(n19734), .X(n54630) );
  inv_x4_sg U41784 ( .A(n19127), .X(n54422) );
  inv_x4_sg U41785 ( .A(n17582), .X(n53857) );
  inv_x4_sg U41786 ( .A(n14462), .X(n52737) );
  inv_x4_sg U41787 ( .A(n41593), .X(n41594) );
  nor_x2_sg U41788 ( .A(n44670), .B(n53504), .X(n16636) );
  inv_x4_sg U41789 ( .A(n16638), .X(n53504) );
  nor_x2_sg U41790 ( .A(n44672), .B(n52946), .X(n15070) );
  inv_x4_sg U41791 ( .A(n15072), .X(n52946) );
  nor_x2_sg U41792 ( .A(n44674), .B(n52112), .X(n12737) );
  inv_x4_sg U41793 ( .A(n12739), .X(n52112) );
  nor_x2_sg U41794 ( .A(n44676), .B(n51555), .X(n11176) );
  inv_x4_sg U41795 ( .A(n11178), .X(n51555) );
  inv_x4_sg U41796 ( .A(n41595), .X(n41596) );
  inv_x4_sg U41797 ( .A(n41597), .X(n41598) );
  inv_x4_sg U41798 ( .A(n41599), .X(n41600) );
  inv_x4_sg U41799 ( .A(n41601), .X(n41602) );
  inv_x4_sg U41800 ( .A(n27435), .X(n41603) );
  inv_x4_sg U41801 ( .A(n26038), .X(n41605) );
  inv_x4_sg U41802 ( .A(n25760), .X(n41607) );
  inv_x4_sg U41803 ( .A(n24345), .X(n41609) );
  inv_x4_sg U41804 ( .A(n31992), .X(n41611) );
  inv_x4_sg U41805 ( .A(n32011), .X(n41613) );
  inv_x4_sg U41806 ( .A(n24326), .X(n41615) );
  nor_x8_sg U41807 ( .A(n27410), .B(n53319), .X(n27417) );
  nor_x8_sg U41808 ( .A(n26013), .B(n51931), .X(n26020) );
  nor_x8_sg U41809 ( .A(n25735), .B(n51650), .X(n25742) );
  nor_x8_sg U41810 ( .A(n29397), .B(n55386), .X(n29404) );
  nor_x8_sg U41811 ( .A(n29115), .B(n55101), .X(n29122) );
  nor_x8_sg U41812 ( .A(n28836), .B(n54818), .X(n28843) );
  nor_x8_sg U41813 ( .A(n28556), .B(n54533), .X(n28563) );
  nor_x8_sg U41814 ( .A(n28278), .B(n54250), .X(n28285) );
  nor_x8_sg U41815 ( .A(n27998), .B(n53968), .X(n28005) );
  nor_x8_sg U41816 ( .A(n26879), .B(n52848), .X(n26886) );
  inv_x4_sg U41817 ( .A(n41617), .X(n41618) );
  inv_x4_sg U41818 ( .A(n41619), .X(n41620) );
  inv_x4_sg U41819 ( .A(n41621), .X(n41622) );
  inv_x4_sg U41820 ( .A(n41623), .X(n41624) );
  inv_x4_sg U41821 ( .A(n41625), .X(n41626) );
  inv_x4_sg U41822 ( .A(n41627), .X(n41628) );
  inv_x4_sg U41823 ( .A(n41629), .X(n41630) );
  inv_x4_sg U41824 ( .A(n41631), .X(n41632) );
  inv_x4_sg U41825 ( .A(n41633), .X(n41634) );
  inv_x4_sg U41826 ( .A(n41635), .X(n41636) );
  inv_x4_sg U41827 ( .A(n41637), .X(n41638) );
  inv_x4_sg U41828 ( .A(n41639), .X(n41640) );
  inv_x4_sg U41829 ( .A(n41641), .X(n41642) );
  inv_x4_sg U41830 ( .A(n41643), .X(n41644) );
  inv_x4_sg U41831 ( .A(n41645), .X(n41646) );
  inv_x4_sg U41832 ( .A(n41647), .X(n41648) );
  nor_x8_sg U41833 ( .A(n24420), .B(n50272), .X(n10078) );
  inv_x1_sg U41834 ( .A(n10078), .X(n50273) );
  nor_x8_sg U41835 ( .A(n32086), .B(n49413), .X(n25186) );
  inv_x1_sg U41836 ( .A(n25186), .X(n49414) );
  inv_x1_sg U41837 ( .A(n10616), .X(n41649) );
  nand_x4_sg U41838 ( .A(n51379), .B(n10617), .X(n10616) );
  inv_x1_sg U41839 ( .A(n21488), .X(n41650) );
  nand_x4_sg U41840 ( .A(n55301), .B(n21489), .X(n21488) );
  inv_x1_sg U41841 ( .A(n19943), .X(n41651) );
  nand_x4_sg U41842 ( .A(n54733), .B(n19944), .X(n19943) );
  inv_x1_sg U41843 ( .A(n16542), .X(n41977) );
  inv_x1_sg U41844 ( .A(n15760), .X(n41981) );
  inv_x1_sg U41845 ( .A(n14976), .X(n41985) );
  inv_x1_sg U41846 ( .A(n13427), .X(n41991) );
  inv_x1_sg U41847 ( .A(n12643), .X(n41995) );
  inv_x1_sg U41848 ( .A(n11865), .X(n41999) );
  inv_x1_sg U41849 ( .A(n11082), .X(n42003) );
  inv_x1_sg U41850 ( .A(n16582), .X(n42009) );
  inv_x1_sg U41851 ( .A(n15016), .X(n42013) );
  inv_x1_sg U41852 ( .A(n13467), .X(n42017) );
  inv_x1_sg U41853 ( .A(n12683), .X(n42021) );
  inv_x1_sg U41854 ( .A(n11905), .X(n42025) );
  inv_x2_sg U41855 ( .A(n31436), .X(n43443) );
  inv_x1_sg U41856 ( .A(n30511), .X(n42950) );
  inv_x1_sg U41857 ( .A(n21802), .X(n42954) );
  inv_x1_sg U41858 ( .A(n21031), .X(n42958) );
  inv_x1_sg U41859 ( .A(n20257), .X(n42962) );
  inv_x1_sg U41860 ( .A(n19487), .X(n42966) );
  inv_x1_sg U41861 ( .A(n18711), .X(n42970) );
  inv_x1_sg U41862 ( .A(n17942), .X(n42974) );
  inv_x1_sg U41863 ( .A(n17169), .X(n42978) );
  inv_x1_sg U41864 ( .A(n15603), .X(n42986) );
  inv_x1_sg U41865 ( .A(n14821), .X(n42990) );
  inv_x1_sg U41866 ( .A(n14050), .X(n42994) );
  inv_x1_sg U41867 ( .A(n13270), .X(n42998) );
  inv_x1_sg U41868 ( .A(n12489), .X(n43002) );
  inv_x1_sg U41869 ( .A(n11709), .X(n43006) );
  inv_x1_sg U41870 ( .A(n22845), .X(n43014) );
  inv_x2_sg U41871 ( .A(n23770), .X(n43445) );
  inv_x2_sg U41872 ( .A(n30191), .X(n42464) );
  inv_x1_sg U41873 ( .A(n24361), .X(n42199) );
  inv_x1_sg U41874 ( .A(n24376), .X(n42203) );
  inv_x1_sg U41875 ( .A(n24158), .X(n42209) );
  inv_x1_sg U41876 ( .A(n23861), .X(n42215) );
  inv_x1_sg U41877 ( .A(n23500), .X(n42221) );
  inv_x2_sg U41878 ( .A(n22525), .X(n42466) );
  inv_x1_sg U41879 ( .A(n30455), .X(n43184) );
  inv_x1_sg U41880 ( .A(n22789), .X(n43188) );
  inv_x1_sg U41881 ( .A(n32027), .X(n42233) );
  inv_x1_sg U41882 ( .A(n32042), .X(n42237) );
  inv_x1_sg U41883 ( .A(n31824), .X(n42243) );
  inv_x1_sg U41884 ( .A(n31527), .X(n42247) );
  inv_x1_sg U41885 ( .A(n31166), .X(n42251) );
  inv_x1_sg U41886 ( .A(n13990), .X(n42076) );
  inv_x1_sg U41887 ( .A(n17069), .X(n42102) );
  nor_x2_sg U41888 ( .A(n53253), .B(n53365), .X(n16160) );
  inv_x4_sg U41889 ( .A(n42311), .X(n53365) );
  inv_x1_sg U41890 ( .A(n16159), .X(n43306) );
  inv_x1_sg U41891 ( .A(n15503), .X(n42104) );
  inv_x1_sg U41892 ( .A(n13950), .X(n42106) );
  inv_x1_sg U41893 ( .A(n13170), .X(n42108) );
  inv_x2_sg U41894 ( .A(n30471), .X(n42500) );
  nor_x2_sg U41895 ( .A(n46513), .B(n51976), .X(n12265) );
  inv_x4_sg U41896 ( .A(n42313), .X(n51976) );
  inv_x1_sg U41897 ( .A(n12264), .X(n43312) );
  inv_x2_sg U41898 ( .A(n22805), .X(n42504) );
  inv_x1_sg U41899 ( .A(n10703), .X(n43316) );
  nor_x2_sg U41900 ( .A(n51306), .B(n51421), .X(n10704) );
  inv_x4_sg U41901 ( .A(n42323), .X(n51421) );
  inv_x1_sg U41902 ( .A(n21575), .X(n43320) );
  nor_x2_sg U41903 ( .A(n55228), .B(n55348), .X(n21576) );
  inv_x4_sg U41904 ( .A(n42325), .X(n55348) );
  inv_x1_sg U41905 ( .A(n20030), .X(n43324) );
  nor_x2_sg U41906 ( .A(n54660), .B(n54780), .X(n20031) );
  inv_x4_sg U41907 ( .A(n42327), .X(n54780) );
  inv_x1_sg U41908 ( .A(n18803), .X(n42124) );
  inv_x1_sg U41909 ( .A(n17256), .X(n42126) );
  inv_x1_sg U41910 ( .A(n15690), .X(n42128) );
  inv_x1_sg U41911 ( .A(n14137), .X(n42130) );
  inv_x1_sg U41912 ( .A(n13357), .X(n42132) );
  inv_x1_sg U41913 ( .A(n12575), .X(n42134) );
  nor_x2_sg U41914 ( .A(n46266), .B(n55064), .X(n20806) );
  inv_x4_sg U41915 ( .A(n42329), .X(n55064) );
  inv_x1_sg U41916 ( .A(n20805), .X(n43328) );
  nor_x2_sg U41917 ( .A(n46311), .B(n54496), .X(n19262) );
  inv_x4_sg U41918 ( .A(n42331), .X(n54496) );
  inv_x1_sg U41919 ( .A(n19261), .X(n43332) );
  nor_x2_sg U41920 ( .A(n46358), .B(n53931), .X(n17717) );
  inv_x4_sg U41921 ( .A(n42333), .X(n53931) );
  inv_x1_sg U41922 ( .A(n17716), .X(n43336) );
  inv_x1_sg U41923 ( .A(n14595), .X(n43340) );
  nor_x2_sg U41924 ( .A(n52695), .B(n52811), .X(n14596) );
  inv_x4_sg U41925 ( .A(n42335), .X(n52811) );
  inv_x2_sg U41926 ( .A(n11803), .X(n43551) );
  inv_x1_sg U41927 ( .A(n10783), .X(n43343) );
  inv_x1_sg U41928 ( .A(n10740), .X(n43101) );
  inv_x2_sg U41929 ( .A(n10733), .X(n42458) );
  inv_x2_sg U41930 ( .A(n17021), .X(n43473) );
  inv_x2_sg U41931 ( .A(n15455), .X(n43475) );
  inv_x2_sg U41932 ( .A(n13122), .X(n43479) );
  inv_x2_sg U41933 ( .A(n11561), .X(n43481) );
  nor_x2_sg U41934 ( .A(n18346), .B(n42138), .X(n18383) );
  inv_x2_sg U41935 ( .A(n18559), .X(n42468) );
  nor_x2_sg U41936 ( .A(n20665), .B(n42140), .X(n20703) );
  nor_x2_sg U41937 ( .A(n19121), .B(n42142), .X(n19159) );
  nor_x2_sg U41938 ( .A(n17576), .B(n42144), .X(n17614) );
  nor_x2_sg U41939 ( .A(n14456), .B(n42146), .X(n14493) );
  inv_x2_sg U41940 ( .A(n20887), .X(n43346) );
  inv_x2_sg U41941 ( .A(n19343), .X(n43348) );
  inv_x2_sg U41942 ( .A(n17798), .X(n43350) );
  inv_x1_sg U41943 ( .A(n26689), .X(n42149) );
  inv_x2_sg U41944 ( .A(n10440), .X(n43260) );
  inv_x1_sg U41945 ( .A(n21325), .X(n43132) );
  inv_x1_sg U41946 ( .A(n19780), .X(n43136) );
  inv_x1_sg U41947 ( .A(n27527), .X(n42169) );
  inv_x1_sg U41948 ( .A(n25571), .X(n42173) );
  inv_x1_sg U41949 ( .A(n29484), .X(n42177) );
  inv_x2_sg U41950 ( .A(n20400), .X(n42436) );
  inv_x1_sg U41951 ( .A(n28923), .X(n42181) );
  inv_x2_sg U41952 ( .A(n18856), .X(n42438) );
  inv_x2_sg U41953 ( .A(n17311), .X(n42440) );
  inv_x1_sg U41954 ( .A(n26132), .X(n42185) );
  inv_x4_sg U41955 ( .A(n41652), .X(n41653) );
  inv_x4_sg U41956 ( .A(n41654), .X(n41655) );
  inv_x4_sg U41957 ( .A(n41656), .X(n41657) );
  inv_x4_sg U41958 ( .A(n41658), .X(n41659) );
  inv_x4_sg U41959 ( .A(n41660), .X(n41661) );
  inv_x4_sg U41960 ( .A(n41662), .X(n41663) );
  inv_x2_sg U41961 ( .A(n41664), .X(n41665) );
  inv_x4_sg U41962 ( .A(n41666), .X(n41667) );
  inv_x2_sg U41963 ( .A(n41668), .X(n41669) );
  inv_x4_sg U41964 ( .A(n41670), .X(n41671) );
  nor_x2_sg U41965 ( .A(n40753), .B(n49822), .X(n31326) );
  inv_x4_sg U41966 ( .A(n41672), .X(n41673) );
  inv_x2_sg U41967 ( .A(n41674), .X(n41675) );
  inv_x4_sg U41968 ( .A(n41676), .X(n41677) );
  inv_x2_sg U41969 ( .A(n41678), .X(n41679) );
  inv_x4_sg U41970 ( .A(n41680), .X(n41681) );
  nor_x2_sg U41971 ( .A(n40754), .B(n50681), .X(n23660) );
  nor_x1_sg U41972 ( .A(n55433), .B(n21734), .X(n21235) );
  nor_x2_sg U41973 ( .A(n43055), .B(n21736), .X(n21734) );
  nor_x1_sg U41974 ( .A(n55148), .B(n20965), .X(n20463) );
  nor_x2_sg U41975 ( .A(n43057), .B(n20967), .X(n20965) );
  nor_x1_sg U41976 ( .A(n54865), .B(n20189), .X(n19690) );
  nor_x2_sg U41977 ( .A(n43063), .B(n20191), .X(n20189) );
  nor_x1_sg U41978 ( .A(n54580), .B(n19421), .X(n18919) );
  nor_x2_sg U41979 ( .A(n43065), .B(n19423), .X(n19421) );
  nor_x1_sg U41980 ( .A(n54297), .B(n18643), .X(n18145) );
  nor_x2_sg U41981 ( .A(n43071), .B(n18645), .X(n18643) );
  nor_x1_sg U41982 ( .A(n54015), .B(n17876), .X(n17374) );
  nor_x2_sg U41983 ( .A(n43073), .B(n17878), .X(n17876) );
  nor_x1_sg U41984 ( .A(n53455), .B(n16318), .X(n15810) );
  nor_x2_sg U41985 ( .A(n42064), .B(n16320), .X(n16318) );
  nor_x1_sg U41986 ( .A(n52895), .B(n14755), .X(n14255) );
  nor_x2_sg U41987 ( .A(n43081), .B(n14757), .X(n14755) );
  nor_x1_sg U41988 ( .A(n51785), .B(n11643), .X(n11131) );
  nor_x2_sg U41989 ( .A(n43093), .B(n11645), .X(n11643) );
  nor_x1_sg U41990 ( .A(n51505), .B(n10863), .X(n10364) );
  nor_x2_sg U41991 ( .A(n43095), .B(n10865), .X(n10863) );
  inv_x4_sg U41992 ( .A(n41682), .X(n41683) );
  inv_x2_sg U41993 ( .A(n41684), .X(n41685) );
  nor_x2_sg U41994 ( .A(n42287), .B(n17120), .X(n17117) );
  inv_x4_sg U41995 ( .A(n41686), .X(n41687) );
  inv_x2_sg U41996 ( .A(n41688), .X(n41689) );
  nor_x2_sg U41997 ( .A(n42290), .B(n15554), .X(n15551) );
  inv_x4_sg U41998 ( .A(n41690), .X(n41691) );
  inv_x2_sg U41999 ( .A(n41692), .X(n41693) );
  nor_x2_sg U42000 ( .A(n42293), .B(n14001), .X(n13998) );
  inv_x4_sg U42001 ( .A(n41694), .X(n41695) );
  inv_x2_sg U42002 ( .A(n41696), .X(n41697) );
  nor_x2_sg U42003 ( .A(n42296), .B(n13221), .X(n13218) );
  inv_x4_sg U42004 ( .A(n41698), .X(n41699) );
  inv_x2_sg U42005 ( .A(n41700), .X(n41701) );
  nor_x2_sg U42006 ( .A(n42299), .B(n12440), .X(n12437) );
  nor_x8_sg U42007 ( .A(n46274), .B(n46281), .X(n20386) );
  nor_x8_sg U42008 ( .A(n46319), .B(n46326), .X(n18842) );
  nor_x8_sg U42009 ( .A(n46366), .B(n46373), .X(n17297) );
  inv_x4_sg U42010 ( .A(n18516), .X(n54186) );
  nand_x2_sg U42011 ( .A(n18478), .B(n18514), .X(n18516) );
  nor_x4_sg U42012 ( .A(n53509), .B(n53556), .X(n16775) );
  nor_x4_sg U42013 ( .A(n52951), .B(n52998), .X(n15209) );
  nor_x4_sg U42014 ( .A(n52117), .B(n52164), .X(n12876) );
  inv_x4_sg U42015 ( .A(n41702), .X(n41703) );
  inv_x4_sg U42016 ( .A(n41704), .X(n41705) );
  inv_x4_sg U42017 ( .A(n41706), .X(n41707) );
  inv_x4_sg U42018 ( .A(n41708), .X(n41709) );
  inv_x4_sg U42019 ( .A(n18239), .X(n41710) );
  inv_x4_sg U42020 ( .A(n41710), .X(n41711) );
  nor_x2_sg U42021 ( .A(n43161), .B(n28383), .X(n28380) );
  inv_x4_sg U42022 ( .A(n41712), .X(n41713) );
  inv_x2_sg U42023 ( .A(n41714), .X(n41715) );
  inv_x4_sg U42024 ( .A(n41716), .X(n41717) );
  inv_x2_sg U42025 ( .A(n41718), .X(n41719) );
  inv_x4_sg U42026 ( .A(n41720), .X(n41721) );
  inv_x2_sg U42027 ( .A(n41722), .X(n41723) );
  inv_x4_sg U42028 ( .A(n41724), .X(n41725) );
  inv_x2_sg U42029 ( .A(n41726), .X(n41727) );
  inv_x4_sg U42030 ( .A(n17223), .X(n53687) );
  nand_x2_sg U42031 ( .A(n17224), .B(n17167), .X(n17223) );
  inv_x4_sg U42032 ( .A(n15657), .X(n53129) );
  nand_x2_sg U42033 ( .A(n15658), .B(n15601), .X(n15657) );
  inv_x4_sg U42034 ( .A(n13324), .X(n52295) );
  nand_x2_sg U42035 ( .A(n13325), .B(n13268), .X(n13324) );
  inv_x4_sg U42036 ( .A(n12543), .X(n52019) );
  nand_x2_sg U42037 ( .A(n12544), .B(n12487), .X(n12543) );
  inv_x4_sg U42038 ( .A(n10329), .X(n41728) );
  inv_x4_sg U42039 ( .A(n18112), .X(n41730) );
  inv_x4_sg U42040 ( .A(n18224), .X(n41732) );
  nor_x8_sg U42041 ( .A(n46340), .B(n46346), .X(n18224) );
  inv_x2_sg U42042 ( .A(n18224), .X(n54063) );
  nor_x2_sg U42043 ( .A(n54053), .B(n54046), .X(n28449) );
  nor_x2_sg U42044 ( .A(n55456), .B(n55408), .X(n29411) );
  nor_x2_sg U42045 ( .A(n55408), .B(n55403), .X(n29421) );
  inv_x4_sg U42046 ( .A(n21796), .X(n55408) );
  nor_x2_sg U42047 ( .A(n55172), .B(n55123), .X(n29129) );
  nor_x2_sg U42048 ( .A(n55123), .B(n55118), .X(n29139) );
  inv_x4_sg U42049 ( .A(n21025), .X(n55123) );
  nor_x2_sg U42050 ( .A(n54888), .B(n54840), .X(n28850) );
  nor_x2_sg U42051 ( .A(n54840), .B(n54835), .X(n28860) );
  inv_x4_sg U42052 ( .A(n20251), .X(n54840) );
  nor_x2_sg U42053 ( .A(n54604), .B(n54555), .X(n28570) );
  nor_x2_sg U42054 ( .A(n54555), .B(n54550), .X(n28580) );
  inv_x4_sg U42055 ( .A(n19481), .X(n54555) );
  nor_x2_sg U42056 ( .A(n54320), .B(n54273), .X(n28292) );
  nor_x2_sg U42057 ( .A(n54273), .B(n54268), .X(n28302) );
  inv_x4_sg U42058 ( .A(n18705), .X(n54273) );
  nor_x2_sg U42059 ( .A(n54039), .B(n53990), .X(n28012) );
  nor_x2_sg U42060 ( .A(n53990), .B(n53985), .X(n28022) );
  inv_x4_sg U42061 ( .A(n17936), .X(n53990) );
  nor_x2_sg U42062 ( .A(n52919), .B(n52870), .X(n26893) );
  nor_x2_sg U42063 ( .A(n52870), .B(n52865), .X(n26903) );
  inv_x4_sg U42064 ( .A(n14815), .X(n52870) );
  nor_x2_sg U42065 ( .A(n55437), .B(n55424), .X(n21634) );
  nor_x2_sg U42066 ( .A(n21242), .B(n55424), .X(n21241) );
  inv_x4_sg U42067 ( .A(n21636), .X(n55424) );
  nor_x2_sg U42068 ( .A(n54869), .B(n54856), .X(n20089) );
  nor_x2_sg U42069 ( .A(n19697), .B(n54856), .X(n19696) );
  inv_x4_sg U42070 ( .A(n20091), .X(n54856) );
  nor_x2_sg U42071 ( .A(n54301), .B(n54288), .X(n18544) );
  nor_x2_sg U42072 ( .A(n18152), .B(n54288), .X(n18151) );
  inv_x4_sg U42073 ( .A(n18546), .X(n54288) );
  nor_x2_sg U42074 ( .A(n53737), .B(n53725), .X(n17005) );
  nor_x2_sg U42075 ( .A(n16598), .B(n53725), .X(n16597) );
  inv_x4_sg U42076 ( .A(n17007), .X(n53725) );
  nor_x2_sg U42077 ( .A(n53179), .B(n53167), .X(n15439) );
  nor_x2_sg U42078 ( .A(n15032), .B(n53167), .X(n15031) );
  inv_x4_sg U42079 ( .A(n15441), .X(n53167) );
  nor_x2_sg U42080 ( .A(n52620), .B(n52608), .X(n13886) );
  nor_x2_sg U42081 ( .A(n13483), .B(n52608), .X(n13482) );
  inv_x4_sg U42082 ( .A(n13888), .X(n52608) );
  nor_x2_sg U42083 ( .A(n52345), .B(n52333), .X(n13106) );
  nor_x2_sg U42084 ( .A(n12699), .B(n52333), .X(n12698) );
  inv_x4_sg U42085 ( .A(n13108), .X(n52333) );
  nor_x2_sg U42086 ( .A(n52068), .B(n52056), .X(n12325) );
  nor_x2_sg U42087 ( .A(n11921), .B(n52056), .X(n11920) );
  inv_x4_sg U42088 ( .A(n12327), .X(n52056) );
  nor_x2_sg U42089 ( .A(n51789), .B(n51776), .X(n11545) );
  nor_x2_sg U42090 ( .A(n11138), .B(n51776), .X(n11137) );
  inv_x4_sg U42091 ( .A(n11547), .X(n51776) );
  inv_x4_sg U42092 ( .A(n41733), .X(n41734) );
  nor_x2_sg U42093 ( .A(n43171), .B(n46473), .X(n13619) );
  inv_x4_sg U42094 ( .A(n41735), .X(n41736) );
  inv_x4_sg U42095 ( .A(n41737), .X(n41738) );
  inv_x4_sg U42096 ( .A(n41739), .X(n41740) );
  inv_x4_sg U42097 ( .A(n41741), .X(n41742) );
  nor_x2_sg U42098 ( .A(n51392), .B(n11006), .X(n11005) );
  inv_x4_sg U42099 ( .A(n41743), .X(n41744) );
  inv_x4_sg U42100 ( .A(n41745), .X(n41746) );
  inv_x4_sg U42101 ( .A(n41747), .X(n41748) );
  inv_x4_sg U42102 ( .A(n41749), .X(n41750) );
  inv_x4_sg U42103 ( .A(n41751), .X(n41752) );
  inv_x4_sg U42104 ( .A(n41753), .X(n41754) );
  inv_x4_sg U42105 ( .A(n41755), .X(n41756) );
  inv_x4_sg U42106 ( .A(n41757), .X(n41758) );
  inv_x4_sg U42107 ( .A(n41759), .X(n41760) );
  inv_x4_sg U42108 ( .A(n41761), .X(n41762) );
  nor_x2_sg U42109 ( .A(n21703), .B(n21701), .X(n21880) );
  nor_x2_sg U42110 ( .A(n55316), .B(n21882), .X(n21881) );
  inv_x4_sg U42111 ( .A(n41763), .X(n41764) );
  nor_x2_sg U42112 ( .A(n20158), .B(n20156), .X(n20335) );
  nor_x2_sg U42113 ( .A(n54748), .B(n20337), .X(n20336) );
  inv_x4_sg U42114 ( .A(n41765), .X(n41766) );
  nor_x2_sg U42115 ( .A(n18612), .B(n18610), .X(n18791) );
  nor_x2_sg U42116 ( .A(n54181), .B(n18793), .X(n18792) );
  inv_x4_sg U42117 ( .A(n41767), .X(n41768) );
  inv_x4_sg U42118 ( .A(n41769), .X(n41770) );
  inv_x4_sg U42119 ( .A(n41771), .X(n41772) );
  inv_x4_sg U42120 ( .A(n41773), .X(n41774) );
  inv_x4_sg U42121 ( .A(n41775), .X(n41776) );
  inv_x4_sg U42122 ( .A(n41777), .X(n41778) );
  inv_x4_sg U42123 ( .A(n41779), .X(n41780) );
  nor_x2_sg U42124 ( .A(n21111), .B(n21112), .X(n21110) );
  inv_x4_sg U42125 ( .A(n41781), .X(n41782) );
  nor_x2_sg U42126 ( .A(n19567), .B(n19568), .X(n19566) );
  inv_x4_sg U42127 ( .A(n41783), .X(n41784) );
  nor_x2_sg U42128 ( .A(n18022), .B(n18023), .X(n18021) );
  inv_x4_sg U42129 ( .A(n41785), .X(n41786) );
  inv_x4_sg U42130 ( .A(n41787), .X(n41788) );
  inv_x4_sg U42131 ( .A(n41789), .X(n41790) );
  inv_x4_sg U42132 ( .A(n41791), .X(n41792) );
  inv_x4_sg U42133 ( .A(n41793), .X(n41794) );
  inv_x4_sg U42134 ( .A(n41795), .X(n41796) );
  inv_x4_sg U42135 ( .A(n41797), .X(n41798) );
  inv_x4_sg U42136 ( .A(n41799), .X(n41800) );
  inv_x4_sg U42137 ( .A(n41801), .X(n41802) );
  inv_x4_sg U42138 ( .A(n41803), .X(n41804) );
  inv_x4_sg U42139 ( .A(n15974), .X(n53288) );
  nand_x2_sg U42140 ( .A(n15975), .B(n53287), .X(n15974) );
  inv_x4_sg U42141 ( .A(n41805), .X(n41806) );
  inv_x4_sg U42142 ( .A(n13640), .X(n52455) );
  nand_x2_sg U42143 ( .A(n13641), .B(n52454), .X(n13640) );
  inv_x4_sg U42144 ( .A(n41807), .X(n41808) );
  inv_x4_sg U42145 ( .A(n12079), .X(n51903) );
  nand_x2_sg U42146 ( .A(n12080), .B(n51902), .X(n12079) );
  inv_x4_sg U42147 ( .A(n41809), .X(n41810) );
  inv_x4_sg U42148 ( .A(n11299), .X(n51621) );
  nand_x2_sg U42149 ( .A(n11300), .B(n51620), .X(n11299) );
  nor_x4_sg U42150 ( .A(n13618), .B(n52443), .X(n13614) );
  nor_x4_sg U42151 ( .A(n41806), .B(n52455), .X(n13618) );
  inv_x4_sg U42152 ( .A(n41811), .X(n41812) );
  inv_x4_sg U42153 ( .A(n41813), .X(n41814) );
  inv_x4_sg U42154 ( .A(n41815), .X(n41816) );
  inv_x4_sg U42155 ( .A(n41817), .X(n41818) );
  inv_x4_sg U42156 ( .A(n41819), .X(n41820) );
  inv_x4_sg U42157 ( .A(n41821), .X(n41822) );
  nand_x8_sg U42158 ( .A(n10919), .B(n25505), .X(n25520) );
  nand_x8_sg U42159 ( .A(n17162), .B(n27739), .X(n27755) );
  nand_x8_sg U42160 ( .A(n16378), .B(n27458), .X(n27474) );
  nand_x8_sg U42161 ( .A(n15596), .B(n27179), .X(n27197) );
  nand_x8_sg U42162 ( .A(n14043), .B(n26622), .X(n26638) );
  nand_x8_sg U42163 ( .A(n13263), .B(n26343), .X(n26360) );
  nand_x8_sg U42164 ( .A(n12482), .B(n26062), .X(n26081) );
  nand_x8_sg U42165 ( .A(n11703), .B(n25783), .X(n25799) );
  inv_x8_sg U42166 ( .A(n31415), .X(n49492) );
  nand_x4_sg U42167 ( .A(n8357), .B(n31416), .X(n31415) );
  nor_x8_sg U42168 ( .A(n25140), .B(n31279), .X(n31414) );
  inv_x8_sg U42169 ( .A(n31406), .X(n49632) );
  nand_x4_sg U42170 ( .A(n8354), .B(n31407), .X(n31406) );
  nor_x8_sg U42171 ( .A(n24995), .B(n31297), .X(n31405) );
  inv_x8_sg U42172 ( .A(n23749), .X(n50351) );
  nand_x4_sg U42173 ( .A(n8657), .B(n23750), .X(n23749) );
  nor_x8_sg U42174 ( .A(n10032), .B(n23613), .X(n23748) );
  inv_x8_sg U42175 ( .A(n23740), .X(n50491) );
  nand_x4_sg U42176 ( .A(n8654), .B(n23741), .X(n23740) );
  nor_x8_sg U42177 ( .A(n9887), .B(n23631), .X(n23739) );
  inv_x4_sg U42178 ( .A(n41823), .X(n41824) );
  inv_x4_sg U42179 ( .A(n41825), .X(n41826) );
  inv_x4_sg U42180 ( .A(n41827), .X(n41828) );
  inv_x4_sg U42181 ( .A(n41829), .X(n41830) );
  nand_x8_sg U42182 ( .A(n49249), .B(n32067), .X(n25379) );
  nand_x2_sg U42183 ( .A(n8482), .B(n40725), .X(n32067) );
  nand_x8_sg U42184 ( .A(n50108), .B(n24401), .X(n10273) );
  nand_x2_sg U42185 ( .A(n8782), .B(n40726), .X(n24401) );
  inv_x8_sg U42186 ( .A(n42630), .X(n42631) );
  inv_x8_sg U42187 ( .A(n42632), .X(n42633) );
  inv_x8_sg U42188 ( .A(n42634), .X(n42635) );
  inv_x8_sg U42189 ( .A(n42636), .X(n42637) );
  inv_x8_sg U42190 ( .A(n42638), .X(n42639) );
  inv_x8_sg U42191 ( .A(n42640), .X(n42641) );
  inv_x8_sg U42192 ( .A(n42642), .X(n42643) );
  inv_x8_sg U42193 ( .A(n42644), .X(n42645) );
  inv_x8_sg U42194 ( .A(n42646), .X(n42647) );
  inv_x8_sg U42195 ( .A(n42648), .X(n42649) );
  inv_x8_sg U42196 ( .A(n42650), .X(n42651) );
  inv_x8_sg U42197 ( .A(n42652), .X(n42653) );
  inv_x8_sg U42198 ( .A(n42654), .X(n42655) );
  inv_x8_sg U42199 ( .A(n42656), .X(n42657) );
  inv_x8_sg U42200 ( .A(n42658), .X(n42659) );
  inv_x8_sg U42201 ( .A(n42660), .X(n42661) );
  inv_x8_sg U42202 ( .A(n42662), .X(n42663) );
  inv_x8_sg U42203 ( .A(n42664), .X(n42665) );
  inv_x8_sg U42204 ( .A(n42666), .X(n42667) );
  inv_x8_sg U42205 ( .A(n42668), .X(n42669) );
  inv_x8_sg U42206 ( .A(n42670), .X(n42671) );
  inv_x8_sg U42207 ( .A(n42674), .X(n42675) );
  inv_x8_sg U42208 ( .A(n42678), .X(n42679) );
  inv_x8_sg U42209 ( .A(n42702), .X(n42703) );
  inv_x8_sg U42210 ( .A(n42704), .X(n42705) );
  inv_x8_sg U42211 ( .A(n42706), .X(n42707) );
  inv_x8_sg U42212 ( .A(n42708), .X(n42709) );
  inv_x8_sg U42213 ( .A(n42710), .X(n42711) );
  inv_x8_sg U42214 ( .A(n42712), .X(n42713) );
  inv_x8_sg U42215 ( .A(n42714), .X(n42715) );
  inv_x8_sg U42216 ( .A(n42716), .X(n42717) );
  inv_x8_sg U42217 ( .A(n42718), .X(n42719) );
  inv_x8_sg U42218 ( .A(n42720), .X(n42721) );
  inv_x8_sg U42219 ( .A(n42722), .X(n42723) );
  inv_x8_sg U42220 ( .A(n42724), .X(n42725) );
  inv_x8_sg U42221 ( .A(n42726), .X(n42727) );
  inv_x8_sg U42222 ( .A(n42728), .X(n42729) );
  inv_x8_sg U42223 ( .A(n42730), .X(n42731) );
  inv_x8_sg U42224 ( .A(n42732), .X(n42733) );
  inv_x8_sg U42225 ( .A(n42734), .X(n42735) );
  inv_x8_sg U42226 ( .A(n42736), .X(n42737) );
  inv_x8_sg U42227 ( .A(n42738), .X(n42739) );
  inv_x8_sg U42228 ( .A(n42740), .X(n42741) );
  inv_x8_sg U42229 ( .A(n42742), .X(n42743) );
  inv_x8_sg U42230 ( .A(n42746), .X(n42747) );
  inv_x8_sg U42231 ( .A(n42750), .X(n42751) );
  inv_x8_sg U42232 ( .A(n42772), .X(n42773) );
  inv_x8_sg U42233 ( .A(n42774), .X(n42775) );
  inv_x8_sg U42234 ( .A(n42776), .X(n42777) );
  inv_x8_sg U42235 ( .A(n42778), .X(n42779) );
  inv_x8_sg U42236 ( .A(n42782), .X(n42783) );
  inv_x8_sg U42237 ( .A(n42784), .X(n42785) );
  inv_x8_sg U42238 ( .A(n42786), .X(n42787) );
  inv_x8_sg U42239 ( .A(n42788), .X(n42789) );
  inv_x8_sg U42240 ( .A(n44656), .X(n44657) );
  inv_x4_sg U42241 ( .A(n24134), .X(n44656) );
  nor_x2_sg U42242 ( .A(n24136), .B(n50544), .X(n24134) );
  inv_x8_sg U42243 ( .A(n45508), .X(n45509) );
  inv_x4_sg U42244 ( .A(n24141), .X(n45508) );
  nor_x2_sg U42245 ( .A(n24170), .B(n50591), .X(n24141) );
  inv_x8_sg U42246 ( .A(n45500), .X(n45501) );
  inv_x4_sg U42247 ( .A(n23997), .X(n45500) );
  nor_x2_sg U42248 ( .A(n24026), .B(n50603), .X(n23997) );
  inv_x8_sg U42249 ( .A(n45506), .X(n45507) );
  inv_x4_sg U42250 ( .A(n23844), .X(n45506) );
  nor_x2_sg U42251 ( .A(n23873), .B(n50649), .X(n23844) );
  inv_x8_sg U42252 ( .A(n45498), .X(n45499) );
  inv_x4_sg U42253 ( .A(n23673), .X(n45498) );
  nor_x2_sg U42254 ( .A(n23702), .B(n50694), .X(n23673) );
  inv_x8_sg U42255 ( .A(n45504), .X(n45505) );
  inv_x4_sg U42256 ( .A(n23483), .X(n45504) );
  nor_x2_sg U42257 ( .A(n23512), .B(n50740), .X(n23483) );
  inv_x8_sg U42258 ( .A(n45496), .X(n45497) );
  inv_x4_sg U42259 ( .A(n23278), .X(n45496) );
  nor_x2_sg U42260 ( .A(n23307), .B(n50786), .X(n23278) );
  inv_x8_sg U42261 ( .A(n45502), .X(n45503) );
  inv_x4_sg U42262 ( .A(n23052), .X(n45502) );
  nor_x2_sg U42263 ( .A(n23081), .B(n50830), .X(n23052) );
  inv_x8_sg U42264 ( .A(n44665), .X(n44666) );
  inv_x4_sg U42265 ( .A(n31800), .X(n44665) );
  nor_x2_sg U42266 ( .A(n31802), .B(n49685), .X(n31800) );
  inv_x8_sg U42267 ( .A(n45522), .X(n45523) );
  inv_x4_sg U42268 ( .A(n31807), .X(n45522) );
  nor_x2_sg U42269 ( .A(n31836), .B(n49732), .X(n31807) );
  inv_x8_sg U42270 ( .A(n45520), .X(n45521) );
  inv_x4_sg U42271 ( .A(n31510), .X(n45520) );
  nor_x2_sg U42272 ( .A(n31539), .B(n49790), .X(n31510) );
  inv_x8_sg U42273 ( .A(n45518), .X(n45519) );
  inv_x4_sg U42274 ( .A(n31149), .X(n45518) );
  nor_x2_sg U42275 ( .A(n31178), .B(n49881), .X(n31149) );
  inv_x8_sg U42276 ( .A(n45516), .X(n45517) );
  inv_x4_sg U42277 ( .A(n30718), .X(n45516) );
  nor_x2_sg U42278 ( .A(n30747), .B(n49971), .X(n30718) );
  inv_x8_sg U42279 ( .A(n45512), .X(n45513) );
  inv_x4_sg U42280 ( .A(n31339), .X(n45512) );
  nor_x2_sg U42281 ( .A(n31368), .B(n49835), .X(n31339) );
  inv_x8_sg U42282 ( .A(n45510), .X(n45511) );
  inv_x4_sg U42283 ( .A(n30944), .X(n45510) );
  nor_x2_sg U42284 ( .A(n30973), .B(n49927), .X(n30944) );
  inv_x8_sg U42285 ( .A(n45514), .X(n45515) );
  inv_x4_sg U42286 ( .A(n31663), .X(n45514) );
  nor_x2_sg U42287 ( .A(n31692), .B(n49744), .X(n31663) );
  inv_x8_sg U42288 ( .A(n45526), .X(n45527) );
  inv_x4_sg U42289 ( .A(n30463), .X(n45526) );
  nor_x2_sg U42290 ( .A(n30492), .B(n50015), .X(n30463) );
  inv_x8_sg U42291 ( .A(n45524), .X(n45525) );
  inv_x4_sg U42292 ( .A(n22797), .X(n45524) );
  nor_x2_sg U42293 ( .A(n22826), .B(n50874), .X(n22797) );
  inv_x4_sg U42294 ( .A(n41831), .X(n41832) );
  nor_x4_sg U42295 ( .A(n41832), .B(n55244), .X(n21368) );
  inv_x4_sg U42296 ( .A(n21378), .X(n55244) );
  nand_x2_sg U42297 ( .A(n42691), .B(n41514), .X(n21378) );
  inv_x4_sg U42298 ( .A(n41833), .X(n41834) );
  nor_x4_sg U42299 ( .A(n41834), .B(n54972), .X(n20597) );
  inv_x4_sg U42300 ( .A(n20607), .X(n54972) );
  nand_x2_sg U42301 ( .A(n42693), .B(n41183), .X(n20607) );
  inv_x4_sg U42302 ( .A(n41835), .X(n41836) );
  nor_x4_sg U42303 ( .A(n41836), .B(n54676), .X(n19823) );
  inv_x4_sg U42304 ( .A(n19833), .X(n54676) );
  nand_x2_sg U42305 ( .A(n42695), .B(n41518), .X(n19833) );
  inv_x4_sg U42306 ( .A(n41837), .X(n41838) );
  nor_x4_sg U42307 ( .A(n41838), .B(n54404), .X(n19053) );
  inv_x4_sg U42308 ( .A(n19063), .X(n54404) );
  nand_x2_sg U42309 ( .A(n42697), .B(n41185), .X(n19063) );
  inv_x4_sg U42310 ( .A(n41839), .X(n41840) );
  nor_x4_sg U42311 ( .A(n41840), .B(n53839), .X(n17508) );
  inv_x4_sg U42312 ( .A(n17518), .X(n53839) );
  nand_x2_sg U42313 ( .A(n42699), .B(n41187), .X(n17518) );
  inv_x4_sg U42314 ( .A(n41841), .X(n41842) );
  nor_x4_sg U42315 ( .A(n41842), .B(n52712), .X(n14387) );
  inv_x4_sg U42316 ( .A(n14397), .X(n52712) );
  nand_x2_sg U42317 ( .A(n42701), .B(n41189), .X(n14397) );
  inv_x4_sg U42318 ( .A(n41843), .X(n41844) );
  nor_x4_sg U42319 ( .A(n41844), .B(n51322), .X(n10496) );
  inv_x4_sg U42320 ( .A(n10506), .X(n51322) );
  nand_x2_sg U42321 ( .A(n41215), .B(n41147), .X(n10506) );
  nor_x4_sg U42322 ( .A(n18277), .B(n18280), .X(n18281) );
  inv_x4_sg U42323 ( .A(n13829), .X(n41845) );
  inv_x4_sg U42324 ( .A(n41845), .X(n41846) );
  inv_x4_sg U42325 ( .A(n41847), .X(n41848) );
  nor_x4_sg U42326 ( .A(n50101), .B(n41848), .X(n29611) );
  inv_x4_sg U42327 ( .A(n30175), .X(n50101) );
  nand_x2_sg U42328 ( .A(n30174), .B(n41484), .X(n30175) );
  inv_x4_sg U42329 ( .A(n41849), .X(n41850) );
  nor_x4_sg U42330 ( .A(n50105), .B(n41850), .X(n29602) );
  inv_x4_sg U42331 ( .A(n29646), .X(n50105) );
  nand_x2_sg U42332 ( .A(n29645), .B(n41482), .X(n29646) );
  inv_x4_sg U42333 ( .A(n41851), .X(n41852) );
  nor_x4_sg U42334 ( .A(n50960), .B(n41852), .X(n21955) );
  inv_x4_sg U42335 ( .A(n22509), .X(n50960) );
  nand_x2_sg U42336 ( .A(n22508), .B(n41488), .X(n22509) );
  inv_x4_sg U42337 ( .A(n41853), .X(n41854) );
  nor_x4_sg U42338 ( .A(n50964), .B(n41854), .X(n21948) );
  inv_x4_sg U42339 ( .A(n21981), .X(n50964) );
  nand_x2_sg U42340 ( .A(n21980), .B(n41486), .X(n21981) );
  nor_x4_sg U42341 ( .A(n15952), .B(n53279), .X(n15948) );
  nor_x4_sg U42342 ( .A(n41804), .B(n53288), .X(n15952) );
  nor_x4_sg U42343 ( .A(n16738), .B(n53561), .X(n16734) );
  nor_x4_sg U42344 ( .A(n15172), .B(n53003), .X(n15168) );
  nor_x4_sg U42345 ( .A(n12839), .B(n52169), .X(n12835) );
  nor_x4_sg U42346 ( .A(n12057), .B(n51892), .X(n12053) );
  nor_x4_sg U42347 ( .A(n41808), .B(n51903), .X(n12057) );
  nor_x4_sg U42348 ( .A(n11278), .B(n51611), .X(n11274) );
  nor_x4_sg U42349 ( .A(n41810), .B(n51621), .X(n11278) );
  nor_x4_sg U42350 ( .A(n50073), .B(n30446), .X(n24502) );
  inv_x4_sg U42351 ( .A(n30448), .X(n50073) );
  nand_x2_sg U42352 ( .A(n30447), .B(n24499), .X(n30448) );
  nor_x4_sg U42353 ( .A(n24499), .B(n30447), .X(n30446) );
  nor_x4_sg U42354 ( .A(n50083), .B(n29841), .X(n24495) );
  inv_x4_sg U42355 ( .A(n29843), .X(n50083) );
  nand_x2_sg U42356 ( .A(n29842), .B(n24523), .X(n29843) );
  nor_x4_sg U42357 ( .A(n24523), .B(n29842), .X(n29841) );
  nor_x4_sg U42358 ( .A(n50932), .B(n22780), .X(n9388) );
  inv_x4_sg U42359 ( .A(n22782), .X(n50932) );
  nand_x2_sg U42360 ( .A(n22781), .B(n9384), .X(n22782) );
  nor_x4_sg U42361 ( .A(n9384), .B(n22781), .X(n22780) );
  nor_x4_sg U42362 ( .A(n50942), .B(n22176), .X(n9380) );
  inv_x4_sg U42363 ( .A(n22178), .X(n50942) );
  nand_x2_sg U42364 ( .A(n22177), .B(n9414), .X(n22178) );
  nor_x4_sg U42365 ( .A(n9414), .B(n22177), .X(n22176) );
  inv_x4_sg U42366 ( .A(n24649), .X(n49941) );
  inv_x4_sg U42367 ( .A(n24600), .X(n49986) );
  inv_x4_sg U42368 ( .A(n24551), .X(n50031) );
  inv_x4_sg U42369 ( .A(n9541), .X(n50800) );
  inv_x4_sg U42370 ( .A(n9492), .X(n50845) );
  inv_x4_sg U42371 ( .A(n9443), .X(n50890) );
  nand_x4_sg U42372 ( .A(n53458), .B(n15808), .X(n16222) );
  nand_x4_sg U42373 ( .A(n42849), .B(n16277), .X(n15808) );
  nor_x1_sg U42374 ( .A(n53387), .B(n16133), .X(n16127) );
  inv_x4_sg U42375 ( .A(n16431), .X(n41865) );
  nor_x1_sg U42376 ( .A(n53666), .B(n16918), .X(n16912) );
  nor_x1_sg U42377 ( .A(n53108), .B(n15352), .X(n15346) );
  nor_x1_sg U42378 ( .A(n52549), .B(n13799), .X(n13793) );
  nor_x1_sg U42379 ( .A(n52274), .B(n13019), .X(n13013) );
  nor_x1_sg U42380 ( .A(n51998), .B(n12238), .X(n12232) );
  nor_x1_sg U42381 ( .A(n51720), .B(n11458), .X(n11452) );
  inv_x4_sg U42382 ( .A(n11757), .X(n41867) );
  nand_x4_sg U42383 ( .A(n14190), .B(n14280), .X(n14197) );
  inv_x4_sg U42384 ( .A(n10443), .X(n41870) );
  nor_x8_sg U42385 ( .A(n46565), .B(n46570), .X(n10443) );
  inv_x2_sg U42386 ( .A(n10443), .X(n51277) );
  inv_x4_sg U42387 ( .A(n18204), .X(n41871) );
  nor_x8_sg U42388 ( .A(n46340), .B(n46341), .X(n18204) );
  inv_x2_sg U42389 ( .A(n18204), .X(n54064) );
  inv_x2_sg U42390 ( .A(n50183), .X(n41872) );
  inv_x8_sg U42391 ( .A(n24320), .X(n50183) );
  inv_x2_sg U42392 ( .A(n49324), .X(n41873) );
  inv_x8_sg U42393 ( .A(n31986), .X(n49324) );
  inv_x4_sg U42394 ( .A(n41874), .X(n41875) );
  inv_x4_sg U42395 ( .A(n41876), .X(n41877) );
  inv_x4_sg U42396 ( .A(n41878), .X(n41879) );
  inv_x4_sg U42397 ( .A(n41880), .X(n41881) );
  inv_x4_sg U42398 ( .A(n41882), .X(n41883) );
  nand_x4_sg U42399 ( .A(n10447), .B(n42853), .X(n10444) );
  inv_x1_sg U42400 ( .A(n21262), .X(n41884) );
  nand_x4_sg U42401 ( .A(n42627), .B(n41884), .X(n21173) );
  inv_x1_sg U42402 ( .A(n21262), .X(n55197) );
  nand_x4_sg U42403 ( .A(n18228), .B(n43139), .X(n18225) );
  nand_x4_sg U42404 ( .A(n42855), .B(n14339), .X(n14336) );
  nand_x4_sg U42405 ( .A(n55310), .B(n21195), .X(n9111) );
  nand_x4_sg U42406 ( .A(n55028), .B(n20422), .X(n9146) );
  nand_x4_sg U42407 ( .A(n54742), .B(n19650), .X(n9201) );
  nand_x4_sg U42408 ( .A(n54460), .B(n18878), .X(n9222) );
  nand_x4_sg U42409 ( .A(n53895), .B(n17333), .X(n9260) );
  nand_x4_sg U42410 ( .A(n53604), .B(n16550), .X(n9298) );
  nand_x4_sg U42411 ( .A(n53514), .B(n16527), .X(n9292) );
  nand_x4_sg U42412 ( .A(n53325), .B(n15768), .X(n9341) );
  nand_x4_sg U42413 ( .A(n53046), .B(n14984), .X(n8981) );
  nand_x4_sg U42414 ( .A(n52956), .B(n14961), .X(n8975) );
  nand_x4_sg U42415 ( .A(n52775), .B(n14214), .X(n8956) );
  nand_x4_sg U42416 ( .A(n14190), .B(n52675), .X(n8950) );
  nand_x4_sg U42417 ( .A(n43147), .B(n14192), .X(n14190) );
  nand_x4_sg U42418 ( .A(n52489), .B(n13435), .X(n8797) );
  nand_x4_sg U42419 ( .A(n52212), .B(n12651), .X(n8842) );
  nand_x4_sg U42420 ( .A(n51937), .B(n11873), .X(n8917) );
  nand_x4_sg U42421 ( .A(n51656), .B(n11090), .X(n8880) );
  nor_x2_sg U42422 ( .A(n25513), .B(n10907), .X(n25512) );
  nor_x4_sg U42423 ( .A(n46231), .B(n25508), .X(n25513) );
  inv_x4_sg U42424 ( .A(n41885), .X(n41886) );
  inv_x4_sg U42425 ( .A(n41887), .X(n41888) );
  inv_x1_sg U42426 ( .A(n21815), .X(n41889) );
  nand_x4_sg U42427 ( .A(n21816), .B(n21817), .X(n21815) );
  inv_x4_sg U42428 ( .A(n55434), .X(n41890) );
  inv_x4_sg U42429 ( .A(n41890), .X(n41891) );
  inv_x4_sg U42430 ( .A(n55149), .X(n41892) );
  inv_x4_sg U42431 ( .A(n41892), .X(n41893) );
  inv_x1_sg U42432 ( .A(n21044), .X(n41894) );
  nand_x4_sg U42433 ( .A(n21045), .B(n21046), .X(n21044) );
  inv_x1_sg U42434 ( .A(n20270), .X(n41895) );
  nand_x4_sg U42435 ( .A(n20271), .B(n20272), .X(n20270) );
  inv_x4_sg U42436 ( .A(n54866), .X(n41896) );
  inv_x4_sg U42437 ( .A(n41896), .X(n41897) );
  inv_x4_sg U42438 ( .A(n54581), .X(n41898) );
  inv_x4_sg U42439 ( .A(n41898), .X(n41899) );
  inv_x1_sg U42440 ( .A(n19500), .X(n41900) );
  nand_x4_sg U42441 ( .A(n19501), .B(n19502), .X(n19500) );
  inv_x1_sg U42442 ( .A(n18724), .X(n41901) );
  nand_x4_sg U42443 ( .A(n18725), .B(n18726), .X(n18724) );
  inv_x4_sg U42444 ( .A(n54298), .X(n41902) );
  inv_x4_sg U42445 ( .A(n41902), .X(n41903) );
  inv_x4_sg U42446 ( .A(n41904), .X(n41905) );
  inv_x4_sg U42447 ( .A(n54016), .X(n41906) );
  inv_x4_sg U42448 ( .A(n41906), .X(n41907) );
  inv_x1_sg U42449 ( .A(n17955), .X(n41908) );
  nand_x4_sg U42450 ( .A(n17956), .B(n17957), .X(n17955) );
  inv_x1_sg U42451 ( .A(n17182), .X(n41909) );
  nand_x4_sg U42452 ( .A(n17183), .B(n17184), .X(n17182) );
  inv_x1_sg U42453 ( .A(n15616), .X(n41910) );
  nand_x4_sg U42454 ( .A(n15617), .B(n15618), .X(n15616) );
  inv_x4_sg U42455 ( .A(n52896), .X(n41911) );
  inv_x4_sg U42456 ( .A(n41911), .X(n41912) );
  inv_x1_sg U42457 ( .A(n14834), .X(n41913) );
  nand_x4_sg U42458 ( .A(n14835), .B(n14836), .X(n14834) );
  inv_x1_sg U42459 ( .A(n14063), .X(n41914) );
  nand_x4_sg U42460 ( .A(n14064), .B(n14065), .X(n14063) );
  inv_x1_sg U42461 ( .A(n13283), .X(n41915) );
  nand_x4_sg U42462 ( .A(n13284), .B(n13285), .X(n13283) );
  inv_x1_sg U42463 ( .A(n12502), .X(n41916) );
  nand_x4_sg U42464 ( .A(n12503), .B(n12504), .X(n12502) );
  inv_x1_sg U42465 ( .A(n11722), .X(n41917) );
  nand_x4_sg U42466 ( .A(n11723), .B(n11724), .X(n11722) );
  inv_x4_sg U42467 ( .A(n51786), .X(n41918) );
  inv_x4_sg U42468 ( .A(n41918), .X(n41919) );
  inv_x4_sg U42469 ( .A(n51506), .X(n41920) );
  inv_x4_sg U42470 ( .A(n41920), .X(n41921) );
  inv_x4_sg U42471 ( .A(n41922), .X(n41923) );
  inv_x1_sg U42472 ( .A(n16397), .X(n41924) );
  nand_x4_sg U42473 ( .A(n16398), .B(n16399), .X(n16397) );
  inv_x1_sg U42474 ( .A(n10939), .X(n41925) );
  nand_x4_sg U42475 ( .A(n10940), .B(n10941), .X(n10939) );
  inv_x4_sg U42476 ( .A(n41926), .X(n41927) );
  inv_x4_sg U42477 ( .A(n41928), .X(n41929) );
  inv_x4_sg U42478 ( .A(n41930), .X(n41931) );
  inv_x4_sg U42479 ( .A(n41932), .X(n41933) );
  inv_x4_sg U42480 ( .A(n41934), .X(n41935) );
  inv_x4_sg U42481 ( .A(n21703), .X(n55331) );
  inv_x4_sg U42482 ( .A(n20158), .X(n54763) );
  inv_x4_sg U42483 ( .A(n18612), .X(n54196) );
  nor_x2_sg U42484 ( .A(n51413), .B(n51393), .X(n11004) );
  inv_x4_sg U42485 ( .A(n10832), .X(n51393) );
  inv_x4_sg U42486 ( .A(n16187), .X(n53342) );
  nor_x4_sg U42487 ( .A(n16190), .B(n46416), .X(n16187) );
  inv_x1_sg U42488 ( .A(n16709), .X(n41936) );
  nand_x4_sg U42489 ( .A(n16710), .B(n16708), .X(n16709) );
  inv_x1_sg U42490 ( .A(n15143), .X(n41937) );
  nand_x4_sg U42491 ( .A(n15144), .B(n15142), .X(n15143) );
  inv_x1_sg U42492 ( .A(n12810), .X(n41938) );
  nand_x4_sg U42493 ( .A(n12811), .B(n12809), .X(n12810) );
  inv_x4_sg U42494 ( .A(n11512), .X(n51673) );
  nor_x4_sg U42495 ( .A(n11515), .B(n46552), .X(n11512) );
  inv_x1_sg U42496 ( .A(n11249), .X(n41939) );
  nand_x4_sg U42497 ( .A(n11250), .B(n11248), .X(n11249) );
  inv_x4_sg U42498 ( .A(n20834), .X(n55038) );
  nor_x4_sg U42499 ( .A(n20837), .B(n46281), .X(n20834) );
  inv_x1_sg U42500 ( .A(n20576), .X(n41940) );
  nand_x4_sg U42501 ( .A(n20577), .B(n20575), .X(n20576) );
  inv_x4_sg U42502 ( .A(n19290), .X(n54470) );
  nor_x4_sg U42503 ( .A(n19293), .B(n46326), .X(n19290) );
  inv_x1_sg U42504 ( .A(n19032), .X(n41941) );
  nand_x4_sg U42505 ( .A(n19033), .B(n19031), .X(n19032) );
  inv_x4_sg U42506 ( .A(n17745), .X(n53905) );
  nor_x4_sg U42507 ( .A(n17748), .B(n46373), .X(n17745) );
  inv_x1_sg U42508 ( .A(n17487), .X(n41942) );
  nand_x4_sg U42509 ( .A(n17488), .B(n17486), .X(n17487) );
  inv_x4_sg U42510 ( .A(n14624), .X(n52785) );
  nor_x4_sg U42511 ( .A(n14627), .B(n46463), .X(n14624) );
  nand_x4_sg U42512 ( .A(n13898), .B(n13899), .X(n13845) );
  nand_x4_sg U42513 ( .A(n13907), .B(n13906), .X(n13899) );
  inv_x4_sg U42514 ( .A(n30688), .X(n41943) );
  inv_x4_sg U42515 ( .A(n30694), .X(n41945) );
  inv_x4_sg U42516 ( .A(n30700), .X(n41947) );
  inv_x4_sg U42517 ( .A(n23022), .X(n41949) );
  inv_x4_sg U42518 ( .A(n23028), .X(n41951) );
  inv_x4_sg U42519 ( .A(n23034), .X(n41953) );
  inv_x4_sg U42520 ( .A(n41955), .X(n41956) );
  inv_x4_sg U42521 ( .A(n41957), .X(n41958) );
  inv_x2_sg U42522 ( .A(n25235), .X(n41959) );
  inv_x2_sg U42523 ( .A(n10127), .X(n41960) );
  inv_x4_sg U42524 ( .A(n41961), .X(n41962) );
  inv_x4_sg U42525 ( .A(n41963), .X(n41964) );
  inv_x1_sg U42526 ( .A(n21227), .X(n42896) );
  inv_x1_sg U42527 ( .A(n20454), .X(n42900) );
  inv_x1_sg U42528 ( .A(n19682), .X(n42904) );
  inv_x1_sg U42529 ( .A(n18910), .X(n42908) );
  inv_x1_sg U42530 ( .A(n18137), .X(n42912) );
  inv_x1_sg U42531 ( .A(n17365), .X(n42916) );
  inv_x1_sg U42532 ( .A(n15801), .X(n42920) );
  inv_x1_sg U42533 ( .A(n14246), .X(n42924) );
  inv_x1_sg U42534 ( .A(n11122), .X(n42928) );
  inv_x1_sg U42535 ( .A(n10355), .X(n42932) );
  inv_x1_sg U42536 ( .A(n16344), .X(n42982) );
  inv_x1_sg U42537 ( .A(n10889), .X(n43010) );
  inv_x1_sg U42538 ( .A(n16366), .X(n43038) );
  inv_x1_sg U42539 ( .A(n21785), .X(n43052) );
  inv_x1_sg U42540 ( .A(n21014), .X(n43058) );
  inv_x1_sg U42541 ( .A(n20240), .X(n43060) );
  inv_x1_sg U42542 ( .A(n19470), .X(n43066) );
  inv_x1_sg U42543 ( .A(n18694), .X(n43068) );
  inv_x1_sg U42544 ( .A(n17925), .X(n43074) );
  inv_x1_sg U42545 ( .A(n17151), .X(n43076) );
  inv_x1_sg U42546 ( .A(n15585), .X(n43078) );
  inv_x1_sg U42547 ( .A(n14804), .X(n43082) );
  inv_x1_sg U42548 ( .A(n14032), .X(n43084) );
  inv_x1_sg U42549 ( .A(n13252), .X(n43086) );
  inv_x1_sg U42550 ( .A(n12471), .X(n43088) );
  inv_x1_sg U42551 ( .A(n11692), .X(n43090) );
  inv_x2_sg U42552 ( .A(n12366), .X(n43469) );
  inv_x2_sg U42553 ( .A(n13902), .X(n43477) );
  inv_x1_sg U42554 ( .A(n10404), .X(n43112) );
  inv_x1_sg U42555 ( .A(n21276), .X(n43116) );
  inv_x1_sg U42556 ( .A(n19731), .X(n43120) );
  inv_x1_sg U42557 ( .A(n15843), .X(n43144) );
  inv_x1_sg U42558 ( .A(n19725), .X(n43150) );
  inv_x1_sg U42559 ( .A(n13510), .X(n43154) );
  inv_x1_sg U42560 ( .A(n11948), .X(n43158) );
  inv_x1_sg U42561 ( .A(n26968), .X(n43164) );
  inv_x2_sg U42562 ( .A(reg_num[0]), .X(n43264) );
  inv_x4_sg U42563 ( .A(n41965), .X(n41966) );
  nor_x2_sg U42564 ( .A(n21189), .B(n55251), .X(n21187) );
  inv_x4_sg U42565 ( .A(n21190), .X(n55251) );
  inv_x4_sg U42566 ( .A(n41967), .X(n41968) );
  nor_x2_sg U42567 ( .A(n20416), .B(n54966), .X(n20414) );
  inv_x4_sg U42568 ( .A(n20417), .X(n54966) );
  inv_x4_sg U42569 ( .A(n41969), .X(n41970) );
  nor_x2_sg U42570 ( .A(n19644), .B(n54683), .X(n19642) );
  inv_x4_sg U42571 ( .A(n19645), .X(n54683) );
  inv_x4_sg U42572 ( .A(n41971), .X(n41972) );
  nor_x2_sg U42573 ( .A(n18872), .B(n54398), .X(n18870) );
  inv_x4_sg U42574 ( .A(n18873), .X(n54398) );
  inv_x4_sg U42575 ( .A(n41973), .X(n41974) );
  nor_x2_sg U42576 ( .A(n17327), .B(n53833), .X(n17325) );
  inv_x4_sg U42577 ( .A(n17328), .X(n53833) );
  inv_x4_sg U42578 ( .A(n41975), .X(n41976) );
  inv_x2_sg U42579 ( .A(n41977), .X(n41978) );
  inv_x4_sg U42580 ( .A(n41979), .X(n41980) );
  inv_x2_sg U42581 ( .A(n41981), .X(n41982) );
  inv_x4_sg U42582 ( .A(n41983), .X(n41984) );
  inv_x2_sg U42583 ( .A(n41985), .X(n41986) );
  inv_x4_sg U42584 ( .A(n41987), .X(n41988) );
  nor_x2_sg U42585 ( .A(n14208), .B(n52719), .X(n14206) );
  inv_x4_sg U42586 ( .A(n14209), .X(n52719) );
  inv_x4_sg U42587 ( .A(n41989), .X(n41990) );
  inv_x2_sg U42588 ( .A(n41991), .X(n41992) );
  inv_x4_sg U42589 ( .A(n41993), .X(n41994) );
  inv_x2_sg U42590 ( .A(n41995), .X(n41996) );
  inv_x4_sg U42591 ( .A(n41997), .X(n41998) );
  inv_x2_sg U42592 ( .A(n41999), .X(n42000) );
  inv_x4_sg U42593 ( .A(n42001), .X(n42002) );
  inv_x2_sg U42594 ( .A(n42003), .X(n42004) );
  inv_x4_sg U42595 ( .A(n42005), .X(n42006) );
  nor_x2_sg U42596 ( .A(n10316), .B(n51329), .X(n10314) );
  inv_x4_sg U42597 ( .A(n10317), .X(n51329) );
  inv_x4_sg U42598 ( .A(n42007), .X(n42008) );
  inv_x2_sg U42599 ( .A(n42009), .X(n42010) );
  inv_x4_sg U42600 ( .A(n42011), .X(n42012) );
  inv_x2_sg U42601 ( .A(n42013), .X(n42014) );
  inv_x4_sg U42602 ( .A(n42015), .X(n42016) );
  inv_x2_sg U42603 ( .A(n42017), .X(n42018) );
  inv_x4_sg U42604 ( .A(n42019), .X(n42020) );
  inv_x2_sg U42605 ( .A(n42021), .X(n42022) );
  inv_x4_sg U42606 ( .A(n42023), .X(n42024) );
  inv_x2_sg U42607 ( .A(n42025), .X(n42026) );
  inv_x4_sg U42608 ( .A(n42027), .X(n42028) );
  nor_x2_sg U42609 ( .A(n42953), .B(n21759), .X(n21757) );
  inv_x4_sg U42610 ( .A(n42029), .X(n42030) );
  nor_x2_sg U42611 ( .A(n42957), .B(n20989), .X(n20987) );
  inv_x4_sg U42612 ( .A(n42031), .X(n42032) );
  nor_x2_sg U42613 ( .A(n42961), .B(n20214), .X(n20212) );
  inv_x4_sg U42614 ( .A(n42033), .X(n42034) );
  nor_x2_sg U42615 ( .A(n42965), .B(n19445), .X(n19443) );
  inv_x4_sg U42616 ( .A(n42035), .X(n42036) );
  nor_x2_sg U42617 ( .A(n42969), .B(n18669), .X(n18667) );
  inv_x4_sg U42618 ( .A(n42037), .X(n42038) );
  nor_x2_sg U42619 ( .A(n42973), .B(n17900), .X(n17898) );
  inv_x4_sg U42620 ( .A(n42039), .X(n42040) );
  nor_x2_sg U42621 ( .A(n42977), .B(n17127), .X(n17125) );
  inv_x4_sg U42622 ( .A(n42041), .X(n42042) );
  nor_x2_sg U42623 ( .A(n42985), .B(n15561), .X(n15559) );
  inv_x4_sg U42624 ( .A(n42043), .X(n42044) );
  nor_x2_sg U42625 ( .A(n42989), .B(n14779), .X(n14777) );
  inv_x4_sg U42626 ( .A(n42045), .X(n42046) );
  nor_x2_sg U42627 ( .A(n42993), .B(n14008), .X(n14006) );
  inv_x4_sg U42628 ( .A(n42047), .X(n42048) );
  nor_x2_sg U42629 ( .A(n42997), .B(n13228), .X(n13226) );
  inv_x4_sg U42630 ( .A(n42049), .X(n42050) );
  nor_x2_sg U42631 ( .A(n43001), .B(n12447), .X(n12445) );
  inv_x4_sg U42632 ( .A(n42051), .X(n42052) );
  nor_x2_sg U42633 ( .A(n43005), .B(n11667), .X(n11665) );
  inv_x4_sg U42634 ( .A(n10973), .X(n42053) );
  inv_x2_sg U42635 ( .A(n42055), .X(n42056) );
  inv_x4_sg U42636 ( .A(n21079), .X(n42057) );
  inv_x4_sg U42637 ( .A(n19535), .X(n42059) );
  inv_x4_sg U42638 ( .A(n17990), .X(n42061) );
  inv_x4_sg U42639 ( .A(n42063), .X(n42064) );
  inv_x2_sg U42640 ( .A(n42065), .X(n42066) );
  nor_x2_sg U42641 ( .A(n43173), .B(n16335), .X(n16333) );
  inv_x4_sg U42642 ( .A(n14869), .X(n42067) );
  inv_x4_sg U42643 ( .A(n17108), .X(n42069) );
  nor_x2_sg U42644 ( .A(n17112), .B(n17111), .X(n17109) );
  nor_x4_sg U42645 ( .A(n17099), .B(n46385), .X(n17111) );
  inv_x4_sg U42646 ( .A(n15542), .X(n42073) );
  nor_x2_sg U42647 ( .A(n15546), .B(n15545), .X(n15543) );
  nor_x4_sg U42648 ( .A(n15533), .B(n46429), .X(n15545) );
  inv_x4_sg U42649 ( .A(n13209), .X(n42077) );
  nor_x2_sg U42650 ( .A(n13213), .B(n13212), .X(n13210) );
  nor_x4_sg U42651 ( .A(n13200), .B(n46497), .X(n13212) );
  inv_x4_sg U42652 ( .A(n12428), .X(n42079) );
  nor_x2_sg U42653 ( .A(n12432), .B(n12431), .X(n12429) );
  nor_x4_sg U42654 ( .A(n46518), .B(n12344), .X(n12431) );
  inv_x4_sg U42655 ( .A(n20970), .X(n42081) );
  inv_x4_sg U42656 ( .A(n19426), .X(n42083) );
  inv_x4_sg U42657 ( .A(n17881), .X(n42085) );
  inv_x4_sg U42658 ( .A(n16323), .X(n42087) );
  nor_x2_sg U42659 ( .A(n16327), .B(n16326), .X(n16324) );
  nor_x4_sg U42660 ( .A(n46406), .B(n16239), .X(n16326) );
  inv_x4_sg U42661 ( .A(n14760), .X(n42089) );
  inv_x4_sg U42662 ( .A(n11648), .X(n42091) );
  inv_x4_sg U42663 ( .A(n10868), .X(n42093) );
  inv_x4_sg U42664 ( .A(n21740), .X(n42095) );
  nor_x2_sg U42665 ( .A(n21744), .B(n21743), .X(n21741) );
  nor_x4_sg U42666 ( .A(n46250), .B(n21653), .X(n21743) );
  inv_x4_sg U42667 ( .A(n20195), .X(n42097) );
  nor_x2_sg U42668 ( .A(n20199), .B(n20198), .X(n20196) );
  nor_x4_sg U42669 ( .A(n46295), .B(n20108), .X(n20198) );
  inv_x4_sg U42670 ( .A(n16274), .X(n42119) );
  nor_x2_sg U42671 ( .A(n43177), .B(n16477), .X(n16475) );
  inv_x4_sg U42672 ( .A(n42137), .X(n42138) );
  nor_x2_sg U42673 ( .A(n54111), .B(n18387), .X(n18384) );
  inv_x2_sg U42674 ( .A(n18387), .X(n54172) );
  nor_x8_sg U42675 ( .A(n18442), .B(n46353), .X(n18387) );
  inv_x4_sg U42676 ( .A(n42139), .X(n42140) );
  nor_x2_sg U42677 ( .A(n54970), .B(n20707), .X(n20704) );
  inv_x2_sg U42678 ( .A(n20707), .X(n55024) );
  nor_x8_sg U42679 ( .A(n20762), .B(n46281), .X(n20707) );
  inv_x4_sg U42680 ( .A(n42141), .X(n42142) );
  nor_x2_sg U42681 ( .A(n54402), .B(n19163), .X(n19160) );
  inv_x2_sg U42682 ( .A(n19163), .X(n54456) );
  nor_x8_sg U42683 ( .A(n19218), .B(n46326), .X(n19163) );
  inv_x4_sg U42684 ( .A(n42143), .X(n42144) );
  nor_x2_sg U42685 ( .A(n53837), .B(n17618), .X(n17615) );
  inv_x2_sg U42686 ( .A(n17618), .X(n53891) );
  nor_x8_sg U42687 ( .A(n17673), .B(n46373), .X(n17618) );
  inv_x4_sg U42688 ( .A(n42145), .X(n42146) );
  nor_x2_sg U42689 ( .A(n52710), .B(n14497), .X(n14494) );
  inv_x2_sg U42690 ( .A(n14497), .X(n52771) );
  nor_x8_sg U42691 ( .A(n14552), .B(n46463), .X(n14497) );
  inv_x4_sg U42692 ( .A(n42147), .X(n42148) );
  inv_x2_sg U42693 ( .A(n42149), .X(n42150) );
  inv_x4_sg U42694 ( .A(n42151), .X(n42152) );
  nor_x2_sg U42695 ( .A(n10427), .B(n44369), .X(n10426) );
  inv_x4_sg U42696 ( .A(n42153), .X(n42154) );
  inv_x4_sg U42697 ( .A(n42155), .X(n42156) );
  inv_x4_sg U42698 ( .A(n42157), .X(n42158) );
  inv_x4_sg U42699 ( .A(n42159), .X(n42160) );
  inv_x4_sg U42700 ( .A(n42161), .X(n42162) );
  nor_x2_sg U42701 ( .A(n20531), .B(n44363), .X(n20530) );
  inv_x4_sg U42702 ( .A(n42163), .X(n42164) );
  nor_x2_sg U42703 ( .A(n18987), .B(n44365), .X(n18986) );
  inv_x4_sg U42704 ( .A(n42165), .X(n42166) );
  nor_x2_sg U42705 ( .A(n17442), .B(n44367), .X(n17441) );
  inv_x4_sg U42706 ( .A(n42167), .X(n42168) );
  inv_x2_sg U42707 ( .A(n42169), .X(n42170) );
  inv_x4_sg U42708 ( .A(n42171), .X(n42172) );
  inv_x2_sg U42709 ( .A(n42173), .X(n42174) );
  inv_x4_sg U42710 ( .A(n42175), .X(n42176) );
  inv_x2_sg U42711 ( .A(n42177), .X(n42178) );
  inv_x4_sg U42712 ( .A(n42179), .X(n42180) );
  inv_x2_sg U42713 ( .A(n42181), .X(n42182) );
  inv_x4_sg U42714 ( .A(n42183), .X(n42184) );
  inv_x2_sg U42715 ( .A(n42185), .X(n42186) );
  inv_x4_sg U42716 ( .A(n42187), .X(n42188) );
  inv_x4_sg U42717 ( .A(n42189), .X(n42190) );
  inv_x4_sg U42718 ( .A(n42191), .X(n42192) );
  inv_x4_sg U42719 ( .A(n42193), .X(n42194) );
  inv_x4_sg U42720 ( .A(n42195), .X(n42196) );
  inv_x4_sg U42721 ( .A(n42197), .X(n42198) );
  inv_x2_sg U42722 ( .A(n42199), .X(n42200) );
  inv_x4_sg U42723 ( .A(n42201), .X(n42202) );
  inv_x2_sg U42724 ( .A(n42203), .X(n42204) );
  inv_x4_sg U42725 ( .A(n42205), .X(n42206) );
  inv_x4_sg U42726 ( .A(n42207), .X(n42208) );
  inv_x2_sg U42727 ( .A(n42209), .X(n42210) );
  inv_x4_sg U42728 ( .A(n42211), .X(n42212) );
  inv_x4_sg U42729 ( .A(n42213), .X(n42214) );
  inv_x2_sg U42730 ( .A(n42215), .X(n42216) );
  inv_x4_sg U42731 ( .A(n42217), .X(n42218) );
  inv_x4_sg U42732 ( .A(n42219), .X(n42220) );
  inv_x2_sg U42733 ( .A(n42221), .X(n42222) );
  inv_x4_sg U42734 ( .A(n42223), .X(n42224) );
  inv_x4_sg U42735 ( .A(n42225), .X(n42226) );
  inv_x4_sg U42736 ( .A(n42227), .X(n42228) );
  inv_x4_sg U42737 ( .A(n42229), .X(n42230) );
  inv_x4_sg U42738 ( .A(n42231), .X(n42232) );
  inv_x2_sg U42739 ( .A(n42233), .X(n42234) );
  inv_x4_sg U42740 ( .A(n42235), .X(n42236) );
  inv_x2_sg U42741 ( .A(n42237), .X(n42238) );
  inv_x4_sg U42742 ( .A(n42239), .X(n42240) );
  inv_x4_sg U42743 ( .A(n42241), .X(n42242) );
  inv_x2_sg U42744 ( .A(n42243), .X(n42244) );
  inv_x4_sg U42745 ( .A(n42245), .X(n42246) );
  inv_x2_sg U42746 ( .A(n42247), .X(n42248) );
  inv_x4_sg U42747 ( .A(n42249), .X(n42250) );
  inv_x2_sg U42748 ( .A(n42251), .X(n42252) );
  inv_x4_sg U42749 ( .A(n42253), .X(n42254) );
  inv_x4_sg U42750 ( .A(n42255), .X(n42256) );
  inv_x4_sg U42751 ( .A(n42257), .X(n42258) );
  inv_x4_sg U42752 ( .A(n42259), .X(n42260) );
  inv_x2_sg U42753 ( .A(n42261), .X(n42262) );
  inv_x4_sg U42754 ( .A(n42263), .X(n42264) );
  inv_x2_sg U42755 ( .A(n42265), .X(n42266) );
  inv_x4_sg U42756 ( .A(n42267), .X(n42268) );
  inv_x2_sg U42757 ( .A(n42269), .X(n42270) );
  inv_x4_sg U42758 ( .A(n42271), .X(n42272) );
  inv_x2_sg U42759 ( .A(n42273), .X(n42274) );
  inv_x4_sg U42760 ( .A(n42275), .X(n42276) );
  inv_x2_sg U42761 ( .A(n42277), .X(n42278) );
  inv_x4_sg U42762 ( .A(n42279), .X(n42280) );
  inv_x4_sg U42763 ( .A(n42281), .X(n42282) );
  inv_x4_sg U42764 ( .A(n15890), .X(n53222) );
  nor_x2_sg U42765 ( .A(n16661), .B(n16662), .X(n16660) );
  nor_x4_sg U42766 ( .A(n16678), .B(n46385), .X(n16662) );
  nand_x4_sg U42767 ( .A(n46391), .B(n16635), .X(n16678) );
  nor_x2_sg U42768 ( .A(n15095), .B(n15096), .X(n15094) );
  nor_x4_sg U42769 ( .A(n15112), .B(n46429), .X(n15096) );
  nand_x4_sg U42770 ( .A(n46435), .B(n15069), .X(n15112) );
  nor_x2_sg U42771 ( .A(n12762), .B(n12763), .X(n12761) );
  nor_x4_sg U42772 ( .A(n12779), .B(n46497), .X(n12763) );
  nand_x4_sg U42773 ( .A(n46503), .B(n12736), .X(n12779) );
  inv_x4_sg U42774 ( .A(n11995), .X(n51834) );
  nor_x2_sg U42775 ( .A(n11201), .B(n11202), .X(n11200) );
  nor_x4_sg U42776 ( .A(n11218), .B(n46541), .X(n11202) );
  nand_x4_sg U42777 ( .A(n46547), .B(n11175), .X(n11218) );
  inv_x4_sg U42778 ( .A(n42283), .X(n42284) );
  inv_x4_sg U42779 ( .A(n42285), .X(n42286) );
  nor_x8_sg U42780 ( .A(n16109), .B(n46407), .X(n16029) );
  nor_x8_sg U42781 ( .A(n11434), .B(n46546), .X(n11354) );
  inv_x4_sg U42782 ( .A(n10330), .X(n42302) );
  inv_x4_sg U42783 ( .A(n18113), .X(n42304) );
  nor_x4_sg U42784 ( .A(n10619), .B(n10618), .X(n10636) );
  nor_x4_sg U42785 ( .A(n21491), .B(n21490), .X(n21508) );
  nor_x4_sg U42786 ( .A(n19946), .B(n19945), .X(n19963) );
  nor_x4_sg U42787 ( .A(n18401), .B(n18400), .X(n18418) );
  nor_x4_sg U42788 ( .A(n44699), .B(n15981), .X(n15775) );
  inv_x4_sg U42789 ( .A(n21202), .X(n42306) );
  nor_x4_sg U42790 ( .A(n20721), .B(n20720), .X(n20738) );
  inv_x4_sg U42791 ( .A(n19657), .X(n42308) );
  nor_x4_sg U42792 ( .A(n19177), .B(n19176), .X(n19194) );
  nor_x4_sg U42793 ( .A(n17632), .B(n17631), .X(n17649) );
  nor_x4_sg U42794 ( .A(n44697), .B(n16766), .X(n16557) );
  inv_x4_sg U42795 ( .A(n42310), .X(n42311) );
  nor_x4_sg U42796 ( .A(n44701), .B(n15200), .X(n14991) );
  nor_x4_sg U42797 ( .A(n14511), .B(n14510), .X(n14528) );
  nor_x4_sg U42798 ( .A(n44703), .B(n13647), .X(n13442) );
  nor_x4_sg U42799 ( .A(n44705), .B(n12867), .X(n12658) );
  nor_x4_sg U42800 ( .A(n44707), .B(n12086), .X(n11880) );
  nor_x4_sg U42801 ( .A(n44709), .B(n11306), .X(n11097) );
  inv_x4_sg U42802 ( .A(n42312), .X(n42313) );
  inv_x4_sg U42803 ( .A(n20429), .X(n42314) );
  inv_x4_sg U42804 ( .A(n18885), .X(n42316) );
  inv_x4_sg U42805 ( .A(n17340), .X(n42318) );
  inv_x4_sg U42806 ( .A(n14221), .X(n42320) );
  inv_x4_sg U42807 ( .A(n42322), .X(n42323) );
  inv_x4_sg U42808 ( .A(n42324), .X(n42325) );
  inv_x4_sg U42809 ( .A(n42326), .X(n42327) );
  inv_x4_sg U42810 ( .A(n42328), .X(n42329) );
  inv_x4_sg U42811 ( .A(n42330), .X(n42331) );
  inv_x4_sg U42812 ( .A(n42332), .X(n42333) );
  inv_x4_sg U42813 ( .A(n42334), .X(n42335) );
  inv_x4_sg U42814 ( .A(n14335), .X(n42336) );
  nor_x8_sg U42815 ( .A(n46451), .B(n46456), .X(n14335) );
  inv_x2_sg U42816 ( .A(n14335), .X(n52666) );
  inv_x4_sg U42817 ( .A(n20547), .X(n42337) );
  nor_x8_sg U42818 ( .A(n46270), .B(n46274), .X(n20547) );
  inv_x2_sg U42819 ( .A(n20547), .X(n54915) );
  inv_x4_sg U42820 ( .A(n19003), .X(n42338) );
  nor_x8_sg U42821 ( .A(n46315), .B(n46319), .X(n19003) );
  inv_x2_sg U42822 ( .A(n19003), .X(n54347) );
  inv_x4_sg U42823 ( .A(n17458), .X(n42339) );
  nor_x8_sg U42824 ( .A(n46362), .B(n46366), .X(n17458) );
  inv_x2_sg U42825 ( .A(n17458), .X(n53782) );
  nor_x2_sg U42826 ( .A(n53755), .B(n53710), .X(n27733) );
  nor_x2_sg U42827 ( .A(n53710), .B(n53707), .X(n27743) );
  inv_x4_sg U42828 ( .A(n17162), .X(n53710) );
  nor_x2_sg U42829 ( .A(n53477), .B(n53430), .X(n27452) );
  nor_x2_sg U42830 ( .A(n53430), .B(n53425), .X(n27462) );
  inv_x4_sg U42831 ( .A(n16378), .X(n53430) );
  nor_x2_sg U42832 ( .A(n53197), .B(n53152), .X(n27173) );
  nor_x2_sg U42833 ( .A(n53152), .B(n53149), .X(n27183) );
  inv_x4_sg U42834 ( .A(n15596), .X(n53152) );
  nor_x2_sg U42835 ( .A(n52638), .B(n52593), .X(n26616) );
  nor_x2_sg U42836 ( .A(n52593), .B(n52590), .X(n26626) );
  inv_x4_sg U42837 ( .A(n14043), .X(n52593) );
  nor_x2_sg U42838 ( .A(n52363), .B(n52318), .X(n26337) );
  nor_x2_sg U42839 ( .A(n52318), .B(n52315), .X(n26347) );
  inv_x4_sg U42840 ( .A(n13263), .X(n52318) );
  nor_x2_sg U42841 ( .A(n52085), .B(n52042), .X(n26056) );
  nor_x2_sg U42842 ( .A(n52042), .B(n52039), .X(n26066) );
  inv_x4_sg U42843 ( .A(n12482), .X(n52042) );
  nor_x2_sg U42844 ( .A(n51809), .B(n51761), .X(n25777) );
  nor_x2_sg U42845 ( .A(n51761), .B(n51756), .X(n25787) );
  inv_x4_sg U42846 ( .A(n11703), .X(n51761) );
  nor_x2_sg U42847 ( .A(n21117), .B(n55090), .X(n21116) );
  nor_x2_sg U42848 ( .A(n55090), .B(n55104), .X(n21108) );
  inv_x4_sg U42849 ( .A(n41816), .X(n55090) );
  nor_x2_sg U42850 ( .A(n19573), .B(n54522), .X(n19572) );
  nor_x2_sg U42851 ( .A(n54522), .B(n54536), .X(n19564) );
  inv_x4_sg U42852 ( .A(n41818), .X(n54522) );
  nor_x2_sg U42853 ( .A(n18028), .B(n53957), .X(n18027) );
  nor_x2_sg U42854 ( .A(n53957), .B(n53971), .X(n18019) );
  inv_x4_sg U42855 ( .A(n41820), .X(n53957) );
  nor_x2_sg U42856 ( .A(n14907), .B(n52837), .X(n14906) );
  nor_x2_sg U42857 ( .A(n52837), .B(n52851), .X(n14898) );
  inv_x4_sg U42858 ( .A(n41822), .X(n52837) );
  inv_x4_sg U42859 ( .A(n42340), .X(n42341) );
  inv_x4_sg U42860 ( .A(n42342), .X(n42343) );
  inv_x4_sg U42861 ( .A(n42344), .X(n42345) );
  inv_x4_sg U42862 ( .A(n42346), .X(n42347) );
  inv_x4_sg U42863 ( .A(n15946), .X(n42348) );
  inv_x4_sg U42864 ( .A(n10498), .X(n51342) );
  inv_x4_sg U42865 ( .A(n21370), .X(n55264) );
  inv_x4_sg U42866 ( .A(n19825), .X(n54696) );
  inv_x4_sg U42867 ( .A(n16732), .X(n42349) );
  inv_x4_sg U42868 ( .A(n15166), .X(n42350) );
  inv_x4_sg U42869 ( .A(n12833), .X(n42351) );
  inv_x4_sg U42870 ( .A(n12051), .X(n42352) );
  inv_x4_sg U42871 ( .A(n11272), .X(n42353) );
  inv_x4_sg U42872 ( .A(n20599), .X(n54985) );
  inv_x4_sg U42873 ( .A(n19055), .X(n54417) );
  inv_x4_sg U42874 ( .A(n17510), .X(n53852) );
  inv_x4_sg U42875 ( .A(n14389), .X(n52732) );
  inv_x4_sg U42876 ( .A(n42354), .X(n42355) );
  nor_x2_sg U42877 ( .A(n46248), .B(n21380), .X(n21414) );
  inv_x4_sg U42878 ( .A(n42356), .X(n42357) );
  nor_x2_sg U42879 ( .A(n46293), .B(n19835), .X(n19869) );
  inv_x4_sg U42880 ( .A(n42358), .X(n42359) );
  nor_x2_sg U42881 ( .A(n54921), .B(n20609), .X(n20643) );
  inv_x4_sg U42882 ( .A(n42360), .X(n42361) );
  nor_x2_sg U42883 ( .A(n54353), .B(n19065), .X(n19099) );
  inv_x4_sg U42884 ( .A(n42362), .X(n42363) );
  nor_x2_sg U42885 ( .A(n53788), .B(n17520), .X(n17554) );
  nor_x4_sg U42886 ( .A(n53537), .B(n16775), .X(n16773) );
  inv_x4_sg U42887 ( .A(n16744), .X(n53537) );
  nor_x4_sg U42888 ( .A(n52979), .B(n15209), .X(n15207) );
  inv_x4_sg U42889 ( .A(n15178), .X(n52979) );
  inv_x4_sg U42890 ( .A(n42364), .X(n42365) );
  nor_x2_sg U42891 ( .A(n46449), .B(n14399), .X(n14435) );
  nor_x4_sg U42892 ( .A(n52145), .B(n12876), .X(n12874) );
  inv_x4_sg U42893 ( .A(n12845), .X(n52145) );
  nor_x4_sg U42894 ( .A(n43195), .B(n53724), .X(n16576) );
  nor_x4_sg U42895 ( .A(n43197), .B(n53166), .X(n15010) );
  nor_x4_sg U42896 ( .A(n43199), .B(n52607), .X(n13461) );
  nor_x4_sg U42897 ( .A(n43201), .B(n52332), .X(n12677) );
  nor_x4_sg U42898 ( .A(n43203), .B(n51775), .X(n11116) );
  inv_x4_sg U42899 ( .A(n12419), .X(n42366) );
  inv_x4_sg U42900 ( .A(n42366), .X(n42367) );
  nor_x4_sg U42901 ( .A(n16764), .B(n43237), .X(n16766) );
  nor_x4_sg U42902 ( .A(n16763), .B(n16762), .X(n16764) );
  nor_x4_sg U42903 ( .A(n15198), .B(n43239), .X(n15200) );
  nor_x4_sg U42904 ( .A(n15197), .B(n15196), .X(n15198) );
  nor_x4_sg U42905 ( .A(n13645), .B(n13649), .X(n13647) );
  nor_x4_sg U42906 ( .A(n13644), .B(n13643), .X(n13645) );
  nor_x4_sg U42907 ( .A(n12865), .B(n43241), .X(n12867) );
  nor_x4_sg U42908 ( .A(n12864), .B(n12863), .X(n12865) );
  inv_x4_sg U42909 ( .A(n10531), .X(n42368) );
  inv_x4_sg U42910 ( .A(n42368), .X(n42369) );
  inv_x4_sg U42911 ( .A(n18313), .X(n42370) );
  inv_x4_sg U42912 ( .A(n42370), .X(n42371) );
  inv_x4_sg U42913 ( .A(n13556), .X(n52386) );
  nand_x8_sg U42914 ( .A(n54184), .B(n46352), .X(n18514) );
  nand_x8_sg U42915 ( .A(n21796), .B(n29417), .X(n29433) );
  nand_x8_sg U42916 ( .A(n21025), .B(n29135), .X(n29153) );
  nand_x8_sg U42917 ( .A(n20251), .B(n28856), .X(n28872) );
  nand_x8_sg U42918 ( .A(n19481), .B(n28576), .X(n28592) );
  nand_x8_sg U42919 ( .A(n18705), .B(n28298), .X(n28315) );
  nand_x8_sg U42920 ( .A(n17936), .B(n28018), .X(n28034) );
  nand_x8_sg U42921 ( .A(n14815), .B(n26899), .X(n26915) );
  inv_x4_sg U42922 ( .A(n21588), .X(n42372) );
  nor_x2_sg U42923 ( .A(n44177), .B(n21633), .X(n21630) );
  inv_x4_sg U42924 ( .A(n20043), .X(n42374) );
  nor_x2_sg U42925 ( .A(n44179), .B(n20088), .X(n20085) );
  inv_x4_sg U42926 ( .A(n18498), .X(n42376) );
  nor_x2_sg U42927 ( .A(n44181), .B(n18543), .X(n18540) );
  inv_x4_sg U42928 ( .A(n12277), .X(n42378) );
  nor_x2_sg U42929 ( .A(n44191), .B(n12324), .X(n12321) );
  inv_x4_sg U42930 ( .A(n42394), .X(n42395) );
  inv_x4_sg U42931 ( .A(n42396), .X(n42397) );
  nor_x4_sg U42932 ( .A(n42395), .B(n42397), .X(n16142) );
  inv_x4_sg U42933 ( .A(n16164), .X(n42398) );
  nor_x2_sg U42934 ( .A(n16241), .B(n16242), .X(n16240) );
  inv_x4_sg U42935 ( .A(n42400), .X(n42401) );
  inv_x4_sg U42936 ( .A(n42402), .X(n42403) );
  nor_x4_sg U42937 ( .A(n42401), .B(n42403), .X(n12247) );
  inv_x4_sg U42938 ( .A(n42404), .X(n42405) );
  nor_x4_sg U42939 ( .A(n10699), .B(n42405), .X(n10686) );
  nor_x4_sg U42940 ( .A(n10702), .B(n41277), .X(n10699) );
  inv_x4_sg U42941 ( .A(n42406), .X(n42407) );
  nor_x4_sg U42942 ( .A(n21571), .B(n42407), .X(n21558) );
  nor_x4_sg U42943 ( .A(n21574), .B(n41572), .X(n21571) );
  inv_x4_sg U42944 ( .A(n42408), .X(n42409) );
  nor_x4_sg U42945 ( .A(n20026), .B(n42409), .X(n20013) );
  nor_x4_sg U42946 ( .A(n20029), .B(n41574), .X(n20026) );
  inv_x4_sg U42947 ( .A(n42410), .X(n42411) );
  inv_x4_sg U42948 ( .A(n42412), .X(n42413) );
  nor_x4_sg U42949 ( .A(n42411), .B(n42413), .X(n20788) );
  inv_x4_sg U42950 ( .A(n42414), .X(n42415) );
  inv_x4_sg U42951 ( .A(n42416), .X(n42417) );
  nor_x4_sg U42952 ( .A(n42415), .B(n42417), .X(n19244) );
  inv_x4_sg U42953 ( .A(n42418), .X(n42419) );
  inv_x4_sg U42954 ( .A(n42420), .X(n42421) );
  nor_x4_sg U42955 ( .A(n42419), .B(n42421), .X(n17699) );
  inv_x4_sg U42956 ( .A(n42422), .X(n42423) );
  inv_x4_sg U42957 ( .A(n42424), .X(n42425) );
  nor_x4_sg U42958 ( .A(n42423), .B(n42425), .X(n14578) );
  inv_x4_sg U42959 ( .A(n21580), .X(n42426) );
  nor_x2_sg U42960 ( .A(n21655), .B(n21656), .X(n21654) );
  inv_x4_sg U42961 ( .A(n20035), .X(n42428) );
  nor_x2_sg U42962 ( .A(n20110), .B(n20111), .X(n20109) );
  inv_x4_sg U42963 ( .A(n20810), .X(n42430) );
  nor_x2_sg U42964 ( .A(n20886), .B(n43347), .X(n20885) );
  inv_x4_sg U42965 ( .A(n19266), .X(n42432) );
  nor_x2_sg U42966 ( .A(n19342), .B(n43349), .X(n19341) );
  inv_x4_sg U42967 ( .A(n17721), .X(n42434) );
  nor_x2_sg U42968 ( .A(n17797), .B(n43351), .X(n17796) );
  inv_x4_sg U42969 ( .A(n42436), .X(n42437) );
  nor_x4_sg U42970 ( .A(n20397), .B(n20396), .X(n20398) );
  inv_x4_sg U42971 ( .A(n42438), .X(n42439) );
  nor_x4_sg U42972 ( .A(n18853), .B(n18852), .X(n18854) );
  inv_x4_sg U42973 ( .A(n42440), .X(n42441) );
  nor_x4_sg U42974 ( .A(n17308), .B(n17307), .X(n17309) );
  nand_x8_sg U42975 ( .A(n49256), .B(n31429), .X(n25382) );
  nand_x2_sg U42976 ( .A(n8382), .B(n25352), .X(n31429) );
  nand_x8_sg U42977 ( .A(n49252), .B(n31868), .X(n25378) );
  nand_x2_sg U42978 ( .A(n8442), .B(n25348), .X(n31868) );
  nand_x8_sg U42979 ( .A(n50111), .B(n24202), .X(n10272) );
  nand_x2_sg U42980 ( .A(n8742), .B(n10245), .X(n24202) );
  nand_x8_sg U42981 ( .A(n50115), .B(n23763), .X(n10276) );
  nand_x2_sg U42982 ( .A(n8682), .B(n10244), .X(n23763) );
  nand_x8_sg U42983 ( .A(n27417), .B(n16190), .X(n27424) );
  nand_x8_sg U42984 ( .A(n26020), .B(n12295), .X(n26027) );
  nand_x8_sg U42985 ( .A(n25742), .B(n11515), .X(n25749) );
  inv_x4_sg U42986 ( .A(n10899), .X(n51498) );
  nor_x4_sg U42987 ( .A(n10919), .B(n46566), .X(n10899) );
  nor_x4_sg U42988 ( .A(n10518), .B(n46565), .X(n10580) );
  nor_x4_sg U42989 ( .A(n46250), .B(n46246), .X(n21452) );
  nor_x4_sg U42990 ( .A(n46295), .B(n46291), .X(n19907) );
  nor_x4_sg U42991 ( .A(n46335), .B(n46340), .X(n18362) );
  nor_x4_sg U42992 ( .A(n20685), .B(n46270), .X(n20681) );
  nor_x4_sg U42993 ( .A(n19141), .B(n46315), .X(n19137) );
  nor_x4_sg U42994 ( .A(n17596), .B(n46362), .X(n17592) );
  nor_x4_sg U42995 ( .A(n46447), .B(n46451), .X(n14472) );
  inv_x8_sg U42996 ( .A(n11522), .X(n51684) );
  inv_x4_sg U42997 ( .A(n42442), .X(n42443) );
  inv_x4_sg U42998 ( .A(n42444), .X(n42445) );
  inv_x4_sg U42999 ( .A(n42446), .X(n42447) );
  inv_x8_sg U43000 ( .A(n44574), .X(n44575) );
  inv_x4_sg U43001 ( .A(n29833), .X(n44574) );
  nor_x2_sg U43002 ( .A(n29835), .B(n49994), .X(n29833) );
  inv_x8_sg U43003 ( .A(n44654), .X(n44655) );
  inv_x4_sg U43004 ( .A(n22168), .X(n44654) );
  nor_x2_sg U43005 ( .A(n22170), .B(n50853), .X(n22168) );
  nor_x4_sg U43006 ( .A(n54200), .B(n18562), .X(n18490) );
  inv_x4_sg U43007 ( .A(n18557), .X(n54200) );
  nor_x4_sg U43008 ( .A(n18563), .B(n18564), .X(n18562) );
  nor_x4_sg U43009 ( .A(n15948), .B(n15947), .X(n15950) );
  nor_x4_sg U43010 ( .A(n44695), .B(n42348), .X(n15947) );
  nor_x4_sg U43011 ( .A(n10500), .B(n10499), .X(n10502) );
  nor_x4_sg U43012 ( .A(n10496), .B(n51342), .X(n10499) );
  nor_x4_sg U43013 ( .A(n21372), .B(n21371), .X(n21374) );
  nor_x4_sg U43014 ( .A(n21368), .B(n55264), .X(n21371) );
  nor_x4_sg U43015 ( .A(n19827), .B(n19826), .X(n19829) );
  nor_x4_sg U43016 ( .A(n19823), .B(n54696), .X(n19826) );
  nor_x4_sg U43017 ( .A(n54133), .B(n18281), .X(n18283) );
  inv_x4_sg U43018 ( .A(n18279), .X(n54133) );
  nor_x4_sg U43019 ( .A(n16734), .B(n16733), .X(n16736) );
  nor_x4_sg U43020 ( .A(n44279), .B(n42349), .X(n16733) );
  nor_x4_sg U43021 ( .A(n15168), .B(n15167), .X(n15170) );
  nor_x4_sg U43022 ( .A(n44281), .B(n42350), .X(n15167) );
  inv_x4_sg U43023 ( .A(n42448), .X(n42449) );
  nor_x4_sg U43024 ( .A(n12835), .B(n12834), .X(n12837) );
  nor_x4_sg U43025 ( .A(n44283), .B(n42351), .X(n12834) );
  nor_x4_sg U43026 ( .A(n12053), .B(n12052), .X(n12055) );
  nor_x4_sg U43027 ( .A(n45529), .B(n42352), .X(n12052) );
  nor_x4_sg U43028 ( .A(n11274), .B(n11273), .X(n11276) );
  nor_x4_sg U43029 ( .A(n44076), .B(n42353), .X(n11273) );
  nor_x4_sg U43030 ( .A(n20601), .B(n20600), .X(n20603) );
  nor_x4_sg U43031 ( .A(n20597), .B(n54985), .X(n20600) );
  nor_x4_sg U43032 ( .A(n19057), .B(n19056), .X(n19059) );
  nor_x4_sg U43033 ( .A(n19053), .B(n54417), .X(n19056) );
  nor_x4_sg U43034 ( .A(n17512), .B(n17511), .X(n17514) );
  nor_x4_sg U43035 ( .A(n17508), .B(n53852), .X(n17511) );
  nor_x4_sg U43036 ( .A(n14391), .B(n14390), .X(n14393) );
  nor_x4_sg U43037 ( .A(n14387), .B(n52732), .X(n14390) );
  inv_x4_sg U43038 ( .A(n16948), .X(n42450) );
  inv_x4_sg U43039 ( .A(n42450), .X(n42451) );
  inv_x4_sg U43040 ( .A(n15382), .X(n42452) );
  inv_x4_sg U43041 ( .A(n42452), .X(n42453) );
  inv_x4_sg U43042 ( .A(n13049), .X(n42454) );
  inv_x4_sg U43043 ( .A(n42454), .X(n42455) );
  inv_x4_sg U43044 ( .A(n11488), .X(n42456) );
  inv_x4_sg U43045 ( .A(n42456), .X(n42457) );
  inv_x4_sg U43046 ( .A(n42458), .X(n42459) );
  nor_x2_sg U43047 ( .A(n10663), .B(n10664), .X(n10661) );
  nor_x4_sg U43048 ( .A(n42459), .B(n51397), .X(n10663) );
  inv_x4_sg U43049 ( .A(n10734), .X(n51397) );
  nand_x2_sg U43050 ( .A(n10696), .B(n51396), .X(n10734) );
  inv_x4_sg U43051 ( .A(n42460), .X(n42461) );
  nor_x2_sg U43052 ( .A(n21535), .B(n21536), .X(n21533) );
  nor_x4_sg U43053 ( .A(n42461), .B(n55321), .X(n21535) );
  inv_x4_sg U43054 ( .A(n21606), .X(n55321) );
  nand_x2_sg U43055 ( .A(n21568), .B(n21604), .X(n21606) );
  inv_x4_sg U43056 ( .A(n42462), .X(n42463) );
  nor_x2_sg U43057 ( .A(n19990), .B(n19991), .X(n19988) );
  nor_x4_sg U43058 ( .A(n42463), .B(n54753), .X(n19990) );
  inv_x4_sg U43059 ( .A(n20061), .X(n54753) );
  nand_x2_sg U43060 ( .A(n20023), .B(n20059), .X(n20061) );
  inv_x4_sg U43061 ( .A(n42464), .X(n42465) );
  nor_x4_sg U43062 ( .A(n50095), .B(n42465), .X(n29625) );
  inv_x4_sg U43063 ( .A(n30193), .X(n50095) );
  nand_x2_sg U43064 ( .A(n30192), .B(n41348), .X(n30193) );
  nand_x4_sg U43065 ( .A(n15889), .B(n16199), .X(n16194) );
  nor_x4_sg U43066 ( .A(n16113), .B(n46402), .X(n16199) );
  inv_x4_sg U43067 ( .A(n42466), .X(n42467) );
  nor_x4_sg U43068 ( .A(n50954), .B(n42467), .X(n21964) );
  inv_x4_sg U43069 ( .A(n22527), .X(n50954) );
  nand_x2_sg U43070 ( .A(n22526), .B(n41350), .X(n22527) );
  nand_x4_sg U43071 ( .A(n13865), .B(n13555), .X(n13860) );
  nor_x4_sg U43072 ( .A(n13779), .B(n46469), .X(n13865) );
  nand_x4_sg U43073 ( .A(n11994), .B(n12304), .X(n12299) );
  nor_x4_sg U43074 ( .A(n12218), .B(n46514), .X(n12304) );
  nor_x2_sg U43075 ( .A(n54899), .B(n54894), .X(n20385) );
  nand_x4_sg U43076 ( .A(n20386), .B(n54894), .X(n20393) );
  inv_x4_sg U43077 ( .A(n20383), .X(n54894) );
  nor_x2_sg U43078 ( .A(n54331), .B(n54326), .X(n18841) );
  nand_x4_sg U43079 ( .A(n18842), .B(n54326), .X(n18849) );
  inv_x4_sg U43080 ( .A(n18839), .X(n54326) );
  nor_x2_sg U43081 ( .A(n53766), .B(n53761), .X(n17296) );
  nand_x4_sg U43082 ( .A(n17297), .B(n53761), .X(n17304) );
  inv_x4_sg U43083 ( .A(n17294), .X(n53761) );
  inv_x4_sg U43084 ( .A(n42468), .X(n42469) );
  nor_x4_sg U43085 ( .A(n42469), .B(n54210), .X(n18487) );
  inv_x4_sg U43086 ( .A(n18560), .X(n54210) );
  nand_x2_sg U43087 ( .A(n18558), .B(n18561), .X(n18560) );
  nor_x2_sg U43088 ( .A(n40755), .B(n31321), .X(n31320) );
  nor_x4_sg U43089 ( .A(n31396), .B(n49775), .X(n31321) );
  inv_x4_sg U43090 ( .A(n31397), .X(n49775) );
  nand_x2_sg U43091 ( .A(n8351), .B(n31398), .X(n31397) );
  nor_x4_sg U43092 ( .A(n24851), .B(n31315), .X(n31396) );
  nor_x2_sg U43093 ( .A(n40756), .B(n23655), .X(n23654) );
  nor_x4_sg U43094 ( .A(n23730), .B(n50634), .X(n23655) );
  inv_x4_sg U43095 ( .A(n23731), .X(n50634) );
  nand_x2_sg U43096 ( .A(n8651), .B(n23732), .X(n23731) );
  nor_x4_sg U43097 ( .A(n9743), .B(n23649), .X(n23730) );
  inv_x4_sg U43098 ( .A(n42470), .X(n42471) );
  inv_x4_sg U43099 ( .A(n42472), .X(n42473) );
  nor_x2_sg U43100 ( .A(n18214), .B(n18215), .X(n18213) );
  nor_x4_sg U43101 ( .A(n42471), .B(n42473), .X(n18214) );
  nor_x2_sg U43102 ( .A(n16514), .B(n53483), .X(n16513) );
  inv_x4_sg U43103 ( .A(n16511), .X(n53483) );
  nor_x2_sg U43104 ( .A(n14948), .B(n52925), .X(n14947) );
  inv_x4_sg U43105 ( .A(n14945), .X(n52925) );
  nor_x2_sg U43106 ( .A(n12615), .B(n52091), .X(n12614) );
  inv_x4_sg U43107 ( .A(n12612), .X(n52091) );
  nor_x2_sg U43108 ( .A(n11054), .B(n51533), .X(n11053) );
  inv_x4_sg U43109 ( .A(n11051), .X(n51533) );
  inv_x4_sg U43110 ( .A(n27725), .X(n42474) );
  inv_x8_sg U43111 ( .A(n42474), .X(n42475) );
  inv_x4_sg U43112 ( .A(n27445), .X(n42476) );
  inv_x8_sg U43113 ( .A(n42476), .X(n42477) );
  inv_x4_sg U43114 ( .A(n27165), .X(n42478) );
  inv_x8_sg U43115 ( .A(n42478), .X(n42479) );
  inv_x4_sg U43116 ( .A(n26608), .X(n42480) );
  inv_x8_sg U43117 ( .A(n42480), .X(n42481) );
  inv_x4_sg U43118 ( .A(n26329), .X(n42482) );
  inv_x8_sg U43119 ( .A(n42482), .X(n42483) );
  inv_x4_sg U43120 ( .A(n26048), .X(n42484) );
  inv_x8_sg U43121 ( .A(n42484), .X(n42485) );
  inv_x4_sg U43122 ( .A(n25770), .X(n42486) );
  inv_x8_sg U43123 ( .A(n42486), .X(n42487) );
  inv_x4_sg U43124 ( .A(n25492), .X(n42488) );
  inv_x8_sg U43125 ( .A(n42488), .X(n42489) );
  inv_x4_sg U43126 ( .A(n42490), .X(n42491) );
  nor_x2_sg U43127 ( .A(n29644), .B(n9415), .X(n29634) );
  nor_x4_sg U43128 ( .A(n42491), .B(n50104), .X(n29644) );
  inv_x4_sg U43129 ( .A(n30165), .X(n50104) );
  nand_x2_sg U43130 ( .A(n41143), .B(n42687), .X(n30165) );
  inv_x4_sg U43131 ( .A(n42492), .X(n42493) );
  nor_x2_sg U43132 ( .A(n29608), .B(n9385), .X(n29604) );
  nor_x4_sg U43133 ( .A(n42493), .B(n50100), .X(n29608) );
  inv_x4_sg U43134 ( .A(n30177), .X(n50100) );
  nand_x2_sg U43135 ( .A(n41179), .B(n42689), .X(n30177) );
  inv_x4_sg U43136 ( .A(n42494), .X(n42495) );
  nor_x2_sg U43137 ( .A(n21979), .B(n9415), .X(n21969) );
  nor_x4_sg U43138 ( .A(n42495), .B(n50963), .X(n21979) );
  inv_x4_sg U43139 ( .A(n22499), .X(n50963) );
  nand_x2_sg U43140 ( .A(n41145), .B(n42759), .X(n22499) );
  inv_x4_sg U43141 ( .A(n42496), .X(n42497) );
  nor_x2_sg U43142 ( .A(n21952), .B(n9385), .X(n21949) );
  nor_x4_sg U43143 ( .A(n42497), .B(n50959), .X(n21952) );
  inv_x4_sg U43144 ( .A(n22511), .X(n50959) );
  nand_x2_sg U43145 ( .A(n41181), .B(n42761), .X(n22511) );
  inv_x4_sg U43146 ( .A(n42498), .X(n42499) );
  inv_x4_sg U43147 ( .A(n42500), .X(n42501) );
  nor_x4_sg U43148 ( .A(n42499), .B(n42501), .X(n24511) );
  inv_x4_sg U43149 ( .A(n42502), .X(n42503) );
  inv_x4_sg U43150 ( .A(n42504), .X(n42505) );
  nor_x4_sg U43151 ( .A(n42503), .B(n42505), .X(n9400) );
  inv_x4_sg U43152 ( .A(n17283), .X(n42506) );
  inv_x8_sg U43153 ( .A(n42506), .X(n42507) );
  inv_x4_sg U43154 ( .A(n15717), .X(n42508) );
  inv_x8_sg U43155 ( .A(n42508), .X(n42509) );
  inv_x4_sg U43156 ( .A(n14164), .X(n42510) );
  inv_x8_sg U43157 ( .A(n42510), .X(n42511) );
  inv_x4_sg U43158 ( .A(n13384), .X(n42512) );
  inv_x8_sg U43159 ( .A(n42512), .X(n42513) );
  inv_x4_sg U43160 ( .A(n12602), .X(n42514) );
  inv_x8_sg U43161 ( .A(n42514), .X(n42515) );
  inv_x4_sg U43162 ( .A(n28449), .X(n42516) );
  inv_x8_sg U43163 ( .A(n42516), .X(n42517) );
  nor_x8_sg U43164 ( .A(n28448), .B(n42517), .X(n28383) );
  nor_x8_sg U43165 ( .A(n28389), .B(n46193), .X(n28448) );
  inv_x4_sg U43166 ( .A(n9981), .X(n50366) );
  inv_x4_sg U43167 ( .A(n25089), .X(n49507) );
  nor_x2_sg U43168 ( .A(n40757), .B(n31291), .X(n31290) );
  inv_x2_sg U43169 ( .A(n31291), .X(n49540) );
  nor_x8_sg U43170 ( .A(n31411), .B(n49539), .X(n31291) );
  inv_x8_sg U43171 ( .A(n31412), .X(n49539) );
  nor_x8_sg U43172 ( .A(n25092), .B(n31285), .X(n31411) );
  nand_x4_sg U43173 ( .A(n8356), .B(n31413), .X(n31412) );
  nor_x2_sg U43174 ( .A(n40758), .B(n31309), .X(n31308) );
  inv_x2_sg U43175 ( .A(n31309), .X(n49680) );
  nor_x8_sg U43176 ( .A(n31402), .B(n49679), .X(n31309) );
  inv_x8_sg U43177 ( .A(n31403), .X(n49679) );
  nor_x8_sg U43178 ( .A(n24947), .B(n31303), .X(n31402) );
  nand_x4_sg U43179 ( .A(n8353), .B(n31404), .X(n31403) );
  nor_x2_sg U43180 ( .A(n40759), .B(n23625), .X(n23624) );
  inv_x2_sg U43181 ( .A(n23625), .X(n50399) );
  nor_x8_sg U43182 ( .A(n23745), .B(n50398), .X(n23625) );
  inv_x8_sg U43183 ( .A(n23746), .X(n50398) );
  nor_x8_sg U43184 ( .A(n9984), .B(n23619), .X(n23745) );
  nand_x4_sg U43185 ( .A(n8656), .B(n23747), .X(n23746) );
  nor_x2_sg U43186 ( .A(n40760), .B(n23643), .X(n23642) );
  inv_x2_sg U43187 ( .A(n23643), .X(n50539) );
  nor_x8_sg U43188 ( .A(n23736), .B(n50538), .X(n23643) );
  inv_x8_sg U43189 ( .A(n23737), .X(n50538) );
  nor_x8_sg U43190 ( .A(n9839), .B(n23637), .X(n23736) );
  nand_x4_sg U43191 ( .A(n8653), .B(n23738), .X(n23737) );
  inv_x2_sg U43192 ( .A(n24423), .X(n50227) );
  inv_x2_sg U43193 ( .A(n32089), .X(n49368) );
  nand_x2_sg U43194 ( .A(n25273), .B(n30847), .X(n31044) );
  nor_x2_sg U43195 ( .A(n25273), .B(n9385), .X(n25270) );
  nor_x8_sg U43196 ( .A(n31057), .B(n49330), .X(n25273) );
  inv_x8_sg U43197 ( .A(n31058), .X(n49330) );
  nor_x8_sg U43198 ( .A(n42631), .B(n25263), .X(n31057) );
  nand_x4_sg U43199 ( .A(n25263), .B(n42631), .X(n31058) );
  nand_x2_sg U43200 ( .A(n25224), .B(n30853), .X(n31041) );
  nor_x2_sg U43201 ( .A(n25224), .B(n9385), .X(n25221) );
  nor_x8_sg U43202 ( .A(n31063), .B(n49374), .X(n25224) );
  inv_x8_sg U43203 ( .A(n31064), .X(n49374) );
  nor_x8_sg U43204 ( .A(n42633), .B(n25214), .X(n31063) );
  nand_x4_sg U43205 ( .A(n25214), .B(n42633), .X(n31064) );
  nand_x2_sg U43206 ( .A(n25175), .B(n30859), .X(n31038) );
  nor_x2_sg U43207 ( .A(n25175), .B(n9385), .X(n25172) );
  nor_x8_sg U43208 ( .A(n31069), .B(n49420), .X(n25175) );
  inv_x8_sg U43209 ( .A(n31070), .X(n49420) );
  nor_x8_sg U43210 ( .A(n42635), .B(n25165), .X(n31069) );
  nand_x4_sg U43211 ( .A(n25165), .B(n42635), .X(n31070) );
  nand_x2_sg U43212 ( .A(n25150), .B(n29939), .X(n30051) );
  nor_x2_sg U43213 ( .A(n25150), .B(n9415), .X(n25141) );
  nor_x8_sg U43214 ( .A(n30091), .B(n49470), .X(n25150) );
  inv_x8_sg U43215 ( .A(n30092), .X(n49470) );
  nor_x8_sg U43216 ( .A(n42637), .B(n25132), .X(n30091) );
  nand_x4_sg U43217 ( .A(n25132), .B(n42637), .X(n30092) );
  nand_x2_sg U43218 ( .A(n25127), .B(n30865), .X(n31035) );
  nor_x2_sg U43219 ( .A(n25127), .B(n9385), .X(n25124) );
  nor_x8_sg U43220 ( .A(n31075), .B(n49466), .X(n25127) );
  inv_x8_sg U43221 ( .A(n31076), .X(n49466) );
  nor_x8_sg U43222 ( .A(n42639), .B(n25117), .X(n31075) );
  nand_x4_sg U43223 ( .A(n25117), .B(n42639), .X(n31076) );
  nand_x2_sg U43224 ( .A(n25078), .B(n30871), .X(n31032) );
  nor_x2_sg U43225 ( .A(n25078), .B(n9385), .X(n25075) );
  nor_x8_sg U43226 ( .A(n31081), .B(n49513), .X(n25078) );
  inv_x8_sg U43227 ( .A(n31082), .X(n49513) );
  nor_x8_sg U43228 ( .A(n42641), .B(n25068), .X(n31081) );
  nand_x4_sg U43229 ( .A(n25068), .B(n42641), .X(n31082) );
  nand_x2_sg U43230 ( .A(n25053), .B(n29951), .X(n30045) );
  nor_x2_sg U43231 ( .A(n25053), .B(n9415), .X(n25044) );
  nor_x8_sg U43232 ( .A(n30103), .B(n49564), .X(n25053) );
  inv_x8_sg U43233 ( .A(n30104), .X(n49564) );
  nor_x8_sg U43234 ( .A(n42643), .B(n25035), .X(n30103) );
  nand_x4_sg U43235 ( .A(n25035), .B(n42643), .X(n30104) );
  nand_x2_sg U43236 ( .A(n25030), .B(n30877), .X(n31029) );
  nor_x2_sg U43237 ( .A(n25030), .B(n9385), .X(n25027) );
  nor_x8_sg U43238 ( .A(n31087), .B(n49560), .X(n25030) );
  inv_x8_sg U43239 ( .A(n31088), .X(n49560) );
  nor_x8_sg U43240 ( .A(n42645), .B(n25020), .X(n31087) );
  nand_x4_sg U43241 ( .A(n25020), .B(n42645), .X(n31088) );
  nand_x2_sg U43242 ( .A(n25005), .B(n29957), .X(n30042) );
  nor_x2_sg U43243 ( .A(n25005), .B(n9415), .X(n24996) );
  nor_x8_sg U43244 ( .A(n30109), .B(n49610), .X(n25005) );
  inv_x8_sg U43245 ( .A(n30110), .X(n49610) );
  nor_x8_sg U43246 ( .A(n42647), .B(n24987), .X(n30109) );
  nand_x4_sg U43247 ( .A(n24987), .B(n42647), .X(n30110) );
  nand_x2_sg U43248 ( .A(n24982), .B(n30883), .X(n31026) );
  nor_x2_sg U43249 ( .A(n24982), .B(n9385), .X(n24979) );
  nor_x8_sg U43250 ( .A(n31093), .B(n49606), .X(n24982) );
  inv_x8_sg U43251 ( .A(n31094), .X(n49606) );
  nor_x8_sg U43252 ( .A(n42649), .B(n24972), .X(n31093) );
  nand_x4_sg U43253 ( .A(n24972), .B(n42649), .X(n31094) );
  nand_x2_sg U43254 ( .A(n24957), .B(n29963), .X(n30039) );
  nor_x2_sg U43255 ( .A(n24957), .B(n9415), .X(n24948) );
  nor_x8_sg U43256 ( .A(n30115), .B(n49657), .X(n24957) );
  inv_x8_sg U43257 ( .A(n30116), .X(n49657) );
  nor_x8_sg U43258 ( .A(n42651), .B(n24939), .X(n30115) );
  nand_x4_sg U43259 ( .A(n24939), .B(n42651), .X(n30116) );
  nand_x2_sg U43260 ( .A(n24934), .B(n30889), .X(n31023) );
  nor_x2_sg U43261 ( .A(n24934), .B(n9385), .X(n24931) );
  nor_x8_sg U43262 ( .A(n31099), .B(n49653), .X(n24934) );
  inv_x8_sg U43263 ( .A(n31100), .X(n49653) );
  nor_x8_sg U43264 ( .A(n42653), .B(n24924), .X(n31099) );
  nand_x4_sg U43265 ( .A(n24924), .B(n42653), .X(n31100) );
  nand_x2_sg U43266 ( .A(n24909), .B(n29969), .X(n30036) );
  nor_x2_sg U43267 ( .A(n24909), .B(n9415), .X(n24900) );
  nor_x8_sg U43268 ( .A(n30121), .B(n49704), .X(n24909) );
  inv_x8_sg U43269 ( .A(n30122), .X(n49704) );
  nor_x8_sg U43270 ( .A(n42655), .B(n24891), .X(n30121) );
  nand_x4_sg U43271 ( .A(n24891), .B(n42655), .X(n30122) );
  nand_x2_sg U43272 ( .A(n24886), .B(n30895), .X(n31020) );
  nor_x2_sg U43273 ( .A(n24886), .B(n9385), .X(n24883) );
  nor_x8_sg U43274 ( .A(n31105), .B(n49700), .X(n24886) );
  inv_x8_sg U43275 ( .A(n31106), .X(n49700) );
  nor_x8_sg U43276 ( .A(n42657), .B(n24876), .X(n31105) );
  nand_x4_sg U43277 ( .A(n24876), .B(n42657), .X(n31106) );
  nand_x2_sg U43278 ( .A(n24861), .B(n29975), .X(n30033) );
  nor_x2_sg U43279 ( .A(n24861), .B(n9415), .X(n24852) );
  nor_x8_sg U43280 ( .A(n30127), .B(n49753), .X(n24861) );
  inv_x8_sg U43281 ( .A(n30128), .X(n49753) );
  nor_x8_sg U43282 ( .A(n42659), .B(n24843), .X(n30127) );
  nand_x4_sg U43283 ( .A(n24843), .B(n42659), .X(n30128) );
  nand_x2_sg U43284 ( .A(n24838), .B(n30901), .X(n31017) );
  nor_x2_sg U43285 ( .A(n24838), .B(n9385), .X(n24835) );
  nor_x8_sg U43286 ( .A(n31111), .B(n49749), .X(n24838) );
  inv_x8_sg U43287 ( .A(n31112), .X(n49749) );
  nor_x8_sg U43288 ( .A(n42661), .B(n24828), .X(n31111) );
  nand_x4_sg U43289 ( .A(n24828), .B(n42661), .X(n31112) );
  nand_x2_sg U43290 ( .A(n24766), .B(n29987), .X(n30027) );
  nor_x2_sg U43291 ( .A(n24766), .B(n9415), .X(n24757) );
  nor_x8_sg U43292 ( .A(n30139), .B(n49848), .X(n24766) );
  inv_x8_sg U43293 ( .A(n30140), .X(n49848) );
  nor_x8_sg U43294 ( .A(n42663), .B(n24748), .X(n30139) );
  nand_x4_sg U43295 ( .A(n24748), .B(n42663), .X(n30140) );
  nand_x2_sg U43296 ( .A(n24743), .B(n30913), .X(n31011) );
  nor_x2_sg U43297 ( .A(n24743), .B(n9385), .X(n24740) );
  nor_x8_sg U43298 ( .A(n31123), .B(n49844), .X(n24743) );
  inv_x8_sg U43299 ( .A(n31124), .X(n49844) );
  nor_x8_sg U43300 ( .A(n42665), .B(n24733), .X(n31123) );
  nand_x4_sg U43301 ( .A(n24733), .B(n42665), .X(n31124) );
  nand_x2_sg U43302 ( .A(n24718), .B(n29993), .X(n30024) );
  nor_x2_sg U43303 ( .A(n24718), .B(n9415), .X(n24709) );
  nor_x8_sg U43304 ( .A(n30145), .B(n49895), .X(n24718) );
  inv_x8_sg U43305 ( .A(n30146), .X(n49895) );
  nor_x8_sg U43306 ( .A(n42667), .B(n24700), .X(n30145) );
  nand_x4_sg U43307 ( .A(n24700), .B(n42667), .X(n30146) );
  nand_x2_sg U43308 ( .A(n24695), .B(n30919), .X(n31008) );
  nor_x2_sg U43309 ( .A(n24695), .B(n9385), .X(n24692) );
  nor_x8_sg U43310 ( .A(n31129), .B(n49891), .X(n24695) );
  inv_x8_sg U43311 ( .A(n31130), .X(n49891) );
  nor_x8_sg U43312 ( .A(n42669), .B(n24685), .X(n31129) );
  nand_x4_sg U43313 ( .A(n24685), .B(n42669), .X(n31130) );
  nand_x2_sg U43314 ( .A(n24670), .B(n29999), .X(n30021) );
  nor_x2_sg U43315 ( .A(n24670), .B(n9415), .X(n24661) );
  nor_x8_sg U43316 ( .A(n30151), .B(n49943), .X(n24670) );
  inv_x8_sg U43317 ( .A(n30152), .X(n49943) );
  nor_x8_sg U43318 ( .A(n42671), .B(n24652), .X(n30151) );
  nand_x4_sg U43319 ( .A(n24652), .B(n42671), .X(n30152) );
  nand_x2_sg U43320 ( .A(n24646), .B(n30925), .X(n31005) );
  nor_x2_sg U43321 ( .A(n24646), .B(n9385), .X(n24643) );
  nor_x8_sg U43322 ( .A(n31135), .B(n49940), .X(n24646) );
  inv_x8_sg U43323 ( .A(n31136), .X(n49940) );
  nor_x8_sg U43324 ( .A(n42673), .B(n24636), .X(n31135) );
  nand_x4_sg U43325 ( .A(n24636), .B(n42673), .X(n31136) );
  nand_x2_sg U43326 ( .A(n24621), .B(n30005), .X(n30018) );
  nor_x2_sg U43327 ( .A(n24621), .B(n9415), .X(n24612) );
  nor_x8_sg U43328 ( .A(n30157), .B(n49988), .X(n24621) );
  inv_x8_sg U43329 ( .A(n30158), .X(n49988) );
  nor_x8_sg U43330 ( .A(n42675), .B(n24603), .X(n30157) );
  nand_x4_sg U43331 ( .A(n24603), .B(n42675), .X(n30158) );
  nand_x2_sg U43332 ( .A(n24597), .B(n30784), .X(n30781) );
  nor_x2_sg U43333 ( .A(n24597), .B(n9385), .X(n24594) );
  nor_x8_sg U43334 ( .A(n30930), .B(n49983), .X(n24597) );
  inv_x8_sg U43335 ( .A(n30931), .X(n49983) );
  nor_x8_sg U43336 ( .A(n42677), .B(n24587), .X(n30930) );
  nand_x4_sg U43337 ( .A(n24587), .B(n42677), .X(n30931) );
  nand_x2_sg U43338 ( .A(n24572), .B(n29855), .X(n29852) );
  nand_x2_sg U43339 ( .A(n30009), .B(n24572), .X(n30007) );
  nor_x2_sg U43340 ( .A(n24572), .B(n9415), .X(n24563) );
  nor_x8_sg U43341 ( .A(n30010), .B(n50035), .X(n24572) );
  inv_x8_sg U43342 ( .A(n30011), .X(n50035) );
  nor_x8_sg U43343 ( .A(n42679), .B(n24554), .X(n30010) );
  nand_x4_sg U43344 ( .A(n24554), .B(n42679), .X(n30011) );
  nand_x2_sg U43345 ( .A(n24548), .B(n30527), .X(n30524) );
  nor_x2_sg U43346 ( .A(n24548), .B(n9385), .X(n24545) );
  nor_x8_sg U43347 ( .A(n30704), .B(n50028), .X(n24548) );
  inv_x8_sg U43348 ( .A(n30705), .X(n50028) );
  nor_x8_sg U43349 ( .A(n42681), .B(n24538), .X(n30704) );
  nand_x4_sg U43350 ( .A(n24538), .B(n42681), .X(n30705) );
  nor_x2_sg U43351 ( .A(n24523), .B(n9415), .X(n24514) );
  nor_x8_sg U43352 ( .A(n29844), .B(n50080), .X(n24523) );
  inv_x8_sg U43353 ( .A(n29845), .X(n50080) );
  nor_x8_sg U43354 ( .A(n42683), .B(n24505), .X(n29844) );
  nand_x4_sg U43355 ( .A(n24505), .B(n42683), .X(n29845) );
  nor_x2_sg U43356 ( .A(n24499), .B(n9385), .X(n24496) );
  nor_x8_sg U43357 ( .A(n30449), .B(n50070), .X(n24499) );
  inv_x8_sg U43358 ( .A(n30450), .X(n50070) );
  nor_x8_sg U43359 ( .A(n42685), .B(n24488), .X(n30449) );
  nand_x4_sg U43360 ( .A(n24488), .B(n42685), .X(n30450) );
  nand_x2_sg U43361 ( .A(n10151), .B(n23936), .X(n24062) );
  nand_x2_sg U43362 ( .A(n23934), .B(n10151), .X(n23932) );
  nor_x2_sg U43363 ( .A(n10151), .B(n9367), .X(n10148) );
  nand_x2_sg U43364 ( .A(n10165), .B(n23181), .X(n23378) );
  nor_x2_sg U43365 ( .A(n10165), .B(n9385), .X(n10162) );
  nor_x8_sg U43366 ( .A(n23391), .B(n50189), .X(n10165) );
  inv_x8_sg U43367 ( .A(n23392), .X(n50189) );
  nor_x8_sg U43368 ( .A(n42703), .B(n10150), .X(n23391) );
  nand_x4_sg U43369 ( .A(n10150), .B(n42703), .X(n23392) );
  nand_x2_sg U43370 ( .A(n10116), .B(n23187), .X(n23375) );
  nor_x2_sg U43371 ( .A(n10116), .B(n9385), .X(n10113) );
  nor_x8_sg U43372 ( .A(n23397), .B(n50233), .X(n10116) );
  inv_x8_sg U43373 ( .A(n23398), .X(n50233) );
  nor_x8_sg U43374 ( .A(n42705), .B(n10101), .X(n23397) );
  nand_x4_sg U43375 ( .A(n10101), .B(n42705), .X(n23398) );
  nand_x2_sg U43376 ( .A(n10067), .B(n23193), .X(n23372) );
  nor_x2_sg U43377 ( .A(n10067), .B(n9385), .X(n10064) );
  nor_x8_sg U43378 ( .A(n23403), .B(n50279), .X(n10067) );
  inv_x8_sg U43379 ( .A(n23404), .X(n50279) );
  nor_x8_sg U43380 ( .A(n42707), .B(n10052), .X(n23403) );
  nand_x4_sg U43381 ( .A(n10052), .B(n42707), .X(n23404) );
  nand_x2_sg U43382 ( .A(n10005), .B(n23954), .X(n24053) );
  nand_x2_sg U43383 ( .A(n23952), .B(n10005), .X(n23950) );
  nor_x2_sg U43384 ( .A(n10005), .B(n9367), .X(n10002) );
  nand_x2_sg U43385 ( .A(n10042), .B(n22274), .X(n22386) );
  nor_x2_sg U43386 ( .A(n10042), .B(n9415), .X(n10033) );
  nor_x8_sg U43387 ( .A(n22426), .B(n50329), .X(n10042) );
  inv_x8_sg U43388 ( .A(n22427), .X(n50329) );
  nor_x8_sg U43389 ( .A(n42709), .B(n10024), .X(n22426) );
  nand_x4_sg U43390 ( .A(n10024), .B(n42709), .X(n22427) );
  nand_x2_sg U43391 ( .A(n10019), .B(n23199), .X(n23369) );
  nor_x2_sg U43392 ( .A(n10019), .B(n9385), .X(n10016) );
  nor_x8_sg U43393 ( .A(n23409), .B(n50325), .X(n10019) );
  inv_x8_sg U43394 ( .A(n23410), .X(n50325) );
  nor_x8_sg U43395 ( .A(n42711), .B(n10004), .X(n23409) );
  nand_x4_sg U43396 ( .A(n10004), .B(n42711), .X(n23410) );
  nand_x2_sg U43397 ( .A(n9956), .B(n23960), .X(n24050) );
  nand_x2_sg U43398 ( .A(n23958), .B(n9956), .X(n23956) );
  nor_x2_sg U43399 ( .A(n9956), .B(n9367), .X(n9953) );
  nand_x2_sg U43400 ( .A(n9970), .B(n23205), .X(n23366) );
  nor_x2_sg U43401 ( .A(n9970), .B(n9385), .X(n9967) );
  nor_x8_sg U43402 ( .A(n23415), .B(n50372), .X(n9970) );
  inv_x8_sg U43403 ( .A(n23416), .X(n50372) );
  nor_x8_sg U43404 ( .A(n42713), .B(n9955), .X(n23415) );
  nand_x4_sg U43405 ( .A(n9955), .B(n42713), .X(n23416) );
  nand_x2_sg U43406 ( .A(n9908), .B(n23966), .X(n24047) );
  nand_x2_sg U43407 ( .A(n23964), .B(n9908), .X(n23962) );
  nor_x2_sg U43408 ( .A(n9908), .B(n9367), .X(n9905) );
  nand_x2_sg U43409 ( .A(n9945), .B(n22286), .X(n22380) );
  nor_x2_sg U43410 ( .A(n9945), .B(n9415), .X(n9936) );
  nor_x8_sg U43411 ( .A(n22438), .B(n50423), .X(n9945) );
  inv_x8_sg U43412 ( .A(n22439), .X(n50423) );
  nor_x8_sg U43413 ( .A(n42715), .B(n9927), .X(n22438) );
  nand_x4_sg U43414 ( .A(n9927), .B(n42715), .X(n22439) );
  nand_x2_sg U43415 ( .A(n9922), .B(n23211), .X(n23363) );
  nor_x2_sg U43416 ( .A(n9922), .B(n9385), .X(n9919) );
  nor_x8_sg U43417 ( .A(n23421), .B(n50419), .X(n9922) );
  inv_x8_sg U43418 ( .A(n23422), .X(n50419) );
  nor_x8_sg U43419 ( .A(n42717), .B(n9907), .X(n23421) );
  nand_x4_sg U43420 ( .A(n9907), .B(n42717), .X(n23422) );
  nand_x2_sg U43421 ( .A(n9860), .B(n23972), .X(n24044) );
  nand_x2_sg U43422 ( .A(n23970), .B(n9860), .X(n23968) );
  nor_x2_sg U43423 ( .A(n9860), .B(n9367), .X(n9857) );
  nand_x2_sg U43424 ( .A(n9897), .B(n22292), .X(n22377) );
  nor_x2_sg U43425 ( .A(n9897), .B(n9415), .X(n9888) );
  nor_x8_sg U43426 ( .A(n22444), .B(n50469), .X(n9897) );
  inv_x8_sg U43427 ( .A(n22445), .X(n50469) );
  nor_x8_sg U43428 ( .A(n42719), .B(n9879), .X(n22444) );
  nand_x4_sg U43429 ( .A(n9879), .B(n42719), .X(n22445) );
  nand_x2_sg U43430 ( .A(n9874), .B(n23217), .X(n23360) );
  nor_x2_sg U43431 ( .A(n9874), .B(n9385), .X(n9871) );
  nor_x8_sg U43432 ( .A(n23427), .B(n50465), .X(n9874) );
  inv_x8_sg U43433 ( .A(n23428), .X(n50465) );
  nor_x8_sg U43434 ( .A(n42721), .B(n9859), .X(n23427) );
  nand_x4_sg U43435 ( .A(n9859), .B(n42721), .X(n23428) );
  nand_x2_sg U43436 ( .A(n9812), .B(n23978), .X(n24041) );
  nand_x2_sg U43437 ( .A(n23976), .B(n9812), .X(n23974) );
  nor_x2_sg U43438 ( .A(n9812), .B(n9367), .X(n9809) );
  nand_x2_sg U43439 ( .A(n9849), .B(n22298), .X(n22374) );
  nor_x2_sg U43440 ( .A(n9849), .B(n9415), .X(n9840) );
  nor_x8_sg U43441 ( .A(n22450), .B(n50516), .X(n9849) );
  inv_x8_sg U43442 ( .A(n22451), .X(n50516) );
  nor_x8_sg U43443 ( .A(n42723), .B(n9831), .X(n22450) );
  nand_x4_sg U43444 ( .A(n9831), .B(n42723), .X(n22451) );
  nand_x2_sg U43445 ( .A(n9826), .B(n23223), .X(n23357) );
  nor_x2_sg U43446 ( .A(n9826), .B(n9385), .X(n9823) );
  nor_x8_sg U43447 ( .A(n23433), .B(n50512), .X(n9826) );
  inv_x8_sg U43448 ( .A(n23434), .X(n50512) );
  nor_x8_sg U43449 ( .A(n42725), .B(n9811), .X(n23433) );
  nand_x4_sg U43450 ( .A(n9811), .B(n42725), .X(n23434) );
  inv_x4_sg U43451 ( .A(n24133), .X(n42536) );
  inv_x8_sg U43452 ( .A(n42536), .X(n42537) );
  nand_x2_sg U43453 ( .A(n9764), .B(n23984), .X(n24038) );
  nand_x2_sg U43454 ( .A(n23982), .B(n9764), .X(n23980) );
  nor_x2_sg U43455 ( .A(n9764), .B(n9367), .X(n9761) );
  nor_x8_sg U43456 ( .A(n24132), .B(n42537), .X(n9764) );
  nor_x8_sg U43457 ( .A(n44657), .B(n24135), .X(n24132) );
  nand_x2_sg U43458 ( .A(n9801), .B(n22304), .X(n22371) );
  nor_x2_sg U43459 ( .A(n9801), .B(n9415), .X(n9792) );
  nor_x8_sg U43460 ( .A(n22456), .B(n50563), .X(n9801) );
  inv_x8_sg U43461 ( .A(n22457), .X(n50563) );
  nor_x8_sg U43462 ( .A(n42727), .B(n9783), .X(n22456) );
  nand_x4_sg U43463 ( .A(n9783), .B(n42727), .X(n22457) );
  nand_x2_sg U43464 ( .A(n9778), .B(n23229), .X(n23354) );
  nor_x2_sg U43465 ( .A(n9778), .B(n9385), .X(n9775) );
  nor_x8_sg U43466 ( .A(n23439), .B(n50559), .X(n9778) );
  inv_x8_sg U43467 ( .A(n23440), .X(n50559) );
  nor_x8_sg U43468 ( .A(n42729), .B(n9763), .X(n23439) );
  nand_x4_sg U43469 ( .A(n9763), .B(n42729), .X(n23440) );
  inv_x4_sg U43470 ( .A(n24140), .X(n42538) );
  inv_x8_sg U43471 ( .A(n42538), .X(n42539) );
  nand_x2_sg U43472 ( .A(n9716), .B(n23990), .X(n24035) );
  nand_x2_sg U43473 ( .A(n23988), .B(n9716), .X(n23986) );
  nor_x2_sg U43474 ( .A(n9716), .B(n9367), .X(n9713) );
  nor_x8_sg U43475 ( .A(n24139), .B(n42539), .X(n9716) );
  nor_x8_sg U43476 ( .A(n45509), .B(n24032), .X(n24139) );
  nand_x2_sg U43477 ( .A(n9753), .B(n22310), .X(n22368) );
  nor_x2_sg U43478 ( .A(n9753), .B(n9415), .X(n9744) );
  nor_x8_sg U43479 ( .A(n22462), .B(n50612), .X(n9753) );
  inv_x8_sg U43480 ( .A(n22463), .X(n50612) );
  nor_x8_sg U43481 ( .A(n42731), .B(n9735), .X(n22462) );
  nand_x4_sg U43482 ( .A(n9735), .B(n42731), .X(n22463) );
  nand_x2_sg U43483 ( .A(n9730), .B(n23235), .X(n23351) );
  nor_x2_sg U43484 ( .A(n9730), .B(n9385), .X(n9727) );
  nor_x8_sg U43485 ( .A(n23445), .B(n50608), .X(n9730) );
  inv_x8_sg U43486 ( .A(n23446), .X(n50608) );
  nor_x8_sg U43487 ( .A(n42733), .B(n9715), .X(n23445) );
  nand_x4_sg U43488 ( .A(n9715), .B(n42733), .X(n23446) );
  inv_x4_sg U43489 ( .A(n23996), .X(n42540) );
  inv_x8_sg U43490 ( .A(n42540), .X(n42541) );
  nand_x2_sg U43491 ( .A(n9669), .B(n23885), .X(n23882) );
  nand_x2_sg U43492 ( .A(n23994), .B(n9669), .X(n23992) );
  nor_x2_sg U43493 ( .A(n9669), .B(n9367), .X(n9666) );
  nor_x8_sg U43494 ( .A(n23995), .B(n42541), .X(n9669) );
  nor_x8_sg U43495 ( .A(n45501), .B(n23879), .X(n23995) );
  inv_x4_sg U43496 ( .A(n23843), .X(n42542) );
  inv_x8_sg U43497 ( .A(n42542), .X(n42543) );
  nand_x2_sg U43498 ( .A(n9621), .B(n23714), .X(n23711) );
  nand_x2_sg U43499 ( .A(n23841), .B(n9621), .X(n23839) );
  nor_x2_sg U43500 ( .A(n9621), .B(n9367), .X(n9618) );
  nor_x8_sg U43501 ( .A(n23842), .B(n42543), .X(n9621) );
  nor_x8_sg U43502 ( .A(n45507), .B(n23708), .X(n23842) );
  nand_x2_sg U43503 ( .A(n9658), .B(n22322), .X(n22362) );
  nor_x2_sg U43504 ( .A(n9658), .B(n9415), .X(n9649) );
  nor_x8_sg U43505 ( .A(n22474), .B(n50707), .X(n9658) );
  inv_x8_sg U43506 ( .A(n22475), .X(n50707) );
  nor_x8_sg U43507 ( .A(n42735), .B(n9640), .X(n22474) );
  nand_x4_sg U43508 ( .A(n9640), .B(n42735), .X(n22475) );
  nand_x2_sg U43509 ( .A(n9635), .B(n23247), .X(n23345) );
  nor_x2_sg U43510 ( .A(n9635), .B(n9385), .X(n9632) );
  nor_x8_sg U43511 ( .A(n23457), .B(n50703), .X(n9635) );
  inv_x8_sg U43512 ( .A(n23458), .X(n50703) );
  nor_x8_sg U43513 ( .A(n42737), .B(n9620), .X(n23457) );
  nand_x4_sg U43514 ( .A(n9620), .B(n42737), .X(n23458) );
  inv_x4_sg U43515 ( .A(n23672), .X(n42544) );
  inv_x8_sg U43516 ( .A(n42544), .X(n42545) );
  nand_x2_sg U43517 ( .A(n9573), .B(n23524), .X(n23521) );
  nand_x2_sg U43518 ( .A(n23670), .B(n9573), .X(n23668) );
  nor_x2_sg U43519 ( .A(n9573), .B(n9367), .X(n9570) );
  nor_x8_sg U43520 ( .A(n23671), .B(n42545), .X(n9573) );
  nor_x8_sg U43521 ( .A(n45499), .B(n23518), .X(n23671) );
  nand_x2_sg U43522 ( .A(n9610), .B(n22328), .X(n22359) );
  nor_x2_sg U43523 ( .A(n9610), .B(n9415), .X(n9601) );
  nor_x8_sg U43524 ( .A(n22480), .B(n50754), .X(n9610) );
  inv_x8_sg U43525 ( .A(n22481), .X(n50754) );
  nor_x8_sg U43526 ( .A(n42739), .B(n9592), .X(n22480) );
  nand_x4_sg U43527 ( .A(n9592), .B(n42739), .X(n22481) );
  nand_x2_sg U43528 ( .A(n9587), .B(n23253), .X(n23342) );
  nor_x2_sg U43529 ( .A(n9587), .B(n9385), .X(n9584) );
  nor_x8_sg U43530 ( .A(n23463), .B(n50750), .X(n9587) );
  inv_x8_sg U43531 ( .A(n23464), .X(n50750) );
  nor_x8_sg U43532 ( .A(n42741), .B(n9572), .X(n23463) );
  nand_x4_sg U43533 ( .A(n9572), .B(n42741), .X(n23464) );
  inv_x4_sg U43534 ( .A(n23482), .X(n42546) );
  inv_x8_sg U43535 ( .A(n42546), .X(n42547) );
  nand_x2_sg U43536 ( .A(n9524), .B(n23319), .X(n23316) );
  nand_x2_sg U43537 ( .A(n23480), .B(n9524), .X(n23478) );
  nor_x2_sg U43538 ( .A(n9524), .B(n9367), .X(n9521) );
  nor_x8_sg U43539 ( .A(n23481), .B(n42547), .X(n9524) );
  nor_x8_sg U43540 ( .A(n45505), .B(n23313), .X(n23481) );
  nand_x2_sg U43541 ( .A(n9562), .B(n22334), .X(n22356) );
  nor_x2_sg U43542 ( .A(n9562), .B(n9415), .X(n9553) );
  nor_x8_sg U43543 ( .A(n22486), .B(n50802), .X(n9562) );
  inv_x8_sg U43544 ( .A(n22487), .X(n50802) );
  nor_x8_sg U43545 ( .A(n42743), .B(n9544), .X(n22486) );
  nand_x4_sg U43546 ( .A(n9544), .B(n42743), .X(n22487) );
  nand_x2_sg U43547 ( .A(n9538), .B(n23259), .X(n23339) );
  nor_x2_sg U43548 ( .A(n9538), .B(n9385), .X(n9535) );
  nor_x8_sg U43549 ( .A(n23469), .B(n50799), .X(n9538) );
  inv_x8_sg U43550 ( .A(n23470), .X(n50799) );
  nor_x8_sg U43551 ( .A(n42745), .B(n9523), .X(n23469) );
  nand_x4_sg U43552 ( .A(n9523), .B(n42745), .X(n23470) );
  inv_x4_sg U43553 ( .A(n23277), .X(n42548) );
  inv_x8_sg U43554 ( .A(n42548), .X(n42549) );
  nand_x2_sg U43555 ( .A(n9475), .B(n23093), .X(n23090) );
  nand_x2_sg U43556 ( .A(n23275), .B(n9475), .X(n23273) );
  nor_x2_sg U43557 ( .A(n9475), .B(n9367), .X(n9472) );
  nor_x8_sg U43558 ( .A(n23276), .B(n42549), .X(n9475) );
  nor_x8_sg U43559 ( .A(n45497), .B(n23087), .X(n23276) );
  nand_x2_sg U43560 ( .A(n9513), .B(n22340), .X(n22353) );
  nor_x2_sg U43561 ( .A(n9513), .B(n9415), .X(n9504) );
  nor_x8_sg U43562 ( .A(n22492), .B(n50847), .X(n9513) );
  inv_x8_sg U43563 ( .A(n22493), .X(n50847) );
  nor_x8_sg U43564 ( .A(n42747), .B(n9495), .X(n22492) );
  nand_x4_sg U43565 ( .A(n9495), .B(n42747), .X(n22493) );
  nand_x2_sg U43566 ( .A(n9489), .B(n23118), .X(n23115) );
  nor_x2_sg U43567 ( .A(n9489), .B(n9385), .X(n9486) );
  nor_x8_sg U43568 ( .A(n23264), .B(n50842), .X(n9489) );
  inv_x8_sg U43569 ( .A(n23265), .X(n50842) );
  nor_x8_sg U43570 ( .A(n42749), .B(n9474), .X(n23264) );
  nand_x4_sg U43571 ( .A(n9474), .B(n42749), .X(n23265) );
  inv_x4_sg U43572 ( .A(n23051), .X(n42550) );
  inv_x8_sg U43573 ( .A(n42550), .X(n42551) );
  nand_x2_sg U43574 ( .A(n9426), .B(n22838), .X(n22835) );
  nand_x2_sg U43575 ( .A(n23049), .B(n9426), .X(n23047) );
  nor_x2_sg U43576 ( .A(n9426), .B(n9367), .X(n9423) );
  nor_x8_sg U43577 ( .A(n23050), .B(n42551), .X(n9426) );
  nor_x8_sg U43578 ( .A(n45503), .B(n22832), .X(n23050) );
  nand_x2_sg U43579 ( .A(n9464), .B(n22190), .X(n22187) );
  nand_x2_sg U43580 ( .A(n22344), .B(n9464), .X(n22342) );
  nor_x2_sg U43581 ( .A(n9464), .B(n9415), .X(n9455) );
  nor_x8_sg U43582 ( .A(n22345), .B(n50894), .X(n9464) );
  inv_x8_sg U43583 ( .A(n22346), .X(n50894) );
  nor_x8_sg U43584 ( .A(n42751), .B(n9446), .X(n22345) );
  nand_x4_sg U43585 ( .A(n9446), .B(n42751), .X(n22346) );
  nand_x2_sg U43586 ( .A(n9440), .B(n22861), .X(n22858) );
  nor_x2_sg U43587 ( .A(n9440), .B(n9385), .X(n9437) );
  nor_x8_sg U43588 ( .A(n23038), .B(n50887), .X(n9440) );
  inv_x8_sg U43589 ( .A(n23039), .X(n50887) );
  nor_x8_sg U43590 ( .A(n42753), .B(n9425), .X(n23038) );
  nand_x4_sg U43591 ( .A(n9425), .B(n42753), .X(n23039) );
  nor_x2_sg U43592 ( .A(n9414), .B(n9415), .X(n9404) );
  nor_x8_sg U43593 ( .A(n22179), .B(n50939), .X(n9414) );
  inv_x8_sg U43594 ( .A(n22180), .X(n50939) );
  nor_x8_sg U43595 ( .A(n42755), .B(n9391), .X(n22179) );
  nand_x4_sg U43596 ( .A(n9391), .B(n42755), .X(n22180) );
  nor_x2_sg U43597 ( .A(n9384), .B(n9385), .X(n9381) );
  nor_x8_sg U43598 ( .A(n22783), .B(n50929), .X(n9384) );
  inv_x8_sg U43599 ( .A(n22784), .X(n50929) );
  nor_x8_sg U43600 ( .A(n42757), .B(n9364), .X(n22783) );
  nand_x4_sg U43601 ( .A(n9364), .B(n42757), .X(n22784) );
  nand_x2_sg U43602 ( .A(n24790), .B(n24811), .X(n29682) );
  nor_x2_sg U43603 ( .A(n24790), .B(n46605), .X(n24789) );
  nand_x2_sg U43604 ( .A(n24797), .B(n30408), .X(n30551) );
  nand_x2_sg U43605 ( .A(n30406), .B(n24797), .X(n30404) );
  nor_x2_sg U43606 ( .A(n24797), .B(n9394), .X(n24794) );
  nand_x2_sg U43607 ( .A(n9682), .B(n9703), .X(n22017) );
  nor_x2_sg U43608 ( .A(n9682), .B(n46603), .X(n9681) );
  nand_x2_sg U43609 ( .A(n9689), .B(n22742), .X(n22885) );
  nand_x2_sg U43610 ( .A(n22740), .B(n9689), .X(n22738) );
  nor_x2_sg U43611 ( .A(n9689), .B(n9394), .X(n9686) );
  nand_x2_sg U43612 ( .A(n25259), .B(n31602), .X(n31728) );
  nand_x2_sg U43613 ( .A(n31600), .B(n25259), .X(n31598) );
  nor_x2_sg U43614 ( .A(n25259), .B(n9367), .X(n25256) );
  nand_x2_sg U43615 ( .A(n25210), .B(n31608), .X(n31725) );
  nand_x2_sg U43616 ( .A(n31606), .B(n25210), .X(n31604) );
  nor_x2_sg U43617 ( .A(n25210), .B(n9367), .X(n25207) );
  nand_x2_sg U43618 ( .A(n25161), .B(n31614), .X(n31722) );
  nand_x2_sg U43619 ( .A(n31612), .B(n25161), .X(n31610) );
  nor_x2_sg U43620 ( .A(n25161), .B(n9367), .X(n25158) );
  nand_x2_sg U43621 ( .A(n25113), .B(n31620), .X(n31719) );
  nand_x2_sg U43622 ( .A(n31618), .B(n25113), .X(n31616) );
  nor_x2_sg U43623 ( .A(n25113), .B(n9367), .X(n25110) );
  nand_x2_sg U43624 ( .A(n25064), .B(n31626), .X(n31716) );
  nand_x2_sg U43625 ( .A(n31624), .B(n25064), .X(n31622) );
  nor_x2_sg U43626 ( .A(n25064), .B(n9367), .X(n25061) );
  nand_x2_sg U43627 ( .A(n25016), .B(n31632), .X(n31713) );
  nand_x2_sg U43628 ( .A(n31630), .B(n25016), .X(n31628) );
  nor_x2_sg U43629 ( .A(n25016), .B(n9367), .X(n25013) );
  nand_x2_sg U43630 ( .A(n24968), .B(n31638), .X(n31710) );
  nand_x2_sg U43631 ( .A(n31636), .B(n24968), .X(n31634) );
  nor_x2_sg U43632 ( .A(n24968), .B(n9367), .X(n24965) );
  nand_x2_sg U43633 ( .A(n24920), .B(n31644), .X(n31707) );
  nand_x2_sg U43634 ( .A(n31642), .B(n24920), .X(n31640) );
  nor_x2_sg U43635 ( .A(n24920), .B(n9367), .X(n24917) );
  inv_x4_sg U43636 ( .A(n31799), .X(n42576) );
  inv_x8_sg U43637 ( .A(n42576), .X(n42577) );
  nand_x2_sg U43638 ( .A(n24872), .B(n31650), .X(n31704) );
  nand_x2_sg U43639 ( .A(n31648), .B(n24872), .X(n31646) );
  nor_x2_sg U43640 ( .A(n24872), .B(n9367), .X(n24869) );
  nor_x8_sg U43641 ( .A(n31798), .B(n42577), .X(n24872) );
  nor_x8_sg U43642 ( .A(n44666), .B(n31801), .X(n31798) );
  inv_x4_sg U43643 ( .A(n31806), .X(n42578) );
  inv_x8_sg U43644 ( .A(n42578), .X(n42579) );
  nand_x2_sg U43645 ( .A(n24824), .B(n31656), .X(n31701) );
  nand_x2_sg U43646 ( .A(n31654), .B(n24824), .X(n31652) );
  nor_x2_sg U43647 ( .A(n24824), .B(n9367), .X(n24821) );
  nor_x8_sg U43648 ( .A(n31805), .B(n42579), .X(n24824) );
  nor_x8_sg U43649 ( .A(n45523), .B(n31698), .X(n31805) );
  inv_x4_sg U43650 ( .A(n31509), .X(n42580) );
  inv_x8_sg U43651 ( .A(n42580), .X(n42581) );
  nand_x2_sg U43652 ( .A(n24729), .B(n31380), .X(n31377) );
  nand_x2_sg U43653 ( .A(n31507), .B(n24729), .X(n31505) );
  nor_x2_sg U43654 ( .A(n24729), .B(n9367), .X(n24726) );
  nor_x8_sg U43655 ( .A(n31508), .B(n42581), .X(n24729) );
  nor_x8_sg U43656 ( .A(n45521), .B(n31374), .X(n31508) );
  inv_x4_sg U43657 ( .A(n31148), .X(n42582) );
  inv_x8_sg U43658 ( .A(n42582), .X(n42583) );
  nand_x2_sg U43659 ( .A(n24632), .B(n30985), .X(n30982) );
  nand_x2_sg U43660 ( .A(n31146), .B(n24632), .X(n31144) );
  nor_x2_sg U43661 ( .A(n24632), .B(n9367), .X(n24629) );
  nor_x8_sg U43662 ( .A(n31147), .B(n42583), .X(n24632) );
  nor_x8_sg U43663 ( .A(n45519), .B(n30979), .X(n31147) );
  inv_x4_sg U43664 ( .A(n30717), .X(n42584) );
  inv_x8_sg U43665 ( .A(n42584), .X(n42585) );
  nand_x2_sg U43666 ( .A(n24534), .B(n30504), .X(n30501) );
  nand_x2_sg U43667 ( .A(n30715), .B(n24534), .X(n30713) );
  nor_x2_sg U43668 ( .A(n24534), .B(n9367), .X(n24531) );
  nor_x8_sg U43669 ( .A(n30716), .B(n42585), .X(n24534) );
  nor_x8_sg U43670 ( .A(n45517), .B(n30498), .X(n30716) );
  nand_x2_sg U43671 ( .A(n10102), .B(n23942), .X(n24059) );
  nand_x2_sg U43672 ( .A(n23940), .B(n10102), .X(n23938) );
  nor_x2_sg U43673 ( .A(n10102), .B(n9367), .X(n10099) );
  nand_x2_sg U43674 ( .A(n10053), .B(n23948), .X(n24056) );
  nand_x2_sg U43675 ( .A(n23946), .B(n10053), .X(n23944) );
  nor_x2_sg U43676 ( .A(n10053), .B(n9367), .X(n10050) );
  inv_x4_sg U43677 ( .A(n31338), .X(n42590) );
  inv_x8_sg U43678 ( .A(n42590), .X(n42591) );
  nand_x2_sg U43679 ( .A(n24681), .B(n31190), .X(n31187) );
  nand_x2_sg U43680 ( .A(n31336), .B(n24681), .X(n31334) );
  nor_x2_sg U43681 ( .A(n24681), .B(n9367), .X(n24678) );
  nor_x8_sg U43682 ( .A(n31337), .B(n42591), .X(n24681) );
  nor_x8_sg U43683 ( .A(n45513), .B(n31184), .X(n31337) );
  inv_x4_sg U43684 ( .A(n30943), .X(n42592) );
  inv_x8_sg U43685 ( .A(n42592), .X(n42593) );
  nand_x2_sg U43686 ( .A(n24583), .B(n30759), .X(n30756) );
  nand_x2_sg U43687 ( .A(n30941), .B(n24583), .X(n30939) );
  nor_x2_sg U43688 ( .A(n24583), .B(n9367), .X(n24580) );
  nor_x8_sg U43689 ( .A(n30942), .B(n42593), .X(n24583) );
  nor_x8_sg U43690 ( .A(n45511), .B(n30753), .X(n30942) );
  nand_x2_sg U43691 ( .A(n25295), .B(n29921), .X(n30060) );
  nor_x2_sg U43692 ( .A(n25295), .B(n9415), .X(n25286) );
  nor_x8_sg U43693 ( .A(n30073), .B(n49334), .X(n25295) );
  inv_x8_sg U43694 ( .A(n30074), .X(n49334) );
  nor_x8_sg U43695 ( .A(n42773), .B(n25278), .X(n30073) );
  nand_x4_sg U43696 ( .A(n25278), .B(n42773), .X(n30074) );
  nand_x2_sg U43697 ( .A(n25248), .B(n29927), .X(n30057) );
  nor_x2_sg U43698 ( .A(n25248), .B(n9415), .X(n25239) );
  nor_x8_sg U43699 ( .A(n30079), .B(n49378), .X(n25248) );
  inv_x8_sg U43700 ( .A(n30080), .X(n49378) );
  nor_x8_sg U43701 ( .A(n42775), .B(n25229), .X(n30079) );
  nand_x4_sg U43702 ( .A(n25229), .B(n42775), .X(n30080) );
  nand_x2_sg U43703 ( .A(n25199), .B(n29933), .X(n30054) );
  nor_x2_sg U43704 ( .A(n25199), .B(n9415), .X(n25190) );
  nor_x8_sg U43705 ( .A(n30085), .B(n49424), .X(n25199) );
  inv_x8_sg U43706 ( .A(n30086), .X(n49424) );
  nor_x8_sg U43707 ( .A(n42777), .B(n25180), .X(n30085) );
  nand_x4_sg U43708 ( .A(n25180), .B(n42777), .X(n30086) );
  nand_x2_sg U43709 ( .A(n25102), .B(n29945), .X(n30048) );
  nor_x2_sg U43710 ( .A(n25102), .B(n9415), .X(n25093) );
  nor_x8_sg U43711 ( .A(n30097), .B(n49517), .X(n25102) );
  inv_x8_sg U43712 ( .A(n30098), .X(n49517) );
  nor_x8_sg U43713 ( .A(n42779), .B(n25083), .X(n30097) );
  nand_x4_sg U43714 ( .A(n25083), .B(n42779), .X(n30098) );
  nand_x2_sg U43715 ( .A(n10187), .B(n22256), .X(n22395) );
  nor_x2_sg U43716 ( .A(n10187), .B(n9415), .X(n10178) );
  nor_x8_sg U43717 ( .A(n22408), .B(n50193), .X(n10187) );
  inv_x8_sg U43718 ( .A(n22409), .X(n50193) );
  nor_x8_sg U43719 ( .A(n42783), .B(n10170), .X(n22408) );
  nand_x4_sg U43720 ( .A(n10170), .B(n42783), .X(n22409) );
  nand_x2_sg U43721 ( .A(n10140), .B(n22262), .X(n22392) );
  nor_x2_sg U43722 ( .A(n10140), .B(n9415), .X(n10131) );
  nor_x8_sg U43723 ( .A(n22414), .B(n50237), .X(n10140) );
  inv_x8_sg U43724 ( .A(n22415), .X(n50237) );
  nor_x8_sg U43725 ( .A(n42785), .B(n10121), .X(n22414) );
  nand_x4_sg U43726 ( .A(n10121), .B(n42785), .X(n22415) );
  nand_x2_sg U43727 ( .A(n10091), .B(n22268), .X(n22389) );
  nor_x2_sg U43728 ( .A(n10091), .B(n9415), .X(n10082) );
  nor_x8_sg U43729 ( .A(n22420), .B(n50283), .X(n10091) );
  inv_x8_sg U43730 ( .A(n22421), .X(n50283) );
  nor_x8_sg U43731 ( .A(n42787), .B(n10072), .X(n22420) );
  nand_x4_sg U43732 ( .A(n10072), .B(n42787), .X(n22421) );
  nand_x2_sg U43733 ( .A(n9994), .B(n22280), .X(n22383) );
  nor_x2_sg U43734 ( .A(n9994), .B(n9415), .X(n9985) );
  nor_x8_sg U43735 ( .A(n22432), .B(n50376), .X(n9994) );
  inv_x8_sg U43736 ( .A(n22433), .X(n50376) );
  nor_x8_sg U43737 ( .A(n42789), .B(n9975), .X(n22432) );
  nand_x4_sg U43738 ( .A(n9975), .B(n42789), .X(n22433) );
  inv_x4_sg U43739 ( .A(n31662), .X(n42594) );
  inv_x8_sg U43740 ( .A(n42594), .X(n42595) );
  nand_x2_sg U43741 ( .A(n24777), .B(n31551), .X(n31548) );
  nand_x2_sg U43742 ( .A(n31660), .B(n24777), .X(n31658) );
  nor_x2_sg U43743 ( .A(n24777), .B(n9367), .X(n24774) );
  nor_x8_sg U43744 ( .A(n31661), .B(n42595), .X(n24777) );
  nor_x8_sg U43745 ( .A(n45515), .B(n31545), .X(n31661) );
  inv_x4_sg U43746 ( .A(n30462), .X(n42596) );
  inv_x8_sg U43747 ( .A(n42596), .X(n42597) );
  nand_x2_sg U43748 ( .A(n30460), .B(n24484), .X(n30458) );
  nor_x2_sg U43749 ( .A(n24484), .B(n9367), .X(n24481) );
  nor_x8_sg U43750 ( .A(n30461), .B(n42597), .X(n24484) );
  nor_x8_sg U43751 ( .A(n45527), .B(n30227), .X(n30461) );
  inv_x4_sg U43752 ( .A(n22796), .X(n42598) );
  inv_x8_sg U43753 ( .A(n42598), .X(n42599) );
  nand_x2_sg U43754 ( .A(n22794), .B(n9366), .X(n22792) );
  nor_x2_sg U43755 ( .A(n9366), .B(n9367), .X(n9362) );
  nor_x8_sg U43756 ( .A(n22795), .B(n42599), .X(n9366) );
  nor_x8_sg U43757 ( .A(n45525), .B(n22561), .X(n22795) );
  inv_x4_sg U43758 ( .A(n18759), .X(n42600) );
  nand_x4_sg U43759 ( .A(n53551), .B(n45469), .X(n16686) );
  nand_x4_sg U43760 ( .A(n52993), .B(n45473), .X(n15120) );
  nand_x4_sg U43761 ( .A(n52159), .B(n45479), .X(n12787) );
  nand_x4_sg U43762 ( .A(n51601), .B(n45483), .X(n11226) );
  nand_x4_sg U43763 ( .A(n54963), .B(n45461), .X(n20555) );
  nand_x4_sg U43764 ( .A(n54395), .B(n45465), .X(n19011) );
  nand_x4_sg U43765 ( .A(n53830), .B(n45467), .X(n17466) );
  inv_x4_sg U43766 ( .A(n54126), .X(n42602) );
  inv_x8_sg U43767 ( .A(n42602), .X(n42603) );
  inv_x4_sg U43768 ( .A(n42604), .X(n42605) );
  inv_x4_sg U43769 ( .A(n42606), .X(n42607) );
  inv_x4_sg U43770 ( .A(n42608), .X(n42609) );
  inv_x4_sg U43771 ( .A(n42610), .X(n42611) );
  inv_x4_sg U43772 ( .A(n42612), .X(n42613) );
  inv_x4_sg U43773 ( .A(n42614), .X(n42615) );
  inv_x4_sg U43774 ( .A(n42616), .X(n42617) );
  inv_x1_sg U43775 ( .A(n10390), .X(n42618) );
  nand_x4_sg U43776 ( .A(n10389), .B(n42618), .X(n10300) );
  inv_x1_sg U43777 ( .A(n10390), .X(n51275) );
  inv_x4_sg U43778 ( .A(n42619), .X(n42620) );
  inv_x4_sg U43779 ( .A(n42621), .X(n42622) );
  inv_x4_sg U43780 ( .A(n42623), .X(n42624) );
  inv_x1_sg U43781 ( .A(n14282), .X(n42625) );
  nand_x4_sg U43782 ( .A(n14281), .B(n42625), .X(n14192) );
  inv_x1_sg U43783 ( .A(n14282), .X(n52664) );
  inv_x4_sg U43784 ( .A(n42626), .X(n42627) );
  inv_x4_sg U43785 ( .A(n42628), .X(n42629) );
  inv_x4_sg U43786 ( .A(n31059), .X(n42630) );
  inv_x4_sg U43787 ( .A(n31065), .X(n42632) );
  inv_x4_sg U43788 ( .A(n31071), .X(n42634) );
  inv_x4_sg U43789 ( .A(n30093), .X(n42636) );
  inv_x4_sg U43790 ( .A(n31077), .X(n42638) );
  inv_x4_sg U43791 ( .A(n31083), .X(n42640) );
  inv_x4_sg U43792 ( .A(n30105), .X(n42642) );
  inv_x4_sg U43793 ( .A(n31089), .X(n42644) );
  inv_x4_sg U43794 ( .A(n30111), .X(n42646) );
  inv_x4_sg U43795 ( .A(n31095), .X(n42648) );
  inv_x4_sg U43796 ( .A(n30117), .X(n42650) );
  inv_x4_sg U43797 ( .A(n31101), .X(n42652) );
  inv_x4_sg U43798 ( .A(n30123), .X(n42654) );
  inv_x4_sg U43799 ( .A(n31107), .X(n42656) );
  inv_x4_sg U43800 ( .A(n30129), .X(n42658) );
  inv_x4_sg U43801 ( .A(n31113), .X(n42660) );
  inv_x4_sg U43802 ( .A(n30141), .X(n42662) );
  inv_x4_sg U43803 ( .A(n31125), .X(n42664) );
  inv_x4_sg U43804 ( .A(n30147), .X(n42666) );
  inv_x4_sg U43805 ( .A(n31131), .X(n42668) );
  inv_x4_sg U43806 ( .A(n30153), .X(n42670) );
  inv_x4_sg U43807 ( .A(n31137), .X(n42672) );
  inv_x4_sg U43808 ( .A(n30159), .X(n42674) );
  inv_x4_sg U43809 ( .A(n30932), .X(n42676) );
  inv_x4_sg U43810 ( .A(n30012), .X(n42678) );
  inv_x4_sg U43811 ( .A(n30706), .X(n42680) );
  inv_x4_sg U43812 ( .A(n29846), .X(n42682) );
  inv_x4_sg U43813 ( .A(n30451), .X(n42684) );
  inv_x4_sg U43814 ( .A(n42686), .X(n42687) );
  inv_x4_sg U43815 ( .A(n42688), .X(n42689) );
  inv_x4_sg U43816 ( .A(n42690), .X(n42691) );
  inv_x4_sg U43817 ( .A(n42692), .X(n42693) );
  inv_x4_sg U43818 ( .A(n42694), .X(n42695) );
  inv_x4_sg U43819 ( .A(n42696), .X(n42697) );
  inv_x4_sg U43820 ( .A(n42698), .X(n42699) );
  inv_x4_sg U43821 ( .A(n42700), .X(n42701) );
  inv_x4_sg U43822 ( .A(n23393), .X(n42702) );
  inv_x4_sg U43823 ( .A(n23399), .X(n42704) );
  inv_x4_sg U43824 ( .A(n23405), .X(n42706) );
  inv_x4_sg U43825 ( .A(n22428), .X(n42708) );
  inv_x4_sg U43826 ( .A(n23411), .X(n42710) );
  inv_x4_sg U43827 ( .A(n23417), .X(n42712) );
  inv_x4_sg U43828 ( .A(n22440), .X(n42714) );
  inv_x4_sg U43829 ( .A(n23423), .X(n42716) );
  inv_x4_sg U43830 ( .A(n22446), .X(n42718) );
  inv_x4_sg U43831 ( .A(n23429), .X(n42720) );
  inv_x4_sg U43832 ( .A(n22452), .X(n42722) );
  inv_x4_sg U43833 ( .A(n23435), .X(n42724) );
  inv_x4_sg U43834 ( .A(n22458), .X(n42726) );
  inv_x4_sg U43835 ( .A(n23441), .X(n42728) );
  inv_x4_sg U43836 ( .A(n22464), .X(n42730) );
  inv_x4_sg U43837 ( .A(n23447), .X(n42732) );
  inv_x4_sg U43838 ( .A(n22476), .X(n42734) );
  inv_x4_sg U43839 ( .A(n23459), .X(n42736) );
  inv_x4_sg U43840 ( .A(n22482), .X(n42738) );
  inv_x4_sg U43841 ( .A(n23465), .X(n42740) );
  inv_x4_sg U43842 ( .A(n22488), .X(n42742) );
  inv_x4_sg U43843 ( .A(n23471), .X(n42744) );
  inv_x4_sg U43844 ( .A(n22494), .X(n42746) );
  inv_x4_sg U43845 ( .A(n23266), .X(n42748) );
  inv_x4_sg U43846 ( .A(n22347), .X(n42750) );
  inv_x4_sg U43847 ( .A(n23040), .X(n42752) );
  inv_x4_sg U43848 ( .A(n22181), .X(n42754) );
  inv_x4_sg U43849 ( .A(n22785), .X(n42756) );
  inv_x4_sg U43850 ( .A(n42758), .X(n42759) );
  inv_x4_sg U43851 ( .A(n42760), .X(n42761) );
  inv_x4_sg U43852 ( .A(n42762), .X(n42763) );
  inv_x4_sg U43853 ( .A(n53456), .X(n42764) );
  inv_x4_sg U43854 ( .A(n42764), .X(n42765) );
  inv_x4_sg U43855 ( .A(n42766), .X(n42767) );
  inv_x4_sg U43856 ( .A(n42768), .X(n42769) );
  inv_x4_sg U43857 ( .A(n42770), .X(n42771) );
  inv_x4_sg U43858 ( .A(n30075), .X(n42772) );
  inv_x4_sg U43859 ( .A(n30081), .X(n42774) );
  inv_x4_sg U43860 ( .A(n30087), .X(n42776) );
  inv_x4_sg U43861 ( .A(n30099), .X(n42778) );
  inv_x4_sg U43862 ( .A(n53388), .X(n42780) );
  inv_x4_sg U43863 ( .A(n42780), .X(n42781) );
  inv_x4_sg U43864 ( .A(n22410), .X(n42782) );
  inv_x4_sg U43865 ( .A(n22416), .X(n42784) );
  inv_x4_sg U43866 ( .A(n22422), .X(n42786) );
  inv_x4_sg U43867 ( .A(n22434), .X(n42788) );
  inv_x4_sg U43868 ( .A(n53667), .X(n42790) );
  inv_x4_sg U43869 ( .A(n42790), .X(n42791) );
  inv_x4_sg U43870 ( .A(n53109), .X(n42792) );
  inv_x4_sg U43871 ( .A(n42792), .X(n42793) );
  inv_x4_sg U43872 ( .A(n52550), .X(n42794) );
  inv_x4_sg U43873 ( .A(n42794), .X(n42795) );
  inv_x4_sg U43874 ( .A(n52275), .X(n42796) );
  inv_x4_sg U43875 ( .A(n42796), .X(n42797) );
  inv_x4_sg U43876 ( .A(n51999), .X(n42798) );
  inv_x4_sg U43877 ( .A(n42798), .X(n42799) );
  inv_x4_sg U43878 ( .A(n51721), .X(n42800) );
  inv_x4_sg U43879 ( .A(n42800), .X(n42801) );
  nor_x2_sg U43880 ( .A(n40795), .B(out_L2[5]), .X(n24430) );
  nor_x2_sg U43881 ( .A(n40796), .B(out_L1[5]), .X(n32096) );
  inv_x4_sg U43882 ( .A(n54212), .X(n42802) );
  inv_x4_sg U43883 ( .A(n42802), .X(n42803) );
  inv_x4_sg U43884 ( .A(n42804), .X(n42805) );
  inv_x4_sg U43885 ( .A(n42806), .X(n42807) );
  inv_x4_sg U43886 ( .A(n42808), .X(n42809) );
  inv_x4_sg U43887 ( .A(n42810), .X(n42811) );
  inv_x4_sg U43888 ( .A(n42812), .X(n42813) );
  inv_x4_sg U43889 ( .A(n42814), .X(n42815) );
  inv_x4_sg U43890 ( .A(n42816), .X(n42817) );
  inv_x4_sg U43891 ( .A(n42818), .X(n42819) );
  inv_x4_sg U43892 ( .A(n42820), .X(n42821) );
  inv_x4_sg U43893 ( .A(n42822), .X(n42823) );
  inv_x4_sg U43894 ( .A(n42824), .X(n42825) );
  inv_x4_sg U43895 ( .A(n42826), .X(n42827) );
  inv_x4_sg U43896 ( .A(n42828), .X(n42829) );
  inv_x4_sg U43897 ( .A(n42830), .X(n42831) );
  inv_x4_sg U43898 ( .A(n42832), .X(n42833) );
  inv_x4_sg U43899 ( .A(n42834), .X(n42835) );
  inv_x4_sg U43900 ( .A(n42836), .X(n42837) );
  inv_x4_sg U43901 ( .A(n42838), .X(n42839) );
  inv_x4_sg U43902 ( .A(n42840), .X(n42841) );
  inv_x2_sg U43903 ( .A(n42842), .X(n42843) );
  inv_x2_sg U43904 ( .A(n42844), .X(n42845) );
  inv_x2_sg U43905 ( .A(n42846), .X(n42847) );
  nor_x4_sg U43906 ( .A(n16525), .B(n44679), .X(n16526) );
  nor_x4_sg U43907 ( .A(n14959), .B(n44681), .X(n14960) );
  nor_x4_sg U43908 ( .A(n12626), .B(n44683), .X(n12627) );
  nor_x4_sg U43909 ( .A(n11065), .B(n44685), .X(n11066) );
  inv_x4_sg U43910 ( .A(n42848), .X(n42849) );
  inv_x4_sg U43911 ( .A(n42850), .X(n42851) );
  nand_x4_sg U43912 ( .A(n18564), .B(n18563), .X(n18557) );
  nor_x4_sg U43913 ( .A(n54199), .B(n54178), .X(n18564) );
  inv_x4_sg U43914 ( .A(n42852), .X(n42853) );
  inv_x4_sg U43915 ( .A(n42854), .X(n42855) );
  inv_x2_sg U43916 ( .A(n16692), .X(n44738) );
  inv_x2_sg U43917 ( .A(n15126), .X(n44740) );
  inv_x2_sg U43918 ( .A(n12793), .X(n44742) );
  inv_x2_sg U43919 ( .A(n11232), .X(n44744) );
  inv_x4_sg U43920 ( .A(n42856), .X(n42857) );
  nor_x2_sg U43921 ( .A(n21206), .B(n55329), .X(n21204) );
  inv_x4_sg U43922 ( .A(n42858), .X(n42859) );
  nor_x2_sg U43923 ( .A(n20433), .B(n55047), .X(n20431) );
  inv_x4_sg U43924 ( .A(n42860), .X(n42861) );
  nor_x2_sg U43925 ( .A(n19661), .B(n54761), .X(n19659) );
  inv_x4_sg U43926 ( .A(n42862), .X(n42863) );
  nor_x2_sg U43927 ( .A(n18889), .B(n54479), .X(n18887) );
  inv_x4_sg U43928 ( .A(n42864), .X(n42865) );
  nor_x2_sg U43929 ( .A(n18116), .B(n54194), .X(n18114) );
  inv_x4_sg U43930 ( .A(n42866), .X(n42867) );
  nor_x2_sg U43931 ( .A(n17344), .B(n53914), .X(n17342) );
  inv_x4_sg U43932 ( .A(n42868), .X(n42869) );
  nor_x2_sg U43933 ( .A(n16561), .B(n53630), .X(n16559) );
  inv_x4_sg U43934 ( .A(n42870), .X(n42871) );
  inv_x4_sg U43935 ( .A(n42872), .X(n42873) );
  nor_x2_sg U43936 ( .A(n15779), .B(n53351), .X(n15777) );
  inv_x4_sg U43937 ( .A(n42874), .X(n42875) );
  nor_x2_sg U43938 ( .A(n14995), .B(n53072), .X(n14993) );
  inv_x4_sg U43939 ( .A(n42876), .X(n42877) );
  inv_x4_sg U43940 ( .A(n42878), .X(n42879) );
  nor_x2_sg U43941 ( .A(n14225), .B(n52794), .X(n14223) );
  inv_x4_sg U43942 ( .A(n42880), .X(n42881) );
  nor_x2_sg U43943 ( .A(n13446), .B(n52515), .X(n13444) );
  inv_x4_sg U43944 ( .A(n42882), .X(n42883) );
  nor_x2_sg U43945 ( .A(n12662), .B(n52238), .X(n12660) );
  inv_x4_sg U43946 ( .A(n42884), .X(n42885) );
  inv_x4_sg U43947 ( .A(n42886), .X(n42887) );
  nor_x2_sg U43948 ( .A(n11884), .B(n51963), .X(n11882) );
  inv_x4_sg U43949 ( .A(n42888), .X(n42889) );
  nor_x2_sg U43950 ( .A(n11101), .B(n51682), .X(n11099) );
  inv_x4_sg U43951 ( .A(n42890), .X(n42891) );
  inv_x4_sg U43952 ( .A(n42892), .X(n42893) );
  nor_x2_sg U43953 ( .A(n10333), .B(n51405), .X(n10331) );
  inv_x4_sg U43954 ( .A(n42894), .X(n42895) );
  inv_x2_sg U43955 ( .A(n42896), .X(n42897) );
  inv_x4_sg U43956 ( .A(n42898), .X(n42899) );
  inv_x2_sg U43957 ( .A(n42900), .X(n42901) );
  inv_x4_sg U43958 ( .A(n42902), .X(n42903) );
  inv_x2_sg U43959 ( .A(n42904), .X(n42905) );
  inv_x4_sg U43960 ( .A(n42906), .X(n42907) );
  inv_x2_sg U43961 ( .A(n42908), .X(n42909) );
  inv_x4_sg U43962 ( .A(n42910), .X(n42911) );
  inv_x2_sg U43963 ( .A(n42912), .X(n42913) );
  inv_x4_sg U43964 ( .A(n42914), .X(n42915) );
  inv_x2_sg U43965 ( .A(n42916), .X(n42917) );
  inv_x4_sg U43966 ( .A(n42918), .X(n42919) );
  inv_x2_sg U43967 ( .A(n42920), .X(n42921) );
  inv_x4_sg U43968 ( .A(n42922), .X(n42923) );
  inv_x2_sg U43969 ( .A(n42924), .X(n42925) );
  inv_x4_sg U43970 ( .A(n42926), .X(n42927) );
  inv_x2_sg U43971 ( .A(n42928), .X(n42929) );
  inv_x4_sg U43972 ( .A(n42930), .X(n42931) );
  inv_x2_sg U43973 ( .A(n42932), .X(n42933) );
  inv_x4_sg U43974 ( .A(n42934), .X(n42935) );
  inv_x2_sg U43975 ( .A(n42936), .X(n42937) );
  inv_x2_sg U43976 ( .A(n31285), .X(n42938) );
  nor_x8_sg U43977 ( .A(n31414), .B(n49492), .X(n31285) );
  inv_x4_sg U43978 ( .A(n42939), .X(n42940) );
  inv_x2_sg U43979 ( .A(n42941), .X(n42942) );
  inv_x2_sg U43980 ( .A(n31303), .X(n42943) );
  nor_x8_sg U43981 ( .A(n31405), .B(n49632), .X(n31303) );
  inv_x4_sg U43982 ( .A(n42944), .X(n42945) );
  nor_x2_sg U43983 ( .A(n40761), .B(n49916), .X(n31198) );
  inv_x4_sg U43984 ( .A(n42946), .X(n42947) );
  nor_x2_sg U43985 ( .A(n40762), .B(n50004), .X(n30767) );
  inv_x4_sg U43986 ( .A(n42948), .X(n42949) );
  inv_x2_sg U43987 ( .A(n42950), .X(n42951) );
  inv_x4_sg U43988 ( .A(n42952), .X(n42953) );
  inv_x2_sg U43989 ( .A(n42954), .X(n42955) );
  inv_x4_sg U43990 ( .A(n42956), .X(n42957) );
  inv_x2_sg U43991 ( .A(n42958), .X(n42959) );
  inv_x4_sg U43992 ( .A(n42960), .X(n42961) );
  inv_x2_sg U43993 ( .A(n42962), .X(n42963) );
  inv_x4_sg U43994 ( .A(n42964), .X(n42965) );
  inv_x2_sg U43995 ( .A(n42966), .X(n42967) );
  inv_x4_sg U43996 ( .A(n42968), .X(n42969) );
  inv_x2_sg U43997 ( .A(n42970), .X(n42971) );
  inv_x4_sg U43998 ( .A(n42972), .X(n42973) );
  inv_x2_sg U43999 ( .A(n42974), .X(n42975) );
  inv_x4_sg U44000 ( .A(n42976), .X(n42977) );
  inv_x2_sg U44001 ( .A(n42978), .X(n42979) );
  inv_x4_sg U44002 ( .A(n42980), .X(n42981) );
  inv_x2_sg U44003 ( .A(n42982), .X(n42983) );
  inv_x4_sg U44004 ( .A(n42984), .X(n42985) );
  inv_x2_sg U44005 ( .A(n42986), .X(n42987) );
  inv_x4_sg U44006 ( .A(n42988), .X(n42989) );
  inv_x2_sg U44007 ( .A(n42990), .X(n42991) );
  inv_x4_sg U44008 ( .A(n42992), .X(n42993) );
  inv_x2_sg U44009 ( .A(n42994), .X(n42995) );
  inv_x4_sg U44010 ( .A(n42996), .X(n42997) );
  inv_x2_sg U44011 ( .A(n42998), .X(n42999) );
  inv_x4_sg U44012 ( .A(n43000), .X(n43001) );
  inv_x2_sg U44013 ( .A(n43002), .X(n43003) );
  inv_x4_sg U44014 ( .A(n43004), .X(n43005) );
  inv_x2_sg U44015 ( .A(n43006), .X(n43007) );
  inv_x4_sg U44016 ( .A(n43008), .X(n43009) );
  inv_x2_sg U44017 ( .A(n43010), .X(n43011) );
  inv_x4_sg U44018 ( .A(n43012), .X(n43013) );
  inv_x2_sg U44019 ( .A(n43014), .X(n43015) );
  inv_x4_sg U44020 ( .A(n43016), .X(n43017) );
  inv_x2_sg U44021 ( .A(n43018), .X(n43019) );
  inv_x2_sg U44022 ( .A(n23619), .X(n43020) );
  nor_x8_sg U44023 ( .A(n23748), .B(n50351), .X(n23619) );
  inv_x4_sg U44024 ( .A(n43021), .X(n43022) );
  inv_x2_sg U44025 ( .A(n43023), .X(n43024) );
  inv_x2_sg U44026 ( .A(n23637), .X(n43025) );
  nor_x8_sg U44027 ( .A(n23739), .B(n50491), .X(n23637) );
  inv_x4_sg U44028 ( .A(n43026), .X(n43027) );
  nor_x2_sg U44029 ( .A(n40763), .B(n50775), .X(n23532) );
  inv_x4_sg U44030 ( .A(n43028), .X(n43029) );
  nor_x2_sg U44031 ( .A(n40764), .B(n50863), .X(n23101) );
  inv_x4_sg U44032 ( .A(n43030), .X(n43031) );
  nor_x2_sg U44033 ( .A(n55086), .B(n55013), .X(n21060) );
  inv_x4_sg U44034 ( .A(n43032), .X(n43033) );
  nor_x2_sg U44035 ( .A(n54518), .B(n54445), .X(n19516) );
  inv_x4_sg U44036 ( .A(n43034), .X(n43035) );
  nor_x2_sg U44037 ( .A(n53953), .B(n53880), .X(n17971) );
  inv_x4_sg U44038 ( .A(n43036), .X(n43037) );
  nor_x2_sg U44039 ( .A(n53680), .B(n53595), .X(n17198) );
  inv_x2_sg U44040 ( .A(n43038), .X(n43039) );
  inv_x4_sg U44041 ( .A(n43040), .X(n43041) );
  nor_x2_sg U44042 ( .A(n53122), .B(n53037), .X(n15632) );
  inv_x4_sg U44043 ( .A(n43042), .X(n43043) );
  nor_x2_sg U44044 ( .A(n52563), .B(n52480), .X(n14079) );
  inv_x4_sg U44045 ( .A(n43044), .X(n43045) );
  nor_x2_sg U44046 ( .A(n52288), .B(n52203), .X(n13299) );
  inv_x4_sg U44047 ( .A(n43046), .X(n43047) );
  nor_x2_sg U44048 ( .A(n52011), .B(n51928), .X(n12518) );
  inv_x4_sg U44049 ( .A(n43048), .X(n43049) );
  nor_x2_sg U44050 ( .A(n51733), .B(n51647), .X(n11738) );
  inv_x4_sg U44051 ( .A(n43050), .X(n43051) );
  nor_x2_sg U44052 ( .A(n53403), .B(n53316), .X(n16412) );
  inv_x2_sg U44053 ( .A(n43052), .X(n43053) );
  inv_x4_sg U44054 ( .A(n43054), .X(n43055) );
  nor_x2_sg U44055 ( .A(n44375), .B(n21752), .X(n21749) );
  inv_x4_sg U44056 ( .A(n43056), .X(n43057) );
  nor_x2_sg U44057 ( .A(n44034), .B(n20982), .X(n20979) );
  inv_x2_sg U44058 ( .A(n43058), .X(n43059) );
  inv_x2_sg U44059 ( .A(n43060), .X(n43061) );
  inv_x4_sg U44060 ( .A(n43062), .X(n43063) );
  nor_x2_sg U44061 ( .A(n44377), .B(n20207), .X(n20204) );
  inv_x4_sg U44062 ( .A(n43064), .X(n43065) );
  nor_x2_sg U44063 ( .A(n44036), .B(n19438), .X(n19435) );
  inv_x2_sg U44064 ( .A(n43066), .X(n43067) );
  inv_x2_sg U44065 ( .A(n43068), .X(n43069) );
  inv_x4_sg U44066 ( .A(n43070), .X(n43071) );
  nor_x2_sg U44067 ( .A(n44213), .B(n18662), .X(n18659) );
  inv_x4_sg U44068 ( .A(n43072), .X(n43073) );
  nor_x2_sg U44069 ( .A(n44038), .B(n17893), .X(n17890) );
  inv_x2_sg U44070 ( .A(n43074), .X(n43075) );
  inv_x2_sg U44071 ( .A(n43076), .X(n43077) );
  inv_x2_sg U44072 ( .A(n43078), .X(n43079) );
  inv_x4_sg U44073 ( .A(n43080), .X(n43081) );
  nor_x2_sg U44074 ( .A(n44215), .B(n14772), .X(n14769) );
  inv_x2_sg U44075 ( .A(n43082), .X(n43083) );
  inv_x2_sg U44076 ( .A(n43084), .X(n43085) );
  inv_x2_sg U44077 ( .A(n43086), .X(n43087) );
  inv_x2_sg U44078 ( .A(n43088), .X(n43089) );
  inv_x2_sg U44079 ( .A(n43090), .X(n43091) );
  inv_x4_sg U44080 ( .A(n43092), .X(n43093) );
  nor_x2_sg U44081 ( .A(n44102), .B(n11659), .X(n11657) );
  inv_x4_sg U44082 ( .A(n43094), .X(n43095) );
  nor_x2_sg U44083 ( .A(n44379), .B(n10879), .X(n10877) );
  inv_x4_sg U44084 ( .A(n21850), .X(n43096) );
  inv_x4_sg U44085 ( .A(n20305), .X(n43098) );
  inv_x4_sg U44086 ( .A(n43102), .X(n43103) );
  inv_x4_sg U44087 ( .A(n43104), .X(n43105) );
  inv_x4_sg U44088 ( .A(n43106), .X(n43107) );
  inv_x4_sg U44089 ( .A(n43108), .X(n43109) );
  inv_x4_sg U44090 ( .A(n43110), .X(n43111) );
  inv_x2_sg U44091 ( .A(n43112), .X(n43113) );
  nor_x2_sg U44092 ( .A(n10406), .B(n10407), .X(n10405) );
  inv_x4_sg U44093 ( .A(n43114), .X(n43115) );
  inv_x2_sg U44094 ( .A(n43116), .X(n43117) );
  nor_x2_sg U44095 ( .A(n21278), .B(n21279), .X(n21277) );
  inv_x4_sg U44096 ( .A(n43118), .X(n43119) );
  inv_x2_sg U44097 ( .A(n43120), .X(n43121) );
  nor_x2_sg U44098 ( .A(n19733), .B(n19734), .X(n19732) );
  inv_x4_sg U44099 ( .A(n43122), .X(n43123) );
  nor_x2_sg U44100 ( .A(n53513), .B(n16638), .X(n16637) );
  inv_x4_sg U44101 ( .A(n44670), .X(n53513) );
  inv_x4_sg U44102 ( .A(n43124), .X(n43125) );
  nor_x2_sg U44103 ( .A(n52955), .B(n15072), .X(n15071) );
  inv_x4_sg U44104 ( .A(n44672), .X(n52955) );
  inv_x4_sg U44105 ( .A(n43126), .X(n43127) );
  nor_x2_sg U44106 ( .A(n52121), .B(n12739), .X(n12738) );
  inv_x4_sg U44107 ( .A(n44674), .X(n52121) );
  inv_x4_sg U44108 ( .A(n43128), .X(n43129) );
  nor_x2_sg U44109 ( .A(n51564), .B(n11178), .X(n11177) );
  inv_x4_sg U44110 ( .A(n44676), .X(n51564) );
  inv_x4_sg U44111 ( .A(n43130), .X(n43131) );
  inv_x2_sg U44112 ( .A(n43132), .X(n43133) );
  inv_x4_sg U44113 ( .A(n43134), .X(n43135) );
  inv_x2_sg U44114 ( .A(n43136), .X(n43137) );
  nor_x2_sg U44115 ( .A(n51162), .B(n46043), .X(n28372) );
  inv_x4_sg U44116 ( .A(n43138), .X(n43139) );
  inv_x4_sg U44117 ( .A(n15850), .X(n43140) );
  nor_x2_sg U44118 ( .A(n15857), .B(n53221), .X(n15854) );
  inv_x4_sg U44119 ( .A(n43142), .X(n43143) );
  inv_x2_sg U44120 ( .A(n43144), .X(n43145) );
  inv_x4_sg U44121 ( .A(n43146), .X(n43147) );
  nor_x2_sg U44122 ( .A(n14298), .B(n14299), .X(n14297) );
  inv_x4_sg U44123 ( .A(n43148), .X(n43149) );
  inv_x2_sg U44124 ( .A(n43150), .X(n43151) );
  inv_x4_sg U44125 ( .A(n43152), .X(n43153) );
  inv_x2_sg U44126 ( .A(n43154), .X(n43155) );
  inv_x4_sg U44127 ( .A(n43156), .X(n43157) );
  inv_x2_sg U44128 ( .A(n43158), .X(n43159) );
  inv_x4_sg U44129 ( .A(n43160), .X(n43161) );
  nor_x2_sg U44130 ( .A(n45270), .B(n46117), .X(n28385) );
  inv_x4_sg U44131 ( .A(n43162), .X(n43163) );
  inv_x2_sg U44132 ( .A(n43164), .X(n43165) );
  inv_x4_sg U44133 ( .A(n27900), .X(n55465) );
  nand_x8_sg U44134 ( .A(n55462), .B(n29612), .X(n27900) );
  inv_x4_sg U44135 ( .A(n43166), .X(n43167) );
  inv_x2_sg U44136 ( .A(n43168), .X(n43169) );
  nor_x2_sg U44137 ( .A(n29426), .B(n55451), .X(n29425) );
  nor_x4_sg U44138 ( .A(n46203), .B(n29420), .X(n29426) );
  nor_x2_sg U44139 ( .A(n29144), .B(n55167), .X(n29143) );
  nor_x4_sg U44140 ( .A(n46205), .B(n29138), .X(n29144) );
  nor_x2_sg U44141 ( .A(n28865), .B(n54883), .X(n28864) );
  nor_x4_sg U44142 ( .A(n46207), .B(n28859), .X(n28865) );
  nor_x2_sg U44143 ( .A(n28585), .B(n54599), .X(n28584) );
  nor_x4_sg U44144 ( .A(n46209), .B(n28579), .X(n28585) );
  nor_x2_sg U44145 ( .A(n28307), .B(n54315), .X(n28306) );
  nor_x4_sg U44146 ( .A(n46211), .B(n28301), .X(n28307) );
  nor_x2_sg U44147 ( .A(n28027), .B(n54034), .X(n28026) );
  nor_x4_sg U44148 ( .A(n46213), .B(n28021), .X(n28027) );
  nor_x2_sg U44149 ( .A(n27748), .B(n53750), .X(n27747) );
  nor_x4_sg U44150 ( .A(n46215), .B(n27742), .X(n27748) );
  nor_x2_sg U44151 ( .A(n27467), .B(n53472), .X(n27466) );
  nor_x4_sg U44152 ( .A(n46217), .B(n27461), .X(n27467) );
  nor_x2_sg U44153 ( .A(n27188), .B(n53192), .X(n27187) );
  nor_x4_sg U44154 ( .A(n46219), .B(n27182), .X(n27188) );
  nor_x2_sg U44155 ( .A(n26908), .B(n52914), .X(n26907) );
  nor_x4_sg U44156 ( .A(n46221), .B(n26902), .X(n26908) );
  nor_x2_sg U44157 ( .A(n26631), .B(n52633), .X(n26630) );
  nor_x4_sg U44158 ( .A(n46223), .B(n26625), .X(n26631) );
  nor_x2_sg U44159 ( .A(n26352), .B(n52358), .X(n26351) );
  nor_x4_sg U44160 ( .A(n46225), .B(n26346), .X(n26352) );
  nor_x2_sg U44161 ( .A(n26071), .B(n52080), .X(n26070) );
  nor_x4_sg U44162 ( .A(n46227), .B(n26065), .X(n26071) );
  nor_x2_sg U44163 ( .A(n25792), .B(n51804), .X(n25791) );
  nor_x4_sg U44164 ( .A(n46229), .B(n25786), .X(n25792) );
  inv_x4_sg U44165 ( .A(n13621), .X(n43170) );
  nor_x2_sg U44166 ( .A(n13624), .B(n13625), .X(n13623) );
  nor_x4_sg U44167 ( .A(n16072), .B(n16071), .X(n16090) );
  inv_x4_sg U44168 ( .A(n16334), .X(n43172) );
  inv_x2_sg U44169 ( .A(n43174), .X(n43175) );
  nor_x2_sg U44170 ( .A(n16357), .B(n16501), .X(n16499) );
  nor_x4_sg U44171 ( .A(n11397), .B(n11396), .X(n11415) );
  nor_x4_sg U44172 ( .A(n10607), .B(n51359), .X(n10599) );
  nor_x4_sg U44173 ( .A(n21479), .B(n55281), .X(n21471) );
  nor_x4_sg U44174 ( .A(n19934), .B(n54713), .X(n19926) );
  nor_x4_sg U44175 ( .A(n18389), .B(n54148), .X(n18381) );
  nor_x4_sg U44176 ( .A(n20709), .B(n55009), .X(n20701) );
  nor_x4_sg U44177 ( .A(n19165), .B(n54441), .X(n19157) );
  nor_x4_sg U44178 ( .A(n17620), .B(n53876), .X(n17612) );
  nor_x4_sg U44179 ( .A(n14499), .B(n52756), .X(n14491) );
  nor_x2_sg U44180 ( .A(n40737), .B(out_L2[4]), .X(n24424) );
  nor_x2_sg U44181 ( .A(n40738), .B(out_L1[4]), .X(n32090) );
  nor_x2_sg U44182 ( .A(n21888), .B(n55375), .X(n21887) );
  nor_x2_sg U44183 ( .A(n55375), .B(n55389), .X(n21879) );
  inv_x4_sg U44184 ( .A(n41812), .X(n55375) );
  nor_x2_sg U44185 ( .A(n20343), .B(n54807), .X(n20342) );
  nor_x2_sg U44186 ( .A(n54807), .B(n54821), .X(n20334) );
  inv_x4_sg U44187 ( .A(n41814), .X(n54807) );
  inv_x4_sg U44188 ( .A(n43176), .X(n43177) );
  inv_x4_sg U44189 ( .A(n43178), .X(n43179) );
  inv_x2_sg U44190 ( .A(n43180), .X(n43181) );
  inv_x4_sg U44191 ( .A(n43182), .X(n43183) );
  inv_x2_sg U44192 ( .A(n43184), .X(n43185) );
  inv_x4_sg U44193 ( .A(n43186), .X(n43187) );
  inv_x2_sg U44194 ( .A(n43188), .X(n43189) );
  inv_x4_sg U44195 ( .A(n43190), .X(n43191) );
  inv_x2_sg U44196 ( .A(n43192), .X(n43193) );
  inv_x4_sg U44197 ( .A(n43194), .X(n43195) );
  inv_x4_sg U44198 ( .A(n43196), .X(n43197) );
  inv_x4_sg U44199 ( .A(n43198), .X(n43199) );
  inv_x4_sg U44200 ( .A(n43200), .X(n43201) );
  inv_x4_sg U44201 ( .A(n43202), .X(n43203) );
  nor_x4_sg U44202 ( .A(n15979), .B(n15983), .X(n15981) );
  nor_x4_sg U44203 ( .A(n15978), .B(n15977), .X(n15979) );
  inv_x4_sg U44204 ( .A(n43204), .X(n43205) );
  nor_x2_sg U44205 ( .A(n10556), .B(n10555), .X(n10553) );
  inv_x4_sg U44206 ( .A(n43206), .X(n43207) );
  nor_x2_sg U44207 ( .A(n21428), .B(n21427), .X(n21425) );
  inv_x4_sg U44208 ( .A(n43208), .X(n43209) );
  nor_x2_sg U44209 ( .A(n19883), .B(n19882), .X(n19880) );
  inv_x4_sg U44210 ( .A(n43210), .X(n43211) );
  nor_x2_sg U44211 ( .A(n18338), .B(n18337), .X(n18335) );
  nor_x4_sg U44212 ( .A(n12084), .B(n12088), .X(n12086) );
  nor_x4_sg U44213 ( .A(n12083), .B(n12082), .X(n12084) );
  nor_x4_sg U44214 ( .A(n11304), .B(n11308), .X(n11306) );
  nor_x4_sg U44215 ( .A(n11303), .B(n11302), .X(n11304) );
  inv_x4_sg U44216 ( .A(n43212), .X(n43213) );
  nor_x2_sg U44217 ( .A(n20657), .B(n20656), .X(n20654) );
  inv_x4_sg U44218 ( .A(n43214), .X(n43215) );
  nor_x2_sg U44219 ( .A(n19113), .B(n19112), .X(n19110) );
  inv_x4_sg U44220 ( .A(n43216), .X(n43217) );
  nor_x2_sg U44221 ( .A(n17568), .B(n17567), .X(n17565) );
  inv_x4_sg U44222 ( .A(n43218), .X(n43219) );
  nor_x2_sg U44223 ( .A(n14448), .B(n14447), .X(n14445) );
  inv_x4_sg U44224 ( .A(n43220), .X(n43221) );
  nor_x2_sg U44225 ( .A(n46563), .B(n10508), .X(n10542) );
  inv_x4_sg U44226 ( .A(n43222), .X(n43223) );
  nor_x4_sg U44227 ( .A(n16060), .B(n53312), .X(n16053) );
  nand_x4_sg U44228 ( .A(n53248), .B(n16029), .X(n16060) );
  nor_x4_sg U44229 ( .A(n11385), .B(n51644), .X(n11378) );
  nand_x4_sg U44230 ( .A(n51581), .B(n11354), .X(n11385) );
  nor_x4_sg U44231 ( .A(n46274), .B(n54905), .X(n20491) );
  nor_x4_sg U44232 ( .A(n46319), .B(n54337), .X(n18947) );
  nor_x4_sg U44233 ( .A(n46366), .B(n53772), .X(n17402) );
  nor_x4_sg U44234 ( .A(n54900), .B(n20491), .X(n20396) );
  inv_x4_sg U44235 ( .A(n20393), .X(n54900) );
  nor_x4_sg U44236 ( .A(n54332), .B(n18947), .X(n18852) );
  inv_x4_sg U44237 ( .A(n18849), .X(n54332) );
  nor_x4_sg U44238 ( .A(n53767), .B(n17402), .X(n17307) );
  inv_x4_sg U44239 ( .A(n17304), .X(n53767) );
  inv_x4_sg U44240 ( .A(n21221), .X(n43224) );
  inv_x4_sg U44241 ( .A(n19676), .X(n43226) );
  inv_x4_sg U44242 ( .A(n18131), .X(n43228) );
  inv_x4_sg U44243 ( .A(n11899), .X(n43230) );
  nor_x4_sg U44244 ( .A(n18285), .B(n18286), .X(n18280) );
  inv_x4_sg U44245 ( .A(n21403), .X(n43232) );
  inv_x4_sg U44246 ( .A(n43232), .X(n43233) );
  inv_x4_sg U44247 ( .A(n19858), .X(n43234) );
  inv_x4_sg U44248 ( .A(n43234), .X(n43235) );
  inv_x4_sg U44249 ( .A(n16768), .X(n43236) );
  inv_x4_sg U44250 ( .A(n43236), .X(n43237) );
  inv_x4_sg U44251 ( .A(n15202), .X(n43238) );
  inv_x4_sg U44252 ( .A(n43238), .X(n43239) );
  nor_x4_sg U44253 ( .A(n13655), .B(n44074), .X(n13649) );
  inv_x4_sg U44254 ( .A(n12869), .X(n43240) );
  inv_x4_sg U44255 ( .A(n43240), .X(n43241) );
  inv_x4_sg U44256 ( .A(n20632), .X(n43242) );
  inv_x4_sg U44257 ( .A(n43242), .X(n43243) );
  inv_x4_sg U44258 ( .A(n19088), .X(n43244) );
  inv_x4_sg U44259 ( .A(n43244), .X(n43245) );
  inv_x4_sg U44260 ( .A(n17543), .X(n43246) );
  inv_x4_sg U44261 ( .A(n43246), .X(n43247) );
  inv_x4_sg U44262 ( .A(n14423), .X(n43248) );
  inv_x4_sg U44263 ( .A(n43248), .X(n43249) );
  inv_x4_sg U44264 ( .A(n43250), .X(n43251) );
  nor_x4_sg U44265 ( .A(n20605), .B(n54974), .X(n20601) );
  nand_x4_sg U44266 ( .A(n54974), .B(n20605), .X(n20599) );
  nor_x4_sg U44267 ( .A(n54984), .B(n43251), .X(n20605) );
  inv_x4_sg U44268 ( .A(n20624), .X(n54984) );
  nand_x2_sg U44269 ( .A(n20622), .B(n20623), .X(n20624) );
  inv_x4_sg U44270 ( .A(n43252), .X(n43253) );
  nor_x4_sg U44271 ( .A(n19061), .B(n54406), .X(n19057) );
  nand_x4_sg U44272 ( .A(n54406), .B(n19061), .X(n19055) );
  nor_x4_sg U44273 ( .A(n54416), .B(n43253), .X(n19061) );
  inv_x4_sg U44274 ( .A(n19080), .X(n54416) );
  nand_x2_sg U44275 ( .A(n19078), .B(n19079), .X(n19080) );
  inv_x4_sg U44276 ( .A(n43254), .X(n43255) );
  nor_x4_sg U44277 ( .A(n17516), .B(n53841), .X(n17512) );
  nand_x4_sg U44278 ( .A(n53841), .B(n17516), .X(n17510) );
  nor_x4_sg U44279 ( .A(n53851), .B(n43255), .X(n17516) );
  inv_x4_sg U44280 ( .A(n17535), .X(n53851) );
  nand_x2_sg U44281 ( .A(n17533), .B(n17534), .X(n17535) );
  inv_x4_sg U44282 ( .A(n43256), .X(n43257) );
  inv_x4_sg U44283 ( .A(n43258), .X(n43259) );
  inv_x4_sg U44284 ( .A(n43260), .X(n43261) );
  inv_x4_sg U44285 ( .A(n43262), .X(n43263) );
  inv_x4_sg U44286 ( .A(n43264), .X(n43265) );
  inv_x4_sg U44287 ( .A(n16172), .X(n43266) );
  nor_x2_sg U44288 ( .A(n44439), .B(n16219), .X(n16216) );
  inv_x4_sg U44289 ( .A(n16957), .X(n43268) );
  nor_x2_sg U44290 ( .A(n44183), .B(n17004), .X(n17001) );
  inv_x4_sg U44291 ( .A(n15391), .X(n43270) );
  nor_x2_sg U44292 ( .A(n44185), .B(n15438), .X(n15435) );
  inv_x4_sg U44293 ( .A(n13838), .X(n43272) );
  nor_x2_sg U44294 ( .A(n44187), .B(n13885), .X(n13882) );
  inv_x4_sg U44295 ( .A(n13058), .X(n43274) );
  nor_x2_sg U44296 ( .A(n44189), .B(n13105), .X(n13102) );
  inv_x4_sg U44297 ( .A(n11497), .X(n43276) );
  nor_x2_sg U44298 ( .A(n44193), .B(n11544), .X(n11541) );
  inv_x4_sg U44299 ( .A(n20818), .X(n43288) );
  nor_x2_sg U44300 ( .A(n44449), .B(n20864), .X(n20861) );
  inv_x4_sg U44301 ( .A(n19274), .X(n43290) );
  nor_x2_sg U44302 ( .A(n44451), .B(n19320), .X(n19317) );
  inv_x4_sg U44303 ( .A(n17729), .X(n43292) );
  nor_x2_sg U44304 ( .A(n44453), .B(n17775), .X(n17772) );
  inv_x4_sg U44305 ( .A(n14608), .X(n43294) );
  nor_x2_sg U44306 ( .A(n44455), .B(n14654), .X(n14651) );
  inv_x4_sg U44307 ( .A(n12331), .X(n43302) );
  inv_x4_sg U44308 ( .A(n16141), .X(n43304) );
  inv_x2_sg U44309 ( .A(n43306), .X(n43307) );
  inv_x4_sg U44310 ( .A(n12269), .X(n43308) );
  nor_x2_sg U44311 ( .A(n12346), .B(n12347), .X(n12345) );
  nor_x4_sg U44312 ( .A(n51964), .B(n51947), .X(n12347) );
  inv_x4_sg U44313 ( .A(n12246), .X(n43310) );
  inv_x2_sg U44314 ( .A(n43312), .X(n43313) );
  inv_x4_sg U44315 ( .A(n10685), .X(n43314) );
  inv_x2_sg U44316 ( .A(n43316), .X(n43317) );
  inv_x4_sg U44317 ( .A(n21557), .X(n43318) );
  inv_x2_sg U44318 ( .A(n43320), .X(n43321) );
  inv_x4_sg U44319 ( .A(n20012), .X(n43322) );
  inv_x2_sg U44320 ( .A(n43324), .X(n43325) );
  inv_x4_sg U44321 ( .A(n20787), .X(n43326) );
  inv_x2_sg U44322 ( .A(n43328), .X(n43329) );
  inv_x4_sg U44323 ( .A(n19243), .X(n43330) );
  inv_x2_sg U44324 ( .A(n43332), .X(n43333) );
  inv_x4_sg U44325 ( .A(n17698), .X(n43334) );
  inv_x2_sg U44326 ( .A(n43336), .X(n43337) );
  inv_x4_sg U44327 ( .A(n14577), .X(n43338) );
  inv_x2_sg U44328 ( .A(n43340), .X(n43341) );
  inv_x4_sg U44329 ( .A(n14600), .X(n43344) );
  nor_x2_sg U44330 ( .A(n14676), .B(n14677), .X(n14675) );
  nor_x4_sg U44331 ( .A(n52778), .B(n52795), .X(n14677) );
  inv_x4_sg U44332 ( .A(n43346), .X(n43347) );
  inv_x4_sg U44333 ( .A(n43348), .X(n43349) );
  inv_x4_sg U44334 ( .A(n43350), .X(n43351) );
  nor_x4_sg U44335 ( .A(n53335), .B(n53353), .X(n16242) );
  inv_x8_sg U44336 ( .A(n16197), .X(n53353) );
  nor_x4_sg U44337 ( .A(n55335), .B(n55313), .X(n21656) );
  inv_x8_sg U44338 ( .A(n21613), .X(n55335) );
  nor_x4_sg U44339 ( .A(n54767), .B(n54745), .X(n20111) );
  inv_x8_sg U44340 ( .A(n20068), .X(n54767) );
  inv_x4_sg U44341 ( .A(n43352), .X(n43353) );
  inv_x4_sg U44342 ( .A(n43354), .X(n43355) );
  inv_x4_sg U44343 ( .A(n43356), .X(n43357) );
  inv_x4_sg U44344 ( .A(n43358), .X(n43359) );
  inv_x4_sg U44345 ( .A(n43360), .X(n43361) );
  inv_x4_sg U44346 ( .A(n43362), .X(n43363) );
  inv_x4_sg U44347 ( .A(n43364), .X(n43365) );
  nor_x4_sg U44348 ( .A(n15951), .B(n15950), .X(n15827) );
  nor_x4_sg U44349 ( .A(n10503), .B(n10502), .X(n10382) );
  nor_x4_sg U44350 ( .A(n21375), .B(n21374), .X(n21254) );
  nor_x4_sg U44351 ( .A(n19830), .B(n19829), .X(n19709) );
  nor_x4_sg U44352 ( .A(n18284), .B(n18283), .X(n18164) );
  nor_x4_sg U44353 ( .A(n16737), .B(n16736), .X(n16609) );
  nor_x4_sg U44354 ( .A(n15171), .B(n15170), .X(n15043) );
  nor_x4_sg U44355 ( .A(n13617), .B(n42449), .X(n13494) );
  nor_x4_sg U44356 ( .A(n12838), .B(n12837), .X(n12710) );
  nor_x4_sg U44357 ( .A(n12056), .B(n12055), .X(n11932) );
  nor_x4_sg U44358 ( .A(n11277), .B(n11276), .X(n11149) );
  nor_x4_sg U44359 ( .A(n20604), .B(n20603), .X(n20482) );
  nor_x4_sg U44360 ( .A(n19060), .B(n19059), .X(n18938) );
  nor_x4_sg U44361 ( .A(n17515), .B(n17514), .X(n17393) );
  nor_x4_sg U44362 ( .A(n14394), .B(n14393), .X(n14274) );
  inv_x4_sg U44363 ( .A(n43366), .X(n43367) );
  inv_x4_sg U44364 ( .A(n43368), .X(n43369) );
  nor_x4_sg U44365 ( .A(n43367), .B(n43369), .X(n21189) );
  inv_x4_sg U44366 ( .A(n43370), .X(n43371) );
  inv_x4_sg U44367 ( .A(n43372), .X(n43373) );
  nor_x4_sg U44368 ( .A(n43371), .B(n43373), .X(n20416) );
  inv_x4_sg U44369 ( .A(n43374), .X(n43375) );
  inv_x4_sg U44370 ( .A(n43376), .X(n43377) );
  nor_x4_sg U44371 ( .A(n43375), .B(n43377), .X(n19644) );
  inv_x4_sg U44372 ( .A(n43378), .X(n43379) );
  inv_x4_sg U44373 ( .A(n43380), .X(n43381) );
  nor_x4_sg U44374 ( .A(n43379), .B(n43381), .X(n18872) );
  inv_x4_sg U44375 ( .A(n43382), .X(n43383) );
  inv_x4_sg U44376 ( .A(n43384), .X(n43385) );
  nor_x4_sg U44377 ( .A(n43383), .B(n43385), .X(n17327) );
  inv_x4_sg U44378 ( .A(n43386), .X(n43387) );
  inv_x4_sg U44379 ( .A(n43388), .X(n43389) );
  nor_x4_sg U44380 ( .A(n43387), .B(n43389), .X(n16544) );
  inv_x4_sg U44381 ( .A(n43390), .X(n43391) );
  inv_x4_sg U44382 ( .A(n43392), .X(n43393) );
  nor_x4_sg U44383 ( .A(n43391), .B(n43393), .X(n15762) );
  inv_x4_sg U44384 ( .A(n43394), .X(n43395) );
  inv_x4_sg U44385 ( .A(n43396), .X(n43397) );
  nor_x4_sg U44386 ( .A(n43395), .B(n43397), .X(n14978) );
  inv_x4_sg U44387 ( .A(n43398), .X(n43399) );
  inv_x4_sg U44388 ( .A(n43400), .X(n43401) );
  nor_x4_sg U44389 ( .A(n43399), .B(n43401), .X(n14208) );
  inv_x4_sg U44390 ( .A(n43402), .X(n43403) );
  inv_x4_sg U44391 ( .A(n43404), .X(n43405) );
  nor_x4_sg U44392 ( .A(n43403), .B(n43405), .X(n13429) );
  inv_x4_sg U44393 ( .A(n43406), .X(n43407) );
  inv_x4_sg U44394 ( .A(n43408), .X(n43409) );
  nor_x4_sg U44395 ( .A(n43407), .B(n43409), .X(n12645) );
  inv_x4_sg U44396 ( .A(n43410), .X(n43411) );
  inv_x4_sg U44397 ( .A(n43412), .X(n43413) );
  nor_x4_sg U44398 ( .A(n43411), .B(n43413), .X(n11867) );
  inv_x4_sg U44399 ( .A(n43414), .X(n43415) );
  inv_x4_sg U44400 ( .A(n43416), .X(n43417) );
  nor_x4_sg U44401 ( .A(n43415), .B(n43417), .X(n11084) );
  inv_x4_sg U44402 ( .A(n43418), .X(n43419) );
  inv_x4_sg U44403 ( .A(n43420), .X(n43421) );
  nor_x4_sg U44404 ( .A(n43419), .B(n43421), .X(n10316) );
  nor_x4_sg U44405 ( .A(n53632), .B(n17024), .X(n16949) );
  inv_x4_sg U44406 ( .A(n17018), .X(n53632) );
  nor_x4_sg U44407 ( .A(n17025), .B(n17026), .X(n17024) );
  nor_x4_sg U44408 ( .A(n53614), .B(n53631), .X(n17026) );
  nor_x4_sg U44409 ( .A(n53074), .B(n15458), .X(n15383) );
  inv_x4_sg U44410 ( .A(n15452), .X(n53074) );
  nor_x4_sg U44411 ( .A(n15459), .B(n15460), .X(n15458) );
  nor_x4_sg U44412 ( .A(n53056), .B(n53073), .X(n15460) );
  inv_x4_sg U44413 ( .A(n13899), .X(n43422) );
  nor_x4_sg U44414 ( .A(n43422), .B(n13905), .X(n13830) );
  nor_x4_sg U44415 ( .A(n13906), .B(n13907), .X(n13905) );
  nor_x4_sg U44416 ( .A(n52499), .B(n52516), .X(n13907) );
  nor_x4_sg U44417 ( .A(n52240), .B(n13125), .X(n13050) );
  inv_x4_sg U44418 ( .A(n13119), .X(n52240) );
  nor_x4_sg U44419 ( .A(n13126), .B(n13127), .X(n13125) );
  nor_x4_sg U44420 ( .A(n52222), .B(n52239), .X(n13127) );
  nor_x4_sg U44421 ( .A(n51685), .B(n11564), .X(n11489) );
  inv_x4_sg U44422 ( .A(n11558), .X(n51685) );
  nor_x4_sg U44423 ( .A(n11565), .B(n11566), .X(n11564) );
  nor_x4_sg U44424 ( .A(n51666), .B(n51684), .X(n11566) );
  inv_x4_sg U44425 ( .A(n43423), .X(n43424) );
  inv_x4_sg U44426 ( .A(n43425), .X(n43426) );
  nor_x2_sg U44427 ( .A(n16926), .B(n16927), .X(n16938) );
  nor_x4_sg U44428 ( .A(n43424), .B(n43426), .X(n16926) );
  inv_x4_sg U44429 ( .A(n43427), .X(n43428) );
  inv_x4_sg U44430 ( .A(n43429), .X(n43430) );
  nor_x2_sg U44431 ( .A(n15360), .B(n15361), .X(n15372) );
  nor_x4_sg U44432 ( .A(n43428), .B(n43430), .X(n15360) );
  inv_x4_sg U44433 ( .A(n43431), .X(n43432) );
  inv_x4_sg U44434 ( .A(n43433), .X(n43434) );
  nor_x2_sg U44435 ( .A(n13807), .B(n13808), .X(n13819) );
  nor_x4_sg U44436 ( .A(n43432), .B(n43434), .X(n13807) );
  inv_x4_sg U44437 ( .A(n43435), .X(n43436) );
  inv_x4_sg U44438 ( .A(n43437), .X(n43438) );
  nor_x2_sg U44439 ( .A(n13027), .B(n13028), .X(n13039) );
  nor_x4_sg U44440 ( .A(n43436), .B(n43438), .X(n13027) );
  inv_x4_sg U44441 ( .A(n43439), .X(n43440) );
  inv_x4_sg U44442 ( .A(n43441), .X(n43442) );
  nor_x2_sg U44443 ( .A(n11466), .B(n11467), .X(n11478) );
  nor_x4_sg U44444 ( .A(n43440), .B(n43442), .X(n11466) );
  inv_x4_sg U44445 ( .A(n43443), .X(n43444) );
  inv_x4_sg U44446 ( .A(n31258), .X(n49329) );
  nor_x4_sg U44447 ( .A(n43444), .B(n49328), .X(n31258) );
  inv_x4_sg U44448 ( .A(n31437), .X(n49328) );
  nand_x2_sg U44449 ( .A(n25262), .B(n41956), .X(n31437) );
  inv_x4_sg U44450 ( .A(n43445), .X(n43446) );
  inv_x4_sg U44451 ( .A(n23592), .X(n50188) );
  nor_x4_sg U44452 ( .A(n43446), .B(n50187), .X(n23592) );
  inv_x4_sg U44453 ( .A(n23771), .X(n50187) );
  nand_x2_sg U44454 ( .A(n10154), .B(n41958), .X(n23771) );
  inv_x4_sg U44455 ( .A(n43447), .X(n43448) );
  nor_x2_sg U44456 ( .A(n16459), .B(n16458), .X(n16492) );
  nor_x4_sg U44457 ( .A(n43448), .B(n53332), .X(n16459) );
  inv_x4_sg U44458 ( .A(n16495), .X(n53332) );
  nand_x2_sg U44459 ( .A(n16457), .B(n16496), .X(n16495) );
  inv_x4_sg U44460 ( .A(n43449), .X(n43450) );
  nor_x2_sg U44461 ( .A(n17236), .B(n17235), .X(n17273) );
  nor_x4_sg U44462 ( .A(n43450), .B(n53611), .X(n17236) );
  inv_x4_sg U44463 ( .A(n17276), .X(n53611) );
  nand_x2_sg U44464 ( .A(n17234), .B(n17277), .X(n17276) );
  inv_x4_sg U44465 ( .A(n43451), .X(n43452) );
  nor_x2_sg U44466 ( .A(n15670), .B(n15669), .X(n15707) );
  nor_x4_sg U44467 ( .A(n43452), .B(n53053), .X(n15670) );
  inv_x4_sg U44468 ( .A(n15710), .X(n53053) );
  nand_x2_sg U44469 ( .A(n15668), .B(n15711), .X(n15710) );
  inv_x4_sg U44470 ( .A(n43453), .X(n43454) );
  nor_x2_sg U44471 ( .A(n14117), .B(n14116), .X(n14154) );
  nor_x4_sg U44472 ( .A(n43454), .B(n52496), .X(n14117) );
  inv_x4_sg U44473 ( .A(n14157), .X(n52496) );
  nand_x2_sg U44474 ( .A(n14115), .B(n14158), .X(n14157) );
  inv_x4_sg U44475 ( .A(n43455), .X(n43456) );
  nor_x2_sg U44476 ( .A(n13337), .B(n13336), .X(n13374) );
  nor_x4_sg U44477 ( .A(n43456), .B(n52219), .X(n13337) );
  inv_x4_sg U44478 ( .A(n13377), .X(n52219) );
  nand_x2_sg U44479 ( .A(n13335), .B(n13378), .X(n13377) );
  inv_x4_sg U44480 ( .A(n43457), .X(n43458) );
  nor_x2_sg U44481 ( .A(n12556), .B(n12555), .X(n12592) );
  nor_x4_sg U44482 ( .A(n43458), .B(n51944), .X(n12556) );
  inv_x4_sg U44483 ( .A(n12595), .X(n51944) );
  nand_x2_sg U44484 ( .A(n12554), .B(n12596), .X(n12595) );
  inv_x4_sg U44485 ( .A(n43459), .X(n43460) );
  nor_x2_sg U44486 ( .A(n21107), .B(n21106), .X(n21139) );
  nor_x4_sg U44487 ( .A(n43460), .B(n55022), .X(n21107) );
  inv_x4_sg U44488 ( .A(n21142), .X(n55022) );
  nand_x2_sg U44489 ( .A(n21105), .B(n21143), .X(n21142) );
  inv_x4_sg U44490 ( .A(n43461), .X(n43462) );
  nor_x2_sg U44491 ( .A(n19563), .B(n19562), .X(n19595) );
  nor_x4_sg U44492 ( .A(n43462), .B(n54454), .X(n19563) );
  inv_x4_sg U44493 ( .A(n19598), .X(n54454) );
  nand_x2_sg U44494 ( .A(n19561), .B(n19599), .X(n19598) );
  inv_x4_sg U44495 ( .A(n43463), .X(n43464) );
  nor_x2_sg U44496 ( .A(n18018), .B(n18017), .X(n18050) );
  nor_x4_sg U44497 ( .A(n43464), .B(n53889), .X(n18018) );
  inv_x4_sg U44498 ( .A(n18053), .X(n53889) );
  nand_x2_sg U44499 ( .A(n18016), .B(n18054), .X(n18053) );
  inv_x4_sg U44500 ( .A(n43465), .X(n43466) );
  nor_x2_sg U44501 ( .A(n14897), .B(n14896), .X(n14929) );
  nor_x4_sg U44502 ( .A(n43466), .B(n52769), .X(n14897) );
  inv_x4_sg U44503 ( .A(n14932), .X(n52769) );
  nand_x2_sg U44504 ( .A(n14895), .B(n14933), .X(n14932) );
  inv_x4_sg U44505 ( .A(n43467), .X(n43468) );
  nor_x2_sg U44506 ( .A(n11784), .B(n11783), .X(n11817) );
  nor_x4_sg U44507 ( .A(n43468), .B(n51663), .X(n11784) );
  inv_x4_sg U44508 ( .A(n11820), .X(n51663) );
  nand_x2_sg U44509 ( .A(n11782), .B(n11821), .X(n11820) );
  inv_x4_sg U44510 ( .A(n43469), .X(n43470) );
  nor_x4_sg U44511 ( .A(n43470), .B(n51986), .X(n12311) );
  inv_x4_sg U44512 ( .A(n12367), .X(n51986) );
  nand_x2_sg U44513 ( .A(n12368), .B(n51893), .X(n12367) );
  inv_x4_sg U44514 ( .A(n18489), .X(n43471) );
  inv_x4_sg U44515 ( .A(n43471), .X(n43472) );
  nor_x4_sg U44516 ( .A(n18487), .B(n54097), .X(n18485) );
  inv_x4_sg U44517 ( .A(n43473), .X(n43474) );
  nor_x2_sg U44518 ( .A(n46377), .B(n16946), .X(n17020) );
  nor_x4_sg U44519 ( .A(n43474), .B(n53642), .X(n16946) );
  inv_x4_sg U44520 ( .A(n17022), .X(n53642) );
  nand_x2_sg U44521 ( .A(n17019), .B(n17023), .X(n17022) );
  inv_x4_sg U44522 ( .A(n43475), .X(n43476) );
  nor_x2_sg U44523 ( .A(n46421), .B(n15380), .X(n15454) );
  nor_x4_sg U44524 ( .A(n43476), .B(n53084), .X(n15380) );
  inv_x4_sg U44525 ( .A(n15456), .X(n53084) );
  nand_x2_sg U44526 ( .A(n15453), .B(n15457), .X(n15456) );
  inv_x4_sg U44527 ( .A(n43477), .X(n43478) );
  nor_x2_sg U44528 ( .A(n46469), .B(n13827), .X(n13901) );
  nor_x4_sg U44529 ( .A(n43478), .B(n52526), .X(n13827) );
  inv_x4_sg U44530 ( .A(n13903), .X(n52526) );
  nand_x2_sg U44531 ( .A(n13900), .B(n13904), .X(n13903) );
  inv_x4_sg U44532 ( .A(n43479), .X(n43480) );
  nor_x2_sg U44533 ( .A(n46489), .B(n13047), .X(n13121) );
  nor_x4_sg U44534 ( .A(n43480), .B(n52250), .X(n13047) );
  inv_x4_sg U44535 ( .A(n13123), .X(n52250) );
  nand_x2_sg U44536 ( .A(n13120), .B(n13124), .X(n13123) );
  inv_x4_sg U44537 ( .A(n43481), .X(n43482) );
  nor_x2_sg U44538 ( .A(n46533), .B(n11486), .X(n11560) );
  nor_x4_sg U44539 ( .A(n43482), .B(n51694), .X(n11486) );
  inv_x4_sg U44540 ( .A(n11562), .X(n51694) );
  nand_x2_sg U44541 ( .A(n11559), .B(n11563), .X(n11562) );
  inv_x4_sg U44542 ( .A(n43483), .X(n43484) );
  nor_x2_sg U44543 ( .A(n10551), .B(n10552), .X(n10549) );
  nor_x4_sg U44544 ( .A(n43484), .B(n51357), .X(n10551) );
  inv_x4_sg U44545 ( .A(n10612), .X(n51357) );
  nand_x2_sg U44546 ( .A(n10613), .B(n10614), .X(n10612) );
  inv_x4_sg U44547 ( .A(n43485), .X(n43486) );
  nor_x2_sg U44548 ( .A(n18333), .B(n18334), .X(n18331) );
  nor_x4_sg U44549 ( .A(n43486), .B(n54146), .X(n18333) );
  inv_x4_sg U44550 ( .A(n18394), .X(n54146) );
  nand_x2_sg U44551 ( .A(n18395), .B(n18396), .X(n18394) );
  inv_x4_sg U44552 ( .A(n43487), .X(n43488) );
  inv_x4_sg U44553 ( .A(n43489), .X(n43490) );
  nor_x4_sg U44554 ( .A(n43490), .B(n43488), .X(n21305) );
  inv_x4_sg U44555 ( .A(n43491), .X(n43492) );
  inv_x4_sg U44556 ( .A(n43493), .X(n43494) );
  nor_x4_sg U44557 ( .A(n43494), .B(n43492), .X(n19760) );
  inv_x4_sg U44558 ( .A(n43495), .X(n43496) );
  nor_x4_sg U44559 ( .A(n13553), .B(n43496), .X(n13546) );
  nor_x4_sg U44560 ( .A(n13556), .B(n13555), .X(n13553) );
  inv_x4_sg U44561 ( .A(n43497), .X(n43498) );
  inv_x4_sg U44562 ( .A(n43499), .X(n43500) );
  nor_x4_sg U44563 ( .A(n43500), .B(n43498), .X(n20537) );
  inv_x4_sg U44564 ( .A(n43501), .X(n43502) );
  inv_x4_sg U44565 ( .A(n43503), .X(n43504) );
  nor_x4_sg U44566 ( .A(n43504), .B(n43502), .X(n18993) );
  inv_x4_sg U44567 ( .A(n43505), .X(n43506) );
  inv_x4_sg U44568 ( .A(n43507), .X(n43508) );
  nor_x4_sg U44569 ( .A(n43508), .B(n43506), .X(n17448) );
  inv_x4_sg U44570 ( .A(n43509), .X(n43510) );
  inv_x4_sg U44571 ( .A(n43511), .X(n43512) );
  nor_x4_sg U44572 ( .A(n43512), .B(n43510), .X(n14325) );
  inv_x4_sg U44573 ( .A(n43513), .X(n43514) );
  nand_x4_sg U44574 ( .A(n43514), .B(n18235), .X(n18233) );
  nor_x2_sg U44575 ( .A(n18235), .B(n18236), .X(n18234) );
  nor_x4_sg U44576 ( .A(n41732), .B(n18223), .X(n18236) );
  inv_x4_sg U44577 ( .A(n43515), .X(n43516) );
  nor_x2_sg U44578 ( .A(n29606), .B(n46603), .X(n29605) );
  nor_x4_sg U44579 ( .A(n50106), .B(n43516), .X(n29606) );
  inv_x4_sg U44580 ( .A(n29642), .X(n50106) );
  nand_x2_sg U44581 ( .A(n29641), .B(n29602), .X(n29642) );
  inv_x4_sg U44582 ( .A(n43517), .X(n43518) );
  nor_x2_sg U44583 ( .A(n29618), .B(n9394), .X(n29613) );
  nor_x4_sg U44584 ( .A(n50102), .B(n43518), .X(n29618) );
  inv_x4_sg U44585 ( .A(n30172), .X(n50102) );
  nand_x2_sg U44586 ( .A(n30171), .B(n29611), .X(n30172) );
  inv_x4_sg U44587 ( .A(n43519), .X(n43520) );
  nor_x2_sg U44588 ( .A(n21951), .B(n46603), .X(n21950) );
  nor_x4_sg U44589 ( .A(n50965), .B(n43520), .X(n21951) );
  inv_x4_sg U44590 ( .A(n21977), .X(n50965) );
  nand_x2_sg U44591 ( .A(n21976), .B(n21948), .X(n21977) );
  inv_x4_sg U44592 ( .A(n43521), .X(n43522) );
  nor_x2_sg U44593 ( .A(n21959), .B(n9394), .X(n21956) );
  nor_x4_sg U44594 ( .A(n50961), .B(n43522), .X(n21959) );
  inv_x4_sg U44595 ( .A(n22506), .X(n50961) );
  nand_x2_sg U44596 ( .A(n22505), .B(n21955), .X(n22506) );
  nor_x2_sg U44597 ( .A(n40721), .B(out_L2[3]), .X(n24418) );
  nor_x4_sg U44598 ( .A(n17186), .B(n53637), .X(n17112) );
  inv_x4_sg U44599 ( .A(n17187), .X(n53637) );
  nor_x4_sg U44600 ( .A(n53616), .B(n17188), .X(n17186) );
  nor_x8_sg U44601 ( .A(n16975), .B(n53509), .X(n17188) );
  nand_x2_sg U44602 ( .A(n17188), .B(n53616), .X(n17187) );
  nor_x2_sg U44603 ( .A(n53359), .B(n16287), .X(n16462) );
  nor_x4_sg U44604 ( .A(n16466), .B(n53331), .X(n16287) );
  inv_x4_sg U44605 ( .A(n16467), .X(n53331) );
  nand_x2_sg U44606 ( .A(n53311), .B(n16464), .X(n16467) );
  nor_x4_sg U44607 ( .A(n16464), .B(n53311), .X(n16466) );
  nand_x8_sg U44608 ( .A(n46405), .B(n53319), .X(n16464) );
  nor_x4_sg U44609 ( .A(n15620), .B(n53079), .X(n15546) );
  inv_x4_sg U44610 ( .A(n15621), .X(n53079) );
  nor_x4_sg U44611 ( .A(n53058), .B(n15622), .X(n15620) );
  nor_x8_sg U44612 ( .A(n15409), .B(n52951), .X(n15622) );
  nand_x2_sg U44613 ( .A(n15622), .B(n53058), .X(n15621) );
  nor_x4_sg U44614 ( .A(n14067), .B(n52521), .X(n13993) );
  inv_x4_sg U44615 ( .A(n14068), .X(n52521) );
  nor_x4_sg U44616 ( .A(n52501), .B(n14069), .X(n14067) );
  nor_x8_sg U44617 ( .A(n13856), .B(n46473), .X(n14069) );
  nand_x2_sg U44618 ( .A(n14069), .B(n52501), .X(n14068) );
  nor_x4_sg U44619 ( .A(n13287), .B(n52245), .X(n13213) );
  inv_x4_sg U44620 ( .A(n13288), .X(n52245) );
  nor_x4_sg U44621 ( .A(n52224), .B(n13289), .X(n13287) );
  nor_x8_sg U44622 ( .A(n13076), .B(n52117), .X(n13289) );
  nand_x2_sg U44623 ( .A(n13289), .B(n52224), .X(n13288) );
  nor_x4_sg U44624 ( .A(n12506), .B(n51970), .X(n12432) );
  inv_x4_sg U44625 ( .A(n12507), .X(n51970) );
  nor_x4_sg U44626 ( .A(n51949), .B(n12508), .X(n12506) );
  nor_x8_sg U44627 ( .A(n12295), .B(n46516), .X(n12508) );
  nand_x2_sg U44628 ( .A(n12508), .B(n51949), .X(n12507) );
  nor_x2_sg U44629 ( .A(n40722), .B(out_L1[3]), .X(n32084) );
  inv_x4_sg U44630 ( .A(n43523), .X(n43524) );
  inv_x4_sg U44631 ( .A(n43525), .X(n43526) );
  nor_x4_sg U44632 ( .A(n43526), .B(n43524), .X(n21701) );
  nor_x4_sg U44633 ( .A(n21048), .B(n55048), .X(n20974) );
  inv_x4_sg U44634 ( .A(n21049), .X(n55048) );
  nor_x4_sg U44635 ( .A(n55033), .B(n21050), .X(n21048) );
  nor_x8_sg U44636 ( .A(n20837), .B(n54921), .X(n21050) );
  nand_x2_sg U44637 ( .A(n21050), .B(n55033), .X(n21049) );
  inv_x4_sg U44638 ( .A(n43527), .X(n43528) );
  inv_x4_sg U44639 ( .A(n43529), .X(n43530) );
  nor_x4_sg U44640 ( .A(n43530), .B(n43528), .X(n20156) );
  nor_x4_sg U44641 ( .A(n19504), .B(n54480), .X(n19430) );
  inv_x4_sg U44642 ( .A(n19505), .X(n54480) );
  nor_x4_sg U44643 ( .A(n54465), .B(n19506), .X(n19504) );
  nor_x8_sg U44644 ( .A(n19293), .B(n54353), .X(n19506) );
  nand_x2_sg U44645 ( .A(n19506), .B(n54465), .X(n19505) );
  inv_x4_sg U44646 ( .A(n43531), .X(n43532) );
  inv_x4_sg U44647 ( .A(n43533), .X(n43534) );
  nor_x4_sg U44648 ( .A(n43534), .B(n43532), .X(n18610) );
  nor_x4_sg U44649 ( .A(n17959), .B(n53915), .X(n17885) );
  inv_x4_sg U44650 ( .A(n17960), .X(n53915) );
  nor_x4_sg U44651 ( .A(n53900), .B(n17961), .X(n17959) );
  nor_x8_sg U44652 ( .A(n17748), .B(n53788), .X(n17961) );
  nand_x2_sg U44653 ( .A(n17961), .B(n53900), .X(n17960) );
  nor_x4_sg U44654 ( .A(n16401), .B(n53352), .X(n16327) );
  inv_x4_sg U44655 ( .A(n16402), .X(n53352) );
  nor_x4_sg U44656 ( .A(n53337), .B(n16403), .X(n16401) );
  nor_x8_sg U44657 ( .A(n16190), .B(n46404), .X(n16403) );
  nand_x2_sg U44658 ( .A(n16403), .B(n53337), .X(n16402) );
  nor_x4_sg U44659 ( .A(n14838), .B(n52802), .X(n14764) );
  inv_x4_sg U44660 ( .A(n14839), .X(n52802) );
  nor_x4_sg U44661 ( .A(n52780), .B(n14840), .X(n14838) );
  nor_x8_sg U44662 ( .A(n14627), .B(n46449), .X(n14840) );
  nand_x2_sg U44663 ( .A(n14840), .B(n52780), .X(n14839) );
  nor_x4_sg U44664 ( .A(n11726), .B(n51683), .X(n11652) );
  inv_x4_sg U44665 ( .A(n11727), .X(n51683) );
  nor_x4_sg U44666 ( .A(n51668), .B(n11728), .X(n11726) );
  nor_x8_sg U44667 ( .A(n11515), .B(n51560), .X(n11728) );
  nand_x2_sg U44668 ( .A(n11728), .B(n51668), .X(n11727) );
  nor_x4_sg U44669 ( .A(n10943), .B(n51407), .X(n10872) );
  inv_x4_sg U44670 ( .A(n10944), .X(n51407) );
  nor_x4_sg U44671 ( .A(n51391), .B(n10945), .X(n10943) );
  nor_x8_sg U44672 ( .A(n46563), .B(n46555), .X(n10945) );
  nand_x2_sg U44673 ( .A(n10945), .B(n51391), .X(n10944) );
  nor_x4_sg U44674 ( .A(n21819), .B(n55334), .X(n21744) );
  inv_x4_sg U44675 ( .A(n21820), .X(n55334) );
  nor_x4_sg U44676 ( .A(n55315), .B(n21821), .X(n21819) );
  nor_x8_sg U44677 ( .A(n21774), .B(n46248), .X(n21821) );
  nand_x2_sg U44678 ( .A(n21821), .B(n55315), .X(n21820) );
  nor_x4_sg U44679 ( .A(n20274), .B(n54766), .X(n20199) );
  inv_x4_sg U44680 ( .A(n20275), .X(n54766) );
  nor_x4_sg U44681 ( .A(n54747), .B(n20276), .X(n20274) );
  nor_x8_sg U44682 ( .A(n20229), .B(n46293), .X(n20276) );
  nand_x2_sg U44683 ( .A(n20276), .B(n54747), .X(n20275) );
  nor_x4_sg U44684 ( .A(n18728), .B(n54206), .X(n18653) );
  inv_x4_sg U44685 ( .A(n18729), .X(n54206) );
  nor_x4_sg U44686 ( .A(n54180), .B(n18730), .X(n18728) );
  nor_x8_sg U44687 ( .A(n18574), .B(n46337), .X(n18730) );
  nand_x2_sg U44688 ( .A(n18730), .B(n54180), .X(n18729) );
  nor_x2_sg U44689 ( .A(n53638), .B(n17071), .X(n17239) );
  nor_x4_sg U44690 ( .A(n17243), .B(n53610), .X(n17071) );
  inv_x4_sg U44691 ( .A(n17244), .X(n53610) );
  nand_x2_sg U44692 ( .A(n53591), .B(n17241), .X(n17244) );
  nor_x4_sg U44693 ( .A(n17241), .B(n53591), .X(n17243) );
  nand_x8_sg U44694 ( .A(n53598), .B(n46384), .X(n17241) );
  nor_x2_sg U44695 ( .A(n53080), .B(n15505), .X(n15673) );
  nor_x4_sg U44696 ( .A(n15677), .B(n53052), .X(n15505) );
  inv_x4_sg U44697 ( .A(n15678), .X(n53052) );
  nand_x2_sg U44698 ( .A(n53033), .B(n15675), .X(n15678) );
  nor_x4_sg U44699 ( .A(n15675), .B(n53033), .X(n15677) );
  nand_x8_sg U44700 ( .A(n53040), .B(n46428), .X(n15675) );
  nor_x2_sg U44701 ( .A(n52522), .B(n13952), .X(n14120) );
  nor_x4_sg U44702 ( .A(n14124), .B(n52495), .X(n13952) );
  inv_x4_sg U44703 ( .A(n14125), .X(n52495) );
  nand_x2_sg U44704 ( .A(n52476), .B(n14122), .X(n14125) );
  nor_x4_sg U44705 ( .A(n14122), .B(n52476), .X(n14124) );
  nand_x8_sg U44706 ( .A(n52483), .B(n46474), .X(n14122) );
  nor_x2_sg U44707 ( .A(n52246), .B(n13172), .X(n13340) );
  nor_x4_sg U44708 ( .A(n13344), .B(n52218), .X(n13172) );
  inv_x4_sg U44709 ( .A(n13345), .X(n52218) );
  nand_x2_sg U44710 ( .A(n52199), .B(n13342), .X(n13345) );
  nor_x4_sg U44711 ( .A(n13342), .B(n52199), .X(n13344) );
  nand_x8_sg U44712 ( .A(n52206), .B(n46496), .X(n13342) );
  nor_x2_sg U44713 ( .A(n51971), .B(n12392), .X(n12558) );
  nor_x4_sg U44714 ( .A(n12562), .B(n51943), .X(n12392) );
  inv_x4_sg U44715 ( .A(n12563), .X(n51943) );
  nand_x2_sg U44716 ( .A(n51923), .B(n12560), .X(n12563) );
  nor_x4_sg U44717 ( .A(n12560), .B(n51923), .X(n12562) );
  nand_x8_sg U44718 ( .A(n51931), .B(n46517), .X(n12560) );
  nor_x2_sg U44719 ( .A(n51690), .B(n11611), .X(n11788) );
  nor_x4_sg U44720 ( .A(n11792), .B(n51662), .X(n11611) );
  inv_x4_sg U44721 ( .A(n11793), .X(n51662) );
  nand_x2_sg U44722 ( .A(n51643), .B(n11790), .X(n11793) );
  nor_x4_sg U44723 ( .A(n11790), .B(n51643), .X(n11792) );
  nand_x8_sg U44724 ( .A(n51650), .B(n46540), .X(n11790) );
  inv_x4_sg U44725 ( .A(n43535), .X(n43536) );
  nor_x4_sg U44726 ( .A(n43536), .B(n53672), .X(n17228) );
  inv_x4_sg U44727 ( .A(n17260), .X(n53672) );
  nand_x2_sg U44728 ( .A(n17230), .B(n17261), .X(n17260) );
  inv_x4_sg U44729 ( .A(n43537), .X(n43538) );
  nor_x4_sg U44730 ( .A(n43538), .B(n53114), .X(n15662) );
  inv_x4_sg U44731 ( .A(n15694), .X(n53114) );
  nand_x2_sg U44732 ( .A(n15664), .B(n15695), .X(n15694) );
  inv_x4_sg U44733 ( .A(n43539), .X(n43540) );
  nor_x4_sg U44734 ( .A(n43540), .B(n52555), .X(n14109) );
  inv_x4_sg U44735 ( .A(n14141), .X(n52555) );
  nand_x2_sg U44736 ( .A(n14111), .B(n14142), .X(n14141) );
  inv_x4_sg U44737 ( .A(n43541), .X(n43542) );
  nor_x4_sg U44738 ( .A(n43542), .B(n52280), .X(n13329) );
  inv_x4_sg U44739 ( .A(n13361), .X(n52280) );
  nand_x2_sg U44740 ( .A(n13331), .B(n13362), .X(n13361) );
  inv_x4_sg U44741 ( .A(n43543), .X(n43544) );
  nor_x4_sg U44742 ( .A(n43544), .B(n52009), .X(n12548) );
  inv_x4_sg U44743 ( .A(n12579), .X(n52009) );
  nand_x2_sg U44744 ( .A(n12550), .B(n12580), .X(n12579) );
  nor_x2_sg U44745 ( .A(n55056), .B(n20933), .X(n21109) );
  nor_x4_sg U44746 ( .A(n21113), .B(n55021), .X(n20933) );
  inv_x4_sg U44747 ( .A(n21114), .X(n55021) );
  nand_x2_sg U44748 ( .A(n55001), .B(n21111), .X(n21114) );
  nor_x4_sg U44749 ( .A(n21111), .B(n55001), .X(n21113) );
  nand_x8_sg U44750 ( .A(n55016), .B(n46269), .X(n21111) );
  nor_x2_sg U44751 ( .A(n54488), .B(n19389), .X(n19565) );
  nor_x4_sg U44752 ( .A(n19569), .B(n54453), .X(n19389) );
  inv_x4_sg U44753 ( .A(n19570), .X(n54453) );
  nand_x2_sg U44754 ( .A(n54433), .B(n19567), .X(n19570) );
  nor_x4_sg U44755 ( .A(n19567), .B(n54433), .X(n19569) );
  nand_x8_sg U44756 ( .A(n54448), .B(n46314), .X(n19567) );
  nor_x2_sg U44757 ( .A(n53923), .B(n17844), .X(n18020) );
  nor_x4_sg U44758 ( .A(n18024), .B(n53888), .X(n17844) );
  inv_x4_sg U44759 ( .A(n18025), .X(n53888) );
  nand_x2_sg U44760 ( .A(n53868), .B(n18022), .X(n18025) );
  nor_x4_sg U44761 ( .A(n18022), .B(n53868), .X(n18024) );
  nand_x8_sg U44762 ( .A(n53883), .B(n46361), .X(n18022) );
  nor_x2_sg U44763 ( .A(n52803), .B(n14723), .X(n14899) );
  nor_x4_sg U44764 ( .A(n14903), .B(n52768), .X(n14723) );
  inv_x4_sg U44765 ( .A(n14904), .X(n52768) );
  nand_x2_sg U44766 ( .A(n52748), .B(n14901), .X(n14904) );
  nor_x4_sg U44767 ( .A(n14901), .B(n52748), .X(n14903) );
  nand_x8_sg U44768 ( .A(n52763), .B(n46450), .X(n14901) );
  nor_x4_sg U44769 ( .A(n16021), .B(n53247), .X(n15975) );
  nor_x4_sg U44770 ( .A(n16019), .B(n53233), .X(n16021) );
  inv_x4_sg U44771 ( .A(n16022), .X(n53247) );
  nand_x2_sg U44772 ( .A(n53233), .B(n16019), .X(n16022) );
  nor_x4_sg U44773 ( .A(n16806), .B(n53530), .X(n16760) );
  nor_x4_sg U44774 ( .A(n16804), .B(n53517), .X(n16806) );
  inv_x4_sg U44775 ( .A(n16807), .X(n53530) );
  nand_x2_sg U44776 ( .A(n53517), .B(n16804), .X(n16807) );
  nor_x4_sg U44777 ( .A(n15240), .B(n52972), .X(n15194) );
  nor_x4_sg U44778 ( .A(n15238), .B(n52959), .X(n15240) );
  inv_x4_sg U44779 ( .A(n15241), .X(n52972) );
  nand_x2_sg U44780 ( .A(n52959), .B(n15238), .X(n15241) );
  nor_x4_sg U44781 ( .A(n13687), .B(n52413), .X(n13641) );
  nor_x4_sg U44782 ( .A(n13685), .B(n52399), .X(n13687) );
  inv_x4_sg U44783 ( .A(n13688), .X(n52413) );
  nand_x2_sg U44784 ( .A(n52399), .B(n13685), .X(n13688) );
  nor_x4_sg U44785 ( .A(n12907), .B(n52138), .X(n12861) );
  nor_x4_sg U44786 ( .A(n12905), .B(n52125), .X(n12907) );
  inv_x4_sg U44787 ( .A(n12908), .X(n52138) );
  nand_x2_sg U44788 ( .A(n52125), .B(n12905), .X(n12908) );
  nor_x4_sg U44789 ( .A(n12126), .B(n51861), .X(n12080) );
  nor_x4_sg U44790 ( .A(n12124), .B(n51847), .X(n12126) );
  inv_x4_sg U44791 ( .A(n12127), .X(n51861) );
  nand_x2_sg U44792 ( .A(n51847), .B(n12124), .X(n12127) );
  nor_x4_sg U44793 ( .A(n11346), .B(n51580), .X(n11300) );
  nor_x4_sg U44794 ( .A(n11344), .B(n51568), .X(n11346) );
  inv_x4_sg U44795 ( .A(n11347), .X(n51580) );
  nand_x2_sg U44796 ( .A(n51568), .B(n11344), .X(n11347) );
  nor_x4_sg U44797 ( .A(n41278), .B(n20383), .X(n20490) );
  nor_x4_sg U44798 ( .A(n41279), .B(n18839), .X(n18946) );
  nor_x4_sg U44799 ( .A(n41280), .B(n17294), .X(n17401) );
  nor_x4_sg U44800 ( .A(n25382), .B(n8362), .X(n31254) );
  nor_x4_sg U44801 ( .A(n25378), .B(n8422), .X(n31741) );
  nor_x4_sg U44802 ( .A(n10272), .B(n8722), .X(n24075) );
  nor_x4_sg U44803 ( .A(n10276), .B(n8662), .X(n23588) );
  nor_x4_sg U44804 ( .A(n40725), .B(n8482), .X(n32070) );
  nor_x4_sg U44805 ( .A(n25379), .B(n8462), .X(n31982) );
  nor_x4_sg U44806 ( .A(n40726), .B(n8782), .X(n24404) );
  nor_x4_sg U44807 ( .A(n10273), .B(n8762), .X(n24316) );
  inv_x4_sg U44808 ( .A(n43545), .X(n43546) );
  nor_x4_sg U44809 ( .A(n50096), .B(n43546), .X(n29588) );
  inv_x4_sg U44810 ( .A(n30190), .X(n50096) );
  nand_x2_sg U44811 ( .A(n30189), .B(n29625), .X(n30190) );
  inv_x4_sg U44812 ( .A(n43547), .X(n43548) );
  nor_x4_sg U44813 ( .A(n50955), .B(n43548), .X(n21937) );
  inv_x4_sg U44814 ( .A(n22524), .X(n50955) );
  nand_x2_sg U44815 ( .A(n22523), .B(n21964), .X(n22524) );
  nor_x4_sg U44816 ( .A(n27424), .B(n53363), .X(n27431) );
  inv_x8_sg U44817 ( .A(n16239), .X(n53363) );
  nor_x4_sg U44818 ( .A(n26027), .B(n51974), .X(n26034) );
  inv_x8_sg U44819 ( .A(n12344), .X(n51974) );
  nor_x4_sg U44820 ( .A(n25749), .B(n51693), .X(n25756) );
  inv_x4_sg U44821 ( .A(n43549), .X(n43550) );
  inv_x4_sg U44822 ( .A(n43551), .X(n43552) );
  nor_x4_sg U44823 ( .A(n43552), .B(n43550), .X(n11776) );
  nor_x8_sg U44824 ( .A(n29433), .B(n55403), .X(n29420) );
  inv_x8_sg U44825 ( .A(n29404), .X(n55403) );
  nor_x8_sg U44826 ( .A(n29153), .B(n55118), .X(n29138) );
  inv_x8_sg U44827 ( .A(n29122), .X(n55118) );
  nor_x8_sg U44828 ( .A(n28872), .B(n54835), .X(n28859) );
  inv_x8_sg U44829 ( .A(n28843), .X(n54835) );
  nor_x8_sg U44830 ( .A(n28592), .B(n54550), .X(n28579) );
  inv_x8_sg U44831 ( .A(n28563), .X(n54550) );
  nor_x8_sg U44832 ( .A(n28315), .B(n54268), .X(n28301) );
  inv_x8_sg U44833 ( .A(n28285), .X(n54268) );
  nor_x8_sg U44834 ( .A(n28034), .B(n53985), .X(n28021) );
  inv_x8_sg U44835 ( .A(n28005), .X(n53985) );
  nor_x8_sg U44836 ( .A(n27755), .B(n53707), .X(n27742) );
  inv_x8_sg U44837 ( .A(n42475), .X(n53707) );
  nor_x8_sg U44838 ( .A(n27474), .B(n53425), .X(n27461) );
  inv_x8_sg U44839 ( .A(n42477), .X(n53425) );
  nor_x8_sg U44840 ( .A(n27197), .B(n53149), .X(n27182) );
  inv_x8_sg U44841 ( .A(n42479), .X(n53149) );
  nor_x8_sg U44842 ( .A(n26915), .B(n52865), .X(n26902) );
  inv_x8_sg U44843 ( .A(n26886), .X(n52865) );
  nor_x8_sg U44844 ( .A(n26638), .B(n52590), .X(n26625) );
  inv_x8_sg U44845 ( .A(n42481), .X(n52590) );
  nor_x8_sg U44846 ( .A(n26360), .B(n52315), .X(n26346) );
  inv_x8_sg U44847 ( .A(n42483), .X(n52315) );
  nor_x8_sg U44848 ( .A(n26081), .B(n52039), .X(n26065) );
  inv_x8_sg U44849 ( .A(n42485), .X(n52039) );
  nor_x8_sg U44850 ( .A(n25799), .B(n51756), .X(n25786) );
  inv_x8_sg U44851 ( .A(n42487), .X(n51756) );
  nor_x8_sg U44852 ( .A(n25520), .B(n51474), .X(n25508) );
  inv_x8_sg U44853 ( .A(n42489), .X(n51474) );
  nand_x4_sg U44854 ( .A(n10580), .B(n10579), .X(n10607) );
  nor_x8_sg U44855 ( .A(n10655), .B(n46566), .X(n10579) );
  nand_x4_sg U44856 ( .A(n21452), .B(n21451), .X(n21479) );
  nor_x8_sg U44857 ( .A(n21527), .B(n46255), .X(n21451) );
  nand_x4_sg U44858 ( .A(n19907), .B(n19906), .X(n19934) );
  nor_x8_sg U44859 ( .A(n19982), .B(n46300), .X(n19906) );
  nand_x4_sg U44860 ( .A(n18362), .B(n18361), .X(n18389) );
  nor_x8_sg U44861 ( .A(n18437), .B(n46341), .X(n18361) );
  nand_x4_sg U44862 ( .A(n20681), .B(n20680), .X(n20709) );
  nor_x8_sg U44863 ( .A(n20757), .B(n46275), .X(n20680) );
  nand_x4_sg U44864 ( .A(n19137), .B(n19136), .X(n19165) );
  nor_x8_sg U44865 ( .A(n19213), .B(n46320), .X(n19136) );
  nand_x4_sg U44866 ( .A(n17592), .B(n17591), .X(n17620) );
  nor_x8_sg U44867 ( .A(n17668), .B(n46367), .X(n17591) );
  nand_x4_sg U44868 ( .A(n14472), .B(n14471), .X(n14499) );
  nor_x8_sg U44869 ( .A(n14547), .B(n46452), .X(n14471) );
  nand_x4_sg U44870 ( .A(n10579), .B(n10696), .X(n10619) );
  nor_x8_sg U44871 ( .A(n51354), .B(n46570), .X(n10696) );
  nand_x4_sg U44872 ( .A(n21451), .B(n21568), .X(n21491) );
  nor_x8_sg U44873 ( .A(n55276), .B(n46254), .X(n21568) );
  nand_x4_sg U44874 ( .A(n19906), .B(n20023), .X(n19946) );
  nor_x8_sg U44875 ( .A(n54708), .B(n46299), .X(n20023) );
  nor_x4_sg U44876 ( .A(n18514), .B(n18478), .X(n18515) );
  nand_x4_sg U44877 ( .A(n18361), .B(n18478), .X(n18401) );
  nor_x8_sg U44878 ( .A(n54143), .B(n46346), .X(n18478) );
  nand_x4_sg U44879 ( .A(n16029), .B(n16152), .X(n16072) );
  nor_x8_sg U44880 ( .A(n16069), .B(n46411), .X(n16152) );
  nand_x4_sg U44881 ( .A(n11354), .B(n11477), .X(n11397) );
  nor_x8_sg U44882 ( .A(n11394), .B(n46545), .X(n11477) );
  nand_x4_sg U44883 ( .A(n20680), .B(n20798), .X(n20721) );
  nor_x8_sg U44884 ( .A(n20717), .B(n46274), .X(n20798) );
  nand_x4_sg U44885 ( .A(n19136), .B(n19254), .X(n19177) );
  nor_x8_sg U44886 ( .A(n19173), .B(n46319), .X(n19254) );
  nand_x4_sg U44887 ( .A(n17591), .B(n17709), .X(n17632) );
  nor_x8_sg U44888 ( .A(n17628), .B(n46366), .X(n17709) );
  nand_x4_sg U44889 ( .A(n14471), .B(n14588), .X(n14511) );
  nor_x8_sg U44890 ( .A(n14507), .B(n46456), .X(n14588) );
  nor_x8_sg U44891 ( .A(n46387), .B(n46389), .X(n16635) );
  nor_x8_sg U44892 ( .A(n46431), .B(n46433), .X(n15069) );
  nor_x8_sg U44893 ( .A(n46499), .B(n46501), .X(n12736) );
  nor_x8_sg U44894 ( .A(n46543), .B(n46545), .X(n11175) );
  inv_x8_sg U44895 ( .A(n28452), .X(n43559) );
  nor_x8_sg U44896 ( .A(n28451), .B(n43559), .X(n28389) );
  nand_x4_sg U44897 ( .A(n44837), .B(n28453), .X(n28452) );
  nor_x8_sg U44898 ( .A(n28394), .B(n46191), .X(n28451) );
  nor_x4_sg U44899 ( .A(n15890), .B(n15889), .X(n15887) );
  inv_x2_sg U44900 ( .A(n15889), .X(n53234) );
  nor_x8_sg U44901 ( .A(n46404), .B(n46407), .X(n15889) );
  inv_x2_sg U44902 ( .A(n13555), .X(n52400) );
  nor_x8_sg U44903 ( .A(n46473), .B(n46480), .X(n13555) );
  nor_x4_sg U44904 ( .A(n11995), .B(n11994), .X(n11992) );
  inv_x2_sg U44905 ( .A(n11994), .X(n51848) );
  nor_x8_sg U44906 ( .A(n46516), .B(n46519), .X(n11994) );
  nor_x2_sg U44907 ( .A(n40765), .B(n31279), .X(n31278) );
  inv_x2_sg U44908 ( .A(n31279), .X(n49446) );
  nor_x2_sg U44909 ( .A(n40766), .B(n31297), .X(n31296) );
  inv_x2_sg U44910 ( .A(n31297), .X(n49586) );
  nor_x2_sg U44911 ( .A(n40767), .B(n31315), .X(n31314) );
  inv_x2_sg U44912 ( .A(n31315), .X(n49726) );
  nor_x2_sg U44913 ( .A(n40768), .B(n23613), .X(n23612) );
  inv_x2_sg U44914 ( .A(n23613), .X(n50305) );
  nor_x2_sg U44915 ( .A(n40769), .B(n23631), .X(n23630) );
  inv_x2_sg U44916 ( .A(n23631), .X(n50445) );
  nor_x2_sg U44917 ( .A(n40770), .B(n23649), .X(n23648) );
  inv_x2_sg U44918 ( .A(n23649), .X(n50585) );
  nand_x2_sg U44919 ( .A(n16640), .B(n16724), .X(n16723) );
  nand_x4_sg U44920 ( .A(n16640), .B(n53483), .X(n16638) );
  nor_x8_sg U44921 ( .A(n46385), .B(n46387), .X(n16640) );
  nand_x2_sg U44922 ( .A(n15074), .B(n15158), .X(n15157) );
  nand_x4_sg U44923 ( .A(n15074), .B(n52925), .X(n15072) );
  nor_x8_sg U44924 ( .A(n46429), .B(n46431), .X(n15074) );
  nand_x2_sg U44925 ( .A(n12741), .B(n12825), .X(n12824) );
  nand_x4_sg U44926 ( .A(n12741), .B(n52091), .X(n12739) );
  nor_x8_sg U44927 ( .A(n46497), .B(n46499), .X(n12741) );
  nand_x2_sg U44928 ( .A(n11180), .B(n11264), .X(n11263) );
  nand_x4_sg U44929 ( .A(n11180), .B(n51533), .X(n11178) );
  nor_x8_sg U44930 ( .A(n46541), .B(n46543), .X(n11180) );
  nand_x2_sg U44931 ( .A(n20510), .B(n20591), .X(n20590) );
  nor_x8_sg U44932 ( .A(n46270), .B(n46272), .X(n20510) );
  nand_x2_sg U44933 ( .A(n18966), .B(n19047), .X(n19046) );
  nor_x8_sg U44934 ( .A(n46315), .B(n46317), .X(n18966) );
  nand_x2_sg U44935 ( .A(n17421), .B(n17502), .X(n17501) );
  nor_x8_sg U44936 ( .A(n46362), .B(n46364), .X(n17421) );
  nand_x2_sg U44937 ( .A(n24791), .B(n30907), .X(n31014) );
  nor_x2_sg U44938 ( .A(n24791), .B(n9385), .X(n24788) );
  nand_x2_sg U44939 ( .A(n9683), .B(n23241), .X(n23348) );
  nor_x2_sg U44940 ( .A(n9683), .B(n9385), .X(n9680) );
  nand_x2_sg U44941 ( .A(n25272), .B(n25293), .X(n29712) );
  nor_x2_sg U44942 ( .A(n25272), .B(n46603), .X(n25271) );
  nand_x2_sg U44943 ( .A(n25223), .B(n25246), .X(n29709) );
  nor_x2_sg U44944 ( .A(n25223), .B(n46603), .X(n25222) );
  nand_x2_sg U44945 ( .A(n25174), .B(n25197), .X(n29706) );
  nor_x2_sg U44946 ( .A(n25174), .B(n46603), .X(n25173) );
  nand_x2_sg U44947 ( .A(n25126), .B(n25148), .X(n29703) );
  nor_x2_sg U44948 ( .A(n25126), .B(n46603), .X(n25125) );
  nand_x2_sg U44949 ( .A(n25133), .B(n30366), .X(n30572) );
  nand_x2_sg U44950 ( .A(n30364), .B(n25133), .X(n30362) );
  nor_x2_sg U44951 ( .A(n25133), .B(n9394), .X(n25130) );
  nand_x2_sg U44952 ( .A(n25077), .B(n25100), .X(n29700) );
  nor_x2_sg U44953 ( .A(n25077), .B(n46603), .X(n25076) );
  nand_x2_sg U44954 ( .A(n25029), .B(n25051), .X(n29697) );
  nor_x2_sg U44955 ( .A(n25029), .B(n46603), .X(n25028) );
  nand_x2_sg U44956 ( .A(n25036), .B(n30378), .X(n30566) );
  nand_x2_sg U44957 ( .A(n30376), .B(n25036), .X(n30374) );
  nor_x2_sg U44958 ( .A(n25036), .B(n9394), .X(n25033) );
  nand_x2_sg U44959 ( .A(n24981), .B(n25003), .X(n29694) );
  nor_x2_sg U44960 ( .A(n24981), .B(n46603), .X(n24980) );
  nand_x2_sg U44961 ( .A(n24988), .B(n30384), .X(n30563) );
  nand_x2_sg U44962 ( .A(n30382), .B(n24988), .X(n30380) );
  nor_x2_sg U44963 ( .A(n24988), .B(n9394), .X(n24985) );
  nand_x2_sg U44964 ( .A(n24933), .B(n24955), .X(n29691) );
  nor_x2_sg U44965 ( .A(n24933), .B(n46603), .X(n24932) );
  nand_x2_sg U44966 ( .A(n24940), .B(n30390), .X(n30560) );
  nand_x2_sg U44967 ( .A(n30388), .B(n24940), .X(n30386) );
  nor_x2_sg U44968 ( .A(n24940), .B(n9394), .X(n24937) );
  nand_x2_sg U44969 ( .A(n24885), .B(n24907), .X(n29688) );
  nor_x2_sg U44970 ( .A(n24885), .B(n46603), .X(n24884) );
  nand_x2_sg U44971 ( .A(n24892), .B(n30396), .X(n30557) );
  nand_x2_sg U44972 ( .A(n30394), .B(n24892), .X(n30392) );
  nor_x2_sg U44973 ( .A(n24892), .B(n9394), .X(n24889) );
  nand_x2_sg U44974 ( .A(n24837), .B(n24859), .X(n29685) );
  nor_x2_sg U44975 ( .A(n24837), .B(n46603), .X(n24836) );
  nand_x2_sg U44976 ( .A(n24844), .B(n30402), .X(n30554) );
  nand_x2_sg U44977 ( .A(n30400), .B(n24844), .X(n30398) );
  nor_x2_sg U44978 ( .A(n24844), .B(n9394), .X(n24841) );
  nand_x2_sg U44979 ( .A(n24742), .B(n24764), .X(n29679) );
  nor_x2_sg U44980 ( .A(n24742), .B(n46603), .X(n24741) );
  nand_x2_sg U44981 ( .A(n24749), .B(n30414), .X(n30548) );
  nand_x2_sg U44982 ( .A(n30412), .B(n24749), .X(n30410) );
  nor_x2_sg U44983 ( .A(n24749), .B(n9394), .X(n24746) );
  nand_x2_sg U44984 ( .A(n24694), .B(n24716), .X(n29676) );
  nor_x2_sg U44985 ( .A(n24694), .B(n46603), .X(n24693) );
  nand_x2_sg U44986 ( .A(n24701), .B(n30420), .X(n30545) );
  nand_x2_sg U44987 ( .A(n30418), .B(n24701), .X(n30416) );
  nor_x2_sg U44988 ( .A(n24701), .B(n9394), .X(n24698) );
  nand_x2_sg U44989 ( .A(n24645), .B(n24668), .X(n29673) );
  nor_x2_sg U44990 ( .A(n24645), .B(n46603), .X(n24644) );
  nand_x2_sg U44991 ( .A(n24653), .B(n30426), .X(n30542) );
  nand_x2_sg U44992 ( .A(n30424), .B(n24653), .X(n30422) );
  nor_x2_sg U44993 ( .A(n24653), .B(n9394), .X(n24650) );
  nand_x2_sg U44994 ( .A(n24596), .B(n24619), .X(n29670) );
  nor_x2_sg U44995 ( .A(n24596), .B(n46603), .X(n24595) );
  nand_x2_sg U44996 ( .A(n24604), .B(n30432), .X(n30539) );
  nand_x2_sg U44997 ( .A(n30430), .B(n24604), .X(n30428) );
  nor_x2_sg U44998 ( .A(n24604), .B(n9394), .X(n24601) );
  inv_x4_sg U44999 ( .A(n29832), .X(n43617) );
  inv_x8_sg U45000 ( .A(n43617), .X(n43618) );
  nand_x2_sg U45001 ( .A(n24547), .B(n24570), .X(n29667) );
  nor_x2_sg U45002 ( .A(n24547), .B(n46603), .X(n24546) );
  nor_x8_sg U45003 ( .A(n29831), .B(n43618), .X(n24547) );
  nor_x8_sg U45004 ( .A(n44575), .B(n29834), .X(n29831) );
  nand_x2_sg U45005 ( .A(n24555), .B(n30438), .X(n30536) );
  nand_x2_sg U45006 ( .A(n30436), .B(n24555), .X(n30434) );
  nor_x2_sg U45007 ( .A(n24555), .B(n9394), .X(n24552) );
  nor_x2_sg U45008 ( .A(n24498), .B(n46603), .X(n24497) );
  nand_x2_sg U45009 ( .A(n30442), .B(n24506), .X(n30440) );
  nor_x2_sg U45010 ( .A(n24506), .B(n9394), .X(n24503) );
  nand_x2_sg U45011 ( .A(n10164), .B(n10185), .X(n22047) );
  nor_x2_sg U45012 ( .A(n10164), .B(n46603), .X(n10163) );
  nand_x2_sg U45013 ( .A(n10115), .B(n10138), .X(n22044) );
  nor_x2_sg U45014 ( .A(n10115), .B(n46603), .X(n10114) );
  nand_x2_sg U45015 ( .A(n10066), .B(n10089), .X(n22041) );
  nor_x2_sg U45016 ( .A(n10066), .B(n46603), .X(n10065) );
  nand_x2_sg U45017 ( .A(n10018), .B(n10040), .X(n22038) );
  nor_x2_sg U45018 ( .A(n10018), .B(n46603), .X(n10017) );
  nand_x2_sg U45019 ( .A(n10025), .B(n22700), .X(n22906) );
  nand_x2_sg U45020 ( .A(n22698), .B(n10025), .X(n22696) );
  nor_x2_sg U45021 ( .A(n10025), .B(n9394), .X(n10022) );
  nand_x2_sg U45022 ( .A(n9969), .B(n9992), .X(n22035) );
  nor_x2_sg U45023 ( .A(n9969), .B(n46603), .X(n9968) );
  nand_x2_sg U45024 ( .A(n9921), .B(n9943), .X(n22032) );
  nor_x2_sg U45025 ( .A(n9921), .B(n46603), .X(n9920) );
  nand_x2_sg U45026 ( .A(n9928), .B(n22712), .X(n22900) );
  nand_x2_sg U45027 ( .A(n22710), .B(n9928), .X(n22708) );
  nor_x2_sg U45028 ( .A(n9928), .B(n9394), .X(n9925) );
  nand_x2_sg U45029 ( .A(n9873), .B(n9895), .X(n22029) );
  nor_x2_sg U45030 ( .A(n9873), .B(n46603), .X(n9872) );
  nand_x2_sg U45031 ( .A(n9880), .B(n22718), .X(n22897) );
  nand_x2_sg U45032 ( .A(n22716), .B(n9880), .X(n22714) );
  nor_x2_sg U45033 ( .A(n9880), .B(n9394), .X(n9877) );
  nand_x2_sg U45034 ( .A(n9825), .B(n9847), .X(n22026) );
  nor_x2_sg U45035 ( .A(n9825), .B(n46603), .X(n9824) );
  nand_x2_sg U45036 ( .A(n9832), .B(n22724), .X(n22894) );
  nand_x2_sg U45037 ( .A(n22722), .B(n9832), .X(n22720) );
  nor_x2_sg U45038 ( .A(n9832), .B(n9394), .X(n9829) );
  nand_x2_sg U45039 ( .A(n9777), .B(n9799), .X(n22023) );
  nor_x2_sg U45040 ( .A(n9777), .B(n46603), .X(n9776) );
  nand_x2_sg U45041 ( .A(n9784), .B(n22730), .X(n22891) );
  nand_x2_sg U45042 ( .A(n22728), .B(n9784), .X(n22726) );
  nor_x2_sg U45043 ( .A(n9784), .B(n9394), .X(n9781) );
  nand_x2_sg U45044 ( .A(n9729), .B(n9751), .X(n22020) );
  nor_x2_sg U45045 ( .A(n9729), .B(n46603), .X(n9728) );
  nand_x2_sg U45046 ( .A(n9736), .B(n22736), .X(n22888) );
  nand_x2_sg U45047 ( .A(n22734), .B(n9736), .X(n22732) );
  nor_x2_sg U45048 ( .A(n9736), .B(n9394), .X(n9733) );
  nand_x2_sg U45049 ( .A(n9634), .B(n9656), .X(n22014) );
  nor_x2_sg U45050 ( .A(n9634), .B(n46603), .X(n9633) );
  nand_x2_sg U45051 ( .A(n9641), .B(n22748), .X(n22882) );
  nand_x2_sg U45052 ( .A(n22746), .B(n9641), .X(n22744) );
  nor_x2_sg U45053 ( .A(n9641), .B(n9394), .X(n9638) );
  nand_x2_sg U45054 ( .A(n9586), .B(n9608), .X(n22011) );
  nor_x2_sg U45055 ( .A(n9586), .B(n46603), .X(n9585) );
  nand_x2_sg U45056 ( .A(n9593), .B(n22754), .X(n22879) );
  nand_x2_sg U45057 ( .A(n22752), .B(n9593), .X(n22750) );
  nor_x2_sg U45058 ( .A(n9593), .B(n9394), .X(n9590) );
  nand_x2_sg U45059 ( .A(n9537), .B(n9560), .X(n22008) );
  nor_x2_sg U45060 ( .A(n9537), .B(n46603), .X(n9536) );
  nand_x2_sg U45061 ( .A(n9545), .B(n22760), .X(n22876) );
  nand_x2_sg U45062 ( .A(n22758), .B(n9545), .X(n22756) );
  nor_x2_sg U45063 ( .A(n9545), .B(n9394), .X(n9542) );
  nand_x2_sg U45064 ( .A(n9488), .B(n9511), .X(n22005) );
  nor_x2_sg U45065 ( .A(n9488), .B(n46603), .X(n9487) );
  nand_x2_sg U45066 ( .A(n9496), .B(n22766), .X(n22873) );
  nand_x2_sg U45067 ( .A(n22764), .B(n9496), .X(n22762) );
  nor_x2_sg U45068 ( .A(n9496), .B(n9394), .X(n9493) );
  inv_x4_sg U45069 ( .A(n22167), .X(n43671) );
  inv_x8_sg U45070 ( .A(n43671), .X(n43672) );
  nand_x2_sg U45071 ( .A(n9439), .B(n9462), .X(n22002) );
  nor_x2_sg U45072 ( .A(n9439), .B(n46603), .X(n9438) );
  nor_x8_sg U45073 ( .A(n22166), .B(n43672), .X(n9439) );
  nor_x8_sg U45074 ( .A(n44655), .B(n22169), .X(n22166) );
  nand_x2_sg U45075 ( .A(n9447), .B(n22772), .X(n22870) );
  nand_x2_sg U45076 ( .A(n22770), .B(n9447), .X(n22768) );
  nor_x2_sg U45077 ( .A(n9447), .B(n9394), .X(n9444) );
  nor_x2_sg U45078 ( .A(n9383), .B(n46603), .X(n9382) );
  nand_x2_sg U45079 ( .A(n22776), .B(n9393), .X(n22774) );
  nor_x2_sg U45080 ( .A(n9393), .B(n9394), .X(n9389) );
  nand_x2_sg U45081 ( .A(n10155), .B(n24214), .X(n24303) );
  nor_x2_sg U45082 ( .A(n10155), .B(n9373), .X(n10152) );
  nand_x2_sg U45083 ( .A(n10009), .B(n24232), .X(n24294) );
  nor_x2_sg U45084 ( .A(n10009), .B(n9373), .X(n10006) );
  nand_x2_sg U45085 ( .A(n9960), .B(n24238), .X(n24291) );
  nor_x2_sg U45086 ( .A(n9960), .B(n9373), .X(n9957) );
  nand_x2_sg U45087 ( .A(n9912), .B(n24244), .X(n24288) );
  nor_x2_sg U45088 ( .A(n9912), .B(n9373), .X(n9909) );
  nand_x2_sg U45089 ( .A(n9864), .B(n24250), .X(n24285) );
  nor_x2_sg U45090 ( .A(n9864), .B(n9373), .X(n9861) );
  nand_x2_sg U45091 ( .A(n9816), .B(n24256), .X(n24282) );
  nor_x2_sg U45092 ( .A(n9816), .B(n9373), .X(n9813) );
  nand_x2_sg U45093 ( .A(n9768), .B(n24169), .X(n24166) );
  nand_x2_sg U45094 ( .A(n24260), .B(n9768), .X(n24258) );
  nor_x2_sg U45095 ( .A(n9768), .B(n9373), .X(n9765) );
  nand_x2_sg U45096 ( .A(n9720), .B(n24025), .X(n24022) );
  nand_x2_sg U45097 ( .A(n24144), .B(n9720), .X(n24142) );
  nor_x2_sg U45098 ( .A(n9720), .B(n9373), .X(n9717) );
  nand_x2_sg U45099 ( .A(n9673), .B(n23872), .X(n23869) );
  nand_x2_sg U45100 ( .A(n24000), .B(n9673), .X(n23998) );
  nor_x2_sg U45101 ( .A(n9673), .B(n9373), .X(n9670) );
  nand_x2_sg U45102 ( .A(n9625), .B(n23701), .X(n23698) );
  nand_x2_sg U45103 ( .A(n23847), .B(n9625), .X(n23845) );
  nor_x2_sg U45104 ( .A(n9625), .B(n9373), .X(n9622) );
  nand_x2_sg U45105 ( .A(n9577), .B(n23511), .X(n23508) );
  nand_x2_sg U45106 ( .A(n23676), .B(n9577), .X(n23674) );
  nor_x2_sg U45107 ( .A(n9577), .B(n9373), .X(n9574) );
  nand_x2_sg U45108 ( .A(n9528), .B(n23306), .X(n23303) );
  nand_x2_sg U45109 ( .A(n23486), .B(n9528), .X(n23484) );
  nor_x2_sg U45110 ( .A(n9528), .B(n9373), .X(n9525) );
  nand_x2_sg U45111 ( .A(n9479), .B(n23080), .X(n23077) );
  nand_x2_sg U45112 ( .A(n23281), .B(n9479), .X(n23279) );
  nor_x2_sg U45113 ( .A(n9479), .B(n9373), .X(n9476) );
  nand_x2_sg U45114 ( .A(n9430), .B(n22825), .X(n22822) );
  nand_x2_sg U45115 ( .A(n23055), .B(n9430), .X(n23053) );
  nor_x2_sg U45116 ( .A(n9430), .B(n9373), .X(n9427) );
  nand_x2_sg U45117 ( .A(n25181), .B(n30360), .X(n30575) );
  nand_x2_sg U45118 ( .A(n30358), .B(n25181), .X(n30356) );
  nor_x2_sg U45119 ( .A(n25181), .B(n9394), .X(n25178) );
  nand_x2_sg U45120 ( .A(n25084), .B(n30372), .X(n30569) );
  nand_x2_sg U45121 ( .A(n30370), .B(n25084), .X(n30368) );
  nor_x2_sg U45122 ( .A(n25084), .B(n9394), .X(n25081) );
  nand_x2_sg U45123 ( .A(n24813), .B(n29981), .X(n30030) );
  nor_x2_sg U45124 ( .A(n24813), .B(n9415), .X(n24804) );
  nand_x2_sg U45125 ( .A(n10073), .B(n22694), .X(n22909) );
  nand_x2_sg U45126 ( .A(n22692), .B(n10073), .X(n22690) );
  nor_x2_sg U45127 ( .A(n10073), .B(n9394), .X(n10070) );
  nand_x2_sg U45128 ( .A(n9976), .B(n22706), .X(n22903) );
  nand_x2_sg U45129 ( .A(n22704), .B(n9976), .X(n22702) );
  nor_x2_sg U45130 ( .A(n9976), .B(n9394), .X(n9973) );
  nand_x2_sg U45131 ( .A(n9705), .B(n22316), .X(n22365) );
  nor_x2_sg U45132 ( .A(n9705), .B(n9415), .X(n9696) );
  nand_x2_sg U45133 ( .A(n25258), .B(n31880), .X(n31969) );
  nor_x2_sg U45134 ( .A(n25258), .B(n9373), .X(n25257) );
  nand_x2_sg U45135 ( .A(n25209), .B(n31886), .X(n31966) );
  nor_x2_sg U45136 ( .A(n25209), .B(n9373), .X(n25208) );
  nand_x2_sg U45137 ( .A(n25160), .B(n31892), .X(n31963) );
  nor_x2_sg U45138 ( .A(n25160), .B(n9373), .X(n25159) );
  nand_x2_sg U45139 ( .A(n25112), .B(n31898), .X(n31960) );
  nor_x2_sg U45140 ( .A(n25112), .B(n9373), .X(n25111) );
  nand_x2_sg U45141 ( .A(n25230), .B(n30354), .X(n30578) );
  nand_x2_sg U45142 ( .A(n30352), .B(n25230), .X(n30350) );
  nor_x2_sg U45143 ( .A(n25230), .B(n9394), .X(n25227) );
  nand_x2_sg U45144 ( .A(n25063), .B(n31904), .X(n31957) );
  nor_x2_sg U45145 ( .A(n25063), .B(n9373), .X(n25062) );
  nand_x2_sg U45146 ( .A(n25015), .B(n31910), .X(n31954) );
  nor_x2_sg U45147 ( .A(n25015), .B(n9373), .X(n25014) );
  nand_x2_sg U45148 ( .A(n24967), .B(n31916), .X(n31951) );
  nor_x2_sg U45149 ( .A(n24967), .B(n9373), .X(n24966) );
  nand_x2_sg U45150 ( .A(n24919), .B(n31922), .X(n31948) );
  nor_x2_sg U45151 ( .A(n24919), .B(n9373), .X(n24918) );
  nand_x2_sg U45152 ( .A(n24871), .B(n31835), .X(n31832) );
  nand_x2_sg U45153 ( .A(n31926), .B(n24871), .X(n31924) );
  nor_x2_sg U45154 ( .A(n24871), .B(n9373), .X(n24870) );
  nand_x2_sg U45155 ( .A(n24823), .B(n31691), .X(n31688) );
  nand_x2_sg U45156 ( .A(n31810), .B(n24823), .X(n31808) );
  nor_x2_sg U45157 ( .A(n24823), .B(n9373), .X(n24822) );
  nand_x2_sg U45158 ( .A(n24728), .B(n31367), .X(n31364) );
  nand_x2_sg U45159 ( .A(n31513), .B(n24728), .X(n31511) );
  nor_x2_sg U45160 ( .A(n24728), .B(n9373), .X(n24727) );
  nand_x2_sg U45161 ( .A(n24631), .B(n30972), .X(n30969) );
  nand_x2_sg U45162 ( .A(n31152), .B(n24631), .X(n31150) );
  nor_x2_sg U45163 ( .A(n24631), .B(n9373), .X(n24630) );
  nand_x2_sg U45164 ( .A(n24533), .B(n30491), .X(n30488) );
  nand_x2_sg U45165 ( .A(n30721), .B(n24533), .X(n30719) );
  nor_x2_sg U45166 ( .A(n24533), .B(n9373), .X(n24532) );
  nand_x2_sg U45167 ( .A(n10106), .B(n24220), .X(n24300) );
  nor_x2_sg U45168 ( .A(n10106), .B(n9373), .X(n10103) );
  nand_x2_sg U45169 ( .A(n10057), .B(n24226), .X(n24297) );
  nor_x2_sg U45170 ( .A(n10057), .B(n9373), .X(n10054) );
  nand_x2_sg U45171 ( .A(n10122), .B(n22688), .X(n22912) );
  nand_x2_sg U45172 ( .A(n22686), .B(n10122), .X(n22684) );
  nor_x2_sg U45173 ( .A(n10122), .B(n9394), .X(n10119) );
  nand_x2_sg U45174 ( .A(n24680), .B(n31177), .X(n31174) );
  nand_x2_sg U45175 ( .A(n31342), .B(n24680), .X(n31340) );
  nor_x2_sg U45176 ( .A(n24680), .B(n9373), .X(n24679) );
  nand_x2_sg U45177 ( .A(n24582), .B(n30746), .X(n30743) );
  nand_x2_sg U45178 ( .A(n30947), .B(n24582), .X(n30945) );
  nor_x2_sg U45179 ( .A(n24582), .B(n9373), .X(n24581) );
  nand_x2_sg U45180 ( .A(n25279), .B(n30348), .X(n30581) );
  nand_x2_sg U45181 ( .A(n30346), .B(n25279), .X(n30344) );
  nor_x2_sg U45182 ( .A(n25279), .B(n9394), .X(n25276) );
  nand_x2_sg U45183 ( .A(n10171), .B(n22682), .X(n22915) );
  nand_x2_sg U45184 ( .A(n22680), .B(n10171), .X(n22678) );
  nor_x2_sg U45185 ( .A(n10171), .B(n9394), .X(n10168) );
  nand_x2_sg U45186 ( .A(n24776), .B(n31538), .X(n31535) );
  nand_x2_sg U45187 ( .A(n31666), .B(n24776), .X(n31664) );
  nor_x2_sg U45188 ( .A(n24776), .B(n9373), .X(n24775) );
  nand_x2_sg U45189 ( .A(n30466), .B(n24483), .X(n30464) );
  nor_x2_sg U45190 ( .A(n24483), .B(n9373), .X(n24482) );
  nand_x2_sg U45191 ( .A(n22800), .B(n9372), .X(n22798) );
  nor_x2_sg U45192 ( .A(n9372), .B(n9373), .X(n9368) );
  inv_x4_sg U45193 ( .A(n25627), .X(n51515) );
  inv_x4_sg U45194 ( .A(n53685), .X(n43735) );
  inv_x8_sg U45195 ( .A(n43735), .X(n43736) );
  nor_x8_sg U45196 ( .A(n43736), .B(n42507), .X(n17167) );
  inv_x4_sg U45197 ( .A(n53127), .X(n43737) );
  inv_x8_sg U45198 ( .A(n43737), .X(n43738) );
  nor_x8_sg U45199 ( .A(n43738), .B(n42509), .X(n15601) );
  inv_x4_sg U45200 ( .A(n52568), .X(n43739) );
  inv_x8_sg U45201 ( .A(n43739), .X(n43740) );
  nor_x8_sg U45202 ( .A(n43740), .B(n42511), .X(n14048) );
  inv_x4_sg U45203 ( .A(n52293), .X(n43741) );
  inv_x8_sg U45204 ( .A(n43741), .X(n43742) );
  nor_x8_sg U45205 ( .A(n43742), .B(n42513), .X(n13268) );
  inv_x4_sg U45206 ( .A(n52017), .X(n43743) );
  inv_x8_sg U45207 ( .A(n43743), .X(n43744) );
  nor_x8_sg U45208 ( .A(n43744), .B(n42515), .X(n12487) );
  nand_x4_sg U45209 ( .A(n11265), .B(n46532), .X(n11777) );
  inv_x2_sg U45210 ( .A(n11777), .X(n51618) );
  nor_x1_sg U45211 ( .A(n14627), .B(n14881), .X(n14878) );
  nor_x1_sg U45212 ( .A(n52844), .B(n14316), .X(n14879) );
  nor_x1_sg U45213 ( .A(n46449), .B(n14552), .X(n14894) );
  nand_x4_sg U45214 ( .A(n46358), .B(n46356), .X(n18011) );
  nor_x1_sg U45215 ( .A(n53964), .B(n46362), .X(n18000) );
  nand_x1_sg U45216 ( .A(n54124), .B(n46339), .X(n18572) );
  nand_x4_sg U45217 ( .A(n54124), .B(n46333), .X(n18780) );
  inv_x2_sg U45218 ( .A(n18780), .X(n54128) );
  nor_x1_sg U45219 ( .A(n18574), .B(n18771), .X(n18768) );
  nand_x4_sg U45220 ( .A(n46311), .B(n46309), .X(n19556) );
  nor_x1_sg U45221 ( .A(n54529), .B(n46315), .X(n19545) );
  nor_x1_sg U45222 ( .A(n54814), .B(n46295), .X(n20315) );
  nand_x4_sg U45223 ( .A(n46266), .B(n46264), .X(n21100) );
  nor_x1_sg U45224 ( .A(n55097), .B(n46270), .X(n21089) );
  nor_x1_sg U45225 ( .A(n55382), .B(n46250), .X(n21860) );
  inv_x1_sg U45226 ( .A(n22867), .X(n50861) );
  inv_x1_sg U45227 ( .A(n22165), .X(n50808) );
  inv_x1_sg U45228 ( .A(n22158), .X(n50760) );
  inv_x1_sg U45229 ( .A(n22151), .X(n50713) );
  inv_x1_sg U45230 ( .A(n22144), .X(n50665) );
  inv_x1_sg U45231 ( .A(n23012), .X(n50674) );
  inv_x1_sg U45232 ( .A(n22137), .X(n50618) );
  inv_x1_sg U45233 ( .A(n23005), .X(n50627) );
  inv_x1_sg U45234 ( .A(n22998), .X(n50578) );
  inv_x1_sg U45235 ( .A(n22130), .X(n50569) );
  inv_x1_sg U45236 ( .A(n22123), .X(n50522) );
  inv_x1_sg U45237 ( .A(n22991), .X(n50531) );
  inv_x1_sg U45238 ( .A(n22116), .X(n50475) );
  inv_x1_sg U45239 ( .A(n22984), .X(n50484) );
  inv_x1_sg U45240 ( .A(n22109), .X(n50429) );
  inv_x1_sg U45241 ( .A(n22977), .X(n50438) );
  inv_x1_sg U45242 ( .A(n22102), .X(n50382) );
  inv_x1_sg U45243 ( .A(n22970), .X(n50391) );
  inv_x1_sg U45244 ( .A(n22095), .X(n50335) );
  inv_x1_sg U45245 ( .A(n22963), .X(n50344) );
  inv_x1_sg U45246 ( .A(n22088), .X(n50289) );
  inv_x1_sg U45247 ( .A(n22081), .X(n50243) );
  inv_x1_sg U45248 ( .A(n22949), .X(n50252) );
  inv_x1_sg U45249 ( .A(n22074), .X(n50199) );
  inv_x1_sg U45250 ( .A(n22067), .X(n50156) );
  nand_x1_sg U45251 ( .A(n46564), .B(n51334), .X(n10793) );
  inv_x2_sg U45252 ( .A(n10949), .X(n43797) );
  nor_x1_sg U45253 ( .A(n10953), .B(n10954), .X(n10949) );
  inv_x1_sg U45254 ( .A(n11590), .X(n51612) );
  nand_x1_sg U45255 ( .A(n46532), .B(n46540), .X(n11574) );
  nor_x1_sg U45256 ( .A(n11438), .B(n51560), .X(n11781) );
  nor_x1_sg U45257 ( .A(n46545), .B(n11623), .X(n11772) );
  nand_x4_sg U45258 ( .A(n11796), .B(n11797), .X(n11787) );
  nand_x1_sg U45259 ( .A(n51740), .B(n11777), .X(n11796) );
  nand_x1_sg U45260 ( .A(n51618), .B(n11778), .X(n11797) );
  inv_x1_sg U45261 ( .A(n11778), .X(n51740) );
  nand_x4_sg U45262 ( .A(n51717), .B(n46547), .X(n11637) );
  nand_x1_sg U45263 ( .A(n51661), .B(n11619), .X(n11625) );
  nand_x1_sg U45264 ( .A(n51672), .B(n11618), .X(n11624) );
  nand_x4_sg U45265 ( .A(n46536), .B(n46532), .X(n11628) );
  nand_x4_sg U45266 ( .A(n11815), .B(n11816), .X(n11627) );
  nand_x1_sg U45267 ( .A(n51744), .B(n11810), .X(n11815) );
  nand_x1_sg U45268 ( .A(n51609), .B(n11811), .X(n11816) );
  nand_x1_sg U45269 ( .A(n11764), .B(n11765), .X(n11763) );
  nand_x1_sg U45270 ( .A(n11769), .B(n51755), .X(n11764) );
  nand_x1_sg U45271 ( .A(n11688), .B(n46551), .X(n11690) );
  nand_x1_sg U45272 ( .A(n51879), .B(n11833), .X(n12100) );
  nand_x1_sg U45273 ( .A(n46517), .B(n51896), .X(n12355) );
  nand_x1_sg U45274 ( .A(n12467), .B(n46529), .X(n12469) );
  inv_x1_sg U45275 ( .A(n13151), .X(n52170) );
  nand_x1_sg U45276 ( .A(n46488), .B(n46496), .X(n13135) );
  inv_x2_sg U45277 ( .A(n13348), .X(n44436) );
  nor_x1_sg U45278 ( .A(n13354), .B(n13198), .X(n13348) );
  nand_x1_sg U45279 ( .A(n52217), .B(n13180), .X(n13186) );
  nand_x1_sg U45280 ( .A(n52228), .B(n13179), .X(n13185) );
  nand_x4_sg U45281 ( .A(n52133), .B(n46488), .X(n13189) );
  nand_x4_sg U45282 ( .A(n13372), .B(n13373), .X(n13188) );
  nand_x1_sg U45283 ( .A(n52301), .B(n13367), .X(n13372) );
  nand_x1_sg U45284 ( .A(n52167), .B(n13368), .X(n13373) );
  nand_x1_sg U45285 ( .A(n13248), .B(n46507), .X(n13250) );
  inv_x1_sg U45286 ( .A(n13931), .X(n52444) );
  nand_x1_sg U45287 ( .A(n52447), .B(n46474), .X(n13915) );
  inv_x2_sg U45288 ( .A(n14128), .X(n44434) );
  nor_x1_sg U45289 ( .A(n14134), .B(n13978), .X(n14128) );
  nand_x1_sg U45290 ( .A(n52494), .B(n13960), .X(n13966) );
  nand_x1_sg U45291 ( .A(n52505), .B(n13959), .X(n13965) );
  nand_x4_sg U45292 ( .A(n52447), .B(n52406), .X(n13969) );
  nand_x4_sg U45293 ( .A(n14152), .B(n14153), .X(n13968) );
  nand_x1_sg U45294 ( .A(n52576), .B(n14147), .X(n14152) );
  nand_x1_sg U45295 ( .A(n52441), .B(n14148), .X(n14153) );
  nand_x1_sg U45296 ( .A(n14028), .B(n46484), .X(n14030) );
  nand_x1_sg U45297 ( .A(n46443), .B(n46450), .X(n14685) );
  inv_x1_sg U45298 ( .A(n14886), .X(n52843) );
  inv_x1_sg U45299 ( .A(n14740), .X(n52728) );
  inv_x1_sg U45300 ( .A(n14920), .X(n52875) );
  nand_x1_sg U45301 ( .A(n14924), .B(n14926), .X(n14925) );
  nand_x1_sg U45302 ( .A(n52713), .B(n52853), .X(n14926) );
  nand_x1_sg U45303 ( .A(n52850), .B(n14890), .X(n14909) );
  inv_x1_sg U45304 ( .A(n14891), .X(n52850) );
  nand_x4_sg U45305 ( .A(n46443), .B(n52683), .X(n14740) );
  nand_x4_sg U45306 ( .A(n14927), .B(n14928), .X(n14739) );
  nand_x1_sg U45307 ( .A(n52713), .B(n14922), .X(n14927) );
  nand_x1_sg U45308 ( .A(n52853), .B(n14923), .X(n14928) );
  nand_x1_sg U45309 ( .A(n14876), .B(n14877), .X(n14875) );
  nand_x1_sg U45310 ( .A(n14878), .B(n14879), .X(n14877) );
  nand_x1_sg U45311 ( .A(n14882), .B(n52864), .X(n14876) );
  nand_x1_sg U45312 ( .A(n14800), .B(n46462), .X(n14802) );
  inv_x1_sg U45313 ( .A(n14897), .X(n52770) );
  nand_x2_sg U45314 ( .A(n14874), .B(n14832), .X(n14873) );
  nand_x1_sg U45315 ( .A(n14884), .B(n14885), .X(n14874) );
  nand_x4_sg U45316 ( .A(n14911), .B(n14912), .X(n14870) );
  nand_x1_sg U45317 ( .A(n52876), .B(n14710), .X(n14912) );
  inv_x1_sg U45318 ( .A(n14711), .X(n52876) );
  inv_x1_sg U45319 ( .A(n15484), .X(n53004) );
  nand_x1_sg U45320 ( .A(n46420), .B(n46428), .X(n15468) );
  inv_x2_sg U45321 ( .A(n15681), .X(n44432) );
  nor_x1_sg U45322 ( .A(n15687), .B(n15531), .X(n15681) );
  nand_x1_sg U45323 ( .A(n53051), .B(n15513), .X(n15519) );
  nand_x1_sg U45324 ( .A(n53062), .B(n15512), .X(n15518) );
  nand_x4_sg U45325 ( .A(n52967), .B(n46420), .X(n15522) );
  nand_x4_sg U45326 ( .A(n15705), .B(n15706), .X(n15521) );
  nand_x1_sg U45327 ( .A(n53135), .B(n15700), .X(n15705) );
  nand_x1_sg U45328 ( .A(n53001), .B(n15701), .X(n15706) );
  nand_x1_sg U45329 ( .A(n15581), .B(n46439), .X(n15583) );
  nand_x1_sg U45330 ( .A(n53266), .B(n46413), .X(n15995) );
  nand_x1_sg U45331 ( .A(n46405), .B(n53282), .X(n16250) );
  nand_x1_sg U45332 ( .A(n53410), .B(n16452), .X(n16471) );
  inv_x1_sg U45333 ( .A(n16453), .X(n53410) );
  nand_x4_sg U45334 ( .A(n53240), .B(n53282), .X(n16304) );
  nand_x4_sg U45335 ( .A(n16490), .B(n16491), .X(n16303) );
  nand_x1_sg U45336 ( .A(n53413), .B(n16485), .X(n16490) );
  nand_x1_sg U45337 ( .A(n53277), .B(n16486), .X(n16491) );
  inv_x1_sg U45338 ( .A(n17050), .X(n53562) );
  nand_x1_sg U45339 ( .A(n46376), .B(n46384), .X(n17034) );
  inv_x2_sg U45340 ( .A(n17247), .X(n44430) );
  nor_x1_sg U45341 ( .A(n17253), .B(n17097), .X(n17247) );
  nand_x1_sg U45342 ( .A(n53609), .B(n17079), .X(n17085) );
  nand_x1_sg U45343 ( .A(n53620), .B(n17078), .X(n17084) );
  nand_x4_sg U45344 ( .A(n53525), .B(n46376), .X(n17088) );
  nand_x4_sg U45345 ( .A(n17271), .B(n17272), .X(n17087) );
  nand_x1_sg U45346 ( .A(n53693), .B(n17266), .X(n17271) );
  nand_x1_sg U45347 ( .A(n53559), .B(n17267), .X(n17272) );
  nand_x1_sg U45348 ( .A(n17147), .B(n46395), .X(n17149) );
  nand_x1_sg U45349 ( .A(n46356), .B(n46361), .X(n17806) );
  inv_x1_sg U45350 ( .A(n18007), .X(n53963) );
  inv_x1_sg U45351 ( .A(n17861), .X(n53848) );
  inv_x1_sg U45352 ( .A(n18041), .X(n53995) );
  nand_x1_sg U45353 ( .A(n18045), .B(n18047), .X(n18046) );
  nand_x1_sg U45354 ( .A(n53840), .B(n53973), .X(n18047) );
  nand_x1_sg U45355 ( .A(n53970), .B(n18011), .X(n18030) );
  inv_x1_sg U45356 ( .A(n18012), .X(n53970) );
  nand_x4_sg U45357 ( .A(n53802), .B(n46356), .X(n17861) );
  nand_x4_sg U45358 ( .A(n18048), .B(n18049), .X(n17860) );
  nand_x1_sg U45359 ( .A(n53840), .B(n18043), .X(n18048) );
  nand_x1_sg U45360 ( .A(n53973), .B(n18044), .X(n18049) );
  nand_x1_sg U45361 ( .A(n17997), .B(n17998), .X(n17996) );
  nand_x1_sg U45362 ( .A(n17999), .B(n18000), .X(n17998) );
  nand_x1_sg U45363 ( .A(n18003), .B(n53984), .X(n17997) );
  nand_x1_sg U45364 ( .A(n17921), .B(n46372), .X(n17923) );
  inv_x1_sg U45365 ( .A(n18018), .X(n53890) );
  nand_x2_sg U45366 ( .A(n17995), .B(n17953), .X(n17994) );
  nand_x1_sg U45367 ( .A(n18005), .B(n18006), .X(n17995) );
  nand_x4_sg U45368 ( .A(n18032), .B(n18033), .X(n17991) );
  nand_x1_sg U45369 ( .A(n53996), .B(n17831), .X(n18033) );
  inv_x1_sg U45370 ( .A(n17832), .X(n53996) );
  nand_x1_sg U45371 ( .A(n18570), .B(n54124), .X(n18569) );
  nor_x1_sg U45372 ( .A(n41710), .B(n18437), .X(n18573) );
  inv_x1_sg U45373 ( .A(n18824), .X(n54170) );
  nor_x1_sg U45374 ( .A(n46346), .B(n18623), .X(n18775) );
  nand_x4_sg U45375 ( .A(n18799), .B(n18800), .X(n18790) );
  nand_x1_sg U45376 ( .A(n54252), .B(n18780), .X(n18799) );
  nand_x1_sg U45377 ( .A(n54128), .B(n18781), .X(n18800) );
  inv_x1_sg U45378 ( .A(n18781), .X(n54252) );
  nand_x4_sg U45379 ( .A(n54229), .B(n46348), .X(n18637) );
  nand_x1_sg U45380 ( .A(n18766), .B(n18767), .X(n18765) );
  nand_x1_sg U45381 ( .A(n18772), .B(n54267), .X(n18766) );
  nand_x1_sg U45382 ( .A(n18768), .B(n18769), .X(n18767) );
  nand_x4_sg U45383 ( .A(n54229), .B(n46343), .X(n18741) );
  nand_x1_sg U45384 ( .A(n18690), .B(n46352), .X(n18692) );
  nand_x1_sg U45385 ( .A(n46309), .B(n46314), .X(n19351) );
  inv_x1_sg U45386 ( .A(n19552), .X(n54528) );
  inv_x1_sg U45387 ( .A(n19406), .X(n54413) );
  inv_x1_sg U45388 ( .A(n19586), .X(n54560) );
  nand_x1_sg U45389 ( .A(n19590), .B(n19592), .X(n19591) );
  nand_x1_sg U45390 ( .A(n54405), .B(n54538), .X(n19592) );
  nand_x1_sg U45391 ( .A(n54535), .B(n19556), .X(n19575) );
  inv_x1_sg U45392 ( .A(n19557), .X(n54535) );
  nand_x4_sg U45393 ( .A(n54367), .B(n46309), .X(n19406) );
  nand_x4_sg U45394 ( .A(n19593), .B(n19594), .X(n19405) );
  nand_x1_sg U45395 ( .A(n54405), .B(n19588), .X(n19593) );
  nand_x1_sg U45396 ( .A(n54538), .B(n19589), .X(n19594) );
  nand_x1_sg U45397 ( .A(n19542), .B(n19543), .X(n19541) );
  nand_x1_sg U45398 ( .A(n19544), .B(n19545), .X(n19543) );
  nand_x1_sg U45399 ( .A(n19548), .B(n54549), .X(n19542) );
  nand_x1_sg U45400 ( .A(n19466), .B(n46325), .X(n19468) );
  inv_x1_sg U45401 ( .A(n19563), .X(n54455) );
  nand_x2_sg U45402 ( .A(n19540), .B(n19498), .X(n19539) );
  nand_x1_sg U45403 ( .A(n19550), .B(n19551), .X(n19540) );
  nand_x4_sg U45404 ( .A(n19577), .B(n19578), .X(n19536) );
  nand_x1_sg U45405 ( .A(n54561), .B(n19376), .X(n19578) );
  inv_x1_sg U45406 ( .A(n19377), .X(n54561) );
  nand_x1_sg U45407 ( .A(n46294), .B(n54688), .X(n20119) );
  inv_x1_sg U45408 ( .A(n20369), .X(n54736) );
  nand_x4_sg U45409 ( .A(n54794), .B(n46296), .X(n20287) );
  nand_x1_sg U45410 ( .A(n54820), .B(n20326), .X(n20345) );
  inv_x1_sg U45411 ( .A(n20327), .X(n54820) );
  nand_x1_sg U45412 ( .A(n20312), .B(n20313), .X(n20311) );
  nand_x1_sg U45413 ( .A(n20314), .B(n20315), .X(n20313) );
  nand_x1_sg U45414 ( .A(n20318), .B(n54834), .X(n20312) );
  nand_x1_sg U45415 ( .A(n20236), .B(n46305), .X(n20238) );
  nand_x1_sg U45416 ( .A(n46264), .B(n46269), .X(n20895) );
  inv_x1_sg U45417 ( .A(n21096), .X(n55096) );
  inv_x1_sg U45418 ( .A(n20950), .X(n54981) );
  inv_x1_sg U45419 ( .A(n21130), .X(n55128) );
  nand_x1_sg U45420 ( .A(n21134), .B(n21136), .X(n21135) );
  nand_x1_sg U45421 ( .A(n54973), .B(n55106), .X(n21136) );
  nand_x1_sg U45422 ( .A(n55103), .B(n21100), .X(n21119) );
  inv_x1_sg U45423 ( .A(n21101), .X(n55103) );
  nand_x4_sg U45424 ( .A(n54935), .B(n46264), .X(n20950) );
  nand_x4_sg U45425 ( .A(n21137), .B(n21138), .X(n20949) );
  nand_x1_sg U45426 ( .A(n54973), .B(n21132), .X(n21137) );
  nand_x1_sg U45427 ( .A(n55106), .B(n21133), .X(n21138) );
  nand_x1_sg U45428 ( .A(n21086), .B(n21087), .X(n21085) );
  nand_x1_sg U45429 ( .A(n21088), .B(n21089), .X(n21087) );
  nand_x1_sg U45430 ( .A(n21092), .B(n55117), .X(n21086) );
  nand_x1_sg U45431 ( .A(n21010), .B(n46280), .X(n21012) );
  inv_x1_sg U45432 ( .A(n21107), .X(n55023) );
  nand_x2_sg U45433 ( .A(n21084), .B(n21042), .X(n21083) );
  nand_x1_sg U45434 ( .A(n21094), .B(n21095), .X(n21084) );
  nand_x4_sg U45435 ( .A(n21121), .B(n21122), .X(n21080) );
  nand_x1_sg U45436 ( .A(n55129), .B(n20920), .X(n21122) );
  inv_x1_sg U45437 ( .A(n20921), .X(n55129) );
  nand_x1_sg U45438 ( .A(n46249), .B(n55256), .X(n21664) );
  inv_x1_sg U45439 ( .A(n21914), .X(n55304) );
  nand_x4_sg U45440 ( .A(n55362), .B(n46251), .X(n21832) );
  nand_x1_sg U45441 ( .A(n55388), .B(n21871), .X(n21890) );
  inv_x1_sg U45442 ( .A(n21872), .X(n55388) );
  nand_x1_sg U45443 ( .A(n21857), .B(n21858), .X(n21856) );
  nand_x1_sg U45444 ( .A(n21859), .B(n21860), .X(n21858) );
  nand_x1_sg U45445 ( .A(n21863), .B(n55402), .X(n21857) );
  nand_x1_sg U45446 ( .A(n21781), .B(n46260), .X(n21783) );
  inv_x1_sg U45447 ( .A(n30533), .X(n50002) );
  inv_x1_sg U45448 ( .A(n29830), .X(n49949) );
  inv_x1_sg U45449 ( .A(n29823), .X(n49901) );
  inv_x1_sg U45450 ( .A(n29816), .X(n49854) );
  inv_x1_sg U45451 ( .A(n29809), .X(n49806) );
  inv_x1_sg U45452 ( .A(n30678), .X(n49815) );
  inv_x1_sg U45453 ( .A(n29802), .X(n49759) );
  inv_x1_sg U45454 ( .A(n30671), .X(n49768) );
  inv_x1_sg U45455 ( .A(n30664), .X(n49719) );
  inv_x1_sg U45456 ( .A(n29795), .X(n49710) );
  inv_x1_sg U45457 ( .A(n29788), .X(n49663) );
  inv_x1_sg U45458 ( .A(n30657), .X(n49672) );
  inv_x1_sg U45459 ( .A(n29781), .X(n49616) );
  inv_x1_sg U45460 ( .A(n30650), .X(n49625) );
  inv_x1_sg U45461 ( .A(n29774), .X(n49570) );
  inv_x1_sg U45462 ( .A(n30643), .X(n49579) );
  inv_x1_sg U45463 ( .A(n29767), .X(n49523) );
  inv_x1_sg U45464 ( .A(n30636), .X(n49532) );
  inv_x1_sg U45465 ( .A(n29760), .X(n49476) );
  inv_x1_sg U45466 ( .A(n30629), .X(n49485) );
  inv_x1_sg U45467 ( .A(n29753), .X(n49430) );
  inv_x1_sg U45468 ( .A(n29746), .X(n49384) );
  inv_x1_sg U45469 ( .A(n30615), .X(n49393) );
  inv_x1_sg U45470 ( .A(n29739), .X(n49340) );
  inv_x1_sg U45471 ( .A(n29732), .X(n49297) );
  inv_x1_sg U45472 ( .A(n22195), .X(n50902) );
  inv_x1_sg U45473 ( .A(n23031), .X(n50817) );
  inv_x1_sg U45474 ( .A(n23025), .X(n50769) );
  inv_x1_sg U45475 ( .A(n23019), .X(n50722) );
  inv_x1_sg U45476 ( .A(n24131), .X(n50496) );
  inv_x1_sg U45477 ( .A(n24124), .X(n50450) );
  inv_x1_sg U45478 ( .A(n24117), .X(n50404) );
  inv_x1_sg U45479 ( .A(n24110), .X(n50356) );
  inv_x1_sg U45480 ( .A(n24348), .X(n50361) );
  inv_x1_sg U45481 ( .A(n22956), .X(n50298) );
  inv_x1_sg U45482 ( .A(n24103), .X(n50310) );
  inv_x1_sg U45483 ( .A(n24096), .X(n50265) );
  inv_x1_sg U45484 ( .A(n24335), .X(n50270) );
  inv_x1_sg U45485 ( .A(n22942), .X(n50208) );
  inv_x1_sg U45486 ( .A(n24089), .X(n50220) );
  inv_x1_sg U45487 ( .A(n22935), .X(n50162) );
  inv_x1_sg U45488 ( .A(n24082), .X(n50172) );
  nand_x1_sg U45489 ( .A(n51306), .B(n46572), .X(n10515) );
  nand_x4_sg U45490 ( .A(n46557), .B(n46574), .X(n10614) );
  inv_x1_sg U45491 ( .A(n10580), .X(n51301) );
  inv_x1_sg U45492 ( .A(n10614), .X(n51356) );
  nand_x1_sg U45493 ( .A(n10615), .B(n46572), .X(n10654) );
  nand_x1_sg U45494 ( .A(n51319), .B(n10646), .X(n10659) );
  nand_x1_sg U45495 ( .A(n51308), .B(n10645), .X(n10658) );
  nand_x4_sg U45496 ( .A(n51306), .B(n46564), .X(n10646) );
  nand_x1_sg U45497 ( .A(n10791), .B(n46564), .X(n10790) );
  nand_x1_sg U45498 ( .A(n10788), .B(n46557), .X(n10787) );
  nand_x4_sg U45499 ( .A(n51306), .B(n51293), .X(n10777) );
  inv_x2_sg U45500 ( .A(n11003), .X(n44502) );
  nor_x1_sg U45501 ( .A(n11012), .B(n11013), .X(n11003) );
  inv_x1_sg U45502 ( .A(n10856), .X(n51446) );
  nor_x1_sg U45503 ( .A(n46570), .B(n10843), .X(n10988) );
  nand_x1_sg U45504 ( .A(n10980), .B(n10981), .X(n10979) );
  nand_x1_sg U45505 ( .A(n10982), .B(n10983), .X(n10981) );
  inv_x1_sg U45506 ( .A(n11037), .X(n51382) );
  inv_x1_sg U45507 ( .A(n11034), .X(n51486) );
  nand_x1_sg U45508 ( .A(n51465), .B(n11030), .X(n11029) );
  nand_x1_sg U45509 ( .A(n51323), .B(n51463), .X(n11030) );
  inv_x1_sg U45510 ( .A(n11021), .X(n51452) );
  inv_x1_sg U45511 ( .A(n10855), .X(n51447) );
  inv_x1_sg U45512 ( .A(n11006), .X(n51373) );
  nand_x1_sg U45513 ( .A(n10974), .B(n42053), .X(n10969) );
  nand_x1_sg U45514 ( .A(n10942), .B(n46564), .X(n10941) );
  nand_x1_sg U45515 ( .A(n10936), .B(n10937), .X(n10938) );
  nand_x1_sg U45516 ( .A(n11265), .B(n11050), .X(n11294) );
  nand_x1_sg U45517 ( .A(n51598), .B(n46547), .X(n11320) );
  nand_x1_sg U45518 ( .A(n51630), .B(n46551), .X(n11392) );
  nand_x1_sg U45519 ( .A(n51630), .B(n46547), .X(n11433) );
  nand_x4_sg U45520 ( .A(n11265), .B(n46540), .X(n11426) );
  nand_x1_sg U45521 ( .A(n51608), .B(n11426), .X(n11440) );
  nand_x1_sg U45522 ( .A(n51595), .B(n11425), .X(n11439) );
  inv_x1_sg U45523 ( .A(n11589), .X(n51708) );
  nand_x1_sg U45524 ( .A(n11572), .B(n46532), .X(n11571) );
  nand_x4_sg U45525 ( .A(n46539), .B(n46532), .X(n11582) );
  nand_x1_sg U45526 ( .A(n11569), .B(n51630), .X(n11568) );
  inv_x1_sg U45527 ( .A(n11628), .X(n51619) );
  inv_x1_sg U45528 ( .A(n11808), .X(n51766) );
  nand_x1_sg U45529 ( .A(n11812), .B(n11814), .X(n11813) );
  inv_x1_sg U45530 ( .A(n11784), .X(n51664) );
  nand_x2_sg U45531 ( .A(n11762), .B(n11720), .X(n11761) );
  nand_x1_sg U45532 ( .A(n11770), .B(n11771), .X(n11762) );
  nand_x4_sg U45533 ( .A(n11798), .B(n11799), .X(n11758) );
  nand_x1_sg U45534 ( .A(n51767), .B(n40531), .X(n11799) );
  nand_x1_sg U45535 ( .A(n11787), .B(n11786), .X(n11795) );
  nand_x4_sg U45536 ( .A(n11634), .B(n11635), .X(n11594) );
  nand_x1_sg U45537 ( .A(n51726), .B(n51713), .X(n11635) );
  nand_x1_sg U45538 ( .A(n11636), .B(n11637), .X(n11634) );
  inv_x1_sg U45539 ( .A(n11636), .X(n51713) );
  nand_x1_sg U45540 ( .A(n11627), .B(n11628), .X(n11629) );
  nand_x1_sg U45541 ( .A(n11719), .B(n11720), .X(n11721) );
  inv_x1_sg U45542 ( .A(n11761), .X(n51758) );
  nand_x1_sg U45543 ( .A(n51598), .B(n51630), .X(n11751) );
  nand_x1_sg U45544 ( .A(n11758), .B(n41867), .X(n11753) );
  nand_x1_sg U45545 ( .A(n11687), .B(n11688), .X(n11686) );
  nand_x1_sg U45546 ( .A(n51911), .B(n46529), .X(n12172) );
  nand_x1_sg U45547 ( .A(n12098), .B(n51879), .X(n12097) );
  nand_x4_sg U45548 ( .A(n51896), .B(n46525), .X(n12134) );
  inv_x2_sg U45549 ( .A(n12046), .X(n51862) );
  nand_x1_sg U45550 ( .A(n51911), .B(n46525), .X(n12213) );
  nand_x4_sg U45551 ( .A(n51826), .B(n51879), .X(n12205) );
  nand_x1_sg U45552 ( .A(n51867), .B(n12205), .X(n12219) );
  nand_x1_sg U45553 ( .A(n51889), .B(n12206), .X(n12220) );
  inv_x1_sg U45554 ( .A(n12294), .X(n51955) );
  nand_x1_sg U45555 ( .A(n12353), .B(n46517), .X(n12352) );
  nand_x4_sg U45556 ( .A(n51896), .B(n51839), .X(n12362) );
  nand_x4_sg U45557 ( .A(n51911), .B(n46517), .X(n12361) );
  nand_x1_sg U45558 ( .A(n12350), .B(n51911), .X(n12349) );
  inv_x1_sg U45559 ( .A(n12311), .X(n51987) );
  inv_x1_sg U45560 ( .A(n12583), .X(n52046) );
  nand_x1_sg U45561 ( .A(n52027), .B(n12589), .X(n12588) );
  nand_x1_sg U45562 ( .A(n51942), .B(n12400), .X(n12406) );
  nand_x1_sg U45563 ( .A(n51953), .B(n12399), .X(n12405) );
  inv_x1_sg U45564 ( .A(n12566), .X(n52021) );
  nand_x4_sg U45565 ( .A(n52004), .B(n12415), .X(n12375) );
  inv_x1_sg U45566 ( .A(n12418), .X(n52004) );
  nand_x1_sg U45567 ( .A(n12416), .B(n12417), .X(n12415) );
  nand_x1_sg U45568 ( .A(n12505), .B(n46517), .X(n12504) );
  nand_x1_sg U45569 ( .A(n12536), .B(n12537), .X(n12533) );
  nand_x1_sg U45570 ( .A(n51911), .B(n51879), .X(n12531) );
  nand_x1_sg U45571 ( .A(n12466), .B(n12467), .X(n12465) );
  nand_x1_sg U45572 ( .A(n52156), .B(n46503), .X(n12881) );
  nand_x1_sg U45573 ( .A(n52187), .B(n46507), .X(n12953) );
  nand_x4_sg U45574 ( .A(n46488), .B(n46503), .X(n12915) );
  inv_x2_sg U45575 ( .A(n12828), .X(n52139) );
  nand_x1_sg U45576 ( .A(n52187), .B(n46503), .X(n12994) );
  nand_x1_sg U45577 ( .A(n52166), .B(n12987), .X(n13001) );
  nand_x1_sg U45578 ( .A(n52153), .B(n12986), .X(n13000) );
  inv_x1_sg U45579 ( .A(n13150), .X(n52264) );
  nand_x1_sg U45580 ( .A(n13133), .B(n46488), .X(n13132) );
  nand_x4_sg U45581 ( .A(n46495), .B(n46488), .X(n13143) );
  nand_x1_sg U45582 ( .A(n13130), .B(n52187), .X(n13129) );
  inv_x1_sg U45583 ( .A(n13189), .X(n52178) );
  inv_x1_sg U45584 ( .A(n13365), .X(n52322) );
  nand_x1_sg U45585 ( .A(n13369), .B(n13371), .X(n13370) );
  nor_x1_sg U45586 ( .A(n12999), .B(n52117), .X(n13334) );
  inv_x1_sg U45587 ( .A(n13346), .X(n52297) );
  inv_x2_sg U45588 ( .A(n52298), .X(n45536) );
  inv_x1_sg U45589 ( .A(n13339), .X(n52298) );
  nand_x1_sg U45590 ( .A(n13188), .B(n13189), .X(n13190) );
  nand_x1_sg U45591 ( .A(n13318), .B(n13317), .X(n13314) );
  nand_x1_sg U45592 ( .A(n52156), .B(n52187), .X(n13312) );
  nand_x1_sg U45593 ( .A(n13247), .B(n13248), .X(n13246) );
  nand_x1_sg U45594 ( .A(n52463), .B(n46484), .X(n13733) );
  nand_x4_sg U45595 ( .A(n52447), .B(n46481), .X(n13695) );
  inv_x2_sg U45596 ( .A(n13607), .X(n52414) );
  nand_x1_sg U45597 ( .A(n52463), .B(n46481), .X(n13774) );
  nand_x4_sg U45598 ( .A(n52430), .B(n52378), .X(n13766) );
  nand_x1_sg U45599 ( .A(n52419), .B(n13766), .X(n13780) );
  nand_x1_sg U45600 ( .A(n52440), .B(n13767), .X(n13781) );
  inv_x1_sg U45601 ( .A(n13855), .X(n52507) );
  inv_x1_sg U45602 ( .A(n13930), .X(n52540) );
  nand_x1_sg U45603 ( .A(n13913), .B(n52447), .X(n13912) );
  nand_x4_sg U45604 ( .A(n52463), .B(n46474), .X(n13922) );
  nand_x4_sg U45605 ( .A(n52447), .B(n52391), .X(n13923) );
  nand_x1_sg U45606 ( .A(n13910), .B(n52463), .X(n13909) );
  inv_x1_sg U45607 ( .A(n13969), .X(n52453) );
  inv_x1_sg U45608 ( .A(n14145), .X(n52597) );
  nand_x1_sg U45609 ( .A(n14149), .B(n14151), .X(n14150) );
  inv_x1_sg U45610 ( .A(n14126), .X(n52572) );
  inv_x2_sg U45611 ( .A(n52573), .X(n45534) );
  inv_x1_sg U45612 ( .A(n14119), .X(n52573) );
  nand_x1_sg U45613 ( .A(n13968), .B(n13969), .X(n13970) );
  nand_x1_sg U45614 ( .A(n14098), .B(n14097), .X(n14094) );
  nand_x1_sg U45615 ( .A(n52463), .B(n52430), .X(n14092) );
  nand_x1_sg U45616 ( .A(n14027), .B(n14028), .X(n14026) );
  nand_x1_sg U45617 ( .A(n52695), .B(n46458), .X(n14407) );
  nand_x1_sg U45618 ( .A(n52689), .B(n14430), .X(n14465) );
  nand_x1_sg U45619 ( .A(n52677), .B(n14429), .X(n14466) );
  inv_x1_sg U45620 ( .A(n14472), .X(n52691) );
  nand_x1_sg U45621 ( .A(n52784), .B(n14730), .X(n14736) );
  nand_x1_sg U45622 ( .A(n52767), .B(n14731), .X(n14737) );
  nand_x1_sg U45623 ( .A(n52747), .B(n14692), .X(n14702) );
  nand_x1_sg U45624 ( .A(n52726), .B(n14691), .X(n14701) );
  nand_x4_sg U45625 ( .A(n52707), .B(n52655), .X(n14537) );
  inv_x1_sg U45626 ( .A(n14626), .X(n52786) );
  nand_x1_sg U45627 ( .A(n14683), .B(n46443), .X(n14682) );
  nand_x4_sg U45628 ( .A(n52695), .B(n52683), .X(n14669) );
  inv_x1_sg U45629 ( .A(n14914), .X(n52845) );
  nand_x4_sg U45630 ( .A(n14911), .B(n14918), .X(n14711) );
  nand_x1_sg U45631 ( .A(n14919), .B(n14920), .X(n14918) );
  inv_x1_sg U45632 ( .A(n14749), .X(n52838) );
  nand_x1_sg U45633 ( .A(n14739), .B(n14740), .X(n14741) );
  nand_x1_sg U45634 ( .A(n14831), .B(n14832), .X(n14833) );
  inv_x1_sg U45635 ( .A(n14873), .X(n52867) );
  inv_x2_sg U45636 ( .A(n14845), .X(n43804) );
  nor_x1_sg U45637 ( .A(n14849), .B(n14850), .X(n14845) );
  nand_x1_sg U45638 ( .A(n14870), .B(n42067), .X(n14865) );
  nand_x1_sg U45639 ( .A(n14799), .B(n14800), .X(n14798) );
  nand_x1_sg U45640 ( .A(n52872), .B(n14873), .X(n14871) );
  inv_x1_sg U45641 ( .A(n14872), .X(n52872) );
  nand_x1_sg U45642 ( .A(n52877), .B(n42067), .X(n14867) );
  nand_x1_sg U45643 ( .A(n42068), .B(n14870), .X(n14868) );
  inv_x1_sg U45644 ( .A(n14870), .X(n52877) );
  nand_x1_sg U45645 ( .A(n52990), .B(n46435), .X(n15214) );
  nand_x1_sg U45646 ( .A(n53021), .B(n46439), .X(n15286) );
  nand_x4_sg U45647 ( .A(n46420), .B(n46435), .X(n15248) );
  inv_x2_sg U45648 ( .A(n15161), .X(n52973) );
  nand_x1_sg U45649 ( .A(n53021), .B(n46435), .X(n15327) );
  nand_x1_sg U45650 ( .A(n53000), .B(n15320), .X(n15334) );
  nand_x1_sg U45651 ( .A(n52987), .B(n15319), .X(n15333) );
  inv_x1_sg U45652 ( .A(n15483), .X(n53098) );
  nand_x1_sg U45653 ( .A(n15466), .B(n46420), .X(n15465) );
  nand_x4_sg U45654 ( .A(n46427), .B(n46420), .X(n15476) );
  nand_x1_sg U45655 ( .A(n15463), .B(n53021), .X(n15462) );
  inv_x1_sg U45656 ( .A(n15522), .X(n53012) );
  inv_x1_sg U45657 ( .A(n15698), .X(n53156) );
  nand_x1_sg U45658 ( .A(n15702), .B(n15704), .X(n15703) );
  nor_x1_sg U45659 ( .A(n15332), .B(n52951), .X(n15667) );
  inv_x1_sg U45660 ( .A(n15679), .X(n53131) );
  inv_x2_sg U45661 ( .A(n53132), .X(n45532) );
  inv_x1_sg U45662 ( .A(n15672), .X(n53132) );
  nand_x1_sg U45663 ( .A(n15521), .B(n15522), .X(n15523) );
  nand_x1_sg U45664 ( .A(n15651), .B(n15650), .X(n15647) );
  nand_x1_sg U45665 ( .A(n52990), .B(n53021), .X(n15645) );
  nand_x1_sg U45666 ( .A(n15580), .B(n15581), .X(n15579) );
  nand_x1_sg U45667 ( .A(n53253), .B(n46413), .X(n15969) );
  nand_x1_sg U45668 ( .A(n15993), .B(n53266), .X(n15992) );
  nand_x4_sg U45669 ( .A(n53266), .B(n53214), .X(n16100) );
  nand_x4_sg U45670 ( .A(n46405), .B(n53253), .X(n16101) );
  nand_x1_sg U45671 ( .A(n53276), .B(n16101), .X(n16115) );
  nand_x1_sg U45672 ( .A(n53254), .B(n16100), .X(n16114) );
  inv_x1_sg U45673 ( .A(n16189), .X(n53343) );
  nand_x1_sg U45674 ( .A(n16248), .B(n46405), .X(n16247) );
  nand_x4_sg U45675 ( .A(n53227), .B(n53282), .X(n16257) );
  nand_x1_sg U45676 ( .A(n16245), .B(n53214), .X(n16244) );
  nand_x4_sg U45677 ( .A(n53240), .B(n53253), .X(n16234) );
  nor_x1_sg U45678 ( .A(n46411), .B(n16299), .X(n16447) );
  nand_x1_sg U45679 ( .A(n16438), .B(n16439), .X(n16437) );
  nand_x1_sg U45680 ( .A(n16440), .B(n16441), .X(n16439) );
  inv_x1_sg U45681 ( .A(n16480), .X(n53400) );
  inv_x1_sg U45682 ( .A(n16304), .X(n53286) );
  inv_x1_sg U45683 ( .A(n16483), .X(n53436) );
  nand_x1_sg U45684 ( .A(n16487), .B(n16489), .X(n16488) );
  nand_x4_sg U45685 ( .A(n16263), .B(n53376), .X(n16206) );
  inv_x1_sg U45686 ( .A(n16264), .X(n53376) );
  nand_x1_sg U45687 ( .A(n16265), .B(n53375), .X(n16263) );
  nand_x1_sg U45688 ( .A(n53330), .B(n16295), .X(n16301) );
  nand_x1_sg U45689 ( .A(n53341), .B(n16294), .X(n16300) );
  nand_x4_sg U45690 ( .A(n16310), .B(n53395), .X(n16269) );
  inv_x1_sg U45691 ( .A(n16311), .X(n53395) );
  nand_x1_sg U45692 ( .A(n16313), .B(n16312), .X(n16310) );
  nand_x1_sg U45693 ( .A(n16303), .B(n16304), .X(n16305) );
  nand_x1_sg U45694 ( .A(n16362), .B(n46417), .X(n16364) );
  nand_x1_sg U45695 ( .A(n16432), .B(n41865), .X(n16427) );
  nand_x1_sg U45696 ( .A(n16400), .B(n46405), .X(n16399) );
  nand_x1_sg U45697 ( .A(n16394), .B(n16395), .X(n16396) );
  nand_x1_sg U45698 ( .A(n53548), .B(n46391), .X(n16780) );
  nand_x1_sg U45699 ( .A(n53579), .B(n46395), .X(n16852) );
  nand_x4_sg U45700 ( .A(n46376), .B(n46391), .X(n16814) );
  inv_x2_sg U45701 ( .A(n16727), .X(n53531) );
  nand_x1_sg U45702 ( .A(n53579), .B(n46391), .X(n16893) );
  nand_x1_sg U45703 ( .A(n53558), .B(n16886), .X(n16900) );
  nand_x1_sg U45704 ( .A(n53545), .B(n16885), .X(n16899) );
  inv_x1_sg U45705 ( .A(n17049), .X(n53656) );
  nand_x1_sg U45706 ( .A(n17032), .B(n46376), .X(n17031) );
  nand_x4_sg U45707 ( .A(n46383), .B(n46376), .X(n17042) );
  nand_x1_sg U45708 ( .A(n17029), .B(n53579), .X(n17028) );
  inv_x1_sg U45709 ( .A(n17088), .X(n53570) );
  inv_x1_sg U45710 ( .A(n17264), .X(n53714) );
  nand_x1_sg U45711 ( .A(n17268), .B(n17270), .X(n17269) );
  nor_x1_sg U45712 ( .A(n16898), .B(n53509), .X(n17233) );
  inv_x1_sg U45713 ( .A(n17245), .X(n53689) );
  inv_x2_sg U45714 ( .A(n53690), .X(n45530) );
  inv_x1_sg U45715 ( .A(n17238), .X(n53690) );
  nand_x1_sg U45716 ( .A(n17087), .B(n17088), .X(n17089) );
  nand_x1_sg U45717 ( .A(n17217), .B(n17216), .X(n17213) );
  nand_x1_sg U45718 ( .A(n53548), .B(n53579), .X(n17211) );
  nand_x1_sg U45719 ( .A(n17146), .B(n17147), .X(n17145) );
  nand_x1_sg U45720 ( .A(n46358), .B(n17293), .X(n17528) );
  nand_x2_sg U45721 ( .A(n53827), .B(n17432), .X(n17531) );
  inv_x1_sg U45722 ( .A(n17592), .X(n53810) );
  nand_x1_sg U45723 ( .A(n53904), .B(n17851), .X(n17857) );
  nand_x1_sg U45724 ( .A(n53887), .B(n17852), .X(n17858) );
  nand_x4_sg U45725 ( .A(n46358), .B(n46361), .X(n17659) );
  nand_x4_sg U45726 ( .A(n53827), .B(n46363), .X(n17658) );
  inv_x1_sg U45727 ( .A(n17747), .X(n53906) );
  nand_x1_sg U45728 ( .A(n17804), .B(n46356), .X(n17803) );
  nand_x4_sg U45729 ( .A(n53802), .B(n46358), .X(n17790) );
  inv_x1_sg U45730 ( .A(n18035), .X(n53965) );
  nand_x4_sg U45731 ( .A(n18032), .B(n18039), .X(n17832) );
  nand_x1_sg U45732 ( .A(n18040), .B(n18041), .X(n18039) );
  inv_x1_sg U45733 ( .A(n17870), .X(n53958) );
  nand_x1_sg U45734 ( .A(n17860), .B(n17861), .X(n17862) );
  nand_x1_sg U45735 ( .A(n17952), .B(n17953), .X(n17954) );
  inv_x1_sg U45736 ( .A(n17994), .X(n53987) );
  nand_x1_sg U45737 ( .A(n17991), .B(n42061), .X(n17986) );
  nand_x1_sg U45738 ( .A(n17920), .B(n17921), .X(n17919) );
  nand_x1_sg U45739 ( .A(n53992), .B(n17994), .X(n17992) );
  inv_x1_sg U45740 ( .A(n17993), .X(n53992) );
  nand_x1_sg U45741 ( .A(n53997), .B(n42061), .X(n17988) );
  nand_x1_sg U45742 ( .A(n42062), .B(n17991), .X(n17989) );
  inv_x1_sg U45743 ( .A(n17991), .X(n53997) );
  nand_x1_sg U45744 ( .A(n46333), .B(n46348), .X(n18297) );
  nand_x4_sg U45745 ( .A(n46329), .B(n46352), .X(n18396) );
  inv_x1_sg U45746 ( .A(n18362), .X(n54093) );
  inv_x1_sg U45747 ( .A(n18396), .X(n54145) );
  nand_x1_sg U45748 ( .A(n18397), .B(n46348), .X(n18436) );
  nand_x1_sg U45749 ( .A(n54169), .B(n18619), .X(n18625) );
  nand_x1_sg U45750 ( .A(n54195), .B(n18618), .X(n18624) );
  nand_x4_sg U45751 ( .A(n54109), .B(n46343), .X(n18427) );
  nand_x4_sg U45752 ( .A(n46333), .B(n46339), .X(n18428) );
  nor_x1_sg U45753 ( .A(n18483), .B(n54159), .X(n18482) );
  nand_x1_sg U45754 ( .A(n18567), .B(n46329), .X(n18566) );
  inv_x1_sg U45755 ( .A(n18821), .X(n54277) );
  nand_x1_sg U45756 ( .A(n54258), .B(n18817), .X(n18816) );
  nand_x1_sg U45757 ( .A(n54114), .B(n54256), .X(n18817) );
  nand_x2_sg U45758 ( .A(n18764), .B(n18722), .X(n18763) );
  nand_x1_sg U45759 ( .A(n18773), .B(n18774), .X(n18764) );
  nand_x4_sg U45760 ( .A(n18801), .B(n18802), .X(n18760) );
  nand_x1_sg U45761 ( .A(n54279), .B(n40537), .X(n18802) );
  nand_x4_sg U45762 ( .A(n18744), .B(n54237), .X(n18657) );
  inv_x1_sg U45763 ( .A(n18745), .X(n54237) );
  nand_x1_sg U45764 ( .A(n54160), .B(n18741), .X(n18744) );
  nand_x1_sg U45765 ( .A(n18790), .B(n18789), .X(n18798) );
  nand_x4_sg U45766 ( .A(n18634), .B(n18635), .X(n18594) );
  nand_x1_sg U45767 ( .A(n54240), .B(n54225), .X(n18635) );
  nand_x1_sg U45768 ( .A(n18636), .B(n18637), .X(n18634) );
  inv_x1_sg U45769 ( .A(n18636), .X(n54225) );
  nand_x4_sg U45770 ( .A(n54270), .B(n18762), .X(n18721) );
  inv_x1_sg U45771 ( .A(n18763), .X(n54270) );
  nand_x1_sg U45772 ( .A(n18721), .B(n18722), .X(n18723) );
  inv_x2_sg U45773 ( .A(n18735), .X(n43942) );
  nor_x1_sg U45774 ( .A(n18739), .B(n18740), .X(n18735) );
  nand_x1_sg U45775 ( .A(n46329), .B(n54109), .X(n18753) );
  nand_x1_sg U45776 ( .A(n18760), .B(n42600), .X(n18755) );
  nand_x1_sg U45777 ( .A(n18689), .B(n18690), .X(n18688) );
  nand_x1_sg U45778 ( .A(n46311), .B(n18838), .X(n19073) );
  nand_x2_sg U45779 ( .A(n54392), .B(n18977), .X(n19076) );
  inv_x1_sg U45780 ( .A(n19137), .X(n54375) );
  nand_x1_sg U45781 ( .A(n54469), .B(n19396), .X(n19402) );
  nand_x1_sg U45782 ( .A(n54452), .B(n19397), .X(n19403) );
  nand_x4_sg U45783 ( .A(n46311), .B(n46314), .X(n19204) );
  nand_x4_sg U45784 ( .A(n54392), .B(n46316), .X(n19203) );
  inv_x1_sg U45785 ( .A(n19292), .X(n54471) );
  nand_x1_sg U45786 ( .A(n19349), .B(n46309), .X(n19348) );
  nand_x4_sg U45787 ( .A(n54367), .B(n46311), .X(n19335) );
  inv_x1_sg U45788 ( .A(n19580), .X(n54530) );
  nand_x4_sg U45789 ( .A(n19577), .B(n19584), .X(n19377) );
  nand_x1_sg U45790 ( .A(n19585), .B(n19586), .X(n19584) );
  inv_x1_sg U45791 ( .A(n19415), .X(n54523) );
  nand_x1_sg U45792 ( .A(n19405), .B(n19406), .X(n19407) );
  nand_x1_sg U45793 ( .A(n19497), .B(n19498), .X(n19499) );
  inv_x1_sg U45794 ( .A(n19539), .X(n54552) );
  nand_x1_sg U45795 ( .A(n19536), .B(n42059), .X(n19531) );
  nand_x1_sg U45796 ( .A(n19465), .B(n19466), .X(n19464) );
  nand_x1_sg U45797 ( .A(n54557), .B(n19539), .X(n19537) );
  inv_x1_sg U45798 ( .A(n19538), .X(n54557) );
  nand_x1_sg U45799 ( .A(n54562), .B(n42059), .X(n19533) );
  nand_x1_sg U45800 ( .A(n42060), .B(n19536), .X(n19534) );
  inv_x1_sg U45801 ( .A(n19536), .X(n54562) );
  nand_x1_sg U45802 ( .A(n54660), .B(n19610), .X(n19842) );
  nand_x1_sg U45803 ( .A(n54653), .B(n19820), .X(n19900) );
  nand_x1_sg U45804 ( .A(n54641), .B(n19864), .X(n19901) );
  nor_x1_sg U45805 ( .A(n19941), .B(n19940), .X(n19938) );
  inv_x1_sg U45806 ( .A(n19907), .X(n54655) );
  inv_x1_sg U45807 ( .A(n19941), .X(n54710) );
  nand_x1_sg U45808 ( .A(n19942), .B(n46301), .X(n19981) );
  nand_x1_sg U45809 ( .A(n54762), .B(n20164), .X(n20170) );
  nand_x1_sg U45810 ( .A(n54735), .B(n20165), .X(n20171) );
  nand_x1_sg U45811 ( .A(n54673), .B(n19973), .X(n19986) );
  nand_x1_sg U45812 ( .A(n54662), .B(n19972), .X(n19985) );
  nand_x4_sg U45813 ( .A(n46294), .B(n54660), .X(n19973) );
  nand_x1_sg U45814 ( .A(n20117), .B(n46294), .X(n20116) );
  nand_x1_sg U45815 ( .A(n20114), .B(n46285), .X(n20113) );
  inv_x1_sg U45816 ( .A(n20322), .X(n54813) );
  inv_x1_sg U45817 ( .A(n20366), .X(n54844) );
  nand_x1_sg U45818 ( .A(n54825), .B(n20362), .X(n20361) );
  nand_x1_sg U45819 ( .A(n54677), .B(n54823), .X(n20362) );
  nand_x2_sg U45820 ( .A(n20310), .B(n20268), .X(n20309) );
  nand_x1_sg U45821 ( .A(n20320), .B(n20321), .X(n20310) );
  nand_x4_sg U45822 ( .A(n20347), .B(n20348), .X(n20306) );
  nand_x1_sg U45823 ( .A(n54846), .B(n20144), .X(n20348) );
  inv_x1_sg U45824 ( .A(n20145), .X(n54846) );
  inv_x1_sg U45825 ( .A(n20291), .X(n54802) );
  nand_x1_sg U45826 ( .A(n54726), .B(n20287), .X(n20290) );
  inv_x1_sg U45827 ( .A(n20183), .X(n54808) );
  nand_x4_sg U45828 ( .A(n54837), .B(n20308), .X(n20267) );
  inv_x1_sg U45829 ( .A(n20309), .X(n54837) );
  nand_x1_sg U45830 ( .A(n20273), .B(n46294), .X(n20272) );
  nand_x1_sg U45831 ( .A(n20267), .B(n20268), .X(n20269) );
  inv_x2_sg U45832 ( .A(n20281), .X(n43846) );
  nor_x1_sg U45833 ( .A(n20285), .B(n20286), .X(n20281) );
  nand_x1_sg U45834 ( .A(n20306), .B(n43098), .X(n20301) );
  nand_x1_sg U45835 ( .A(n20235), .B(n20236), .X(n20234) );
  nand_x1_sg U45836 ( .A(n46266), .B(n20382), .X(n20617) );
  nand_x2_sg U45837 ( .A(n54960), .B(n20521), .X(n20620) );
  inv_x1_sg U45838 ( .A(n20681), .X(n54943) );
  nand_x1_sg U45839 ( .A(n55037), .B(n20940), .X(n20946) );
  nand_x1_sg U45840 ( .A(n55020), .B(n20941), .X(n20947) );
  nand_x4_sg U45841 ( .A(n46266), .B(n46269), .X(n20748) );
  nand_x4_sg U45842 ( .A(n54960), .B(n46271), .X(n20747) );
  inv_x1_sg U45843 ( .A(n20836), .X(n55039) );
  nand_x1_sg U45844 ( .A(n20893), .B(n46264), .X(n20892) );
  nand_x4_sg U45845 ( .A(n54935), .B(n46266), .X(n20879) );
  inv_x1_sg U45846 ( .A(n21124), .X(n55098) );
  nand_x4_sg U45847 ( .A(n21121), .B(n21128), .X(n20921) );
  nand_x1_sg U45848 ( .A(n21129), .B(n21130), .X(n21128) );
  inv_x1_sg U45849 ( .A(n20959), .X(n55091) );
  nand_x1_sg U45850 ( .A(n20949), .B(n20950), .X(n20951) );
  nand_x1_sg U45851 ( .A(n21041), .B(n21042), .X(n21043) );
  inv_x1_sg U45852 ( .A(n21083), .X(n55120) );
  nand_x1_sg U45853 ( .A(n21080), .B(n42057), .X(n21075) );
  nand_x1_sg U45854 ( .A(n21009), .B(n21010), .X(n21008) );
  nand_x1_sg U45855 ( .A(n55125), .B(n21083), .X(n21081) );
  inv_x1_sg U45856 ( .A(n21082), .X(n55125) );
  nand_x1_sg U45857 ( .A(n55130), .B(n42057), .X(n21077) );
  nand_x1_sg U45858 ( .A(n42058), .B(n21080), .X(n21078) );
  inv_x1_sg U45859 ( .A(n21080), .X(n55130) );
  nand_x1_sg U45860 ( .A(n55228), .B(n21155), .X(n21387) );
  nand_x1_sg U45861 ( .A(n55221), .B(n21365), .X(n21445) );
  nand_x1_sg U45862 ( .A(n55209), .B(n21409), .X(n21446) );
  nor_x1_sg U45863 ( .A(n21486), .B(n21485), .X(n21483) );
  inv_x1_sg U45864 ( .A(n21452), .X(n55223) );
  inv_x1_sg U45865 ( .A(n21486), .X(n55278) );
  nand_x1_sg U45866 ( .A(n21487), .B(n46256), .X(n21526) );
  nand_x1_sg U45867 ( .A(n55330), .B(n21709), .X(n21715) );
  nand_x1_sg U45868 ( .A(n55303), .B(n21710), .X(n21716) );
  nand_x1_sg U45869 ( .A(n55241), .B(n21518), .X(n21531) );
  nand_x1_sg U45870 ( .A(n55230), .B(n21517), .X(n21530) );
  nand_x4_sg U45871 ( .A(n46249), .B(n55228), .X(n21518) );
  nand_x1_sg U45872 ( .A(n21662), .B(n46249), .X(n21661) );
  nand_x1_sg U45873 ( .A(n21659), .B(n46240), .X(n21658) );
  inv_x1_sg U45874 ( .A(n21867), .X(n55381) );
  inv_x1_sg U45875 ( .A(n21911), .X(n55412) );
  nand_x1_sg U45876 ( .A(n55393), .B(n21907), .X(n21906) );
  nand_x1_sg U45877 ( .A(n55245), .B(n55391), .X(n21907) );
  nand_x2_sg U45878 ( .A(n21855), .B(n21813), .X(n21854) );
  nand_x1_sg U45879 ( .A(n21865), .B(n21866), .X(n21855) );
  nand_x4_sg U45880 ( .A(n21892), .B(n21893), .X(n21851) );
  nand_x1_sg U45881 ( .A(n55414), .B(n21689), .X(n21893) );
  inv_x1_sg U45882 ( .A(n21690), .X(n55414) );
  inv_x1_sg U45883 ( .A(n21836), .X(n55370) );
  nand_x1_sg U45884 ( .A(n55294), .B(n21832), .X(n21835) );
  inv_x1_sg U45885 ( .A(n21728), .X(n55376) );
  nand_x4_sg U45886 ( .A(n55405), .B(n21853), .X(n21812) );
  inv_x1_sg U45887 ( .A(n21854), .X(n55405) );
  nand_x1_sg U45888 ( .A(n21818), .B(n46249), .X(n21817) );
  nand_x1_sg U45889 ( .A(n21812), .B(n21813), .X(n21814) );
  inv_x2_sg U45890 ( .A(n21826), .X(n43844) );
  nor_x1_sg U45891 ( .A(n21830), .B(n21831), .X(n21826) );
  nand_x1_sg U45892 ( .A(n21851), .B(n43096), .X(n21846) );
  nand_x1_sg U45893 ( .A(n21780), .B(n21781), .X(n21779) );
  inv_x1_sg U45894 ( .A(n29860), .X(n50043) );
  inv_x1_sg U45895 ( .A(n30697), .X(n49958) );
  inv_x1_sg U45896 ( .A(n30691), .X(n49910) );
  inv_x1_sg U45897 ( .A(n30685), .X(n49863) );
  inv_x1_sg U45898 ( .A(n31797), .X(n49637) );
  inv_x1_sg U45899 ( .A(n31790), .X(n49591) );
  inv_x1_sg U45900 ( .A(n31783), .X(n49545) );
  inv_x1_sg U45901 ( .A(n31776), .X(n49497) );
  inv_x1_sg U45902 ( .A(n32014), .X(n49502) );
  inv_x1_sg U45903 ( .A(n30622), .X(n49439) );
  inv_x1_sg U45904 ( .A(n31769), .X(n49451) );
  inv_x1_sg U45905 ( .A(n31762), .X(n49406) );
  inv_x1_sg U45906 ( .A(n32001), .X(n49411) );
  inv_x1_sg U45907 ( .A(n30608), .X(n49349) );
  inv_x1_sg U45908 ( .A(n31755), .X(n49361) );
  inv_x1_sg U45909 ( .A(n30601), .X(n49303) );
  inv_x1_sg U45910 ( .A(n31748), .X(n49313) );
  inv_x1_sg U45911 ( .A(n46077), .X(n43780) );
  inv_x1_sg U45912 ( .A(n46049), .X(n43764) );
  inv_x1_sg U45913 ( .A(n46047), .X(n43762) );
  inv_x1_sg U45914 ( .A(n46045), .X(n43760) );
  inv_x1_sg U45915 ( .A(n46043), .X(n43758) );
  nand_x1_sg U45916 ( .A(n8504), .B(n50944), .X(n21993) );
  inv_x1_sg U45917 ( .A(n21994), .X(n50944) );
  nand_x1_sg U45918 ( .A(n8584), .B(n50934), .X(n22603) );
  inv_x1_sg U45919 ( .A(n22604), .X(n50934) );
  nand_x1_sg U45920 ( .A(n8664), .B(n50922), .X(n22574) );
  nand_x1_sg U45921 ( .A(n9370), .B(n22576), .X(n22573) );
  inv_x1_sg U45922 ( .A(n22575), .X(n50922) );
  nand_x1_sg U45923 ( .A(n8744), .B(n50911), .X(n22545) );
  inv_x1_sg U45924 ( .A(n22546), .X(n50911) );
  nand_x1_sg U45925 ( .A(n8504), .B(n21995), .X(n22192) );
  nand_x1_sg U45926 ( .A(n8584), .B(n22605), .X(n22863) );
  inv_x1_sg U45927 ( .A(n22843), .X(n50879) );
  inv_x1_sg U45928 ( .A(n22824), .X(n50869) );
  inv_x1_sg U45929 ( .A(n22830), .X(n50873) );
  inv_x1_sg U45930 ( .A(n23098), .X(n50835) );
  inv_x1_sg U45931 ( .A(n22355), .X(n50855) );
  nand_x1_sg U45932 ( .A(n8505), .B(n22172), .X(n22171) );
  inv_x1_sg U45933 ( .A(n23079), .X(n50825) );
  inv_x1_sg U45934 ( .A(n23085), .X(n50829) );
  inv_x1_sg U45935 ( .A(n23324), .X(n50791) );
  inv_x1_sg U45936 ( .A(n22358), .X(n50811) );
  nand_x1_sg U45937 ( .A(n8506), .B(n22165), .X(n22164) );
  inv_x1_sg U45938 ( .A(n23305), .X(n50781) );
  inv_x1_sg U45939 ( .A(n23311), .X(n50785) );
  nor_x1_sg U45940 ( .A(n9552), .B(n50775), .X(n23328) );
  nor_x1_sg U45941 ( .A(n23289), .B(out_L2[15]), .X(n23288) );
  inv_x1_sg U45942 ( .A(n23529), .X(n50745) );
  inv_x1_sg U45943 ( .A(n22361), .X(n50763) );
  nand_x1_sg U45944 ( .A(n8507), .B(n22158), .X(n22157) );
  inv_x1_sg U45945 ( .A(n23510), .X(n50735) );
  inv_x1_sg U45946 ( .A(n23516), .X(n50739) );
  inv_x1_sg U45947 ( .A(n23719), .X(n50699) );
  inv_x1_sg U45948 ( .A(n22364), .X(n50716) );
  nand_x1_sg U45949 ( .A(n8508), .B(n22151), .X(n22150) );
  inv_x1_sg U45950 ( .A(n23347), .X(n50725) );
  nand_x1_sg U45951 ( .A(n8588), .B(n23019), .X(n23018) );
  inv_x1_sg U45952 ( .A(n23700), .X(n50689) );
  inv_x1_sg U45953 ( .A(n23706), .X(n50693) );
  nor_x1_sg U45954 ( .A(n9648), .B(n50681), .X(n23723) );
  nor_x1_sg U45955 ( .A(n23684), .B(out_L2[13]), .X(n23683) );
  inv_x1_sg U45956 ( .A(n23890), .X(n50682) );
  inv_x1_sg U45957 ( .A(n22367), .X(n50668) );
  nand_x1_sg U45958 ( .A(n8509), .B(n22144), .X(n22143) );
  inv_x1_sg U45959 ( .A(n23350), .X(n50677) );
  nand_x1_sg U45960 ( .A(n8589), .B(n23012), .X(n23011) );
  inv_x1_sg U45961 ( .A(n23871), .X(n50644) );
  inv_x1_sg U45962 ( .A(n23877), .X(n50648) );
  inv_x1_sg U45963 ( .A(n22370), .X(n50621) );
  inv_x1_sg U45964 ( .A(n23353), .X(n50630) );
  nand_x1_sg U45965 ( .A(n8590), .B(n23005), .X(n23004) );
  nand_x1_sg U45966 ( .A(n8510), .B(n22137), .X(n22136) );
  inv_x1_sg U45967 ( .A(n23893), .X(n50636) );
  inv_x1_sg U45968 ( .A(n22639), .X(n50623) );
  inv_x1_sg U45969 ( .A(n24024), .X(n50598) );
  inv_x1_sg U45970 ( .A(n24030), .X(n50602) );
  nor_x1_sg U45971 ( .A(n24008), .B(out_L2[11]), .X(n24007) );
  inv_x1_sg U45972 ( .A(n23896), .X(n50586) );
  inv_x1_sg U45973 ( .A(n22373), .X(n50572) );
  nand_x1_sg U45974 ( .A(n8511), .B(n22130), .X(n22129) );
  inv_x1_sg U45975 ( .A(n23356), .X(n50581) );
  nand_x1_sg U45976 ( .A(n8591), .B(n22998), .X(n22997) );
  inv_x1_sg U45977 ( .A(n24168), .X(n50552) );
  inv_x1_sg U45978 ( .A(n24174), .X(n50590) );
  inv_x1_sg U45979 ( .A(n23899), .X(n50540) );
  inv_x1_sg U45980 ( .A(n22376), .X(n50525) );
  nand_x1_sg U45981 ( .A(n8512), .B(n22123), .X(n22122) );
  inv_x1_sg U45982 ( .A(n23359), .X(n50534) );
  nand_x1_sg U45983 ( .A(n8592), .B(n22991), .X(n22990) );
  inv_x1_sg U45984 ( .A(n24284), .X(n50546) );
  nor_x1_sg U45985 ( .A(n24268), .B(out_L2[9]), .X(n24267) );
  inv_x1_sg U45986 ( .A(n23902), .X(n50492) );
  inv_x1_sg U45987 ( .A(n22379), .X(n50478) );
  nand_x1_sg U45988 ( .A(n8513), .B(n22116), .X(n22115) );
  inv_x1_sg U45989 ( .A(n23362), .X(n50487) );
  nand_x1_sg U45990 ( .A(n8593), .B(n22984), .X(n22983) );
  inv_x1_sg U45991 ( .A(n24287), .X(n50499) );
  inv_x1_sg U45992 ( .A(n23905), .X(n50446) );
  inv_x1_sg U45993 ( .A(n22382), .X(n50432) );
  nand_x1_sg U45994 ( .A(n8514), .B(n22109), .X(n22108) );
  inv_x1_sg U45995 ( .A(n23365), .X(n50441) );
  nand_x1_sg U45996 ( .A(n8594), .B(n22977), .X(n22976) );
  inv_x1_sg U45997 ( .A(n24290), .X(n50453) );
  inv_x1_sg U45998 ( .A(n24355), .X(n50409) );
  inv_x1_sg U45999 ( .A(n23908), .X(n50400) );
  inv_x1_sg U46000 ( .A(n22385), .X(n50385) );
  nand_x1_sg U46001 ( .A(n8515), .B(n22102), .X(n22101) );
  inv_x1_sg U46002 ( .A(n23368), .X(n50394) );
  nand_x1_sg U46003 ( .A(n8595), .B(n22970), .X(n22969) );
  inv_x1_sg U46004 ( .A(n24293), .X(n50407) );
  nor_x1_sg U46005 ( .A(n24452), .B(out_L2[6]), .X(n24451) );
  inv_x2_sg U46006 ( .A(n24450), .X(n44300) );
  nor_x1_sg U46007 ( .A(n40851), .B(n50363), .X(n24450) );
  inv_x1_sg U46008 ( .A(n23371), .X(n50347) );
  inv_x1_sg U46009 ( .A(n23911), .X(n50352) );
  inv_x1_sg U46010 ( .A(n22657), .X(n50340) );
  inv_x1_sg U46011 ( .A(n22388), .X(n50338) );
  nand_x1_sg U46012 ( .A(n8516), .B(n22095), .X(n22094) );
  inv_x1_sg U46013 ( .A(n24296), .X(n50359) );
  inv_x1_sg U46014 ( .A(n24342), .X(n50315) );
  inv_x1_sg U46015 ( .A(n23914), .X(n50306) );
  inv_x1_sg U46016 ( .A(n22391), .X(n50292) );
  nand_x1_sg U46017 ( .A(n8517), .B(n22088), .X(n22087) );
  inv_x1_sg U46018 ( .A(n23374), .X(n50301) );
  nand_x1_sg U46019 ( .A(n8597), .B(n22956), .X(n22955) );
  inv_x1_sg U46020 ( .A(n24299), .X(n50313) );
  inv_x1_sg U46021 ( .A(n23377), .X(n50255) );
  inv_x1_sg U46022 ( .A(n22663), .X(n50248) );
  inv_x1_sg U46023 ( .A(n22394), .X(n50246) );
  nand_x1_sg U46024 ( .A(n8518), .B(n22081), .X(n22080) );
  inv_x1_sg U46025 ( .A(n23917), .X(n50261) );
  inv_x1_sg U46026 ( .A(n24329), .X(n50225) );
  inv_x1_sg U46027 ( .A(n24302), .X(n50268) );
  inv_x1_sg U46028 ( .A(n23380), .X(n50211) );
  inv_x1_sg U46029 ( .A(n22666), .X(n50204) );
  inv_x1_sg U46030 ( .A(n22397), .X(n50202) );
  nand_x1_sg U46031 ( .A(n8519), .B(n22074), .X(n22073) );
  inv_x1_sg U46032 ( .A(n23920), .X(n50216) );
  inv_x1_sg U46033 ( .A(n23595), .X(n50167) );
  inv_x1_sg U46034 ( .A(n24323), .X(n50176) );
  inv_x1_sg U46035 ( .A(n24305), .X(n50223) );
  nand_x1_sg U46036 ( .A(n8520), .B(n22067), .X(n22066) );
  nand_x2_sg U46037 ( .A(n23388), .B(n23389), .X(n23387) );
  nand_x1_sg U46038 ( .A(n10514), .B(n51306), .X(n10513) );
  inv_x1_sg U46039 ( .A(n10517), .X(n51324) );
  nand_x1_sg U46040 ( .A(n51293), .B(n46572), .X(n10463) );
  nor_x1_sg U46041 ( .A(n10545), .B(n51307), .X(n10544) );
  nand_x4_sg U46042 ( .A(n46567), .B(n51293), .X(n10537) );
  nor_x1_sg U46043 ( .A(n46573), .B(n10492), .X(n10491) );
  inv_x1_sg U46044 ( .A(n10579), .X(n51346) );
  nand_x1_sg U46045 ( .A(n10652), .B(n46557), .X(n10651) );
  inv_x1_sg U46046 ( .A(n10638), .X(n51335) );
  nand_x4_sg U46047 ( .A(n46567), .B(n51334), .X(n10638) );
  inv_x1_sg U46048 ( .A(n10686), .X(n51371) );
  inv_x1_sg U46049 ( .A(n10752), .X(n51436) );
  inv_x2_sg U46050 ( .A(n10746), .X(n44466) );
  nor_x1_sg U46051 ( .A(n51419), .B(n10748), .X(n10746) );
  inv_x2_sg U46052 ( .A(n10647), .X(n44081) );
  nand_x1_sg U46053 ( .A(n10605), .B(n10604), .X(n10647) );
  inv_x1_sg U46054 ( .A(n10709), .X(n51422) );
  inv_x1_sg U46055 ( .A(n10812), .X(n51448) );
  nand_x4_sg U46056 ( .A(n10777), .B(n10778), .X(n10709) );
  nand_x1_sg U46057 ( .A(n51306), .B(n51421), .X(n10778) );
  nand_x4_sg U46058 ( .A(n11014), .B(n11015), .X(n10974) );
  nand_x1_sg U46059 ( .A(n51488), .B(n10818), .X(n11015) );
  nand_x2_sg U46060 ( .A(n10978), .B(n10937), .X(n10977) );
  nand_x1_sg U46061 ( .A(n10986), .B(n10987), .X(n10978) );
  inv_x1_sg U46062 ( .A(n10977), .X(n51478) );
  nand_x1_sg U46063 ( .A(n11023), .B(n51487), .X(n11022) );
  inv_x1_sg U46064 ( .A(n11024), .X(n51487) );
  nand_x4_sg U46065 ( .A(n11016), .B(n11017), .X(n10818) );
  nand_x1_sg U46066 ( .A(n11018), .B(n51453), .X(n11017) );
  nand_x1_sg U46067 ( .A(n10992), .B(n51415), .X(n11016) );
  nand_x1_sg U46068 ( .A(n10800), .B(n10802), .X(n10801) );
  nand_x1_sg U46069 ( .A(n51455), .B(n10840), .X(n10839) );
  inv_x1_sg U46070 ( .A(n10836), .X(n51455) );
  inv_x2_sg U46071 ( .A(n10878), .X(n44378) );
  nor_x1_sg U46072 ( .A(n11041), .B(n11042), .X(n10878) );
  nand_x1_sg U46073 ( .A(n10901), .B(n51293), .X(n10896) );
  nand_x1_sg U46074 ( .A(n10922), .B(n46567), .X(n10921) );
  nand_x1_sg U46075 ( .A(n10966), .B(n46557), .X(n10965) );
  nand_x1_sg U46076 ( .A(n10935), .B(n10936), .X(n10934) );
  nand_x1_sg U46077 ( .A(n11293), .B(n11265), .X(n11292) );
  inv_x1_sg U46078 ( .A(n11297), .X(n51599) );
  nand_x1_sg U46079 ( .A(n11318), .B(n51598), .X(n11317) );
  nand_x1_sg U46080 ( .A(n11265), .B(n46551), .X(n11264) );
  nand_x1_sg U46081 ( .A(n11390), .B(n51630), .X(n11389) );
  nand_x4_sg U46082 ( .A(n11352), .B(n11353), .X(n11339) );
  nand_x1_sg U46083 ( .A(n51581), .B(n51625), .X(n11352) );
  nand_x1_sg U46084 ( .A(n11354), .B(n11267), .X(n11353) );
  inv_x1_sg U46085 ( .A(n11354), .X(n51625) );
  nand_x1_sg U46086 ( .A(n11431), .B(n51630), .X(n11430) );
  inv_x1_sg U46087 ( .A(n11417), .X(n51615) );
  inv_x1_sg U46088 ( .A(n11514), .X(n51674) );
  inv_x1_sg U46089 ( .A(n11443), .X(n51676) );
  inv_x2_sg U46090 ( .A(n11528), .X(n44149) );
  nor_x1_sg U46091 ( .A(n11529), .B(n11530), .X(n11528) );
  inv_x2_sg U46092 ( .A(n11527), .X(n45412) );
  nor_x1_sg U46093 ( .A(n51718), .B(n11533), .X(n11527) );
  nand_x4_sg U46094 ( .A(n11484), .B(n11485), .X(n11467) );
  nand_x1_sg U46095 ( .A(n51695), .B(n11265), .X(n11484) );
  nand_x1_sg U46096 ( .A(n46533), .B(n11486), .X(n11485) );
  inv_x1_sg U46097 ( .A(n11486), .X(n51695) );
  inv_x1_sg U46098 ( .A(n11592), .X(n51727) );
  nand_x1_sg U46099 ( .A(n11594), .B(n11593), .X(n11591) );
  nand_x1_sg U46100 ( .A(n51710), .B(n11584), .X(n11583) );
  nand_x1_sg U46101 ( .A(n51617), .B(n51641), .X(n11584) );
  nand_x1_sg U46102 ( .A(n51763), .B(n11761), .X(n11759) );
  inv_x1_sg U46103 ( .A(n11760), .X(n51763) );
  nand_x1_sg U46104 ( .A(n51768), .B(n41867), .X(n11755) );
  nand_x1_sg U46105 ( .A(n41868), .B(n11758), .X(n11756) );
  inv_x1_sg U46106 ( .A(n11758), .X(n51768) );
  inv_x2_sg U46107 ( .A(n11658), .X(n44101) );
  nor_x1_sg U46108 ( .A(n11825), .B(n11826), .X(n11658) );
  nand_x1_sg U46109 ( .A(n51598), .B(n11594), .X(n11633) );
  nand_x1_sg U46110 ( .A(n51732), .B(n11621), .X(n11620) );
  nand_x1_sg U46111 ( .A(n11718), .B(n11719), .X(n11717) );
  nand_x1_sg U46112 ( .A(n11750), .B(n51598), .X(n11749) );
  inv_x1_sg U46113 ( .A(n12077), .X(n51880) );
  nor_x1_sg U46114 ( .A(n46528), .B(n12045), .X(n12044) );
  nand_x1_sg U46115 ( .A(n12170), .B(n51911), .X(n12169) );
  nand_x4_sg U46116 ( .A(n12132), .B(n12133), .X(n12119) );
  nand_x1_sg U46117 ( .A(n51899), .B(n12046), .X(n12133) );
  nand_x1_sg U46118 ( .A(n51862), .B(n12134), .X(n12132) );
  nand_x1_sg U46119 ( .A(n12211), .B(n51911), .X(n12210) );
  inv_x1_sg U46120 ( .A(n12197), .X(n51897) );
  nand_x4_sg U46121 ( .A(n51826), .B(n51896), .X(n12197) );
  inv_x1_sg U46122 ( .A(n12247), .X(n51927) );
  inv_x1_sg U46123 ( .A(n12223), .X(n51957) );
  nand_x1_sg U46124 ( .A(n51966), .B(n51948), .X(n12297) );
  inv_x1_sg U46125 ( .A(n12298), .X(n51966) );
  inv_x1_sg U46126 ( .A(n12308), .X(n51997) );
  inv_x1_sg U46127 ( .A(n12270), .X(n51977) );
  inv_x1_sg U46128 ( .A(n12373), .X(n52005) );
  nand_x1_sg U46129 ( .A(n12375), .B(n12374), .X(n12372) );
  nand_x1_sg U46130 ( .A(n46513), .B(n51976), .X(n12340) );
  nand_x1_sg U46131 ( .A(n12363), .B(n12365), .X(n12364) );
  nand_x1_sg U46132 ( .A(n51898), .B(n51922), .X(n12365) );
  inv_x1_sg U46133 ( .A(n12556), .X(n51945) );
  nand_x4_sg U46134 ( .A(n42366), .B(n12557), .X(n12537) );
  inv_x1_sg U46135 ( .A(n12536), .X(n52048) );
  nand_x4_sg U46136 ( .A(n12573), .B(n12574), .X(n12536) );
  nand_x1_sg U46137 ( .A(n52047), .B(n40532), .X(n12574) );
  inv_x1_sg U46138 ( .A(n12310), .X(n51989) );
  nand_x4_sg U46139 ( .A(n12313), .B(n51996), .X(n12308) );
  inv_x1_sg U46140 ( .A(n12314), .X(n51996) );
  nand_x1_sg U46141 ( .A(n12316), .B(n12315), .X(n12313) );
  nand_x1_sg U46142 ( .A(n52063), .B(n51896), .X(n12605) );
  nand_x1_sg U46143 ( .A(n51879), .B(n12375), .X(n12414) );
  nand_x1_sg U46144 ( .A(n52010), .B(n12402), .X(n12401) );
  nand_x1_sg U46145 ( .A(n12498), .B(n12499), .X(n12497) );
  nand_x1_sg U46146 ( .A(n12530), .B(n51911), .X(n12529) );
  inv_x1_sg U46147 ( .A(n12858), .X(n52157) );
  nand_x1_sg U46148 ( .A(n12879), .B(n52156), .X(n12878) );
  nand_x1_sg U46149 ( .A(n12951), .B(n52187), .X(n12950) );
  nand_x4_sg U46150 ( .A(n12913), .B(n12914), .X(n12900) );
  nand_x1_sg U46151 ( .A(n52139), .B(n12915), .X(n12913) );
  nand_x1_sg U46152 ( .A(n52176), .B(n12828), .X(n12914) );
  nand_x1_sg U46153 ( .A(n12992), .B(n52187), .X(n12991) );
  inv_x1_sg U46154 ( .A(n12978), .X(n52173) );
  inv_x1_sg U46155 ( .A(n13075), .X(n52230) );
  inv_x1_sg U46156 ( .A(n13004), .X(n52232) );
  inv_x2_sg U46157 ( .A(n13089), .X(n44147) );
  nor_x1_sg U46158 ( .A(n13090), .B(n13091), .X(n13089) );
  inv_x2_sg U46159 ( .A(n13088), .X(n45410) );
  nor_x1_sg U46160 ( .A(n52272), .B(n13094), .X(n13088) );
  nand_x4_sg U46161 ( .A(n13045), .B(n13046), .X(n13028) );
  nand_x1_sg U46162 ( .A(n52251), .B(n12826), .X(n13045) );
  nand_x1_sg U46163 ( .A(n46489), .B(n13047), .X(n13046) );
  inv_x1_sg U46164 ( .A(n13153), .X(n52283) );
  nand_x1_sg U46165 ( .A(n13155), .B(n13154), .X(n13152) );
  nand_x1_sg U46166 ( .A(n52266), .B(n13145), .X(n13144) );
  nand_x1_sg U46167 ( .A(n52175), .B(n52197), .X(n13145) );
  inv_x1_sg U46168 ( .A(n13337), .X(n52220) );
  nand_x1_sg U46169 ( .A(n52340), .B(n46488), .X(n13387) );
  inv_x1_sg U46170 ( .A(n13197), .X(n52282) );
  nand_x1_sg U46171 ( .A(n52281), .B(n13182), .X(n13181) );
  nand_x1_sg U46172 ( .A(n13279), .B(n13280), .X(n13278) );
  nand_x1_sg U46173 ( .A(n13311), .B(n52156), .X(n13310) );
  inv_x1_sg U46174 ( .A(n13638), .X(n52431) );
  nand_x4_sg U46175 ( .A(n13657), .B(n13658), .X(n13624) );
  nand_x1_sg U46176 ( .A(n13660), .B(n13661), .X(n13657) );
  nand_x1_sg U46177 ( .A(n13659), .B(n52430), .X(n13658) );
  nand_x1_sg U46178 ( .A(n52430), .B(n46481), .X(n13661) );
  nor_x1_sg U46179 ( .A(n46485), .B(n13606), .X(n13605) );
  nand_x1_sg U46180 ( .A(n13731), .B(n52463), .X(n13730) );
  nand_x4_sg U46181 ( .A(n13693), .B(n13694), .X(n13680) );
  nand_x1_sg U46182 ( .A(n52451), .B(n13607), .X(n13694) );
  nand_x1_sg U46183 ( .A(n52414), .B(n13695), .X(n13693) );
  nand_x1_sg U46184 ( .A(n13772), .B(n52463), .X(n13771) );
  inv_x1_sg U46185 ( .A(n13758), .X(n52448) );
  inv_x1_sg U46186 ( .A(n13784), .X(n52509) );
  nand_x1_sg U46187 ( .A(n52517), .B(n52500), .X(n13858) );
  inv_x1_sg U46188 ( .A(n13859), .X(n52517) );
  inv_x2_sg U46189 ( .A(n13869), .X(n44145) );
  nor_x1_sg U46190 ( .A(n13870), .B(n13871), .X(n13869) );
  inv_x2_sg U46191 ( .A(n13868), .X(n45408) );
  nor_x1_sg U46192 ( .A(n52547), .B(n13874), .X(n13868) );
  nand_x4_sg U46193 ( .A(n13825), .B(n13826), .X(n13808) );
  nand_x1_sg U46194 ( .A(n52527), .B(n46468), .X(n13825) );
  nand_x1_sg U46195 ( .A(n13604), .B(n13827), .X(n13826) );
  inv_x1_sg U46196 ( .A(n13827), .X(n52527) );
  inv_x1_sg U46197 ( .A(n13933), .X(n52558) );
  nand_x1_sg U46198 ( .A(n13935), .B(n13934), .X(n13932) );
  nand_x1_sg U46199 ( .A(n52542), .B(n13925), .X(n13924) );
  nand_x1_sg U46200 ( .A(n52450), .B(n52474), .X(n13925) );
  inv_x1_sg U46201 ( .A(n14117), .X(n52497) );
  nand_x4_sg U46202 ( .A(n42268), .B(n14101), .X(n14060) );
  nand_x1_sg U46203 ( .A(n52615), .B(n52447), .X(n14167) );
  inv_x1_sg U46204 ( .A(n13977), .X(n52557) );
  nand_x1_sg U46205 ( .A(n52556), .B(n13962), .X(n13961) );
  nand_x1_sg U46206 ( .A(n14059), .B(n14060), .X(n14058) );
  nand_x1_sg U46207 ( .A(n14091), .B(n52463), .X(n14090) );
  inv_x1_sg U46208 ( .A(n14409), .X(n52714) );
  nand_x1_sg U46209 ( .A(n14406), .B(n52695), .X(n14405) );
  nand_x1_sg U46210 ( .A(n52683), .B(n14174), .X(n14355) );
  nor_x1_sg U46211 ( .A(n14438), .B(n52696), .X(n14437) );
  nor_x1_sg U46212 ( .A(n14413), .B(n14414), .X(n14412) );
  nand_x4_sg U46213 ( .A(n52670), .B(n46450), .X(n14430) );
  nand_x4_sg U46214 ( .A(n52683), .B(n52655), .X(n14429) );
  nand_x4_sg U46215 ( .A(n52750), .B(n14503), .X(n14443) );
  inv_x1_sg U46216 ( .A(n14505), .X(n52750) );
  nand_x1_sg U46217 ( .A(n14504), .B(n52749), .X(n14503) );
  inv_x1_sg U46218 ( .A(n14471), .X(n52736) );
  inv_x1_sg U46219 ( .A(n14644), .X(n52825) );
  inv_x2_sg U46220 ( .A(n14638), .X(n44446) );
  nor_x1_sg U46221 ( .A(n52807), .B(n14640), .X(n14638) );
  inv_x1_sg U46222 ( .A(n14530), .X(n52724) );
  nand_x4_sg U46223 ( .A(n46443), .B(n52655), .X(n14530) );
  inv_x1_sg U46224 ( .A(n14578), .X(n52759) );
  inv_x1_sg U46225 ( .A(n14555), .X(n52788) );
  inv_x1_sg U46226 ( .A(n14630), .X(n52797) );
  inv_x1_sg U46227 ( .A(n14601), .X(n52812) );
  nand_x4_sg U46228 ( .A(n46443), .B(n52670), .X(n14692) );
  nand_x1_sg U46229 ( .A(n14705), .B(n14704), .X(n14706) );
  nand_x1_sg U46230 ( .A(n14693), .B(n14695), .X(n14694) );
  nand_x4_sg U46231 ( .A(n14669), .B(n14670), .X(n14601) );
  nand_x1_sg U46232 ( .A(n52695), .B(n52811), .X(n14670) );
  inv_x1_sg U46233 ( .A(n14709), .X(n52881) );
  nand_x1_sg U46234 ( .A(n14710), .B(n14711), .X(n14708) );
  inv_x2_sg U46235 ( .A(n14771), .X(n44214) );
  nor_x1_sg U46236 ( .A(n14937), .B(n14938), .X(n14771) );
  nand_x1_sg U46237 ( .A(n52707), .B(n14705), .X(n14745) );
  nand_x1_sg U46238 ( .A(n52832), .B(n14733), .X(n14732) );
  nand_x1_sg U46239 ( .A(n14830), .B(n14831), .X(n14829) );
  nand_x1_sg U46240 ( .A(n14862), .B(n52707), .X(n14861) );
  inv_x1_sg U46241 ( .A(n14774), .X(n45448) );
  inv_x1_sg U46242 ( .A(n15191), .X(n52991) );
  nand_x1_sg U46243 ( .A(n15212), .B(n52990), .X(n15211) );
  nand_x1_sg U46244 ( .A(n15284), .B(n53021), .X(n15283) );
  nand_x4_sg U46245 ( .A(n15246), .B(n15247), .X(n15233) );
  nand_x1_sg U46246 ( .A(n52973), .B(n15248), .X(n15246) );
  nand_x1_sg U46247 ( .A(n53010), .B(n15161), .X(n15247) );
  nand_x1_sg U46248 ( .A(n15325), .B(n53021), .X(n15324) );
  inv_x1_sg U46249 ( .A(n15311), .X(n53007) );
  inv_x1_sg U46250 ( .A(n15408), .X(n53064) );
  inv_x1_sg U46251 ( .A(n15337), .X(n53066) );
  inv_x2_sg U46252 ( .A(n15422), .X(n44143) );
  nor_x1_sg U46253 ( .A(n15423), .B(n15424), .X(n15422) );
  inv_x2_sg U46254 ( .A(n15421), .X(n45406) );
  nor_x1_sg U46255 ( .A(n53106), .B(n15427), .X(n15421) );
  nand_x4_sg U46256 ( .A(n15378), .B(n15379), .X(n15361) );
  nand_x1_sg U46257 ( .A(n53085), .B(n15159), .X(n15378) );
  nand_x1_sg U46258 ( .A(n46421), .B(n15380), .X(n15379) );
  inv_x1_sg U46259 ( .A(n15486), .X(n53117) );
  nand_x1_sg U46260 ( .A(n15488), .B(n15487), .X(n15485) );
  nand_x1_sg U46261 ( .A(n53100), .B(n15478), .X(n15477) );
  nand_x1_sg U46262 ( .A(n53009), .B(n53031), .X(n15478) );
  inv_x1_sg U46263 ( .A(n15670), .X(n53054) );
  nand_x1_sg U46264 ( .A(n53174), .B(n46420), .X(n15720) );
  inv_x1_sg U46265 ( .A(n15530), .X(n53116) );
  nand_x1_sg U46266 ( .A(n53115), .B(n15515), .X(n15514) );
  nand_x1_sg U46267 ( .A(n15612), .B(n15613), .X(n15611) );
  nand_x1_sg U46268 ( .A(n15644), .B(n52990), .X(n15643) );
  inv_x1_sg U46269 ( .A(n15972), .X(n53267) );
  nand_x1_sg U46270 ( .A(n15968), .B(n53253), .X(n15967) );
  nand_x4_sg U46271 ( .A(n16027), .B(n16028), .X(n16014) );
  nand_x1_sg U46272 ( .A(n53248), .B(n53292), .X(n16027) );
  nand_x1_sg U46273 ( .A(n16029), .B(n15941), .X(n16028) );
  inv_x1_sg U46274 ( .A(n16029), .X(n53292) );
  inv_x1_sg U46275 ( .A(n16092), .X(n53283) );
  nand_x4_sg U46276 ( .A(n53214), .B(n53282), .X(n16092) );
  inv_x1_sg U46277 ( .A(n16142), .X(n53315) );
  inv_x1_sg U46278 ( .A(n16118), .X(n53345) );
  nand_x1_sg U46279 ( .A(n53355), .B(n53336), .X(n16192) );
  inv_x1_sg U46280 ( .A(n16193), .X(n53355) );
  inv_x1_sg U46281 ( .A(n16203), .X(n53386) );
  inv_x1_sg U46282 ( .A(n16165), .X(n53366) );
  nand_x1_sg U46283 ( .A(n16269), .B(n16268), .X(n16270) );
  nand_x4_sg U46284 ( .A(n16234), .B(n16235), .X(n16165) );
  nand_x1_sg U46285 ( .A(n53253), .B(n53365), .X(n16235) );
  nand_x4_sg U46286 ( .A(n16473), .B(n16474), .X(n16432) );
  nand_x1_sg U46287 ( .A(n53437), .B(n42119), .X(n16474) );
  nand_x2_sg U46288 ( .A(n16436), .B(n16395), .X(n16435) );
  nand_x1_sg U46289 ( .A(n16445), .B(n16446), .X(n16436) );
  inv_x1_sg U46290 ( .A(n16459), .X(n53333) );
  inv_x1_sg U46291 ( .A(n16435), .X(n53427) );
  nand_x1_sg U46292 ( .A(n16258), .B(n16260), .X(n16259) );
  nand_x1_sg U46293 ( .A(n53284), .B(n53309), .X(n16260) );
  inv_x1_sg U46294 ( .A(n16205), .X(n53377) );
  nand_x4_sg U46295 ( .A(n16208), .B(n53385), .X(n16203) );
  inv_x1_sg U46296 ( .A(n16209), .X(n53385) );
  nand_x1_sg U46297 ( .A(n16211), .B(n16210), .X(n16208) );
  nand_x1_sg U46298 ( .A(n53266), .B(n16269), .X(n16309) );
  nand_x1_sg U46299 ( .A(n53402), .B(n16297), .X(n16296) );
  nand_x1_sg U46300 ( .A(n53451), .B(n53282), .X(n16503) );
  nand_x1_sg U46301 ( .A(n16361), .B(n16362), .X(n16360) );
  nand_x1_sg U46302 ( .A(n16424), .B(n53266), .X(n16423) );
  nand_x1_sg U46303 ( .A(n16393), .B(n16394), .X(n16392) );
  inv_x1_sg U46304 ( .A(n16757), .X(n53549) );
  nand_x1_sg U46305 ( .A(n16778), .B(n53548), .X(n16777) );
  nand_x1_sg U46306 ( .A(n16850), .B(n53579), .X(n16849) );
  nand_x4_sg U46307 ( .A(n16812), .B(n16813), .X(n16799) );
  nand_x1_sg U46308 ( .A(n53531), .B(n16814), .X(n16812) );
  nand_x1_sg U46309 ( .A(n53568), .B(n16727), .X(n16813) );
  nand_x1_sg U46310 ( .A(n16891), .B(n53579), .X(n16890) );
  inv_x1_sg U46311 ( .A(n16877), .X(n53565) );
  inv_x1_sg U46312 ( .A(n16974), .X(n53622) );
  inv_x1_sg U46313 ( .A(n16903), .X(n53624) );
  inv_x2_sg U46314 ( .A(n16988), .X(n44141) );
  nor_x1_sg U46315 ( .A(n16989), .B(n16990), .X(n16988) );
  inv_x2_sg U46316 ( .A(n16987), .X(n45404) );
  nor_x1_sg U46317 ( .A(n53664), .B(n16993), .X(n16987) );
  nand_x4_sg U46318 ( .A(n16944), .B(n16945), .X(n16927) );
  nand_x1_sg U46319 ( .A(n53643), .B(n16725), .X(n16944) );
  nand_x1_sg U46320 ( .A(n46377), .B(n16946), .X(n16945) );
  inv_x1_sg U46321 ( .A(n17052), .X(n53675) );
  nand_x1_sg U46322 ( .A(n17054), .B(n17053), .X(n17051) );
  nand_x1_sg U46323 ( .A(n53658), .B(n17044), .X(n17043) );
  nand_x1_sg U46324 ( .A(n53567), .B(n53589), .X(n17044) );
  inv_x1_sg U46325 ( .A(n17236), .X(n53612) );
  nand_x1_sg U46326 ( .A(n53732), .B(n46376), .X(n17286) );
  inv_x1_sg U46327 ( .A(n17096), .X(n53674) );
  nand_x1_sg U46328 ( .A(n53673), .B(n17081), .X(n17080) );
  nand_x1_sg U46329 ( .A(n17178), .B(n17179), .X(n17177) );
  nand_x1_sg U46330 ( .A(n17210), .B(n53548), .X(n17209) );
  nand_x1_sg U46331 ( .A(n17527), .B(n43864), .X(n17526) );
  nand_x1_sg U46332 ( .A(n53808), .B(n17531), .X(n17530) );
  nand_x1_sg U46333 ( .A(n53828), .B(n17492), .X(n17529) );
  inv_x1_sg U46334 ( .A(n17531), .X(n53828) );
  nand_x1_sg U46335 ( .A(n53802), .B(n46368), .X(n17478) );
  nor_x1_sg U46336 ( .A(n17557), .B(n53823), .X(n17556) );
  nand_x4_sg U46337 ( .A(n17585), .B(n17586), .X(n17533) );
  nand_x1_sg U46338 ( .A(n53809), .B(n17505), .X(n17585) );
  nand_x1_sg U46339 ( .A(n53796), .B(n17549), .X(n17586) );
  nand_x4_sg U46340 ( .A(n46356), .B(n46372), .X(n17534) );
  nand_x4_sg U46341 ( .A(n53802), .B(n46363), .X(n17549) );
  nand_x1_sg U46342 ( .A(n46358), .B(n46372), .X(n17502) );
  nand_x4_sg U46343 ( .A(n53870), .B(n17624), .X(n17563) );
  inv_x1_sg U46344 ( .A(n17626), .X(n53870) );
  nand_x1_sg U46345 ( .A(n17625), .B(n53869), .X(n17624) );
  inv_x1_sg U46346 ( .A(n17591), .X(n53856) );
  inv_x1_sg U46347 ( .A(n17765), .X(n53945) );
  inv_x2_sg U46348 ( .A(n17759), .X(n44444) );
  nor_x1_sg U46349 ( .A(n53927), .B(n17761), .X(n17759) );
  inv_x1_sg U46350 ( .A(n17651), .X(n53844) );
  inv_x1_sg U46351 ( .A(n17699), .X(n53879) );
  inv_x1_sg U46352 ( .A(n17676), .X(n53908) );
  inv_x1_sg U46353 ( .A(n17751), .X(n53918) );
  inv_x1_sg U46354 ( .A(n17722), .X(n53932) );
  nand_x4_sg U46355 ( .A(n46360), .B(n46356), .X(n17813) );
  nand_x1_sg U46356 ( .A(n17826), .B(n17825), .X(n17827) );
  nand_x1_sg U46357 ( .A(n17814), .B(n17816), .X(n17815) );
  nand_x1_sg U46358 ( .A(n53846), .B(n53867), .X(n17816) );
  nand_x4_sg U46359 ( .A(n17790), .B(n17791), .X(n17722) );
  nand_x1_sg U46360 ( .A(n46358), .B(n53931), .X(n17791) );
  inv_x1_sg U46361 ( .A(n17830), .X(n54001) );
  nand_x1_sg U46362 ( .A(n17831), .B(n17832), .X(n17829) );
  inv_x2_sg U46363 ( .A(n17892), .X(n44037) );
  nor_x1_sg U46364 ( .A(n18058), .B(n18059), .X(n17892) );
  nand_x1_sg U46365 ( .A(n53827), .B(n17826), .X(n17866) );
  nand_x1_sg U46366 ( .A(n53952), .B(n17854), .X(n17853) );
  nand_x1_sg U46367 ( .A(n17951), .B(n17952), .X(n17950) );
  nand_x1_sg U46368 ( .A(n17983), .B(n53827), .X(n17982) );
  inv_x1_sg U46369 ( .A(n17895), .X(n45444) );
  nand_x1_sg U46370 ( .A(n54084), .B(n18065), .X(n18245) );
  inv_x1_sg U46371 ( .A(n18299), .X(n54115) );
  nand_x1_sg U46372 ( .A(n18296), .B(n43811), .X(n18295) );
  nand_x4_sg U46373 ( .A(n54084), .B(n46343), .X(n18320) );
  nand_x4_sg U46374 ( .A(n54070), .B(n46339), .X(n18319) );
  inv_x1_sg U46375 ( .A(n18361), .X(n54136) );
  nand_x1_sg U46376 ( .A(n18434), .B(n46329), .X(n18433) );
  inv_x1_sg U46377 ( .A(n18420), .X(n54125) );
  nand_x4_sg U46378 ( .A(n54124), .B(n46343), .X(n18420) );
  inv_x1_sg U46379 ( .A(n18533), .X(n54230) );
  inv_x2_sg U46380 ( .A(n18527), .X(n44210) );
  nor_x1_sg U46381 ( .A(n54223), .B(n18529), .X(n18527) );
  inv_x1_sg U46382 ( .A(n18514), .X(n54185) );
  inv_x2_sg U46383 ( .A(n18482), .X(n44718) );
  inv_x1_sg U46384 ( .A(n18592), .X(n54241) );
  nand_x1_sg U46385 ( .A(n18594), .B(n18593), .X(n18591) );
  nand_x1_sg U46386 ( .A(n18810), .B(n54278), .X(n18809) );
  inv_x1_sg U46387 ( .A(n18811), .X(n54278) );
  nand_x1_sg U46388 ( .A(n18580), .B(n18582), .X(n18581) );
  nand_x1_sg U46389 ( .A(n54275), .B(n18763), .X(n18761) );
  inv_x1_sg U46390 ( .A(n18762), .X(n54275) );
  nand_x1_sg U46391 ( .A(n54280), .B(n42600), .X(n18757) );
  nand_x1_sg U46392 ( .A(n42601), .B(n18760), .X(n18758) );
  inv_x1_sg U46393 ( .A(n18760), .X(n54280) );
  nand_x1_sg U46394 ( .A(n18657), .B(n18656), .X(n18658) );
  inv_x2_sg U46395 ( .A(n18661), .X(n44212) );
  nor_x1_sg U46396 ( .A(n18830), .B(n18831), .X(n18661) );
  nand_x1_sg U46397 ( .A(n54109), .B(n18594), .X(n18633) );
  nand_x1_sg U46398 ( .A(n54247), .B(n18621), .X(n18620) );
  inv_x1_sg U46399 ( .A(n18611), .X(n54197) );
  nand_x1_sg U46400 ( .A(n18720), .B(n18721), .X(n18719) );
  nand_x1_sg U46401 ( .A(n18752), .B(n46329), .X(n18751) );
  nand_x1_sg U46402 ( .A(n19072), .B(n43862), .X(n19071) );
  nand_x1_sg U46403 ( .A(n54373), .B(n19076), .X(n19075) );
  nand_x1_sg U46404 ( .A(n54393), .B(n19037), .X(n19074) );
  inv_x1_sg U46405 ( .A(n19076), .X(n54393) );
  nand_x1_sg U46406 ( .A(n54367), .B(n46321), .X(n19023) );
  nor_x1_sg U46407 ( .A(n19102), .B(n54388), .X(n19101) );
  nand_x4_sg U46408 ( .A(n19130), .B(n19131), .X(n19078) );
  nand_x1_sg U46409 ( .A(n54374), .B(n19050), .X(n19130) );
  nand_x1_sg U46410 ( .A(n54361), .B(n19094), .X(n19131) );
  nand_x4_sg U46411 ( .A(n46309), .B(n46325), .X(n19079) );
  nand_x4_sg U46412 ( .A(n54367), .B(n46316), .X(n19094) );
  nand_x1_sg U46413 ( .A(n46311), .B(n46325), .X(n19047) );
  nand_x4_sg U46414 ( .A(n54435), .B(n19169), .X(n19108) );
  inv_x1_sg U46415 ( .A(n19171), .X(n54435) );
  nand_x1_sg U46416 ( .A(n19170), .B(n54434), .X(n19169) );
  inv_x1_sg U46417 ( .A(n19136), .X(n54421) );
  inv_x1_sg U46418 ( .A(n19310), .X(n54510) );
  inv_x2_sg U46419 ( .A(n19304), .X(n44442) );
  nor_x1_sg U46420 ( .A(n54492), .B(n19306), .X(n19304) );
  inv_x1_sg U46421 ( .A(n19196), .X(n54409) );
  inv_x1_sg U46422 ( .A(n19244), .X(n54444) );
  inv_x1_sg U46423 ( .A(n19221), .X(n54473) );
  inv_x1_sg U46424 ( .A(n19296), .X(n54483) );
  inv_x1_sg U46425 ( .A(n19267), .X(n54497) );
  nand_x4_sg U46426 ( .A(n46313), .B(n46309), .X(n19358) );
  nand_x1_sg U46427 ( .A(n19371), .B(n19370), .X(n19372) );
  nand_x1_sg U46428 ( .A(n19359), .B(n19361), .X(n19360) );
  nand_x1_sg U46429 ( .A(n54411), .B(n54432), .X(n19361) );
  nand_x4_sg U46430 ( .A(n19335), .B(n19336), .X(n19267) );
  nand_x1_sg U46431 ( .A(n46311), .B(n54496), .X(n19336) );
  inv_x1_sg U46432 ( .A(n19375), .X(n54566) );
  nand_x1_sg U46433 ( .A(n19376), .B(n19377), .X(n19374) );
  inv_x2_sg U46434 ( .A(n19437), .X(n44035) );
  nor_x1_sg U46435 ( .A(n19603), .B(n19604), .X(n19437) );
  nand_x1_sg U46436 ( .A(n54392), .B(n19371), .X(n19411) );
  nand_x1_sg U46437 ( .A(n54517), .B(n19399), .X(n19398) );
  nand_x1_sg U46438 ( .A(n19496), .B(n19497), .X(n19495) );
  nand_x1_sg U46439 ( .A(n19528), .B(n54392), .X(n19527) );
  inv_x1_sg U46440 ( .A(n19440), .X(n45436) );
  nand_x1_sg U46441 ( .A(n19841), .B(n54660), .X(n19840) );
  inv_x1_sg U46442 ( .A(n19844), .X(n54678) );
  nand_x1_sg U46443 ( .A(n54647), .B(n46301), .X(n19790) );
  nor_x1_sg U46444 ( .A(n19848), .B(n19849), .X(n19847) );
  nand_x4_sg U46445 ( .A(n46296), .B(n54647), .X(n19864) );
  inv_x2_sg U46446 ( .A(n19938), .X(n44728) );
  inv_x1_sg U46447 ( .A(n19906), .X(n54700) );
  nand_x1_sg U46448 ( .A(n19979), .B(n46285), .X(n19978) );
  inv_x1_sg U46449 ( .A(n19965), .X(n54689) );
  nand_x4_sg U46450 ( .A(n46296), .B(n54688), .X(n19965) );
  inv_x1_sg U46451 ( .A(n20013), .X(n54725) );
  inv_x1_sg U46452 ( .A(n20078), .X(n54795) );
  inv_x2_sg U46453 ( .A(n20072), .X(n44464) );
  nor_x1_sg U46454 ( .A(n54777), .B(n20074), .X(n20072) );
  inv_x1_sg U46455 ( .A(n20059), .X(n54752) );
  inv_x2_sg U46456 ( .A(n19974), .X(n44079) );
  nand_x1_sg U46457 ( .A(n19932), .B(n19931), .X(n19974) );
  inv_x1_sg U46458 ( .A(n20036), .X(n54781) );
  inv_x1_sg U46459 ( .A(n20137), .X(n44416) );
  nand_x1_sg U46460 ( .A(n54660), .B(n54780), .X(n20104) );
  nand_x1_sg U46461 ( .A(n20126), .B(n20128), .X(n20127) );
  inv_x1_sg U46462 ( .A(n20350), .X(n54815) );
  nand_x4_sg U46463 ( .A(n20347), .B(n20354), .X(n20145) );
  nand_x1_sg U46464 ( .A(n20355), .B(n54845), .X(n20354) );
  inv_x1_sg U46465 ( .A(n20356), .X(n54845) );
  nand_x1_sg U46466 ( .A(n54842), .B(n20309), .X(n20307) );
  inv_x1_sg U46467 ( .A(n20308), .X(n54842) );
  nand_x1_sg U46468 ( .A(n54847), .B(n43098), .X(n20303) );
  nand_x1_sg U46469 ( .A(n43099), .B(n20306), .X(n20304) );
  inv_x1_sg U46470 ( .A(n20306), .X(n54847) );
  inv_x2_sg U46471 ( .A(n20206), .X(n44376) );
  nor_x1_sg U46472 ( .A(n20375), .B(n20376), .X(n20206) );
  nand_x1_sg U46473 ( .A(n54805), .B(n20167), .X(n20166) );
  inv_x1_sg U46474 ( .A(n20157), .X(n54764) );
  nand_x1_sg U46475 ( .A(n20266), .B(n20267), .X(n20265) );
  nand_x1_sg U46476 ( .A(n20298), .B(n46285), .X(n20297) );
  nand_x1_sg U46477 ( .A(n20616), .B(n43860), .X(n20615) );
  nand_x1_sg U46478 ( .A(n54941), .B(n20620), .X(n20619) );
  nand_x1_sg U46479 ( .A(n54961), .B(n20581), .X(n20618) );
  inv_x1_sg U46480 ( .A(n20620), .X(n54961) );
  nand_x1_sg U46481 ( .A(n54935), .B(n46276), .X(n20567) );
  nor_x1_sg U46482 ( .A(n20646), .B(n54956), .X(n20645) );
  nand_x4_sg U46483 ( .A(n20674), .B(n20675), .X(n20622) );
  nand_x1_sg U46484 ( .A(n54942), .B(n20594), .X(n20674) );
  nand_x1_sg U46485 ( .A(n54929), .B(n20638), .X(n20675) );
  nand_x4_sg U46486 ( .A(n46264), .B(n46280), .X(n20623) );
  nand_x4_sg U46487 ( .A(n54935), .B(n46271), .X(n20638) );
  nand_x1_sg U46488 ( .A(n46266), .B(n46280), .X(n20591) );
  nand_x4_sg U46489 ( .A(n55003), .B(n20713), .X(n20652) );
  inv_x1_sg U46490 ( .A(n20715), .X(n55003) );
  nand_x1_sg U46491 ( .A(n20714), .B(n55002), .X(n20713) );
  inv_x1_sg U46492 ( .A(n20680), .X(n54989) );
  inv_x1_sg U46493 ( .A(n20854), .X(n55078) );
  inv_x2_sg U46494 ( .A(n20848), .X(n44440) );
  nor_x1_sg U46495 ( .A(n55060), .B(n20850), .X(n20848) );
  inv_x1_sg U46496 ( .A(n20740), .X(n54977) );
  inv_x1_sg U46497 ( .A(n20788), .X(n55012) );
  inv_x1_sg U46498 ( .A(n20765), .X(n55041) );
  inv_x1_sg U46499 ( .A(n20840), .X(n55051) );
  inv_x1_sg U46500 ( .A(n20811), .X(n55065) );
  nand_x4_sg U46501 ( .A(n46268), .B(n46264), .X(n20902) );
  nand_x1_sg U46502 ( .A(n20915), .B(n20914), .X(n20916) );
  nand_x1_sg U46503 ( .A(n20903), .B(n20905), .X(n20904) );
  nand_x1_sg U46504 ( .A(n54979), .B(n55000), .X(n20905) );
  nand_x4_sg U46505 ( .A(n20879), .B(n20880), .X(n20811) );
  nand_x1_sg U46506 ( .A(n46266), .B(n55064), .X(n20880) );
  inv_x1_sg U46507 ( .A(n20919), .X(n55134) );
  nand_x1_sg U46508 ( .A(n20920), .B(n20921), .X(n20918) );
  inv_x2_sg U46509 ( .A(n20981), .X(n44033) );
  nor_x1_sg U46510 ( .A(n21147), .B(n21148), .X(n20981) );
  nand_x1_sg U46511 ( .A(n54960), .B(n20915), .X(n20955) );
  nand_x1_sg U46512 ( .A(n55085), .B(n20943), .X(n20942) );
  nand_x1_sg U46513 ( .A(n21040), .B(n21041), .X(n21039) );
  nand_x1_sg U46514 ( .A(n21072), .B(n54960), .X(n21071) );
  inv_x1_sg U46515 ( .A(n20984), .X(n45428) );
  nand_x1_sg U46516 ( .A(n21386), .B(n55228), .X(n21385) );
  inv_x1_sg U46517 ( .A(n21389), .X(n55246) );
  nand_x1_sg U46518 ( .A(n55215), .B(n46256), .X(n21335) );
  nor_x1_sg U46519 ( .A(n21393), .B(n21394), .X(n21392) );
  nand_x4_sg U46520 ( .A(n46251), .B(n55215), .X(n21409) );
  inv_x2_sg U46521 ( .A(n21483), .X(n44726) );
  inv_x1_sg U46522 ( .A(n21451), .X(n55268) );
  nand_x1_sg U46523 ( .A(n21524), .B(n46240), .X(n21523) );
  inv_x1_sg U46524 ( .A(n21510), .X(n55257) );
  nand_x4_sg U46525 ( .A(n46251), .B(n55256), .X(n21510) );
  inv_x1_sg U46526 ( .A(n21558), .X(n55293) );
  inv_x1_sg U46527 ( .A(n21623), .X(n55363) );
  inv_x2_sg U46528 ( .A(n21617), .X(n44462) );
  nor_x1_sg U46529 ( .A(n55345), .B(n21619), .X(n21617) );
  inv_x1_sg U46530 ( .A(n21604), .X(n55320) );
  inv_x2_sg U46531 ( .A(n21519), .X(n44077) );
  nand_x1_sg U46532 ( .A(n21477), .B(n21476), .X(n21519) );
  inv_x1_sg U46533 ( .A(n21581), .X(n55349) );
  inv_x1_sg U46534 ( .A(n21682), .X(n44414) );
  nand_x1_sg U46535 ( .A(n55228), .B(n55348), .X(n21649) );
  nand_x1_sg U46536 ( .A(n21671), .B(n21673), .X(n21672) );
  inv_x1_sg U46537 ( .A(n21895), .X(n55383) );
  nand_x4_sg U46538 ( .A(n21892), .B(n21899), .X(n21690) );
  nand_x1_sg U46539 ( .A(n21900), .B(n55413), .X(n21899) );
  inv_x1_sg U46540 ( .A(n21901), .X(n55413) );
  nand_x1_sg U46541 ( .A(n55410), .B(n21854), .X(n21852) );
  inv_x1_sg U46542 ( .A(n21853), .X(n55410) );
  nand_x1_sg U46543 ( .A(n55415), .B(n43096), .X(n21848) );
  nand_x1_sg U46544 ( .A(n43097), .B(n21851), .X(n21849) );
  inv_x1_sg U46545 ( .A(n21851), .X(n55415) );
  inv_x2_sg U46546 ( .A(n21751), .X(n44374) );
  nor_x1_sg U46547 ( .A(n21920), .B(n21921), .X(n21751) );
  nand_x1_sg U46548 ( .A(n55373), .B(n21712), .X(n21711) );
  inv_x1_sg U46549 ( .A(n21702), .X(n55332) );
  nand_x1_sg U46550 ( .A(n21811), .B(n21812), .X(n21810) );
  nand_x1_sg U46551 ( .A(n21843), .B(n46240), .X(n21842) );
  nand_x1_sg U46552 ( .A(n8204), .B(n50085), .X(n29658) );
  inv_x1_sg U46553 ( .A(n29659), .X(n50085) );
  nand_x1_sg U46554 ( .A(n8284), .B(n50075), .X(n30269) );
  inv_x1_sg U46555 ( .A(n30270), .X(n50075) );
  nand_x1_sg U46556 ( .A(n8364), .B(n50063), .X(n30240) );
  nand_x1_sg U46557 ( .A(n24487), .B(n30242), .X(n30239) );
  inv_x1_sg U46558 ( .A(n30241), .X(n50063) );
  nand_x1_sg U46559 ( .A(n8444), .B(n50052), .X(n30211) );
  inv_x1_sg U46560 ( .A(n30212), .X(n50052) );
  nand_x1_sg U46561 ( .A(n8204), .B(n29660), .X(n29857) );
  nand_x1_sg U46562 ( .A(n8284), .B(n30271), .X(n30529) );
  inv_x1_sg U46563 ( .A(n30509), .X(n50020) );
  inv_x1_sg U46564 ( .A(n30490), .X(n50010) );
  inv_x1_sg U46565 ( .A(n30496), .X(n50014) );
  inv_x1_sg U46566 ( .A(n30020), .X(n49996) );
  nand_x1_sg U46567 ( .A(n8205), .B(n29837), .X(n29836) );
  inv_x1_sg U46568 ( .A(n30764), .X(n49976) );
  inv_x1_sg U46569 ( .A(n30745), .X(n49966) );
  inv_x1_sg U46570 ( .A(n30751), .X(n49970) );
  inv_x1_sg U46571 ( .A(n30990), .X(n49932) );
  inv_x1_sg U46572 ( .A(n30023), .X(n49952) );
  nand_x1_sg U46573 ( .A(n8206), .B(n29830), .X(n29829) );
  inv_x1_sg U46574 ( .A(n30971), .X(n49922) );
  inv_x1_sg U46575 ( .A(n30977), .X(n49926) );
  nor_x1_sg U46576 ( .A(n30955), .B(out_L1[15]), .X(n30954) );
  inv_x1_sg U46577 ( .A(n30026), .X(n49904) );
  nand_x1_sg U46578 ( .A(n8207), .B(n29823), .X(n29822) );
  inv_x1_sg U46579 ( .A(n31195), .X(n49886) );
  inv_x1_sg U46580 ( .A(n31176), .X(n49876) );
  inv_x1_sg U46581 ( .A(n31182), .X(n49880) );
  inv_x1_sg U46582 ( .A(n31385), .X(n49840) );
  inv_x1_sg U46583 ( .A(n30029), .X(n49857) );
  nand_x1_sg U46584 ( .A(n8208), .B(n29816), .X(n29815) );
  inv_x1_sg U46585 ( .A(n31013), .X(n49866) );
  nand_x1_sg U46586 ( .A(n8288), .B(n30685), .X(n30684) );
  inv_x1_sg U46587 ( .A(n31366), .X(n49830) );
  inv_x1_sg U46588 ( .A(n31372), .X(n49834) );
  nor_x1_sg U46589 ( .A(n31350), .B(out_L1[13]), .X(n31349) );
  inv_x1_sg U46590 ( .A(n30032), .X(n49809) );
  nand_x1_sg U46591 ( .A(n8209), .B(n29809), .X(n29808) );
  inv_x1_sg U46592 ( .A(n31016), .X(n49818) );
  nand_x1_sg U46593 ( .A(n8289), .B(n30678), .X(n30677) );
  inv_x1_sg U46594 ( .A(n31556), .X(n49823) );
  inv_x1_sg U46595 ( .A(n31537), .X(n49785) );
  inv_x1_sg U46596 ( .A(n31543), .X(n49789) );
  inv_x1_sg U46597 ( .A(n30035), .X(n49762) );
  inv_x1_sg U46598 ( .A(n31019), .X(n49771) );
  nand_x1_sg U46599 ( .A(n8290), .B(n30671), .X(n30670) );
  nand_x1_sg U46600 ( .A(n8210), .B(n29802), .X(n29801) );
  inv_x1_sg U46601 ( .A(n30305), .X(n49764) );
  inv_x1_sg U46602 ( .A(n31559), .X(n49777) );
  inv_x1_sg U46603 ( .A(n31690), .X(n49739) );
  inv_x1_sg U46604 ( .A(n31696), .X(n49743) );
  nor_x1_sg U46605 ( .A(n31674), .B(out_L1[11]), .X(n31673) );
  inv_x1_sg U46606 ( .A(n30038), .X(n49713) );
  nand_x1_sg U46607 ( .A(n8211), .B(n29795), .X(n29794) );
  inv_x1_sg U46608 ( .A(n31022), .X(n49722) );
  nand_x1_sg U46609 ( .A(n8291), .B(n30664), .X(n30663) );
  inv_x1_sg U46610 ( .A(n31562), .X(n49727) );
  inv_x1_sg U46611 ( .A(n31834), .X(n49693) );
  inv_x1_sg U46612 ( .A(n31840), .X(n49731) );
  inv_x1_sg U46613 ( .A(n30041), .X(n49666) );
  nand_x1_sg U46614 ( .A(n8212), .B(n29788), .X(n29787) );
  inv_x1_sg U46615 ( .A(n31025), .X(n49675) );
  nand_x1_sg U46616 ( .A(n8292), .B(n30657), .X(n30656) );
  inv_x1_sg U46617 ( .A(n31565), .X(n49681) );
  inv_x1_sg U46618 ( .A(n31950), .X(n49687) );
  nor_x1_sg U46619 ( .A(n31934), .B(out_L1[9]), .X(n31933) );
  inv_x1_sg U46620 ( .A(n30044), .X(n49619) );
  nand_x1_sg U46621 ( .A(n8213), .B(n29781), .X(n29780) );
  inv_x1_sg U46622 ( .A(n31028), .X(n49628) );
  nand_x1_sg U46623 ( .A(n8293), .B(n30650), .X(n30649) );
  inv_x1_sg U46624 ( .A(n31568), .X(n49633) );
  inv_x1_sg U46625 ( .A(n31953), .X(n49640) );
  inv_x1_sg U46626 ( .A(n30047), .X(n49573) );
  nand_x1_sg U46627 ( .A(n8214), .B(n29774), .X(n29773) );
  inv_x1_sg U46628 ( .A(n31031), .X(n49582) );
  nand_x1_sg U46629 ( .A(n8294), .B(n30643), .X(n30642) );
  inv_x1_sg U46630 ( .A(n31571), .X(n49587) );
  inv_x1_sg U46631 ( .A(n31956), .X(n49594) );
  inv_x1_sg U46632 ( .A(n32021), .X(n49550) );
  inv_x1_sg U46633 ( .A(n30050), .X(n49526) );
  nand_x1_sg U46634 ( .A(n8215), .B(n29767), .X(n29766) );
  inv_x1_sg U46635 ( .A(n31034), .X(n49535) );
  nand_x1_sg U46636 ( .A(n8295), .B(n30636), .X(n30635) );
  inv_x1_sg U46637 ( .A(n31574), .X(n49541) );
  inv_x1_sg U46638 ( .A(n31959), .X(n49548) );
  nor_x1_sg U46639 ( .A(n32118), .B(out_L1[6]), .X(n32117) );
  inv_x2_sg U46640 ( .A(n32116), .X(n44296) );
  nor_x1_sg U46641 ( .A(n40852), .B(n49504), .X(n32116) );
  inv_x1_sg U46642 ( .A(n31037), .X(n49488) );
  inv_x1_sg U46643 ( .A(n30323), .X(n49481) );
  inv_x1_sg U46644 ( .A(n30053), .X(n49479) );
  nand_x1_sg U46645 ( .A(n8216), .B(n29760), .X(n29759) );
  inv_x1_sg U46646 ( .A(n31577), .X(n49493) );
  inv_x1_sg U46647 ( .A(n31962), .X(n49500) );
  inv_x1_sg U46648 ( .A(n32008), .X(n49456) );
  inv_x1_sg U46649 ( .A(n30056), .X(n49433) );
  nand_x1_sg U46650 ( .A(n8217), .B(n29753), .X(n29752) );
  inv_x1_sg U46651 ( .A(n31040), .X(n49442) );
  nand_x1_sg U46652 ( .A(n8297), .B(n30622), .X(n30621) );
  inv_x1_sg U46653 ( .A(n31580), .X(n49447) );
  inv_x1_sg U46654 ( .A(n31965), .X(n49454) );
  inv_x1_sg U46655 ( .A(n31043), .X(n49396) );
  inv_x1_sg U46656 ( .A(n30329), .X(n49389) );
  inv_x1_sg U46657 ( .A(n30059), .X(n49387) );
  nand_x1_sg U46658 ( .A(n8218), .B(n29746), .X(n29745) );
  inv_x1_sg U46659 ( .A(n31583), .X(n49402) );
  inv_x1_sg U46660 ( .A(n31995), .X(n49366) );
  inv_x1_sg U46661 ( .A(n31968), .X(n49409) );
  inv_x1_sg U46662 ( .A(n31046), .X(n49352) );
  inv_x1_sg U46663 ( .A(n30332), .X(n49345) );
  inv_x1_sg U46664 ( .A(n30062), .X(n49343) );
  nand_x1_sg U46665 ( .A(n8219), .B(n29739), .X(n29738) );
  inv_x1_sg U46666 ( .A(n31586), .X(n49357) );
  inv_x1_sg U46667 ( .A(n31261), .X(n49308) );
  inv_x1_sg U46668 ( .A(n31989), .X(n49317) );
  inv_x1_sg U46669 ( .A(n31971), .X(n49364) );
  nand_x1_sg U46670 ( .A(n8220), .B(n29732), .X(n29731) );
  inv_x1_sg U46671 ( .A(n10266), .X(n55461) );
  nand_x2_sg U46672 ( .A(n51265), .B(n25595), .X(n25593) );
  inv_x1_sg U46673 ( .A(n25596), .X(n51265) );
  inv_x1_sg U46674 ( .A(n25593), .X(n51266) );
  nand_x2_sg U46675 ( .A(n51541), .B(n25876), .X(n25874) );
  inv_x1_sg U46676 ( .A(n25877), .X(n51541) );
  inv_x1_sg U46677 ( .A(n25874), .X(n51542) );
  nand_x1_sg U46678 ( .A(n25875), .B(n50988), .X(n25934) );
  nand_x2_sg U46679 ( .A(n51550), .B(n25870), .X(n25868) );
  inv_x1_sg U46680 ( .A(n25871), .X(n51550) );
  inv_x1_sg U46681 ( .A(n25868), .X(n51551) );
  inv_x1_sg U46682 ( .A(n25859), .X(n51574) );
  nor_x1_sg U46683 ( .A(n25849), .B(n25850), .X(n25848) );
  inv_x1_sg U46684 ( .A(n46035), .X(n43756) );
  inv_x1_sg U46685 ( .A(n25930), .X(n51549) );
  inv_x1_sg U46686 ( .A(n25857), .X(n51557) );
  nand_x2_sg U46687 ( .A(n51824), .B(n26156), .X(n26154) );
  inv_x1_sg U46688 ( .A(n26157), .X(n51824) );
  inv_x1_sg U46689 ( .A(n26154), .X(n51825) );
  nand_x2_sg U46690 ( .A(n52098), .B(n26435), .X(n26433) );
  inv_x1_sg U46691 ( .A(n26436), .X(n52098) );
  inv_x1_sg U46692 ( .A(n26433), .X(n52099) );
  nand_x1_sg U46693 ( .A(n26434), .B(n51026), .X(n26493) );
  nand_x2_sg U46694 ( .A(n52107), .B(n26429), .X(n26427) );
  inv_x1_sg U46695 ( .A(n26430), .X(n52107) );
  inv_x1_sg U46696 ( .A(n26427), .X(n52108) );
  inv_x1_sg U46697 ( .A(n26418), .X(n52131) );
  nor_x1_sg U46698 ( .A(n26408), .B(n26409), .X(n26407) );
  nand_x1_sg U46699 ( .A(n26408), .B(n26409), .X(n26410) );
  inv_x1_sg U46700 ( .A(n26416), .X(n52114) );
  inv_x1_sg U46701 ( .A(n45225), .X(n43752) );
  inv_x1_sg U46702 ( .A(n26489), .X(n52106) );
  nand_x2_sg U46703 ( .A(n52376), .B(n26713), .X(n26711) );
  inv_x1_sg U46704 ( .A(n26714), .X(n52376) );
  inv_x1_sg U46705 ( .A(n26711), .X(n52377) );
  nand_x2_sg U46706 ( .A(n52653), .B(n26992), .X(n26990) );
  inv_x1_sg U46707 ( .A(n26993), .X(n52653) );
  inv_x1_sg U46708 ( .A(n26990), .X(n52654) );
  inv_x1_sg U46709 ( .A(n27042), .X(n44322) );
  nand_x2_sg U46710 ( .A(n52932), .B(n27272), .X(n27270) );
  inv_x1_sg U46711 ( .A(n27273), .X(n52932) );
  inv_x1_sg U46712 ( .A(n27270), .X(n52933) );
  nand_x1_sg U46713 ( .A(n27271), .B(n51084), .X(n27330) );
  nand_x2_sg U46714 ( .A(n52941), .B(n27266), .X(n27264) );
  inv_x1_sg U46715 ( .A(n27267), .X(n52941) );
  inv_x1_sg U46716 ( .A(n27264), .X(n52942) );
  inv_x1_sg U46717 ( .A(n27255), .X(n52965) );
  nor_x1_sg U46718 ( .A(n27245), .B(n27246), .X(n27244) );
  nand_x1_sg U46719 ( .A(n27245), .B(n27246), .X(n27247) );
  inv_x1_sg U46720 ( .A(n27253), .X(n52948) );
  inv_x1_sg U46721 ( .A(n45223), .X(n43750) );
  inv_x1_sg U46722 ( .A(n27326), .X(n52940) );
  nand_x2_sg U46723 ( .A(n53212), .B(n27551), .X(n27549) );
  inv_x1_sg U46724 ( .A(n27552), .X(n53212) );
  inv_x1_sg U46725 ( .A(n27549), .X(n53213) );
  nand_x2_sg U46726 ( .A(n53490), .B(n27830), .X(n27828) );
  inv_x1_sg U46727 ( .A(n27831), .X(n53490) );
  inv_x1_sg U46728 ( .A(n27828), .X(n53491) );
  nand_x1_sg U46729 ( .A(n27829), .B(n51122), .X(n27888) );
  nand_x2_sg U46730 ( .A(n53499), .B(n27824), .X(n27822) );
  inv_x1_sg U46731 ( .A(n27825), .X(n53499) );
  inv_x1_sg U46732 ( .A(n27822), .X(n53500) );
  inv_x1_sg U46733 ( .A(n27813), .X(n53523) );
  nor_x1_sg U46734 ( .A(n27803), .B(n27804), .X(n27802) );
  nand_x1_sg U46735 ( .A(n27803), .B(n27804), .X(n27805) );
  inv_x1_sg U46736 ( .A(n27811), .X(n53506) );
  inv_x1_sg U46737 ( .A(n45221), .X(n43748) );
  inv_x1_sg U46738 ( .A(n27884), .X(n53498) );
  nand_x2_sg U46739 ( .A(n53770), .B(n28111), .X(n28109) );
  inv_x1_sg U46740 ( .A(n28112), .X(n53770) );
  inv_x1_sg U46741 ( .A(n28109), .X(n53771) );
  nand_x2_sg U46742 ( .A(n53777), .B(n28105), .X(n28103) );
  inv_x1_sg U46743 ( .A(n28106), .X(n53777) );
  inv_x1_sg U46744 ( .A(n28103), .X(n53778) );
  nand_x1_sg U46745 ( .A(n28110), .B(n51141), .X(n28169) );
  nand_x1_sg U46746 ( .A(n28084), .B(n28085), .X(n28086) );
  inv_x1_sg U46747 ( .A(n28092), .X(n53785) );
  nand_x1_sg U46748 ( .A(n45219), .B(n28444), .X(n28443) );
  nand_x1_sg U46749 ( .A(n28377), .B(n51161), .X(n28442) );
  nand_x1_sg U46750 ( .A(n28363), .B(n28364), .X(n28365) );
  inv_x1_sg U46751 ( .A(n28364), .X(n54081) );
  nand_x2_sg U46752 ( .A(n54335), .B(n28669), .X(n28667) );
  inv_x1_sg U46753 ( .A(n28670), .X(n54335) );
  inv_x1_sg U46754 ( .A(n28667), .X(n54336) );
  nand_x2_sg U46755 ( .A(n54342), .B(n28663), .X(n28661) );
  inv_x1_sg U46756 ( .A(n28664), .X(n54342) );
  inv_x1_sg U46757 ( .A(n28661), .X(n54343) );
  nand_x1_sg U46758 ( .A(n28668), .B(n51178), .X(n28727) );
  nand_x1_sg U46759 ( .A(n28642), .B(n28643), .X(n28644) );
  inv_x1_sg U46760 ( .A(n28650), .X(n54350) );
  nand_x2_sg U46761 ( .A(n54619), .B(n28947), .X(n28945) );
  inv_x1_sg U46762 ( .A(n28948), .X(n54619) );
  inv_x1_sg U46763 ( .A(n28945), .X(n54620) );
  nand_x2_sg U46764 ( .A(n54903), .B(n29230), .X(n29228) );
  inv_x1_sg U46765 ( .A(n29231), .X(n54903) );
  inv_x1_sg U46766 ( .A(n29228), .X(n54904) );
  nand_x2_sg U46767 ( .A(n54910), .B(n29224), .X(n29222) );
  inv_x1_sg U46768 ( .A(n29225), .X(n54910) );
  inv_x1_sg U46769 ( .A(n29222), .X(n54911) );
  nand_x1_sg U46770 ( .A(n29229), .B(n51216), .X(n29288) );
  nand_x1_sg U46771 ( .A(n29203), .B(n29204), .X(n29205) );
  inv_x1_sg U46772 ( .A(n29211), .X(n54918) );
  nand_x2_sg U46773 ( .A(n55187), .B(n29508), .X(n29506) );
  inv_x1_sg U46774 ( .A(n29509), .X(n55187) );
  inv_x1_sg U46775 ( .A(n29506), .X(n55188) );
  inv_x2_sg U46776 ( .A(n39307), .X(n43784) );
  nor_x1_sg U46777 ( .A(n39303), .B(n39300), .X(n39307) );
  nand_x1_sg U46778 ( .A(n8484), .B(n50947), .X(n22000) );
  inv_x1_sg U46779 ( .A(n22001), .X(n50947) );
  nand_x1_sg U46780 ( .A(n8544), .B(n50949), .X(n22617) );
  nand_x1_sg U46781 ( .A(n9391), .B(n22184), .X(n22616) );
  inv_x1_sg U46782 ( .A(n22618), .X(n50949) );
  nand_x1_sg U46783 ( .A(n8624), .B(n50927), .X(n22589) );
  nand_x1_sg U46784 ( .A(n9364), .B(n22591), .X(n22588) );
  inv_x1_sg U46785 ( .A(n22590), .X(n50927) );
  nand_x1_sg U46786 ( .A(n8524), .B(n50940), .X(n21986) );
  inv_x1_sg U46787 ( .A(n21987), .X(n50940) );
  inv_x1_sg U46788 ( .A(n21991), .X(n50945) );
  nand_x1_sg U46789 ( .A(n8503), .B(n21990), .X(n21989) );
  nand_x1_sg U46790 ( .A(n8564), .B(n50936), .X(n22610) );
  inv_x1_sg U46791 ( .A(n22611), .X(n50936) );
  nand_x1_sg U46792 ( .A(n8604), .B(n50930), .X(n22596) );
  inv_x1_sg U46793 ( .A(n22597), .X(n50930) );
  inv_x1_sg U46794 ( .A(n22601), .X(n50935) );
  nand_x1_sg U46795 ( .A(n8583), .B(n22600), .X(n22599) );
  nand_x1_sg U46796 ( .A(n8724), .B(n50913), .X(n22552) );
  inv_x1_sg U46797 ( .A(n22553), .X(n50913) );
  nand_x1_sg U46798 ( .A(n8663), .B(n22572), .X(n22571) );
  nand_x1_sg U46799 ( .A(n8644), .B(n22582), .X(n22581) );
  nand_x1_sg U46800 ( .A(n8704), .B(n50917), .X(n22559) );
  nand_x1_sg U46801 ( .A(n22561), .B(n22562), .X(n22558) );
  inv_x1_sg U46802 ( .A(n22560), .X(n50917) );
  inv_x1_sg U46803 ( .A(n22543), .X(n50912) );
  nand_x1_sg U46804 ( .A(n8743), .B(n22542), .X(n22541) );
  nand_x1_sg U46805 ( .A(n8684), .B(n50919), .X(n22567) );
  inv_x1_sg U46806 ( .A(n22568), .X(n50919) );
  inv_x1_sg U46807 ( .A(n22004), .X(n50900) );
  inv_x1_sg U46808 ( .A(n22621), .X(n50905) );
  inv_x1_sg U46809 ( .A(n22854), .X(n50885) );
  inv_x1_sg U46810 ( .A(n22189), .X(n50895) );
  inv_x2_sg U46811 ( .A(n22175), .X(n44652) );
  nor_x1_sg U46812 ( .A(n22191), .B(n50903), .X(n22175) );
  inv_x1_sg U46813 ( .A(n22872), .X(n50907) );
  inv_x1_sg U46814 ( .A(n22860), .X(n50888) );
  inv_x2_sg U46815 ( .A(n22779), .X(n44632) );
  nor_x1_sg U46816 ( .A(n22862), .B(n50891), .X(n22779) );
  nor_x1_sg U46817 ( .A(n22808), .B(out_L2[17]), .X(n22807) );
  nor_x1_sg U46818 ( .A(n9454), .B(n50863), .X(n22847) );
  nand_x1_sg U46819 ( .A(n8664), .B(n22576), .X(n22840) );
  nand_x1_sg U46820 ( .A(n8744), .B(n22547), .X(n22814) );
  inv_x1_sg U46821 ( .A(n22837), .X(n50876) );
  inv_x1_sg U46822 ( .A(n22821), .X(n50870) );
  nand_x1_sg U46823 ( .A(n8724), .B(n22554), .X(n22820) );
  nand_x1_sg U46824 ( .A(n8704), .B(n22562), .X(n22827) );
  inv_x1_sg U46825 ( .A(n22007), .X(n50851) );
  inv_x1_sg U46826 ( .A(n22624), .X(n50857) );
  nand_x1_sg U46827 ( .A(n8665), .B(n22844), .X(n23095) );
  inv_x1_sg U46828 ( .A(n22875), .X(n50859) );
  inv_x1_sg U46829 ( .A(n23117), .X(n50843) );
  nand_x1_sg U46830 ( .A(n8585), .B(n22867), .X(n23120) );
  inv_x1_sg U46831 ( .A(n23111), .X(n50840) );
  inv_x1_sg U46832 ( .A(n22352), .X(n50856) );
  nand_x1_sg U46833 ( .A(n8525), .B(n22190), .X(n22351) );
  inv_x1_sg U46834 ( .A(n23076), .X(n50826) );
  nand_x1_sg U46835 ( .A(n8725), .B(n22825), .X(n23075) );
  nand_x1_sg U46836 ( .A(n8705), .B(n22831), .X(n23082) );
  nand_x1_sg U46837 ( .A(n8646), .B(n23105), .X(n23104) );
  inv_x1_sg U46838 ( .A(n23067), .X(n50864) );
  inv_x1_sg U46839 ( .A(n22010), .X(n50806) );
  inv_x1_sg U46840 ( .A(n22627), .X(n50813) );
  nand_x1_sg U46841 ( .A(n8666), .B(n23099), .X(n23321) );
  inv_x1_sg U46842 ( .A(n22878), .X(n50815) );
  inv_x1_sg U46843 ( .A(n23341), .X(n50819) );
  nand_x1_sg U46844 ( .A(n8586), .B(n23031), .X(n23030) );
  inv_x1_sg U46845 ( .A(n23335), .X(n50797) );
  inv_x1_sg U46846 ( .A(n22341), .X(n50812) );
  nand_x1_sg U46847 ( .A(n8526), .B(n22340), .X(n22339) );
  inv_x2_sg U46848 ( .A(n22161), .X(n44618) );
  nor_x1_sg U46849 ( .A(n22163), .B(n50809), .X(n22161) );
  inv_x1_sg U46850 ( .A(n23302), .X(n50782) );
  nand_x1_sg U46851 ( .A(n8726), .B(n23080), .X(n23301) );
  nand_x1_sg U46852 ( .A(n8706), .B(n23086), .X(n23308) );
  inv_x2_sg U46853 ( .A(n23328), .X(n44288) );
  nand_x2_sg U46854 ( .A(n23292), .B(n23293), .X(n23287) );
  inv_x2_sg U46855 ( .A(n23288), .X(n44304) );
  inv_x1_sg U46856 ( .A(n22013), .X(n50758) );
  inv_x1_sg U46857 ( .A(n22630), .X(n50765) );
  nand_x1_sg U46858 ( .A(n8667), .B(n23325), .X(n23526) );
  inv_x1_sg U46859 ( .A(n22881), .X(n50767) );
  inv_x1_sg U46860 ( .A(n23344), .X(n50771) );
  nand_x1_sg U46861 ( .A(n8587), .B(n23025), .X(n23024) );
  inv_x1_sg U46862 ( .A(n23542), .X(n50773) );
  inv_x1_sg U46863 ( .A(n22335), .X(n50764) );
  nand_x1_sg U46864 ( .A(n8527), .B(n22334), .X(n22333) );
  inv_x2_sg U46865 ( .A(n22154), .X(n44616) );
  nor_x1_sg U46866 ( .A(n22156), .B(n50761), .X(n22154) );
  inv_x1_sg U46867 ( .A(n23507), .X(n50736) );
  nand_x1_sg U46868 ( .A(n8727), .B(n23306), .X(n23506) );
  nand_x1_sg U46869 ( .A(n8707), .B(n23312), .X(n23513) );
  nand_x1_sg U46870 ( .A(n8648), .B(n23536), .X(n23535) );
  nand_x1_sg U46871 ( .A(n23504), .B(n23505), .X(n23501) );
  nand_x1_sg U46872 ( .A(n8748), .B(n23503), .X(n23502) );
  inv_x1_sg U46873 ( .A(n23498), .X(n50777) );
  inv_x1_sg U46874 ( .A(n22016), .X(n50711) );
  inv_x1_sg U46875 ( .A(n22633), .X(n50718) );
  nand_x1_sg U46876 ( .A(n8668), .B(n23530), .X(n23716) );
  inv_x1_sg U46877 ( .A(n23545), .X(n50727) );
  inv_x1_sg U46878 ( .A(n22329), .X(n50717) );
  nand_x1_sg U46879 ( .A(n8528), .B(n22328), .X(n22327) );
  inv_x2_sg U46880 ( .A(n22147), .X(n44612) );
  nor_x1_sg U46881 ( .A(n22149), .B(n50714), .X(n22147) );
  inv_x1_sg U46882 ( .A(n22884), .X(n50720) );
  inv_x1_sg U46883 ( .A(n23254), .X(n50726) );
  nand_x1_sg U46884 ( .A(n8608), .B(n23253), .X(n23252) );
  inv_x2_sg U46885 ( .A(n23015), .X(n44614) );
  nor_x1_sg U46886 ( .A(n23017), .B(n50723), .X(n23015) );
  inv_x1_sg U46887 ( .A(n23697), .X(n50690) );
  nand_x1_sg U46888 ( .A(n8728), .B(n23511), .X(n23696) );
  nand_x1_sg U46889 ( .A(n8708), .B(n23517), .X(n23703) );
  inv_x2_sg U46890 ( .A(n23723), .X(n44286) );
  nand_x2_sg U46891 ( .A(n23687), .B(n23688), .X(n23682) );
  inv_x2_sg U46892 ( .A(n23683), .X(n45584) );
  inv_x1_sg U46893 ( .A(n22019), .X(n50663) );
  inv_x1_sg U46894 ( .A(n22636), .X(n50670) );
  nand_x1_sg U46895 ( .A(n8669), .B(n23720), .X(n23887) );
  inv_x1_sg U46896 ( .A(n23548), .X(n50679) );
  inv_x1_sg U46897 ( .A(n22323), .X(n50669) );
  nand_x1_sg U46898 ( .A(n8529), .B(n22322), .X(n22321) );
  inv_x2_sg U46899 ( .A(n22140), .X(n44608) );
  nor_x1_sg U46900 ( .A(n22142), .B(n50666), .X(n22140) );
  inv_x1_sg U46901 ( .A(n22887), .X(n50672) );
  inv_x1_sg U46902 ( .A(n23248), .X(n50678) );
  nand_x1_sg U46903 ( .A(n8609), .B(n23247), .X(n23246) );
  inv_x2_sg U46904 ( .A(n23008), .X(n44610) );
  nor_x1_sg U46905 ( .A(n23010), .B(n50675), .X(n23008) );
  inv_x1_sg U46906 ( .A(n23868), .X(n50645) );
  nand_x1_sg U46907 ( .A(n8729), .B(n23701), .X(n23867) );
  nand_x1_sg U46908 ( .A(n8709), .B(n23707), .X(n23874) );
  nand_x1_sg U46909 ( .A(n8650), .B(n23728), .X(n23727) );
  nand_x1_sg U46910 ( .A(n23865), .B(n23866), .X(n23862) );
  nand_x1_sg U46911 ( .A(n8750), .B(n23864), .X(n23863) );
  inv_x1_sg U46912 ( .A(n23859), .X(n50685) );
  inv_x1_sg U46913 ( .A(n23551), .X(n50632) );
  inv_x1_sg U46914 ( .A(n22317), .X(n50622) );
  nand_x1_sg U46915 ( .A(n8530), .B(n22316), .X(n22315) );
  inv_x1_sg U46916 ( .A(n22890), .X(n50625) );
  inv_x1_sg U46917 ( .A(n23242), .X(n50631) );
  nand_x1_sg U46918 ( .A(n8610), .B(n23241), .X(n23240) );
  inv_x2_sg U46919 ( .A(n23001), .X(n44644) );
  nor_x1_sg U46920 ( .A(n23003), .B(n50628), .X(n23001) );
  inv_x2_sg U46921 ( .A(n22133), .X(n44606) );
  nor_x1_sg U46922 ( .A(n22135), .B(n50619), .X(n22133) );
  inv_x1_sg U46923 ( .A(n22022), .X(n50616) );
  nand_x1_sg U46924 ( .A(n8670), .B(n23835), .X(n23834) );
  nand_x1_sg U46925 ( .A(n8550), .B(n22473), .X(n22472) );
  inv_x1_sg U46926 ( .A(n24021), .X(n50599) );
  nand_x1_sg U46927 ( .A(n8730), .B(n23872), .X(n24020) );
  nand_x1_sg U46928 ( .A(n8710), .B(n23878), .X(n24027) );
  nand_x2_sg U46929 ( .A(n24011), .B(n24012), .X(n24006) );
  inv_x2_sg U46930 ( .A(n24007), .X(n44724) );
  inv_x1_sg U46931 ( .A(n22025), .X(n50567) );
  inv_x1_sg U46932 ( .A(n22642), .X(n50574) );
  nand_x1_sg U46933 ( .A(n8671), .B(n23829), .X(n23828) );
  inv_x1_sg U46934 ( .A(n23554), .X(n50583) );
  inv_x1_sg U46935 ( .A(n22311), .X(n50573) );
  nand_x1_sg U46936 ( .A(n8531), .B(n22310), .X(n22309) );
  inv_x2_sg U46937 ( .A(n22126), .X(n44602) );
  nor_x1_sg U46938 ( .A(n22128), .B(n50570), .X(n22126) );
  inv_x1_sg U46939 ( .A(n22893), .X(n50576) );
  inv_x1_sg U46940 ( .A(n23236), .X(n50582) );
  nand_x1_sg U46941 ( .A(n8611), .B(n23235), .X(n23234) );
  inv_x2_sg U46942 ( .A(n22994), .X(n44604) );
  nor_x1_sg U46943 ( .A(n22996), .B(n50579), .X(n22994) );
  inv_x1_sg U46944 ( .A(n24165), .X(n50553) );
  nand_x1_sg U46945 ( .A(n8731), .B(n24025), .X(n24164) );
  nand_x1_sg U46946 ( .A(n8711), .B(n24031), .X(n24171) );
  nand_x1_sg U46947 ( .A(n24162), .B(n24163), .X(n24159) );
  nand_x1_sg U46948 ( .A(n8752), .B(n24161), .X(n24160) );
  inv_x1_sg U46949 ( .A(n24156), .X(n50594) );
  inv_x1_sg U46950 ( .A(n22028), .X(n50520) );
  inv_x1_sg U46951 ( .A(n22645), .X(n50527) );
  nand_x1_sg U46952 ( .A(n8672), .B(n23823), .X(n23822) );
  inv_x1_sg U46953 ( .A(n23557), .X(n50536) );
  inv_x1_sg U46954 ( .A(n22305), .X(n50526) );
  nand_x1_sg U46955 ( .A(n8532), .B(n22304), .X(n22303) );
  inv_x2_sg U46956 ( .A(n22119), .X(n44598) );
  nor_x1_sg U46957 ( .A(n22121), .B(n50523), .X(n22119) );
  inv_x1_sg U46958 ( .A(n22896), .X(n50529) );
  inv_x1_sg U46959 ( .A(n23230), .X(n50535) );
  nand_x1_sg U46960 ( .A(n8612), .B(n23229), .X(n23228) );
  inv_x2_sg U46961 ( .A(n22987), .X(n44600) );
  nor_x1_sg U46962 ( .A(n22989), .B(n50532), .X(n22987) );
  inv_x1_sg U46963 ( .A(n24281), .X(n50547) );
  nand_x1_sg U46964 ( .A(n8732), .B(n24169), .X(n24280) );
  nand_x1_sg U46965 ( .A(n8712), .B(n24138), .X(n24137) );
  nand_x2_sg U46966 ( .A(n24271), .B(n24272), .X(n24266) );
  inv_x2_sg U46967 ( .A(n24267), .X(n45588) );
  inv_x1_sg U46968 ( .A(n22031), .X(n50473) );
  inv_x1_sg U46969 ( .A(n22648), .X(n50480) );
  nand_x1_sg U46970 ( .A(n8673), .B(n23817), .X(n23816) );
  inv_x1_sg U46971 ( .A(n23560), .X(n50489) );
  inv_x1_sg U46972 ( .A(n22299), .X(n50479) );
  nand_x1_sg U46973 ( .A(n8533), .B(n22298), .X(n22297) );
  inv_x2_sg U46974 ( .A(n22112), .X(n44594) );
  nor_x1_sg U46975 ( .A(n22114), .B(n50476), .X(n22112) );
  inv_x1_sg U46976 ( .A(n22899), .X(n50482) );
  inv_x1_sg U46977 ( .A(n23224), .X(n50488) );
  nand_x1_sg U46978 ( .A(n8613), .B(n23223), .X(n23222) );
  inv_x2_sg U46979 ( .A(n22980), .X(n44596) );
  nor_x1_sg U46980 ( .A(n22982), .B(n50485), .X(n22980) );
  inv_x1_sg U46981 ( .A(n24257), .X(n50500) );
  nand_x1_sg U46982 ( .A(n8733), .B(n24256), .X(n24255) );
  nand_x1_sg U46983 ( .A(n8713), .B(n24131), .X(n24130) );
  nand_x1_sg U46984 ( .A(n8754), .B(n24379), .X(n24378) );
  nand_x1_sg U46985 ( .A(n24358), .B(n24362), .X(n24377) );
  inv_x1_sg U46986 ( .A(n24374), .X(n50503) );
  inv_x1_sg U46987 ( .A(n22034), .X(n50427) );
  inv_x1_sg U46988 ( .A(n22651), .X(n50434) );
  nand_x1_sg U46989 ( .A(n8674), .B(n23811), .X(n23810) );
  inv_x1_sg U46990 ( .A(n23563), .X(n50443) );
  inv_x1_sg U46991 ( .A(n22293), .X(n50433) );
  nand_x1_sg U46992 ( .A(n8534), .B(n22292), .X(n22291) );
  inv_x2_sg U46993 ( .A(n22105), .X(n44590) );
  nor_x1_sg U46994 ( .A(n22107), .B(n50430), .X(n22105) );
  inv_x1_sg U46995 ( .A(n22902), .X(n50436) );
  inv_x1_sg U46996 ( .A(n23218), .X(n50442) );
  nand_x1_sg U46997 ( .A(n8614), .B(n23217), .X(n23216) );
  inv_x2_sg U46998 ( .A(n22973), .X(n44592) );
  nor_x1_sg U46999 ( .A(n22975), .B(n50439), .X(n22973) );
  inv_x1_sg U47000 ( .A(n24251), .X(n50454) );
  nand_x1_sg U47001 ( .A(n8734), .B(n24250), .X(n24249) );
  nand_x1_sg U47002 ( .A(n8714), .B(n24124), .X(n24123) );
  nand_x1_sg U47003 ( .A(n8755), .B(n24382), .X(n24381) );
  nand_x1_sg U47004 ( .A(n8774), .B(n40799), .X(n24468) );
  nand_x1_sg U47005 ( .A(out_L2[8]), .B(n40800), .X(n24469) );
  inv_x1_sg U47006 ( .A(n22037), .X(n50380) );
  inv_x1_sg U47007 ( .A(n22654), .X(n50387) );
  nand_x1_sg U47008 ( .A(n8675), .B(n23805), .X(n23804) );
  inv_x1_sg U47009 ( .A(n23566), .X(n50396) );
  inv_x1_sg U47010 ( .A(n22287), .X(n50386) );
  nand_x1_sg U47011 ( .A(n8535), .B(n22286), .X(n22285) );
  inv_x2_sg U47012 ( .A(n22098), .X(n44586) );
  nor_x1_sg U47013 ( .A(n22100), .B(n50383), .X(n22098) );
  inv_x1_sg U47014 ( .A(n22905), .X(n50389) );
  inv_x1_sg U47015 ( .A(n23212), .X(n50395) );
  nand_x1_sg U47016 ( .A(n8615), .B(n23211), .X(n23210) );
  inv_x2_sg U47017 ( .A(n22966), .X(n44588) );
  nor_x1_sg U47018 ( .A(n22968), .B(n50392), .X(n22966) );
  inv_x1_sg U47019 ( .A(n24245), .X(n50408) );
  nand_x1_sg U47020 ( .A(n8735), .B(n24244), .X(n24243) );
  nand_x1_sg U47021 ( .A(n8715), .B(n24117), .X(n24116) );
  inv_x2_sg U47022 ( .A(n24451), .X(n44298) );
  nand_x1_sg U47023 ( .A(n8755), .B(n24355), .X(n24354) );
  inv_x1_sg U47024 ( .A(n23206), .X(n50348) );
  nand_x1_sg U47025 ( .A(n8616), .B(n23205), .X(n23204) );
  nand_x1_sg U47026 ( .A(n8596), .B(n22963), .X(n22962) );
  inv_x1_sg U47027 ( .A(n22908), .X(n50342) );
  nand_x1_sg U47028 ( .A(n8676), .B(n23799), .X(n23798) );
  inv_x1_sg U47029 ( .A(n22040), .X(n50333) );
  nand_x1_sg U47030 ( .A(n8556), .B(n22437), .X(n22436) );
  inv_x1_sg U47031 ( .A(n23569), .X(n50349) );
  inv_x1_sg U47032 ( .A(n22281), .X(n50339) );
  nand_x1_sg U47033 ( .A(n8536), .B(n22280), .X(n22279) );
  inv_x2_sg U47034 ( .A(n22091), .X(n44584) );
  nor_x1_sg U47035 ( .A(n22093), .B(n50336), .X(n22091) );
  inv_x1_sg U47036 ( .A(n24239), .X(n50360) );
  nand_x1_sg U47037 ( .A(n8736), .B(n24238), .X(n24237) );
  nand_x1_sg U47038 ( .A(n8716), .B(n24110), .X(n24109) );
  inv_x1_sg U47039 ( .A(n22043), .X(n50287) );
  inv_x1_sg U47040 ( .A(n22660), .X(n50294) );
  nand_x1_sg U47041 ( .A(n8677), .B(n23793), .X(n23792) );
  inv_x1_sg U47042 ( .A(n23572), .X(n50303) );
  inv_x1_sg U47043 ( .A(n22275), .X(n50293) );
  nand_x1_sg U47044 ( .A(n8537), .B(n22274), .X(n22273) );
  inv_x2_sg U47045 ( .A(n22084), .X(n44580) );
  nor_x1_sg U47046 ( .A(n22086), .B(n50290), .X(n22084) );
  inv_x1_sg U47047 ( .A(n22911), .X(n50296) );
  inv_x1_sg U47048 ( .A(n23200), .X(n50302) );
  nand_x1_sg U47049 ( .A(n8617), .B(n23199), .X(n23198) );
  inv_x2_sg U47050 ( .A(n22952), .X(n44582) );
  nor_x1_sg U47051 ( .A(n22954), .B(n50299), .X(n22952) );
  inv_x1_sg U47052 ( .A(n24233), .X(n50314) );
  nand_x1_sg U47053 ( .A(n8737), .B(n24232), .X(n24231) );
  nand_x1_sg U47054 ( .A(n8717), .B(n24103), .X(n24102) );
  nand_x1_sg U47055 ( .A(n8757), .B(n24342), .X(n24341) );
  inv_x1_sg U47056 ( .A(n23194), .X(n50256) );
  nand_x1_sg U47057 ( .A(n8618), .B(n23193), .X(n23192) );
  nand_x1_sg U47058 ( .A(n8598), .B(n22949), .X(n22948) );
  inv_x1_sg U47059 ( .A(n22914), .X(n50250) );
  inv_x1_sg U47060 ( .A(n22046), .X(n50241) );
  nand_x1_sg U47061 ( .A(n8558), .B(n22425), .X(n22424) );
  inv_x1_sg U47062 ( .A(n23575), .X(n50257) );
  inv_x1_sg U47063 ( .A(n22269), .X(n50247) );
  nand_x1_sg U47064 ( .A(n8538), .B(n22268), .X(n22267) );
  inv_x2_sg U47065 ( .A(n22077), .X(n44578) );
  nor_x1_sg U47066 ( .A(n22079), .B(n50244), .X(n22077) );
  nand_x1_sg U47067 ( .A(n8678), .B(n23787), .X(n23786) );
  inv_x1_sg U47068 ( .A(n24061), .X(n50263) );
  inv_x1_sg U47069 ( .A(n24227), .X(n50269) );
  nand_x1_sg U47070 ( .A(n8738), .B(n24226), .X(n24225) );
  nand_x1_sg U47071 ( .A(n8718), .B(n24096), .X(n24095) );
  inv_x1_sg U47072 ( .A(n23188), .X(n50212) );
  nand_x1_sg U47073 ( .A(n8619), .B(n23187), .X(n23186) );
  nand_x1_sg U47074 ( .A(n8599), .B(n22942), .X(n22941) );
  inv_x1_sg U47075 ( .A(n22917), .X(n50206) );
  inv_x1_sg U47076 ( .A(n22049), .X(n50197) );
  nand_x1_sg U47077 ( .A(n8559), .B(n22419), .X(n22418) );
  inv_x1_sg U47078 ( .A(n23578), .X(n50213) );
  inv_x1_sg U47079 ( .A(n22263), .X(n50203) );
  nand_x1_sg U47080 ( .A(n8539), .B(n22262), .X(n22261) );
  inv_x2_sg U47081 ( .A(n22070), .X(n44576) );
  nor_x1_sg U47082 ( .A(n22072), .B(n50200), .X(n22070) );
  nand_x1_sg U47083 ( .A(n8679), .B(n23781), .X(n23780) );
  nand_x1_sg U47084 ( .A(n8660), .B(n23759), .X(n23758) );
  inv_x1_sg U47085 ( .A(n24064), .X(n50218) );
  inv_x1_sg U47086 ( .A(n24221), .X(n50224) );
  nand_x1_sg U47087 ( .A(n8739), .B(n24220), .X(n24219) );
  nand_x1_sg U47088 ( .A(n8719), .B(n24089), .X(n24088) );
  inv_x1_sg U47089 ( .A(n23182), .X(n50165) );
  nand_x1_sg U47090 ( .A(n8620), .B(n23181), .X(n23180) );
  nand_x1_sg U47091 ( .A(n8600), .B(n22935), .X(n22934) );
  nand_x1_sg U47092 ( .A(n8560), .B(n22413), .X(n22412) );
  inv_x1_sg U47093 ( .A(n22257), .X(n50159) );
  nand_x1_sg U47094 ( .A(n8540), .B(n22256), .X(n22255) );
  inv_x2_sg U47095 ( .A(n22063), .X(n44069) );
  nor_x1_sg U47096 ( .A(n22065), .B(n50157), .X(n22063) );
  inv_x1_sg U47097 ( .A(n24215), .X(n50175) );
  nand_x1_sg U47098 ( .A(n8740), .B(n24214), .X(n24213) );
  nand_x1_sg U47099 ( .A(n8720), .B(n24082), .X(n24081) );
  nand_x1_sg U47100 ( .A(n8680), .B(n23775), .X(n23774) );
  nand_x2_sg U47101 ( .A(n50181), .B(n24412), .X(n24410) );
  inv_x1_sg U47102 ( .A(n24413), .X(n50181) );
  nand_x1_sg U47103 ( .A(n8760), .B(n24323), .X(n24322) );
  nand_x2_sg U47104 ( .A(n23174), .B(n23175), .X(n23173) );
  nand_x2_sg U47105 ( .A(n22926), .B(n22927), .X(n22925) );
  nand_x2_sg U47106 ( .A(n24406), .B(n24407), .X(n24405) );
  nand_x2_sg U47107 ( .A(n22405), .B(n22406), .X(n22404) );
  nand_x2_sg U47108 ( .A(n22058), .B(n22059), .X(n22057) );
  nand_x2_sg U47109 ( .A(n22249), .B(n22250), .X(n22248) );
  nand_x1_sg U47110 ( .A(n10197), .B(n50133), .X(n23386) );
  nand_x1_sg U47111 ( .A(n23387), .B(n50147), .X(n23385) );
  inv_x1_sg U47112 ( .A(n23387), .X(n50133) );
  nand_x2_sg U47113 ( .A(n24207), .B(n24208), .X(n24206) );
  nand_x2_sg U47114 ( .A(n24314), .B(n24315), .X(n24313) );
  nand_x1_sg U47115 ( .A(n25663), .B(n51254), .X(n25662) );
  inv_x2_sg U47116 ( .A(n25600), .X(n44256) );
  nor_x1_sg U47117 ( .A(n25601), .B(n25602), .X(n25600) );
  nand_x1_sg U47118 ( .A(n51309), .B(n10397), .X(n10477) );
  nand_x1_sg U47119 ( .A(n10461), .B(n51293), .X(n10460) );
  inv_x2_sg U47120 ( .A(n10544), .X(n44306) );
  inv_x1_sg U47121 ( .A(n10576), .X(n51348) );
  nand_x1_sg U47122 ( .A(n10538), .B(n10572), .X(n10571) );
  nand_x1_sg U47123 ( .A(n51287), .B(n51299), .X(n10572) );
  nand_x1_sg U47124 ( .A(n10488), .B(n46567), .X(n10487) );
  nand_x1_sg U47125 ( .A(n10491), .B(n51306), .X(n10486) );
  inv_x2_sg U47126 ( .A(n10563), .X(n44426) );
  nor_x1_sg U47127 ( .A(n10602), .B(n10603), .X(n10563) );
  inv_x1_sg U47128 ( .A(n10583), .X(n51367) );
  inv_x1_sg U47129 ( .A(n10745), .X(n51437) );
  nand_x1_sg U47130 ( .A(n51390), .B(n40541), .X(n10729) );
  inv_x1_sg U47131 ( .A(n10663), .X(n51398) );
  inv_x1_sg U47132 ( .A(n10643), .X(n51400) );
  nand_x1_sg U47133 ( .A(n40542), .B(n10709), .X(n10706) );
  nand_x2_sg U47134 ( .A(n10774), .B(n10795), .X(n10722) );
  nand_x1_sg U47135 ( .A(n10796), .B(n51449), .X(n10795) );
  inv_x1_sg U47136 ( .A(n10797), .X(n51449) );
  inv_x1_sg U47137 ( .A(n10722), .X(n51450) );
  nand_x4_sg U47138 ( .A(n10971), .B(n10972), .X(n10883) );
  nand_x1_sg U47139 ( .A(n51489), .B(n42053), .X(n10971) );
  nand_x1_sg U47140 ( .A(n42054), .B(n10974), .X(n10972) );
  inv_x1_sg U47141 ( .A(n10974), .X(n51489) );
  nand_x1_sg U47142 ( .A(n51483), .B(n10977), .X(n10975) );
  inv_x1_sg U47143 ( .A(n10976), .X(n51483) );
  nand_x1_sg U47144 ( .A(n10818), .B(n10819), .X(n10816) );
  inv_x1_sg U47145 ( .A(n10818), .X(n51454) );
  inv_x1_sg U47146 ( .A(n10773), .X(n51468) );
  nand_x1_sg U47147 ( .A(n10757), .B(n10758), .X(n10755) );
  inv_x1_sg U47148 ( .A(n10757), .X(n51414) );
  nand_x1_sg U47149 ( .A(n51438), .B(n10682), .X(n10728) );
  nand_x4_sg U47150 ( .A(n10827), .B(n10828), .X(n10773) );
  nand_x1_sg U47151 ( .A(n51467), .B(n10757), .X(n10828) );
  inv_x1_sg U47152 ( .A(n10959), .X(n51443) );
  inv_x1_sg U47153 ( .A(n10361), .X(n51445) );
  inv_x1_sg U47154 ( .A(n10894), .X(n51518) );
  inv_x1_sg U47155 ( .A(n10962), .X(n51513) );
  inv_x2_sg U47156 ( .A(n10927), .X(n44332) );
  nor_x1_sg U47157 ( .A(n10929), .B(n10930), .X(n10927) );
  nand_x1_sg U47158 ( .A(n25942), .B(n51530), .X(n25941) );
  inv_x2_sg U47159 ( .A(n25881), .X(n44258) );
  nor_x1_sg U47160 ( .A(n25882), .B(n25883), .X(n25881) );
  nand_x1_sg U47161 ( .A(n46540), .B(n46547), .X(n11195) );
  nor_x1_sg U47162 ( .A(n51543), .B(n51562), .X(n11196) );
  nand_x4_sg U47163 ( .A(n46539), .B(n46547), .X(n11216) );
  inv_x2_sg U47164 ( .A(n11311), .X(n44420) );
  nor_x1_sg U47165 ( .A(n11348), .B(n11349), .X(n11311) );
  inv_x1_sg U47166 ( .A(n11323), .X(n51631) );
  inv_x2_sg U47167 ( .A(n11359), .X(n45550) );
  nor_x1_sg U47168 ( .A(n51651), .B(n11380), .X(n11359) );
  inv_x1_sg U47169 ( .A(n11357), .X(n51638) );
  nand_x1_sg U47170 ( .A(n11421), .B(n51677), .X(n11420) );
  inv_x1_sg U47171 ( .A(n11422), .X(n51677) );
  nand_x4_sg U47172 ( .A(n46532), .B(n51543), .X(n11417) );
  inv_x1_sg U47173 ( .A(n11414), .X(n51698) );
  nand_x1_sg U47174 ( .A(n51686), .B(n51667), .X(n11517) );
  inv_x1_sg U47175 ( .A(n11518), .X(n51686) );
  nand_x1_sg U47176 ( .A(n51665), .B(n11436), .X(n11435) );
  inv_x1_sg U47177 ( .A(n11423), .X(n51665) );
  inv_x1_sg U47178 ( .A(n11490), .X(n51705) );
  inv_x1_sg U47179 ( .A(n11467), .X(n51696) );
  nand_x2_sg U47180 ( .A(n11556), .B(n11576), .X(n11503) );
  nand_x1_sg U47181 ( .A(n11577), .B(n51728), .X(n11576) );
  inv_x1_sg U47182 ( .A(n11578), .X(n51728) );
  inv_x1_sg U47183 ( .A(n11503), .X(n51729) );
  inv_x1_sg U47184 ( .A(n11662), .X(n45452) );
  inv_x1_sg U47185 ( .A(n11552), .X(n51748) );
  nand_x1_sg U47186 ( .A(n51719), .B(n51711), .X(n11508) );
  inv_x1_sg U47187 ( .A(n11128), .X(n51735) );
  nand_x4_sg U47188 ( .A(n11607), .B(n11608), .X(n11552) );
  nand_x1_sg U47189 ( .A(n51747), .B(n40543), .X(n11608) );
  inv_x1_sg U47190 ( .A(n11714), .X(n51782) );
  inv_x1_sg U47191 ( .A(n11696), .X(n51762) );
  inv_x2_sg U47192 ( .A(n11671), .X(n44340) );
  nor_x1_sg U47193 ( .A(n51799), .B(n11673), .X(n11671) );
  nand_x1_sg U47194 ( .A(n26222), .B(n51812), .X(n26221) );
  inv_x2_sg U47195 ( .A(n26161), .X(n44276) );
  nor_x1_sg U47196 ( .A(n26162), .B(n26163), .X(n26161) );
  nor_x1_sg U47197 ( .A(n51826), .B(n51840), .X(n11975) );
  nand_x1_sg U47198 ( .A(n51868), .B(n11947), .X(n12031) );
  nand_x1_sg U47199 ( .A(n12029), .B(n51846), .X(n12028) );
  nand_x2_sg U47200 ( .A(n51854), .B(n11833), .X(n12015) );
  inv_x2_sg U47201 ( .A(n12091), .X(n44151) );
  nor_x1_sg U47202 ( .A(n12128), .B(n12129), .X(n12091) );
  nand_x1_sg U47203 ( .A(n12041), .B(n51826), .X(n12040) );
  inv_x1_sg U47204 ( .A(n12103), .X(n51912) );
  inv_x2_sg U47205 ( .A(n12139), .X(n45548) );
  nor_x1_sg U47206 ( .A(n51932), .B(n12160), .X(n12139) );
  inv_x1_sg U47207 ( .A(n12137), .X(n51919) );
  nand_x1_sg U47208 ( .A(n12201), .B(n51958), .X(n12200) );
  inv_x1_sg U47209 ( .A(n12202), .X(n51958) );
  nand_x1_sg U47210 ( .A(n51946), .B(n12216), .X(n12215) );
  inv_x1_sg U47211 ( .A(n12203), .X(n51946) );
  nand_x4_sg U47212 ( .A(n12225), .B(n51967), .X(n12190) );
  inv_x1_sg U47213 ( .A(n12226), .X(n51967) );
  nand_x1_sg U47214 ( .A(n12308), .B(n51990), .X(n12305) );
  nand_x1_sg U47215 ( .A(n12307), .B(n51997), .X(n12306) );
  inv_x1_sg U47216 ( .A(n12307), .X(n51990) );
  nand_x1_sg U47217 ( .A(n43308), .B(n12270), .X(n12267) );
  nand_x2_sg U47218 ( .A(n12336), .B(n12357), .X(n12283) );
  nand_x1_sg U47219 ( .A(n12358), .B(n52006), .X(n12357) );
  inv_x1_sg U47220 ( .A(n12359), .X(n52006) );
  inv_x1_sg U47221 ( .A(n12283), .X(n52007) );
  inv_x1_sg U47222 ( .A(n11915), .X(n52031) );
  nand_x1_sg U47223 ( .A(n52023), .B(n12536), .X(n12535) );
  nand_x1_sg U47224 ( .A(n52048), .B(n12537), .X(n12534) );
  inv_x1_sg U47225 ( .A(n12537), .X(n52023) );
  inv_x1_sg U47226 ( .A(n12332), .X(n52030) );
  nand_x1_sg U47227 ( .A(n12308), .B(n12307), .X(n12288) );
  inv_x1_sg U47228 ( .A(n11911), .X(n52013) );
  nand_x4_sg U47229 ( .A(n12388), .B(n12389), .X(n12332) );
  nand_x1_sg U47230 ( .A(n52029), .B(n40544), .X(n12389) );
  inv_x1_sg U47231 ( .A(n12494), .X(n52062) );
  inv_x1_sg U47232 ( .A(n12475), .X(n52043) );
  inv_x2_sg U47233 ( .A(n12451), .X(n44338) );
  nor_x1_sg U47234 ( .A(n52075), .B(n12453), .X(n12451) );
  nand_x1_sg U47235 ( .A(n26501), .B(n52088), .X(n26500) );
  inv_x2_sg U47236 ( .A(n26440), .X(n44274) );
  nor_x1_sg U47237 ( .A(n26441), .B(n26442), .X(n26440) );
  nand_x1_sg U47238 ( .A(n46496), .B(n46503), .X(n12756) );
  nor_x1_sg U47239 ( .A(n52100), .B(n52119), .X(n12757) );
  nand_x4_sg U47240 ( .A(n46495), .B(n46503), .X(n12777) );
  inv_x1_sg U47241 ( .A(n12884), .X(n52188) );
  inv_x2_sg U47242 ( .A(n12920), .X(n45546) );
  nor_x1_sg U47243 ( .A(n52207), .B(n12941), .X(n12920) );
  inv_x1_sg U47244 ( .A(n12918), .X(n52194) );
  nand_x1_sg U47245 ( .A(n12982), .B(n52233), .X(n12981) );
  inv_x1_sg U47246 ( .A(n12983), .X(n52233) );
  nand_x4_sg U47247 ( .A(n46488), .B(n52100), .X(n12978) );
  inv_x1_sg U47248 ( .A(n12975), .X(n52254) );
  nand_x1_sg U47249 ( .A(n52241), .B(n52223), .X(n13078) );
  inv_x1_sg U47250 ( .A(n13079), .X(n52241) );
  nand_x1_sg U47251 ( .A(n52221), .B(n12997), .X(n12996) );
  inv_x1_sg U47252 ( .A(n12984), .X(n52221) );
  inv_x1_sg U47253 ( .A(n13051), .X(n52261) );
  inv_x1_sg U47254 ( .A(n13028), .X(n52252) );
  nand_x2_sg U47255 ( .A(n13117), .B(n13137), .X(n13064) );
  nand_x1_sg U47256 ( .A(n13138), .B(n52284), .X(n13137) );
  inv_x1_sg U47257 ( .A(n13139), .X(n52284) );
  inv_x1_sg U47258 ( .A(n13064), .X(n52285) );
  nand_x1_sg U47259 ( .A(n40533), .B(n13160), .X(n13157) );
  inv_x1_sg U47260 ( .A(n12693), .X(n52306) );
  inv_x1_sg U47261 ( .A(n13316), .X(n52325) );
  nand_x1_sg U47262 ( .A(n52273), .B(n52267), .X(n13069) );
  inv_x1_sg U47263 ( .A(n12689), .X(n52290) );
  nand_x4_sg U47264 ( .A(n13156), .B(n13195), .X(n13193) );
  nand_x1_sg U47265 ( .A(n52156), .B(n13155), .X(n13195) );
  inv_x2_sg U47266 ( .A(n13113), .X(n44412) );
  nor_x1_sg U47267 ( .A(n13191), .B(n13192), .X(n13113) );
  nand_x4_sg U47268 ( .A(n13168), .B(n13169), .X(n13112) );
  nand_x1_sg U47269 ( .A(n52304), .B(n40546), .X(n13169) );
  inv_x1_sg U47270 ( .A(n13275), .X(n52339) );
  inv_x1_sg U47271 ( .A(n13256), .X(n52319) );
  inv_x2_sg U47272 ( .A(n13232), .X(n43970) );
  nor_x1_sg U47273 ( .A(n52353), .B(n13234), .X(n13232) );
  nand_x1_sg U47274 ( .A(n26779), .B(n52365), .X(n26778) );
  inv_x2_sg U47275 ( .A(n26718), .X(n44268) );
  nor_x1_sg U47276 ( .A(n26719), .B(n26720), .X(n26718) );
  nor_x1_sg U47277 ( .A(n52378), .B(n52392), .X(n13536) );
  nand_x1_sg U47278 ( .A(n46474), .B(n46481), .X(n13535) );
  nand_x1_sg U47279 ( .A(n52420), .B(n46477), .X(n13596) );
  nand_x1_sg U47280 ( .A(n13594), .B(n52398), .X(n13593) );
  nand_x2_sg U47281 ( .A(n52406), .B(n46481), .X(n13576) );
  nand_x1_sg U47282 ( .A(n13602), .B(n46474), .X(n13601) );
  inv_x1_sg U47283 ( .A(n13664), .X(n52464) );
  inv_x2_sg U47284 ( .A(n13654), .X(n44073) );
  nor_x1_sg U47285 ( .A(n13625), .B(n13656), .X(n13654) );
  inv_x2_sg U47286 ( .A(n13700), .X(n45544) );
  nor_x1_sg U47287 ( .A(n52484), .B(n13721), .X(n13700) );
  inv_x1_sg U47288 ( .A(n13698), .X(n52471) );
  nand_x1_sg U47289 ( .A(n13762), .B(n52510), .X(n13761) );
  inv_x1_sg U47290 ( .A(n13763), .X(n52510) );
  nand_x4_sg U47291 ( .A(n52447), .B(n52378), .X(n13758) );
  inv_x1_sg U47292 ( .A(n13755), .X(n52530) );
  nand_x1_sg U47293 ( .A(n52498), .B(n13777), .X(n13776) );
  inv_x1_sg U47294 ( .A(n13764), .X(n52498) );
  nand_x4_sg U47295 ( .A(n13786), .B(n52518), .X(n13751) );
  inv_x1_sg U47296 ( .A(n13787), .X(n52518) );
  inv_x1_sg U47297 ( .A(n13831), .X(n52537) );
  inv_x1_sg U47298 ( .A(n13808), .X(n52528) );
  nand_x2_sg U47299 ( .A(n13897), .B(n13917), .X(n13844) );
  nand_x1_sg U47300 ( .A(n13918), .B(n52559), .X(n13917) );
  inv_x1_sg U47301 ( .A(n13919), .X(n52559) );
  inv_x1_sg U47302 ( .A(n13844), .X(n52560) );
  nand_x1_sg U47303 ( .A(n40534), .B(n13940), .X(n13937) );
  inv_x1_sg U47304 ( .A(n13477), .X(n52581) );
  inv_x1_sg U47305 ( .A(n14096), .X(n52600) );
  nand_x1_sg U47306 ( .A(n52548), .B(n52543), .X(n13849) );
  inv_x1_sg U47307 ( .A(n13473), .X(n52565) );
  nand_x4_sg U47308 ( .A(n13936), .B(n13975), .X(n13973) );
  nand_x1_sg U47309 ( .A(n52430), .B(n13935), .X(n13975) );
  inv_x2_sg U47310 ( .A(n13893), .X(n44410) );
  nor_x1_sg U47311 ( .A(n13971), .B(n13972), .X(n13893) );
  nand_x4_sg U47312 ( .A(n13948), .B(n13949), .X(n13892) );
  nand_x1_sg U47313 ( .A(n52579), .B(n40548), .X(n13949) );
  inv_x1_sg U47314 ( .A(n14055), .X(n52614) );
  inv_x1_sg U47315 ( .A(n14036), .X(n52594) );
  inv_x2_sg U47316 ( .A(n14012), .X(n43968) );
  nor_x1_sg U47317 ( .A(n52628), .B(n14014), .X(n14012) );
  nand_x1_sg U47318 ( .A(n27058), .B(n52641), .X(n27057) );
  inv_x2_sg U47319 ( .A(n26997), .X(n44264) );
  nor_x1_sg U47320 ( .A(n26998), .B(n26999), .X(n26997) );
  nand_x1_sg U47321 ( .A(n52698), .B(n14289), .X(n14369) );
  nand_x1_sg U47322 ( .A(n14353), .B(n52683), .X(n14352) );
  inv_x2_sg U47323 ( .A(n14437), .X(n44750) );
  inv_x2_sg U47324 ( .A(n14412), .X(n44714) );
  inv_x1_sg U47325 ( .A(n14468), .X(n52738) );
  nand_x1_sg U47326 ( .A(n14431), .B(n14464), .X(n14463) );
  nand_x1_sg U47327 ( .A(n14380), .B(n46450), .X(n14379) );
  nand_x1_sg U47328 ( .A(n14383), .B(n52695), .X(n14378) );
  inv_x1_sg U47329 ( .A(n14475), .X(n52744) );
  nand_x1_sg U47330 ( .A(n14534), .B(n52789), .X(n14533) );
  inv_x1_sg U47331 ( .A(n14535), .X(n52789) );
  inv_x1_sg U47332 ( .A(n14637), .X(n52826) );
  nand_x1_sg U47333 ( .A(n52779), .B(n14630), .X(n14621) );
  nand_x4_sg U47334 ( .A(n14557), .B(n52798), .X(n14523) );
  inv_x1_sg U47335 ( .A(n14558), .X(n52798) );
  nand_x1_sg U47336 ( .A(n43344), .B(n14601), .X(n14598) );
  nand_x2_sg U47337 ( .A(n14666), .B(n14687), .X(n14614) );
  inv_x1_sg U47338 ( .A(n14614), .X(n52841) );
  inv_x1_sg U47339 ( .A(n14662), .X(n52857) );
  nand_x1_sg U47340 ( .A(n52827), .B(n14574), .X(n14620) );
  inv_x1_sg U47341 ( .A(n14252), .X(n52835) );
  nand_x1_sg U47342 ( .A(n52856), .B(n40551), .X(n14720) );
  inv_x1_sg U47343 ( .A(n14826), .X(n52892) );
  inv_x1_sg U47344 ( .A(n14808), .X(n52871) );
  inv_x2_sg U47345 ( .A(n14783), .X(n44336) );
  nor_x1_sg U47346 ( .A(n52909), .B(n14785), .X(n14783) );
  inv_x1_sg U47347 ( .A(n14716), .X(n52897) );
  inv_x2_sg U47348 ( .A(n14713), .X(n45446) );
  nor_x1_sg U47349 ( .A(n14773), .B(n45449), .X(n14713) );
  nand_x1_sg U47350 ( .A(n27338), .B(n52922), .X(n27337) );
  inv_x2_sg U47351 ( .A(n27277), .X(n44272) );
  nor_x1_sg U47352 ( .A(n27278), .B(n27279), .X(n27277) );
  nand_x1_sg U47353 ( .A(n46428), .B(n46435), .X(n15089) );
  nor_x1_sg U47354 ( .A(n52934), .B(n52953), .X(n15090) );
  nand_x4_sg U47355 ( .A(n46427), .B(n46435), .X(n15110) );
  inv_x1_sg U47356 ( .A(n15217), .X(n53022) );
  inv_x2_sg U47357 ( .A(n15253), .X(n45542) );
  nor_x1_sg U47358 ( .A(n53041), .B(n15274), .X(n15253) );
  inv_x1_sg U47359 ( .A(n15251), .X(n53028) );
  nand_x1_sg U47360 ( .A(n15315), .B(n53067), .X(n15314) );
  inv_x1_sg U47361 ( .A(n15316), .X(n53067) );
  nand_x4_sg U47362 ( .A(n46420), .B(n52934), .X(n15311) );
  inv_x1_sg U47363 ( .A(n15308), .X(n53088) );
  nand_x1_sg U47364 ( .A(n53075), .B(n53057), .X(n15411) );
  inv_x1_sg U47365 ( .A(n15412), .X(n53075) );
  nand_x1_sg U47366 ( .A(n53055), .B(n15330), .X(n15329) );
  inv_x1_sg U47367 ( .A(n15317), .X(n53055) );
  inv_x1_sg U47368 ( .A(n15384), .X(n53095) );
  inv_x1_sg U47369 ( .A(n15361), .X(n53086) );
  nand_x2_sg U47370 ( .A(n15450), .B(n15470), .X(n15397) );
  nand_x1_sg U47371 ( .A(n15471), .B(n53118), .X(n15470) );
  inv_x1_sg U47372 ( .A(n15472), .X(n53118) );
  inv_x1_sg U47373 ( .A(n15397), .X(n53119) );
  nand_x1_sg U47374 ( .A(n40535), .B(n15493), .X(n15490) );
  inv_x1_sg U47375 ( .A(n15026), .X(n53140) );
  inv_x1_sg U47376 ( .A(n15649), .X(n53159) );
  nand_x1_sg U47377 ( .A(n53107), .B(n53101), .X(n15402) );
  inv_x1_sg U47378 ( .A(n15022), .X(n53124) );
  nand_x4_sg U47379 ( .A(n15489), .B(n15528), .X(n15526) );
  nand_x1_sg U47380 ( .A(n52990), .B(n15488), .X(n15528) );
  inv_x2_sg U47381 ( .A(n15446), .X(n44408) );
  nor_x1_sg U47382 ( .A(n15524), .B(n15525), .X(n15446) );
  nand_x4_sg U47383 ( .A(n15501), .B(n15502), .X(n15445) );
  nand_x1_sg U47384 ( .A(n53138), .B(n40552), .X(n15502) );
  inv_x1_sg U47385 ( .A(n15608), .X(n53173) );
  inv_x1_sg U47386 ( .A(n15589), .X(n53153) );
  inv_x2_sg U47387 ( .A(n15565), .X(n43966) );
  nor_x1_sg U47388 ( .A(n53187), .B(n15567), .X(n15565) );
  nand_x1_sg U47389 ( .A(n27617), .B(n53200), .X(n27616) );
  inv_x2_sg U47390 ( .A(n27556), .X(n44260) );
  nor_x1_sg U47391 ( .A(n27557), .B(n27558), .X(n27556) );
  nor_x1_sg U47392 ( .A(n53214), .B(n53228), .X(n15870) );
  nand_x1_sg U47393 ( .A(n53255), .B(n15842), .X(n15926) );
  nand_x1_sg U47394 ( .A(n15924), .B(n53232), .X(n15923) );
  nand_x2_sg U47395 ( .A(n53240), .B(n46413), .X(n15910) );
  inv_x2_sg U47396 ( .A(n15986), .X(n44418) );
  nor_x1_sg U47397 ( .A(n16023), .B(n16024), .X(n15986) );
  nand_x1_sg U47398 ( .A(n15936), .B(n46405), .X(n15935) );
  nand_x1_sg U47399 ( .A(n15939), .B(n53253), .X(n15934) );
  nand_x4_sg U47400 ( .A(n46405), .B(n53240), .X(n15941) );
  inv_x1_sg U47401 ( .A(n15998), .X(n53299) );
  inv_x2_sg U47402 ( .A(n16034), .X(n45540) );
  nor_x1_sg U47403 ( .A(n53320), .B(n16055), .X(n16034) );
  inv_x1_sg U47404 ( .A(n16032), .X(n53306) );
  nand_x1_sg U47405 ( .A(n16096), .B(n53346), .X(n16095) );
  inv_x1_sg U47406 ( .A(n16097), .X(n53346) );
  nand_x1_sg U47407 ( .A(n53334), .B(n16111), .X(n16110) );
  inv_x1_sg U47408 ( .A(n16098), .X(n53334) );
  nand_x4_sg U47409 ( .A(n16120), .B(n53356), .X(n16085) );
  inv_x1_sg U47410 ( .A(n16121), .X(n53356) );
  nand_x1_sg U47411 ( .A(n16203), .B(n53378), .X(n16200) );
  nand_x1_sg U47412 ( .A(n16202), .B(n53386), .X(n16201) );
  inv_x1_sg U47413 ( .A(n16202), .X(n53378) );
  nand_x1_sg U47414 ( .A(n42398), .B(n16165), .X(n16162) );
  nand_x2_sg U47415 ( .A(n16231), .B(n16252), .X(n16178) );
  inv_x1_sg U47416 ( .A(n16178), .X(n53398) );
  nand_x4_sg U47417 ( .A(n16429), .B(n16430), .X(n16338) );
  nand_x1_sg U47418 ( .A(n53438), .B(n41865), .X(n16429) );
  nand_x1_sg U47419 ( .A(n41866), .B(n16432), .X(n16430) );
  inv_x1_sg U47420 ( .A(n16432), .X(n53438) );
  nand_x1_sg U47421 ( .A(n53432), .B(n16435), .X(n16433) );
  inv_x1_sg U47422 ( .A(n16434), .X(n53432) );
  inv_x1_sg U47423 ( .A(n16230), .X(n53417) );
  nand_x1_sg U47424 ( .A(n16203), .B(n16202), .X(n16183) );
  nand_x4_sg U47425 ( .A(n16283), .B(n16284), .X(n16230) );
  nand_x1_sg U47426 ( .A(n53416), .B(n40554), .X(n16284) );
  inv_x1_sg U47427 ( .A(n15807), .X(n53405) );
  inv_x1_sg U47428 ( .A(n16349), .X(n53467) );
  inv_x1_sg U47429 ( .A(n16420), .X(n53453) );
  inv_x2_sg U47430 ( .A(n16385), .X(n44330) );
  nor_x1_sg U47431 ( .A(n16387), .B(n16388), .X(n16385) );
  nand_x1_sg U47432 ( .A(n27896), .B(n53480), .X(n27895) );
  inv_x2_sg U47433 ( .A(n27835), .X(n44270) );
  nor_x1_sg U47434 ( .A(n27836), .B(n27837), .X(n27835) );
  nand_x1_sg U47435 ( .A(n46384), .B(n46391), .X(n16655) );
  nor_x1_sg U47436 ( .A(n53492), .B(n53511), .X(n16656) );
  nand_x4_sg U47437 ( .A(n46383), .B(n46391), .X(n16676) );
  inv_x1_sg U47438 ( .A(n16783), .X(n53580) );
  inv_x2_sg U47439 ( .A(n16819), .X(n45538) );
  nor_x1_sg U47440 ( .A(n53599), .B(n16840), .X(n16819) );
  inv_x1_sg U47441 ( .A(n16817), .X(n53586) );
  nand_x1_sg U47442 ( .A(n16881), .B(n53625), .X(n16880) );
  inv_x1_sg U47443 ( .A(n16882), .X(n53625) );
  nand_x4_sg U47444 ( .A(n46376), .B(n53492), .X(n16877) );
  inv_x1_sg U47445 ( .A(n16874), .X(n53646) );
  nand_x1_sg U47446 ( .A(n53633), .B(n53615), .X(n16977) );
  inv_x1_sg U47447 ( .A(n16978), .X(n53633) );
  nand_x1_sg U47448 ( .A(n53613), .B(n16896), .X(n16895) );
  inv_x1_sg U47449 ( .A(n16883), .X(n53613) );
  inv_x1_sg U47450 ( .A(n16950), .X(n53653) );
  inv_x1_sg U47451 ( .A(n16927), .X(n53644) );
  nand_x2_sg U47452 ( .A(n17016), .B(n17036), .X(n16963) );
  nand_x1_sg U47453 ( .A(n17037), .B(n53676), .X(n17036) );
  inv_x1_sg U47454 ( .A(n17038), .X(n53676) );
  inv_x1_sg U47455 ( .A(n16963), .X(n53677) );
  nand_x1_sg U47456 ( .A(n40536), .B(n17059), .X(n17056) );
  inv_x1_sg U47457 ( .A(n16592), .X(n53698) );
  inv_x1_sg U47458 ( .A(n17215), .X(n53717) );
  nand_x1_sg U47459 ( .A(n53665), .B(n53659), .X(n16968) );
  inv_x1_sg U47460 ( .A(n16588), .X(n53682) );
  nand_x4_sg U47461 ( .A(n17055), .B(n17094), .X(n17092) );
  nand_x1_sg U47462 ( .A(n53548), .B(n17054), .X(n17094) );
  inv_x2_sg U47463 ( .A(n17012), .X(n44406) );
  nor_x1_sg U47464 ( .A(n17090), .B(n17091), .X(n17012) );
  nand_x4_sg U47465 ( .A(n17067), .B(n17068), .X(n17011) );
  nand_x1_sg U47466 ( .A(n53696), .B(n40555), .X(n17068) );
  inv_x1_sg U47467 ( .A(n17174), .X(n53731) );
  inv_x1_sg U47468 ( .A(n17155), .X(n53711) );
  inv_x2_sg U47469 ( .A(n17131), .X(n43964) );
  nor_x1_sg U47470 ( .A(n53745), .B(n17133), .X(n17131) );
  nand_x1_sg U47471 ( .A(n28177), .B(n53758), .X(n28176) );
  inv_x2_sg U47472 ( .A(n28116), .X(n44254) );
  nor_x1_sg U47473 ( .A(n28117), .B(n28118), .X(n28116) );
  nand_x1_sg U47474 ( .A(n17476), .B(n53802), .X(n17475) );
  inv_x2_sg U47475 ( .A(n17556), .X(n44756) );
  inv_x1_sg U47476 ( .A(n17588), .X(n53858) );
  nand_x1_sg U47477 ( .A(n17550), .B(n17584), .X(n17583) );
  nand_x1_sg U47478 ( .A(n53796), .B(n53809), .X(n17584) );
  inv_x1_sg U47479 ( .A(n17595), .X(n53864) );
  nand_x1_sg U47480 ( .A(n17655), .B(n53909), .X(n17654) );
  inv_x1_sg U47481 ( .A(n17656), .X(n53909) );
  inv_x1_sg U47482 ( .A(n17758), .X(n53946) );
  nand_x1_sg U47483 ( .A(n53899), .B(n17751), .X(n17742) );
  nand_x4_sg U47484 ( .A(n17678), .B(n53919), .X(n17644) );
  inv_x1_sg U47485 ( .A(n17679), .X(n53919) );
  nand_x1_sg U47486 ( .A(n42434), .B(n17722), .X(n17719) );
  nand_x2_sg U47487 ( .A(n17787), .B(n17808), .X(n17735) );
  inv_x1_sg U47488 ( .A(n17735), .X(n53961) );
  inv_x1_sg U47489 ( .A(n17783), .X(n53977) );
  nand_x1_sg U47490 ( .A(n53947), .B(n17695), .X(n17741) );
  inv_x1_sg U47491 ( .A(n17371), .X(n53955) );
  nand_x1_sg U47492 ( .A(n53976), .B(n40557), .X(n17841) );
  inv_x1_sg U47493 ( .A(n17947), .X(n54012) );
  inv_x1_sg U47494 ( .A(n17929), .X(n53991) );
  inv_x2_sg U47495 ( .A(n17904), .X(n43962) );
  nor_x1_sg U47496 ( .A(n54029), .B(n17906), .X(n17904) );
  inv_x1_sg U47497 ( .A(n17837), .X(n54017) );
  inv_x2_sg U47498 ( .A(n17834), .X(n45442) );
  nor_x1_sg U47499 ( .A(n17894), .B(n45445), .X(n17834) );
  inv_x1_sg U47500 ( .A(n28397), .X(n54048) );
  nand_x1_sg U47501 ( .A(n18243), .B(n54084), .X(n18242) );
  nand_x1_sg U47502 ( .A(n46339), .B(n18258), .X(n18257) );
  nand_x1_sg U47503 ( .A(n54099), .B(n46342), .X(n18258) );
  nand_x1_sg U47504 ( .A(n18304), .B(n18305), .X(n18302) );
  inv_x1_sg U47505 ( .A(n18304), .X(n54092) );
  nand_x1_sg U47506 ( .A(n18293), .B(n54109), .X(n18292) );
  inv_x1_sg U47507 ( .A(n18358), .X(n54138) );
  nand_x1_sg U47508 ( .A(n54091), .B(n54077), .X(n18354) );
  inv_x1_sg U47509 ( .A(n18280), .X(n54132) );
  nand_x1_sg U47510 ( .A(n18272), .B(n46333), .X(n18268) );
  nand_x1_sg U47511 ( .A(n18270), .B(n41711), .X(n18269) );
  inv_x1_sg U47512 ( .A(n18365), .X(n54156) );
  inv_x1_sg U47513 ( .A(n18480), .X(n54213) );
  inv_x1_sg U47514 ( .A(n18526), .X(n54231) );
  nand_x1_sg U47515 ( .A(n54179), .B(n18519), .X(n18511) );
  inv_x1_sg U47516 ( .A(n18445), .X(n54187) );
  inv_x1_sg U47517 ( .A(n18519), .X(n54201) );
  nand_x1_sg U47518 ( .A(n54106), .B(n54110), .X(n18439) );
  inv_x1_sg U47519 ( .A(n18491), .X(n54221) );
  nand_x2_sg U47520 ( .A(n18555), .B(n18575), .X(n18504) );
  nand_x1_sg U47521 ( .A(n18576), .B(n54242), .X(n18575) );
  inv_x1_sg U47522 ( .A(n18577), .X(n54242) );
  inv_x1_sg U47523 ( .A(n18504), .X(n54243) );
  inv_x1_sg U47524 ( .A(n18664), .X(n45440) );
  inv_x1_sg U47525 ( .A(n18551), .X(n54261) );
  nand_x1_sg U47526 ( .A(n18538), .B(n18539), .X(n18536) );
  inv_x1_sg U47527 ( .A(n18538), .X(n54198) );
  nand_x1_sg U47528 ( .A(n54232), .B(n18464), .X(n18510) );
  inv_x2_sg U47529 ( .A(n18648), .X(n44328) );
  nor_x1_sg U47530 ( .A(n54238), .B(n18655), .X(n18648) );
  nand_x4_sg U47531 ( .A(n18607), .B(n18608), .X(n18551) );
  nand_x1_sg U47532 ( .A(n54260), .B(n18538), .X(n18608) );
  inv_x1_sg U47533 ( .A(n18716), .X(n54294) );
  inv_x1_sg U47534 ( .A(n18698), .X(n54274) );
  inv_x2_sg U47535 ( .A(n18673), .X(n44334) );
  nor_x1_sg U47536 ( .A(n54310), .B(n18675), .X(n18673) );
  nand_x1_sg U47537 ( .A(n28735), .B(n54323), .X(n28734) );
  inv_x2_sg U47538 ( .A(n28674), .X(n44252) );
  nor_x1_sg U47539 ( .A(n28675), .B(n28676), .X(n28674) );
  nand_x1_sg U47540 ( .A(n19021), .B(n54367), .X(n19020) );
  inv_x2_sg U47541 ( .A(n19101), .X(n44754) );
  inv_x1_sg U47542 ( .A(n19133), .X(n54423) );
  nand_x1_sg U47543 ( .A(n19095), .B(n19129), .X(n19128) );
  nand_x1_sg U47544 ( .A(n54361), .B(n54374), .X(n19129) );
  inv_x1_sg U47545 ( .A(n19140), .X(n54429) );
  nand_x1_sg U47546 ( .A(n19200), .B(n54474), .X(n19199) );
  inv_x1_sg U47547 ( .A(n19201), .X(n54474) );
  inv_x1_sg U47548 ( .A(n19303), .X(n54511) );
  nand_x1_sg U47549 ( .A(n54464), .B(n19296), .X(n19287) );
  nand_x4_sg U47550 ( .A(n19223), .B(n54484), .X(n19189) );
  inv_x1_sg U47551 ( .A(n19224), .X(n54484) );
  nand_x1_sg U47552 ( .A(n42432), .B(n19267), .X(n19264) );
  nand_x2_sg U47553 ( .A(n19332), .B(n19353), .X(n19280) );
  inv_x1_sg U47554 ( .A(n19280), .X(n54526) );
  inv_x1_sg U47555 ( .A(n19328), .X(n54542) );
  nand_x1_sg U47556 ( .A(n54512), .B(n19240), .X(n19286) );
  inv_x1_sg U47557 ( .A(n18916), .X(n54520) );
  nand_x1_sg U47558 ( .A(n54541), .B(n40559), .X(n19386) );
  inv_x1_sg U47559 ( .A(n19492), .X(n54577) );
  inv_x1_sg U47560 ( .A(n19474), .X(n54556) );
  inv_x2_sg U47561 ( .A(n19449), .X(n43960) );
  nor_x1_sg U47562 ( .A(n54594), .B(n19451), .X(n19449) );
  inv_x1_sg U47563 ( .A(n19382), .X(n54582) );
  inv_x2_sg U47564 ( .A(n19379), .X(n45434) );
  nor_x1_sg U47565 ( .A(n19439), .B(n45437), .X(n19379) );
  nand_x1_sg U47566 ( .A(n29013), .B(n54607), .X(n29012) );
  inv_x2_sg U47567 ( .A(n28952), .X(n44262) );
  nor_x1_sg U47568 ( .A(n28953), .B(n28954), .X(n28952) );
  nand_x1_sg U47569 ( .A(n54663), .B(n46297), .X(n19804) );
  nand_x1_sg U47570 ( .A(n19788), .B(n54647), .X(n19787) );
  inv_x2_sg U47571 ( .A(n19847), .X(n44712) );
  inv_x1_sg U47572 ( .A(n19903), .X(n54702) );
  nand_x1_sg U47573 ( .A(n19865), .B(n19899), .X(n19898) );
  nand_x1_sg U47574 ( .A(n19815), .B(n46296), .X(n19814) );
  nand_x1_sg U47575 ( .A(n19818), .B(n54660), .X(n19813) );
  inv_x2_sg U47576 ( .A(n19890), .X(n44424) );
  nor_x1_sg U47577 ( .A(n19929), .B(n19930), .X(n19890) );
  inv_x1_sg U47578 ( .A(n19910), .X(n54721) );
  inv_x1_sg U47579 ( .A(n20071), .X(n54796) );
  nand_x1_sg U47580 ( .A(n54746), .B(n20064), .X(n20056) );
  inv_x1_sg U47581 ( .A(n19990), .X(n54754) );
  inv_x1_sg U47582 ( .A(n20064), .X(n54769) );
  inv_x1_sg U47583 ( .A(n19970), .X(n54756) );
  nand_x1_sg U47584 ( .A(n42428), .B(n20036), .X(n20033) );
  nand_x2_sg U47585 ( .A(n20100), .B(n20121), .X(n20049) );
  inv_x1_sg U47586 ( .A(n20049), .X(n54811) );
  inv_x1_sg U47587 ( .A(n20143), .X(n54851) );
  nand_x1_sg U47588 ( .A(n20144), .B(n20145), .X(n20142) );
  inv_x1_sg U47589 ( .A(n20209), .X(n45432) );
  inv_x1_sg U47590 ( .A(n20096), .X(n54828) );
  nand_x1_sg U47591 ( .A(n20083), .B(n20084), .X(n20081) );
  inv_x1_sg U47592 ( .A(n20083), .X(n54765) );
  nand_x1_sg U47593 ( .A(n54797), .B(n20009), .X(n20055) );
  inv_x2_sg U47594 ( .A(n20194), .X(n45416) );
  nor_x1_sg U47595 ( .A(n54803), .B(n20200), .X(n20194) );
  nand_x4_sg U47596 ( .A(n20153), .B(n20154), .X(n20096) );
  nand_x1_sg U47597 ( .A(n54827), .B(n20083), .X(n20154) );
  inv_x1_sg U47598 ( .A(n20262), .X(n54862) );
  inv_x1_sg U47599 ( .A(n20244), .X(n54841) );
  inv_x2_sg U47600 ( .A(n20218), .X(n43958) );
  nor_x1_sg U47601 ( .A(n54878), .B(n20220), .X(n20218) );
  nand_x1_sg U47602 ( .A(n29296), .B(n54891), .X(n29295) );
  inv_x2_sg U47603 ( .A(n29235), .X(n44250) );
  nor_x1_sg U47604 ( .A(n29236), .B(n29237), .X(n29235) );
  nand_x1_sg U47605 ( .A(n20565), .B(n54935), .X(n20564) );
  inv_x2_sg U47606 ( .A(n20645), .X(n44752) );
  inv_x1_sg U47607 ( .A(n20677), .X(n54991) );
  nand_x1_sg U47608 ( .A(n20639), .B(n20673), .X(n20672) );
  nand_x1_sg U47609 ( .A(n54929), .B(n54942), .X(n20673) );
  inv_x1_sg U47610 ( .A(n20684), .X(n54997) );
  nand_x1_sg U47611 ( .A(n20744), .B(n55042), .X(n20743) );
  inv_x1_sg U47612 ( .A(n20745), .X(n55042) );
  inv_x1_sg U47613 ( .A(n20847), .X(n55079) );
  nand_x1_sg U47614 ( .A(n55032), .B(n20840), .X(n20831) );
  nand_x4_sg U47615 ( .A(n20767), .B(n55052), .X(n20733) );
  inv_x1_sg U47616 ( .A(n20768), .X(n55052) );
  nand_x1_sg U47617 ( .A(n42430), .B(n20811), .X(n20808) );
  nand_x2_sg U47618 ( .A(n20876), .B(n20897), .X(n20824) );
  inv_x1_sg U47619 ( .A(n20824), .X(n55094) );
  inv_x1_sg U47620 ( .A(n20872), .X(n55110) );
  nand_x1_sg U47621 ( .A(n55080), .B(n20784), .X(n20830) );
  inv_x1_sg U47622 ( .A(n20460), .X(n55088) );
  nand_x1_sg U47623 ( .A(n55109), .B(n40560), .X(n20930) );
  inv_x1_sg U47624 ( .A(n21036), .X(n55145) );
  inv_x1_sg U47625 ( .A(n21018), .X(n55124) );
  inv_x2_sg U47626 ( .A(n20993), .X(n43956) );
  nor_x1_sg U47627 ( .A(n55162), .B(n20995), .X(n20993) );
  inv_x1_sg U47628 ( .A(n20926), .X(n55150) );
  inv_x2_sg U47629 ( .A(n20923), .X(n45426) );
  nor_x1_sg U47630 ( .A(n20983), .B(n45429), .X(n20923) );
  nand_x1_sg U47631 ( .A(n29574), .B(n55175), .X(n29573) );
  inv_x2_sg U47632 ( .A(n29513), .X(n44266) );
  nor_x1_sg U47633 ( .A(n29514), .B(n29515), .X(n29513) );
  nand_x1_sg U47634 ( .A(n55231), .B(n21269), .X(n21349) );
  nand_x1_sg U47635 ( .A(n21333), .B(n55215), .X(n21332) );
  inv_x2_sg U47636 ( .A(n21392), .X(n44710) );
  inv_x1_sg U47637 ( .A(n21448), .X(n55270) );
  nand_x1_sg U47638 ( .A(n21410), .B(n21444), .X(n21443) );
  nand_x1_sg U47639 ( .A(n21360), .B(n46251), .X(n21359) );
  nand_x1_sg U47640 ( .A(n21363), .B(n55228), .X(n21358) );
  inv_x2_sg U47641 ( .A(n21435), .X(n44422) );
  nor_x1_sg U47642 ( .A(n21474), .B(n21475), .X(n21435) );
  inv_x1_sg U47643 ( .A(n21455), .X(n55289) );
  inv_x1_sg U47644 ( .A(n21616), .X(n55364) );
  nand_x1_sg U47645 ( .A(n55314), .B(n21609), .X(n21601) );
  inv_x1_sg U47646 ( .A(n21535), .X(n55322) );
  inv_x1_sg U47647 ( .A(n21609), .X(n55337) );
  inv_x1_sg U47648 ( .A(n21515), .X(n55324) );
  nand_x1_sg U47649 ( .A(n42426), .B(n21581), .X(n21578) );
  nand_x2_sg U47650 ( .A(n21645), .B(n21666), .X(n21594) );
  inv_x1_sg U47651 ( .A(n21594), .X(n55379) );
  inv_x1_sg U47652 ( .A(n21688), .X(n55419) );
  nand_x1_sg U47653 ( .A(n21689), .B(n21690), .X(n21687) );
  inv_x1_sg U47654 ( .A(n21754), .X(n45424) );
  inv_x1_sg U47655 ( .A(n21641), .X(n55396) );
  nand_x1_sg U47656 ( .A(n21628), .B(n21629), .X(n21626) );
  inv_x1_sg U47657 ( .A(n21628), .X(n55333) );
  nand_x1_sg U47658 ( .A(n55365), .B(n21554), .X(n21600) );
  inv_x2_sg U47659 ( .A(n21739), .X(n45414) );
  nor_x1_sg U47660 ( .A(n55371), .B(n21745), .X(n21739) );
  nand_x4_sg U47661 ( .A(n21698), .B(n21699), .X(n21641) );
  nand_x1_sg U47662 ( .A(n55395), .B(n21628), .X(n21699) );
  inv_x1_sg U47663 ( .A(n21807), .X(n55430) );
  inv_x1_sg U47664 ( .A(n21789), .X(n55409) );
  inv_x2_sg U47665 ( .A(n21763), .X(n43954) );
  nor_x1_sg U47666 ( .A(n55446), .B(n21765), .X(n21763) );
  nand_x1_sg U47667 ( .A(n8184), .B(n50088), .X(n29665) );
  inv_x1_sg U47668 ( .A(n29666), .X(n50088) );
  nand_x1_sg U47669 ( .A(n8244), .B(n50090), .X(n30283) );
  nand_x1_sg U47670 ( .A(n24505), .B(n29849), .X(n30282) );
  inv_x1_sg U47671 ( .A(n30284), .X(n50090) );
  nand_x1_sg U47672 ( .A(n8324), .B(n50068), .X(n30255) );
  nand_x1_sg U47673 ( .A(n24488), .B(n30257), .X(n30254) );
  inv_x1_sg U47674 ( .A(n30256), .X(n50068) );
  nand_x1_sg U47675 ( .A(n8224), .B(n50081), .X(n29651) );
  inv_x1_sg U47676 ( .A(n29652), .X(n50081) );
  inv_x1_sg U47677 ( .A(n29656), .X(n50086) );
  nand_x1_sg U47678 ( .A(n8203), .B(n29655), .X(n29654) );
  nand_x1_sg U47679 ( .A(n8264), .B(n50077), .X(n30276) );
  inv_x1_sg U47680 ( .A(n30277), .X(n50077) );
  nand_x1_sg U47681 ( .A(n8304), .B(n50071), .X(n30262) );
  inv_x1_sg U47682 ( .A(n30263), .X(n50071) );
  inv_x1_sg U47683 ( .A(n30267), .X(n50076) );
  nand_x1_sg U47684 ( .A(n8283), .B(n30266), .X(n30265) );
  nand_x1_sg U47685 ( .A(n8424), .B(n50054), .X(n30218) );
  inv_x1_sg U47686 ( .A(n30219), .X(n50054) );
  nand_x1_sg U47687 ( .A(n8363), .B(n30238), .X(n30237) );
  nand_x1_sg U47688 ( .A(n8344), .B(n30248), .X(n30247) );
  nand_x1_sg U47689 ( .A(n8404), .B(n50058), .X(n30225) );
  nand_x1_sg U47690 ( .A(n30227), .B(n30228), .X(n30224) );
  inv_x1_sg U47691 ( .A(n30226), .X(n50058) );
  inv_x1_sg U47692 ( .A(n30209), .X(n50053) );
  nand_x1_sg U47693 ( .A(n8443), .B(n30208), .X(n30207) );
  nand_x1_sg U47694 ( .A(n8384), .B(n50060), .X(n30233) );
  inv_x1_sg U47695 ( .A(n30234), .X(n50060) );
  inv_x1_sg U47696 ( .A(n29669), .X(n50041) );
  inv_x1_sg U47697 ( .A(n30287), .X(n50046) );
  inv_x1_sg U47698 ( .A(n30520), .X(n50026) );
  inv_x1_sg U47699 ( .A(n29854), .X(n50036) );
  inv_x2_sg U47700 ( .A(n29840), .X(n44528) );
  nor_x1_sg U47701 ( .A(n29856), .B(n50044), .X(n29840) );
  inv_x1_sg U47702 ( .A(n30538), .X(n50048) );
  inv_x1_sg U47703 ( .A(n30526), .X(n50029) );
  inv_x2_sg U47704 ( .A(n30445), .X(n44630) );
  nor_x1_sg U47705 ( .A(n30528), .B(n50032), .X(n30445) );
  nor_x1_sg U47706 ( .A(n30474), .B(out_L1[17]), .X(n30473) );
  nor_x1_sg U47707 ( .A(n24562), .B(n50004), .X(n30513) );
  nand_x1_sg U47708 ( .A(n8364), .B(n30242), .X(n30506) );
  nand_x1_sg U47709 ( .A(n8444), .B(n30213), .X(n30480) );
  inv_x1_sg U47710 ( .A(n30487), .X(n50011) );
  nand_x1_sg U47711 ( .A(n8424), .B(n30220), .X(n30486) );
  nand_x1_sg U47712 ( .A(n8404), .B(n30228), .X(n30493) );
  inv_x1_sg U47713 ( .A(n30503), .X(n50017) );
  inv_x1_sg U47714 ( .A(n29672), .X(n49992) );
  inv_x1_sg U47715 ( .A(n30290), .X(n49998) );
  inv_x1_sg U47716 ( .A(n30541), .X(n50000) );
  inv_x1_sg U47717 ( .A(n30783), .X(n49984) );
  nand_x1_sg U47718 ( .A(n8285), .B(n30533), .X(n30786) );
  inv_x1_sg U47719 ( .A(n30777), .X(n49981) );
  inv_x1_sg U47720 ( .A(n30017), .X(n49997) );
  nand_x1_sg U47721 ( .A(n8225), .B(n29855), .X(n30016) );
  nand_x1_sg U47722 ( .A(n8365), .B(n30510), .X(n30761) );
  inv_x1_sg U47723 ( .A(n30742), .X(n49967) );
  nand_x1_sg U47724 ( .A(n8425), .B(n30491), .X(n30741) );
  nand_x1_sg U47725 ( .A(n8405), .B(n30497), .X(n30748) );
  inv_x1_sg U47726 ( .A(n30733), .X(n50005) );
  inv_x1_sg U47727 ( .A(n30758), .X(n49973) );
  inv_x1_sg U47728 ( .A(n29675), .X(n49947) );
  inv_x1_sg U47729 ( .A(n30293), .X(n49954) );
  nand_x1_sg U47730 ( .A(n8366), .B(n30765), .X(n30987) );
  inv_x1_sg U47731 ( .A(n30544), .X(n49956) );
  inv_x1_sg U47732 ( .A(n31007), .X(n49960) );
  nand_x1_sg U47733 ( .A(n8286), .B(n30697), .X(n30696) );
  inv_x1_sg U47734 ( .A(n31001), .X(n49938) );
  inv_x1_sg U47735 ( .A(n30006), .X(n49953) );
  nand_x1_sg U47736 ( .A(n8226), .B(n30005), .X(n30004) );
  inv_x2_sg U47737 ( .A(n29826), .X(n44572) );
  nor_x1_sg U47738 ( .A(n29828), .B(n49950), .X(n29826) );
  nor_x1_sg U47739 ( .A(n24660), .B(n49916), .X(n30994) );
  inv_x1_sg U47740 ( .A(n30968), .X(n49923) );
  nand_x1_sg U47741 ( .A(n8426), .B(n30746), .X(n30967) );
  nand_x1_sg U47742 ( .A(n8406), .B(n30752), .X(n30974) );
  nand_x2_sg U47743 ( .A(n30958), .B(n30959), .X(n30953) );
  inv_x2_sg U47744 ( .A(n30954), .X(n44302) );
  inv_x1_sg U47745 ( .A(n30984), .X(n49929) );
  inv_x1_sg U47746 ( .A(n29678), .X(n49899) );
  inv_x1_sg U47747 ( .A(n30296), .X(n49906) );
  inv_x1_sg U47748 ( .A(n30547), .X(n49908) );
  inv_x1_sg U47749 ( .A(n31010), .X(n49912) );
  nand_x1_sg U47750 ( .A(n8287), .B(n30691), .X(n30690) );
  inv_x1_sg U47751 ( .A(n31208), .X(n49914) );
  inv_x1_sg U47752 ( .A(n30000), .X(n49905) );
  nand_x1_sg U47753 ( .A(n8227), .B(n29999), .X(n29998) );
  inv_x2_sg U47754 ( .A(n29819), .X(n44570) );
  nor_x1_sg U47755 ( .A(n29821), .B(n49902), .X(n29819) );
  nand_x1_sg U47756 ( .A(n8367), .B(n30991), .X(n31192) );
  inv_x1_sg U47757 ( .A(n31173), .X(n49877) );
  nand_x1_sg U47758 ( .A(n8427), .B(n30972), .X(n31172) );
  nand_x1_sg U47759 ( .A(n8407), .B(n30978), .X(n31179) );
  nand_x1_sg U47760 ( .A(n31170), .B(n31171), .X(n31167) );
  nand_x1_sg U47761 ( .A(n8448), .B(n31169), .X(n31168) );
  inv_x1_sg U47762 ( .A(n31164), .X(n49918) );
  inv_x1_sg U47763 ( .A(n31189), .X(n49883) );
  inv_x1_sg U47764 ( .A(n29681), .X(n49852) );
  inv_x1_sg U47765 ( .A(n30299), .X(n49859) );
  nand_x1_sg U47766 ( .A(n8368), .B(n31196), .X(n31382) );
  inv_x1_sg U47767 ( .A(n31211), .X(n49868) );
  inv_x1_sg U47768 ( .A(n29994), .X(n49858) );
  nand_x1_sg U47769 ( .A(n8228), .B(n29993), .X(n29992) );
  inv_x2_sg U47770 ( .A(n29812), .X(n44566) );
  nor_x1_sg U47771 ( .A(n29814), .B(n49855), .X(n29812) );
  inv_x1_sg U47772 ( .A(n30550), .X(n49861) );
  inv_x1_sg U47773 ( .A(n30920), .X(n49867) );
  nand_x1_sg U47774 ( .A(n8308), .B(n30919), .X(n30918) );
  inv_x2_sg U47775 ( .A(n30681), .X(n44568) );
  nor_x1_sg U47776 ( .A(n30683), .B(n49864), .X(n30681) );
  nor_x1_sg U47777 ( .A(n24756), .B(n49822), .X(n31389) );
  inv_x1_sg U47778 ( .A(n31363), .X(n49831) );
  nand_x1_sg U47779 ( .A(n8428), .B(n31177), .X(n31362) );
  nand_x1_sg U47780 ( .A(n8408), .B(n31183), .X(n31369) );
  nand_x2_sg U47781 ( .A(n31353), .B(n31354), .X(n31348) );
  inv_x2_sg U47782 ( .A(n31349), .X(n45582) );
  inv_x1_sg U47783 ( .A(n31379), .X(n49837) );
  inv_x1_sg U47784 ( .A(n29684), .X(n49804) );
  inv_x1_sg U47785 ( .A(n30302), .X(n49811) );
  inv_x1_sg U47786 ( .A(n31214), .X(n49820) );
  inv_x1_sg U47787 ( .A(n29988), .X(n49810) );
  nand_x1_sg U47788 ( .A(n8229), .B(n29987), .X(n29986) );
  inv_x2_sg U47789 ( .A(n29805), .X(n44562) );
  nor_x1_sg U47790 ( .A(n29807), .B(n49807), .X(n29805) );
  inv_x1_sg U47791 ( .A(n30553), .X(n49813) );
  inv_x1_sg U47792 ( .A(n30914), .X(n49819) );
  nand_x1_sg U47793 ( .A(n8309), .B(n30913), .X(n30912) );
  inv_x2_sg U47794 ( .A(n30674), .X(n44564) );
  nor_x1_sg U47795 ( .A(n30676), .B(n49816), .X(n30674) );
  nand_x1_sg U47796 ( .A(n8369), .B(n31386), .X(n31553) );
  inv_x1_sg U47797 ( .A(n31534), .X(n49786) );
  nand_x1_sg U47798 ( .A(n8429), .B(n31367), .X(n31533) );
  nand_x1_sg U47799 ( .A(n8409), .B(n31373), .X(n31540) );
  nand_x1_sg U47800 ( .A(n31531), .B(n31532), .X(n31528) );
  nand_x1_sg U47801 ( .A(n8450), .B(n31530), .X(n31529) );
  inv_x1_sg U47802 ( .A(n31525), .X(n49826) );
  inv_x1_sg U47803 ( .A(n31550), .X(n49792) );
  inv_x1_sg U47804 ( .A(n31217), .X(n49773) );
  inv_x1_sg U47805 ( .A(n29982), .X(n49763) );
  nand_x1_sg U47806 ( .A(n8230), .B(n29981), .X(n29980) );
  inv_x1_sg U47807 ( .A(n30556), .X(n49766) );
  inv_x1_sg U47808 ( .A(n30908), .X(n49772) );
  nand_x1_sg U47809 ( .A(n8310), .B(n30907), .X(n30906) );
  inv_x2_sg U47810 ( .A(n30667), .X(n44638) );
  nor_x1_sg U47811 ( .A(n30669), .B(n49769), .X(n30667) );
  inv_x2_sg U47812 ( .A(n29798), .X(n44560) );
  nor_x1_sg U47813 ( .A(n29800), .B(n49760), .X(n29798) );
  inv_x1_sg U47814 ( .A(n29687), .X(n49757) );
  nand_x1_sg U47815 ( .A(n8250), .B(n30138), .X(n30137) );
  nand_x1_sg U47816 ( .A(n8370), .B(n31501), .X(n31500) );
  inv_x1_sg U47817 ( .A(n31687), .X(n49740) );
  nand_x1_sg U47818 ( .A(n8430), .B(n31538), .X(n31686) );
  nand_x1_sg U47819 ( .A(n8410), .B(n31544), .X(n31693) );
  nand_x2_sg U47820 ( .A(n31677), .B(n31678), .X(n31672) );
  inv_x2_sg U47821 ( .A(n31673), .X(n44722) );
  inv_x1_sg U47822 ( .A(n31703), .X(n49779) );
  inv_x1_sg U47823 ( .A(n29690), .X(n49708) );
  inv_x1_sg U47824 ( .A(n30308), .X(n49715) );
  inv_x1_sg U47825 ( .A(n31220), .X(n49724) );
  inv_x1_sg U47826 ( .A(n29976), .X(n49714) );
  nand_x1_sg U47827 ( .A(n8231), .B(n29975), .X(n29974) );
  inv_x2_sg U47828 ( .A(n29791), .X(n44556) );
  nor_x1_sg U47829 ( .A(n29793), .B(n49711), .X(n29791) );
  inv_x1_sg U47830 ( .A(n30559), .X(n49717) );
  inv_x1_sg U47831 ( .A(n30902), .X(n49723) );
  nand_x1_sg U47832 ( .A(n8311), .B(n30901), .X(n30900) );
  inv_x2_sg U47833 ( .A(n30660), .X(n44558) );
  nor_x1_sg U47834 ( .A(n30662), .B(n49720), .X(n30660) );
  nand_x1_sg U47835 ( .A(n8371), .B(n31495), .X(n31494) );
  inv_x1_sg U47836 ( .A(n31831), .X(n49694) );
  nand_x1_sg U47837 ( .A(n8431), .B(n31691), .X(n31830) );
  nand_x1_sg U47838 ( .A(n8411), .B(n31697), .X(n31837) );
  nand_x1_sg U47839 ( .A(n31828), .B(n31829), .X(n31825) );
  nand_x1_sg U47840 ( .A(n8452), .B(n31827), .X(n31826) );
  inv_x1_sg U47841 ( .A(n31822), .X(n49735) );
  inv_x1_sg U47842 ( .A(n31706), .X(n49729) );
  inv_x1_sg U47843 ( .A(n29693), .X(n49661) );
  inv_x1_sg U47844 ( .A(n30311), .X(n49668) );
  inv_x1_sg U47845 ( .A(n31223), .X(n49677) );
  inv_x1_sg U47846 ( .A(n29970), .X(n49667) );
  nand_x1_sg U47847 ( .A(n8232), .B(n29969), .X(n29968) );
  inv_x2_sg U47848 ( .A(n29784), .X(n44552) );
  nor_x1_sg U47849 ( .A(n29786), .B(n49664), .X(n29784) );
  inv_x1_sg U47850 ( .A(n30562), .X(n49670) );
  inv_x1_sg U47851 ( .A(n30896), .X(n49676) );
  nand_x1_sg U47852 ( .A(n8312), .B(n30895), .X(n30894) );
  inv_x2_sg U47853 ( .A(n30653), .X(n44554) );
  nor_x1_sg U47854 ( .A(n30655), .B(n49673), .X(n30653) );
  nand_x1_sg U47855 ( .A(n8372), .B(n31489), .X(n31488) );
  inv_x1_sg U47856 ( .A(n31947), .X(n49688) );
  nand_x1_sg U47857 ( .A(n8432), .B(n31835), .X(n31946) );
  nand_x1_sg U47858 ( .A(n8412), .B(n31804), .X(n31803) );
  nand_x2_sg U47859 ( .A(n31937), .B(n31938), .X(n31932) );
  inv_x2_sg U47860 ( .A(n31933), .X(n45586) );
  inv_x1_sg U47861 ( .A(n31709), .X(n49683) );
  inv_x1_sg U47862 ( .A(n29696), .X(n49614) );
  inv_x1_sg U47863 ( .A(n30314), .X(n49621) );
  inv_x1_sg U47864 ( .A(n31226), .X(n49630) );
  inv_x1_sg U47865 ( .A(n29964), .X(n49620) );
  nand_x1_sg U47866 ( .A(n8233), .B(n29963), .X(n29962) );
  inv_x2_sg U47867 ( .A(n29777), .X(n44548) );
  nor_x1_sg U47868 ( .A(n29779), .B(n49617), .X(n29777) );
  inv_x1_sg U47869 ( .A(n30565), .X(n49623) );
  inv_x1_sg U47870 ( .A(n30890), .X(n49629) );
  nand_x1_sg U47871 ( .A(n8313), .B(n30889), .X(n30888) );
  inv_x2_sg U47872 ( .A(n30646), .X(n44550) );
  nor_x1_sg U47873 ( .A(n30648), .B(n49626), .X(n30646) );
  nand_x1_sg U47874 ( .A(n8373), .B(n31483), .X(n31482) );
  inv_x1_sg U47875 ( .A(n31923), .X(n49641) );
  nand_x1_sg U47876 ( .A(n8433), .B(n31922), .X(n31921) );
  nand_x1_sg U47877 ( .A(n8413), .B(n31797), .X(n31796) );
  nand_x1_sg U47878 ( .A(n8454), .B(n32045), .X(n32044) );
  nand_x1_sg U47879 ( .A(n32024), .B(n32028), .X(n32043) );
  inv_x1_sg U47880 ( .A(n32040), .X(n49644) );
  inv_x1_sg U47881 ( .A(n31712), .X(n49635) );
  inv_x1_sg U47882 ( .A(n29699), .X(n49568) );
  inv_x1_sg U47883 ( .A(n30317), .X(n49575) );
  inv_x1_sg U47884 ( .A(n31229), .X(n49584) );
  inv_x1_sg U47885 ( .A(n29958), .X(n49574) );
  nand_x1_sg U47886 ( .A(n8234), .B(n29957), .X(n29956) );
  inv_x2_sg U47887 ( .A(n29770), .X(n44544) );
  nor_x1_sg U47888 ( .A(n29772), .B(n49571), .X(n29770) );
  inv_x1_sg U47889 ( .A(n30568), .X(n49577) );
  inv_x1_sg U47890 ( .A(n30884), .X(n49583) );
  nand_x1_sg U47891 ( .A(n8314), .B(n30883), .X(n30882) );
  inv_x2_sg U47892 ( .A(n30639), .X(n44546) );
  nor_x1_sg U47893 ( .A(n30641), .B(n49580), .X(n30639) );
  nand_x1_sg U47894 ( .A(n8374), .B(n31477), .X(n31476) );
  inv_x1_sg U47895 ( .A(n31917), .X(n49595) );
  nand_x1_sg U47896 ( .A(n8434), .B(n31916), .X(n31915) );
  nand_x1_sg U47897 ( .A(n8414), .B(n31790), .X(n31789) );
  nand_x1_sg U47898 ( .A(n8455), .B(n32048), .X(n32047) );
  nand_x1_sg U47899 ( .A(n8474), .B(n40801), .X(n32134) );
  nand_x1_sg U47900 ( .A(out_L1[8]), .B(n40802), .X(n32135) );
  inv_x1_sg U47901 ( .A(n31715), .X(n49589) );
  inv_x1_sg U47902 ( .A(n29702), .X(n49521) );
  inv_x1_sg U47903 ( .A(n30320), .X(n49528) );
  inv_x1_sg U47904 ( .A(n31232), .X(n49537) );
  inv_x1_sg U47905 ( .A(n29952), .X(n49527) );
  nand_x1_sg U47906 ( .A(n8235), .B(n29951), .X(n29950) );
  inv_x2_sg U47907 ( .A(n29763), .X(n44540) );
  nor_x1_sg U47908 ( .A(n29765), .B(n49524), .X(n29763) );
  inv_x1_sg U47909 ( .A(n30571), .X(n49530) );
  inv_x1_sg U47910 ( .A(n30878), .X(n49536) );
  nand_x1_sg U47911 ( .A(n8315), .B(n30877), .X(n30876) );
  inv_x2_sg U47912 ( .A(n30632), .X(n44542) );
  nor_x1_sg U47913 ( .A(n30634), .B(n49533), .X(n30632) );
  nand_x1_sg U47914 ( .A(n8375), .B(n31471), .X(n31470) );
  inv_x1_sg U47915 ( .A(n31911), .X(n49549) );
  nand_x1_sg U47916 ( .A(n8435), .B(n31910), .X(n31909) );
  nand_x1_sg U47917 ( .A(n8415), .B(n31783), .X(n31782) );
  inv_x2_sg U47918 ( .A(n32117), .X(n44294) );
  nand_x1_sg U47919 ( .A(n8455), .B(n32021), .X(n32020) );
  inv_x1_sg U47920 ( .A(n31718), .X(n49543) );
  inv_x1_sg U47921 ( .A(n30872), .X(n49489) );
  nand_x1_sg U47922 ( .A(n8316), .B(n30871), .X(n30870) );
  nand_x1_sg U47923 ( .A(n8296), .B(n30629), .X(n30628) );
  inv_x1_sg U47924 ( .A(n30574), .X(n49483) );
  inv_x1_sg U47925 ( .A(n29705), .X(n49474) );
  nand_x1_sg U47926 ( .A(n8256), .B(n30102), .X(n30101) );
  inv_x1_sg U47927 ( .A(n31235), .X(n49490) );
  inv_x1_sg U47928 ( .A(n29946), .X(n49480) );
  nand_x1_sg U47929 ( .A(n8236), .B(n29945), .X(n29944) );
  inv_x2_sg U47930 ( .A(n29756), .X(n44538) );
  nor_x1_sg U47931 ( .A(n29758), .B(n49477), .X(n29756) );
  nand_x1_sg U47932 ( .A(n8376), .B(n31465), .X(n31464) );
  inv_x1_sg U47933 ( .A(n31905), .X(n49501) );
  nand_x1_sg U47934 ( .A(n8436), .B(n31904), .X(n31903) );
  nand_x1_sg U47935 ( .A(n8416), .B(n31776), .X(n31775) );
  inv_x1_sg U47936 ( .A(n31721), .X(n49495) );
  inv_x1_sg U47937 ( .A(n29708), .X(n49428) );
  inv_x1_sg U47938 ( .A(n30326), .X(n49435) );
  inv_x1_sg U47939 ( .A(n31238), .X(n49444) );
  inv_x1_sg U47940 ( .A(n29940), .X(n49434) );
  nand_x1_sg U47941 ( .A(n8237), .B(n29939), .X(n29938) );
  inv_x2_sg U47942 ( .A(n29749), .X(n44534) );
  nor_x1_sg U47943 ( .A(n29751), .B(n49431), .X(n29749) );
  inv_x1_sg U47944 ( .A(n30577), .X(n49437) );
  inv_x1_sg U47945 ( .A(n30866), .X(n49443) );
  nand_x1_sg U47946 ( .A(n8317), .B(n30865), .X(n30864) );
  inv_x2_sg U47947 ( .A(n30618), .X(n44536) );
  nor_x1_sg U47948 ( .A(n30620), .B(n49440), .X(n30618) );
  nand_x1_sg U47949 ( .A(n8377), .B(n31459), .X(n31458) );
  inv_x1_sg U47950 ( .A(n31899), .X(n49455) );
  nand_x1_sg U47951 ( .A(n8437), .B(n31898), .X(n31897) );
  nand_x1_sg U47952 ( .A(n8417), .B(n31769), .X(n31768) );
  nand_x1_sg U47953 ( .A(n8457), .B(n32008), .X(n32007) );
  inv_x1_sg U47954 ( .A(n31724), .X(n49449) );
  inv_x1_sg U47955 ( .A(n30860), .X(n49397) );
  nand_x1_sg U47956 ( .A(n8318), .B(n30859), .X(n30858) );
  nand_x1_sg U47957 ( .A(n8298), .B(n30615), .X(n30614) );
  inv_x1_sg U47958 ( .A(n30580), .X(n49391) );
  inv_x1_sg U47959 ( .A(n29711), .X(n49382) );
  nand_x1_sg U47960 ( .A(n8258), .B(n30090), .X(n30089) );
  inv_x1_sg U47961 ( .A(n31241), .X(n49398) );
  inv_x1_sg U47962 ( .A(n29934), .X(n49388) );
  nand_x1_sg U47963 ( .A(n8238), .B(n29933), .X(n29932) );
  inv_x2_sg U47964 ( .A(n29742), .X(n44532) );
  nor_x1_sg U47965 ( .A(n29744), .B(n49385), .X(n29742) );
  nand_x1_sg U47966 ( .A(n8378), .B(n31453), .X(n31452) );
  inv_x1_sg U47967 ( .A(n31893), .X(n49410) );
  nand_x1_sg U47968 ( .A(n8438), .B(n31892), .X(n31891) );
  nand_x1_sg U47969 ( .A(n8418), .B(n31762), .X(n31761) );
  inv_x1_sg U47970 ( .A(n31727), .X(n49404) );
  inv_x1_sg U47971 ( .A(n30854), .X(n49353) );
  nand_x1_sg U47972 ( .A(n8319), .B(n30853), .X(n30852) );
  nand_x1_sg U47973 ( .A(n8299), .B(n30608), .X(n30607) );
  inv_x1_sg U47974 ( .A(n30583), .X(n49347) );
  inv_x1_sg U47975 ( .A(n29714), .X(n49338) );
  nand_x1_sg U47976 ( .A(n8259), .B(n30084), .X(n30083) );
  inv_x1_sg U47977 ( .A(n31244), .X(n49354) );
  inv_x1_sg U47978 ( .A(n29928), .X(n49344) );
  nand_x1_sg U47979 ( .A(n8239), .B(n29927), .X(n29926) );
  inv_x2_sg U47980 ( .A(n29735), .X(n44530) );
  nor_x1_sg U47981 ( .A(n29737), .B(n49341), .X(n29735) );
  nand_x1_sg U47982 ( .A(n8379), .B(n31447), .X(n31446) );
  nand_x1_sg U47983 ( .A(n8360), .B(n31425), .X(n31424) );
  inv_x1_sg U47984 ( .A(n31887), .X(n49365) );
  nand_x1_sg U47985 ( .A(n8439), .B(n31886), .X(n31885) );
  nand_x1_sg U47986 ( .A(n8419), .B(n31755), .X(n31754) );
  inv_x1_sg U47987 ( .A(n31730), .X(n49359) );
  inv_x1_sg U47988 ( .A(n30848), .X(n49306) );
  nand_x1_sg U47989 ( .A(n8320), .B(n30847), .X(n30846) );
  nand_x1_sg U47990 ( .A(n8300), .B(n30601), .X(n30600) );
  nand_x1_sg U47991 ( .A(n8260), .B(n30078), .X(n30077) );
  inv_x1_sg U47992 ( .A(n29922), .X(n49300) );
  nand_x1_sg U47993 ( .A(n8240), .B(n29921), .X(n29920) );
  inv_x2_sg U47994 ( .A(n29728), .X(n44065) );
  nor_x1_sg U47995 ( .A(n29730), .B(n49298), .X(n29728) );
  inv_x1_sg U47996 ( .A(n31881), .X(n49316) );
  nand_x1_sg U47997 ( .A(n8440), .B(n31880), .X(n31879) );
  nand_x1_sg U47998 ( .A(n8420), .B(n31748), .X(n31747) );
  nand_x2_sg U47999 ( .A(n49322), .B(n32078), .X(n32076) );
  inv_x1_sg U48000 ( .A(n32079), .X(n49322) );
  nand_x1_sg U48001 ( .A(n8460), .B(n31989), .X(n31988) );
  nand_x2_sg U48002 ( .A(n30840), .B(n30841), .X(n30839) );
  nand_x2_sg U48003 ( .A(n30592), .B(n30593), .X(n30591) );
  nand_x2_sg U48004 ( .A(n32072), .B(n32073), .X(n32071) );
  nand_x2_sg U48005 ( .A(n31873), .B(n31874), .X(n31872) );
  nand_x2_sg U48006 ( .A(n30070), .B(n30071), .X(n30069) );
  nand_x2_sg U48007 ( .A(n29723), .B(n29724), .X(n29722) );
  nand_x2_sg U48008 ( .A(n31054), .B(n31055), .X(n31053) );
  nand_x2_sg U48009 ( .A(n29914), .B(n29915), .X(n29913) );
  nand_x2_sg U48010 ( .A(n31980), .B(n31981), .X(n31979) );
  nand_x2_sg U48011 ( .A(n31739), .B(n31740), .X(n31738) );
  nand_x1_sg U48012 ( .A(n51266), .B(n51259), .X(n25592) );
  nand_x1_sg U48013 ( .A(n25593), .B(n25594), .X(n25591) );
  nand_x1_sg U48014 ( .A(n51272), .B(n25588), .X(n25585) );
  nand_x1_sg U48015 ( .A(n45275), .B(n25654), .X(n25653) );
  nand_x1_sg U48016 ( .A(n25588), .B(n50970), .X(n25652) );
  nand_x2_sg U48017 ( .A(n25565), .B(n25566), .X(n25563) );
  inv_x1_sg U48018 ( .A(n25564), .X(n51303) );
  inv_x1_sg U48019 ( .A(n25563), .X(n51318) );
  nand_x2_sg U48020 ( .A(n45125), .B(n51317), .X(n25565) );
  inv_x1_sg U48021 ( .A(n25645), .X(n51302) );
  nand_x1_sg U48022 ( .A(n51542), .B(n51535), .X(n25873) );
  nand_x1_sg U48023 ( .A(n25874), .B(n25875), .X(n25872) );
  nand_x1_sg U48024 ( .A(n25861), .B(n25862), .X(n25863) );
  nand_x1_sg U48025 ( .A(n51551), .B(n51540), .X(n25867) );
  nand_x1_sg U48026 ( .A(n25868), .B(n25869), .X(n25866) );
  inv_x1_sg U48027 ( .A(n25855), .X(n51575) );
  nand_x1_sg U48028 ( .A(n25856), .B(n25857), .X(n25854) );
  inv_x1_sg U48029 ( .A(n25848), .X(n46202) );
  nand_x1_sg U48030 ( .A(n25849), .B(n25850), .X(n25851) );
  nand_x2_sg U48031 ( .A(n25846), .B(n25847), .X(n25844) );
  inv_x1_sg U48032 ( .A(n25845), .X(n51585) );
  inv_x1_sg U48033 ( .A(n25844), .X(n51597) );
  nand_x2_sg U48034 ( .A(n45107), .B(n51669), .X(n25822) );
  nand_x1_sg U48035 ( .A(n51825), .B(n51817), .X(n26153) );
  nand_x1_sg U48036 ( .A(n26154), .B(n26155), .X(n26152) );
  nand_x1_sg U48037 ( .A(n45281), .B(n26213), .X(n26212) );
  nand_x1_sg U48038 ( .A(n26149), .B(n51008), .X(n26211) );
  nand_x1_sg U48039 ( .A(n51832), .B(n26149), .X(n26146) );
  nand_x2_sg U48040 ( .A(n26126), .B(n26127), .X(n26124) );
  inv_x1_sg U48041 ( .A(n26125), .X(n51864) );
  inv_x1_sg U48042 ( .A(n26124), .X(n51878) );
  nand_x2_sg U48043 ( .A(n45091), .B(n51950), .X(n26102) );
  nand_x1_sg U48044 ( .A(n52099), .B(n52093), .X(n26432) );
  nand_x1_sg U48045 ( .A(n26433), .B(n26434), .X(n26431) );
  nand_x1_sg U48046 ( .A(n26420), .B(n26421), .X(n26422) );
  nand_x1_sg U48047 ( .A(n52108), .B(n52097), .X(n26426) );
  nand_x1_sg U48048 ( .A(n26427), .B(n26428), .X(n26425) );
  inv_x1_sg U48049 ( .A(n26414), .X(n52132) );
  nand_x1_sg U48050 ( .A(n26415), .B(n26416), .X(n26413) );
  nand_x4_sg U48051 ( .A(n26410), .B(n46198), .X(n43745) );
  inv_x8_sg U48052 ( .A(n43745), .X(n12826) );
  nand_x2_sg U48053 ( .A(n26405), .B(n26406), .X(n26403) );
  inv_x1_sg U48054 ( .A(n26404), .X(n52143) );
  inv_x1_sg U48055 ( .A(n26403), .X(n52155) );
  nand_x2_sg U48056 ( .A(n45075), .B(n52269), .X(n26369) );
  nand_x1_sg U48057 ( .A(n52377), .B(n52370), .X(n26710) );
  nand_x1_sg U48058 ( .A(n26711), .B(n26712), .X(n26709) );
  nand_x1_sg U48059 ( .A(n45291), .B(n26770), .X(n26769) );
  nand_x1_sg U48060 ( .A(n26706), .B(n51047), .X(n26768) );
  nand_x1_sg U48061 ( .A(n52384), .B(n26706), .X(n26703) );
  inv_x1_sg U48062 ( .A(n26692), .X(n52405) );
  nand_x1_sg U48063 ( .A(n26693), .B(n26694), .X(n26691) );
  nand_x2_sg U48064 ( .A(n26683), .B(n26684), .X(n26681) );
  inv_x1_sg U48065 ( .A(n26682), .X(n52416) );
  inv_x1_sg U48066 ( .A(n26681), .X(n52429) );
  nand_x2_sg U48067 ( .A(n45067), .B(n52428), .X(n26683) );
  inv_x1_sg U48068 ( .A(n26761), .X(n52415) );
  nand_x2_sg U48069 ( .A(n45171), .B(n52445), .X(n26677) );
  nand_x2_sg U48070 ( .A(n45061), .B(n52544), .X(n26647) );
  nand_x1_sg U48071 ( .A(n52654), .B(n52646), .X(n26989) );
  nand_x1_sg U48072 ( .A(n26990), .B(n26991), .X(n26988) );
  nand_x1_sg U48073 ( .A(n45309), .B(n27049), .X(n27048) );
  nand_x1_sg U48074 ( .A(n26985), .B(n51066), .X(n27047) );
  nand_x1_sg U48075 ( .A(n52661), .B(n26985), .X(n26982) );
  inv_x1_sg U48076 ( .A(n26971), .X(n52682) );
  nand_x1_sg U48077 ( .A(n26972), .B(n26973), .X(n26970) );
  nand_x1_sg U48078 ( .A(n52933), .B(n52927), .X(n27269) );
  nand_x1_sg U48079 ( .A(n27270), .B(n27271), .X(n27268) );
  nand_x1_sg U48080 ( .A(n27257), .B(n27258), .X(n27259) );
  nand_x1_sg U48081 ( .A(n52942), .B(n52931), .X(n27263) );
  nand_x1_sg U48082 ( .A(n27264), .B(n27265), .X(n27262) );
  inv_x1_sg U48083 ( .A(n27251), .X(n52966) );
  nand_x1_sg U48084 ( .A(n27252), .B(n27253), .X(n27250) );
  nand_x4_sg U48085 ( .A(n27247), .B(n46197), .X(n43746) );
  inv_x8_sg U48086 ( .A(n43746), .X(n15159) );
  nand_x2_sg U48087 ( .A(n27242), .B(n27243), .X(n27240) );
  inv_x1_sg U48088 ( .A(n27241), .X(n52977) );
  inv_x1_sg U48089 ( .A(n27240), .X(n52989) );
  nand_x2_sg U48090 ( .A(n45033), .B(n53103), .X(n27206) );
  nand_x1_sg U48091 ( .A(n53213), .B(n53205), .X(n27548) );
  nand_x1_sg U48092 ( .A(n27549), .B(n27550), .X(n27547) );
  nand_x1_sg U48093 ( .A(n45285), .B(n27608), .X(n27607) );
  nand_x1_sg U48094 ( .A(n27544), .B(n51104), .X(n27606) );
  nand_x1_sg U48095 ( .A(n53220), .B(n27544), .X(n27541) );
  nand_x2_sg U48096 ( .A(n27521), .B(n27522), .X(n27519) );
  inv_x1_sg U48097 ( .A(n27520), .X(n53250) );
  inv_x1_sg U48098 ( .A(n27519), .X(n53265) );
  nand_x2_sg U48099 ( .A(n45025), .B(n53264), .X(n27521) );
  inv_x1_sg U48100 ( .A(n27599), .X(n53249) );
  nand_x2_sg U48101 ( .A(n45181), .B(n53280), .X(n27515) );
  nand_x2_sg U48102 ( .A(n45019), .B(n53338), .X(n27497) );
  nand_x1_sg U48103 ( .A(n53491), .B(n53485), .X(n27827) );
  nand_x1_sg U48104 ( .A(n27828), .B(n27829), .X(n27826) );
  nand_x1_sg U48105 ( .A(n27815), .B(n27816), .X(n27817) );
  nand_x1_sg U48106 ( .A(n53500), .B(n53489), .X(n27821) );
  nand_x1_sg U48107 ( .A(n27822), .B(n27823), .X(n27820) );
  inv_x1_sg U48108 ( .A(n27809), .X(n53524) );
  nand_x1_sg U48109 ( .A(n27810), .B(n27811), .X(n27808) );
  nand_x4_sg U48110 ( .A(n27805), .B(n46196), .X(n43747) );
  inv_x8_sg U48111 ( .A(n43747), .X(n16725) );
  nand_x2_sg U48112 ( .A(n27800), .B(n27801), .X(n27798) );
  inv_x1_sg U48113 ( .A(n27799), .X(n53535) );
  inv_x1_sg U48114 ( .A(n27798), .X(n53547) );
  nand_x2_sg U48115 ( .A(n45003), .B(n53661), .X(n27764) );
  nand_x1_sg U48116 ( .A(n53771), .B(n53763), .X(n28108) );
  nand_x1_sg U48117 ( .A(n28109), .B(n28110), .X(n28107) );
  nand_x1_sg U48118 ( .A(n28096), .B(n28097), .X(n28098) );
  nand_x1_sg U48119 ( .A(n53778), .B(n53769), .X(n28102) );
  nand_x1_sg U48120 ( .A(n28103), .B(n28104), .X(n28101) );
  inv_x1_sg U48121 ( .A(n46041), .X(n43778) );
  inv_x2_sg U48122 ( .A(n17503), .X(n43863) );
  nor_x1_sg U48123 ( .A(n53813), .B(n28083), .X(n17503) );
  inv_x1_sg U48124 ( .A(n28383), .X(n54057) );
  nand_x2_sg U48125 ( .A(n28378), .B(n28379), .X(n28376) );
  inv_x1_sg U48126 ( .A(n28376), .X(n54069) );
  nand_x1_sg U48127 ( .A(n54083), .B(n28371), .X(n28368) );
  inv_x2_sg U48128 ( .A(n18273), .X(n43810) );
  nor_x1_sg U48129 ( .A(n54096), .B(n28362), .X(n18273) );
  nand_x2_sg U48130 ( .A(n28360), .B(n28361), .X(n28358) );
  inv_x1_sg U48131 ( .A(n28359), .X(n54094) );
  inv_x1_sg U48132 ( .A(n28358), .X(n54108) );
  nand_x2_sg U48133 ( .A(n44981), .B(n54107), .X(n28360) );
  nand_x1_sg U48134 ( .A(n28364), .B(n51163), .X(n28436) );
  nand_x1_sg U48135 ( .A(n45211), .B(n28438), .X(n28437) );
  nand_x1_sg U48136 ( .A(n54336), .B(n54328), .X(n28666) );
  nand_x1_sg U48137 ( .A(n28667), .B(n28668), .X(n28665) );
  nand_x1_sg U48138 ( .A(n28654), .B(n28655), .X(n28656) );
  nand_x1_sg U48139 ( .A(n54343), .B(n54334), .X(n28660) );
  nand_x1_sg U48140 ( .A(n28661), .B(n28662), .X(n28659) );
  inv_x1_sg U48141 ( .A(n46039), .X(n43776) );
  inv_x2_sg U48142 ( .A(n19048), .X(n43861) );
  nor_x1_sg U48143 ( .A(n54378), .B(n28641), .X(n19048) );
  nand_x1_sg U48144 ( .A(n54620), .B(n54612), .X(n28944) );
  nand_x1_sg U48145 ( .A(n28945), .B(n28946), .X(n28943) );
  nand_x1_sg U48146 ( .A(n45289), .B(n29004), .X(n29003) );
  nand_x1_sg U48147 ( .A(n28940), .B(n51198), .X(n29002) );
  nand_x1_sg U48148 ( .A(n54626), .B(n28940), .X(n28937) );
  inv_x1_sg U48149 ( .A(n28926), .X(n54646) );
  nand_x1_sg U48150 ( .A(n28927), .B(n28928), .X(n28925) );
  nand_x2_sg U48151 ( .A(n28917), .B(n28918), .X(n28915) );
  inv_x1_sg U48152 ( .A(n28916), .X(n54657) );
  inv_x1_sg U48153 ( .A(n28915), .X(n54672) );
  nand_x1_sg U48154 ( .A(n54904), .B(n54896), .X(n29227) );
  nand_x1_sg U48155 ( .A(n29228), .B(n29229), .X(n29226) );
  nand_x1_sg U48156 ( .A(n29215), .B(n29216), .X(n29217) );
  nand_x1_sg U48157 ( .A(n54911), .B(n54902), .X(n29221) );
  nand_x1_sg U48158 ( .A(n29222), .B(n29223), .X(n29220) );
  inv_x1_sg U48159 ( .A(n46037), .X(n43774) );
  inv_x2_sg U48160 ( .A(n20592), .X(n43859) );
  nor_x1_sg U48161 ( .A(n54946), .B(n29202), .X(n20592) );
  nand_x1_sg U48162 ( .A(n55188), .B(n55180), .X(n29505) );
  nand_x1_sg U48163 ( .A(n29506), .B(n29507), .X(n29504) );
  nand_x1_sg U48164 ( .A(n45287), .B(n29565), .X(n29564) );
  nand_x1_sg U48165 ( .A(n29501), .B(n51236), .X(n29563) );
  nand_x1_sg U48166 ( .A(n55194), .B(n29501), .X(n29498) );
  nand_x2_sg U48167 ( .A(n29478), .B(n29479), .X(n29476) );
  inv_x1_sg U48168 ( .A(n29477), .X(n55225) );
  inv_x1_sg U48169 ( .A(n29476), .X(n55240) );
  nand_x2_sg U48170 ( .A(n44921), .B(n55239), .X(n29478) );
  inv_x1_sg U48171 ( .A(n29556), .X(n55224) );
  nand_x2_sg U48172 ( .A(n44919), .B(n55273), .X(n29466) );
  nand_x2_sg U48173 ( .A(n44917), .B(n55297), .X(n29462) );
  nand_x2_sg U48174 ( .A(n44915), .B(n55317), .X(n29456) );
  nand_x2_sg U48175 ( .A(n45149), .B(n55342), .X(n29450) );
  inv_x1_sg U48176 ( .A(n21998), .X(n50948) );
  nand_x1_sg U48177 ( .A(n8483), .B(n21997), .X(n21996) );
  nand_x1_sg U48178 ( .A(n8543), .B(n22615), .X(n22614) );
  nand_x1_sg U48179 ( .A(n8623), .B(n22587), .X(n22586) );
  inv_x1_sg U48180 ( .A(n21984), .X(n50941) );
  nand_x1_sg U48181 ( .A(n8523), .B(n21983), .X(n21982) );
  inv_x1_sg U48182 ( .A(n22608), .X(n50937) );
  nand_x1_sg U48183 ( .A(n8563), .B(n22607), .X(n22606) );
  inv_x1_sg U48184 ( .A(n22594), .X(n50931) );
  nand_x1_sg U48185 ( .A(n8603), .B(n22593), .X(n22592) );
  nand_x1_sg U48186 ( .A(n22537), .B(n40739), .X(n22536) );
  nand_x1_sg U48187 ( .A(n8763), .B(n40803), .X(n22539) );
  nand_x1_sg U48188 ( .A(out_L2[19]), .B(n40804), .X(n22540) );
  inv_x1_sg U48189 ( .A(n22550), .X(n50914) );
  nand_x1_sg U48190 ( .A(n8723), .B(n22549), .X(n22548) );
  inv_x2_sg U48191 ( .A(n22517), .X(n45370) );
  nor_x1_sg U48192 ( .A(n22570), .B(n50923), .X(n22517) );
  nand_x1_sg U48193 ( .A(n8643), .B(n22579), .X(n22578) );
  inv_x1_sg U48194 ( .A(n22557), .X(n50918) );
  nand_x1_sg U48195 ( .A(n8703), .B(n22556), .X(n22555) );
  nor_x1_sg U48196 ( .A(n21965), .B(n22529), .X(n22528) );
  inv_x1_sg U48197 ( .A(n22565), .X(n50920) );
  nand_x1_sg U48198 ( .A(n8683), .B(n22564), .X(n22563) );
  inv_x1_sg U48199 ( .A(n9413), .X(n50901) );
  nand_x1_sg U48200 ( .A(n8484), .B(n9412), .X(n9411) );
  nand_x1_sg U48201 ( .A(n8544), .B(n22184), .X(n22183) );
  nand_x1_sg U48202 ( .A(n8624), .B(n22591), .X(n22851) );
  inv_x1_sg U48203 ( .A(n22186), .X(n50896) );
  nand_x1_sg U48204 ( .A(n8524), .B(n21988), .X(n22185) );
  inv_x1_sg U48205 ( .A(n22869), .X(n50908) );
  nand_x1_sg U48206 ( .A(n8564), .B(n22612), .X(n22868) );
  inv_x1_sg U48207 ( .A(n22857), .X(n50889) );
  nand_x1_sg U48208 ( .A(n8604), .B(n22598), .X(n22856) );
  inv_x2_sg U48209 ( .A(n22807), .X(n44730) );
  inv_x2_sg U48210 ( .A(n22847), .X(n44734) );
  inv_x2_sg U48211 ( .A(n22803), .X(n44646) );
  nor_x1_sg U48212 ( .A(n22813), .B(n50867), .X(n22803) );
  inv_x1_sg U48213 ( .A(n22834), .X(n50877) );
  nand_x1_sg U48214 ( .A(n8684), .B(n22569), .X(n22833) );
  inv_x1_sg U48215 ( .A(n9463), .X(n50852) );
  nand_x1_sg U48216 ( .A(n8485), .B(n9462), .X(n9461) );
  nand_x1_sg U48217 ( .A(n8545), .B(n22350), .X(n22349) );
  inv_x2_sg U48218 ( .A(n23045), .X(n45386) );
  nor_x1_sg U48219 ( .A(n23094), .B(n50836), .X(n23045) );
  inv_x1_sg U48220 ( .A(n22773), .X(n50860) );
  nand_x1_sg U48221 ( .A(n8565), .B(n22772), .X(n22771) );
  inv_x1_sg U48222 ( .A(n23114), .X(n50844) );
  nand_x1_sg U48223 ( .A(n8605), .B(n22861), .X(n23113) );
  nand_x1_sg U48224 ( .A(n8625), .B(n22855), .X(n23108) );
  inv_x1_sg U48225 ( .A(n23092), .X(n50832) );
  inv_x1_sg U48226 ( .A(n9512), .X(n50807) );
  nand_x1_sg U48227 ( .A(n8486), .B(n9511), .X(n9510) );
  nand_x1_sg U48228 ( .A(n8546), .B(n22497), .X(n22496) );
  inv_x2_sg U48229 ( .A(n23271), .X(n45334) );
  nor_x1_sg U48230 ( .A(n23320), .B(n50792), .X(n23271) );
  inv_x1_sg U48231 ( .A(n22767), .X(n50816) );
  nand_x1_sg U48232 ( .A(n8566), .B(n22766), .X(n22765) );
  inv_x1_sg U48233 ( .A(n23338), .X(n50820) );
  nand_x1_sg U48234 ( .A(n8606), .B(n23118), .X(n23337) );
  nand_x1_sg U48235 ( .A(n8626), .B(n23112), .X(n23332) );
  inv_x1_sg U48236 ( .A(n22337), .X(n50848) );
  inv_x1_sg U48237 ( .A(n23318), .X(n50788) );
  nand_x1_sg U48238 ( .A(n8646), .B(n50795), .X(n23327) );
  inv_x1_sg U48239 ( .A(n23287), .X(n50822) );
  inv_x1_sg U48240 ( .A(n9561), .X(n50759) );
  nand_x1_sg U48241 ( .A(n8487), .B(n9560), .X(n9559) );
  nand_x1_sg U48242 ( .A(n8547), .B(n22491), .X(n22490) );
  inv_x2_sg U48243 ( .A(n23476), .X(n45384) );
  nor_x1_sg U48244 ( .A(n23525), .B(n50746), .X(n23476) );
  inv_x1_sg U48245 ( .A(n22761), .X(n50768) );
  nand_x1_sg U48246 ( .A(n8567), .B(n22760), .X(n22759) );
  inv_x1_sg U48247 ( .A(n23260), .X(n50772) );
  nand_x1_sg U48248 ( .A(n8607), .B(n23259), .X(n23258) );
  nand_x1_sg U48249 ( .A(n8627), .B(n23336), .X(n23539) );
  inv_x1_sg U48250 ( .A(n22331), .X(n50803) );
  inv_x1_sg U48251 ( .A(n23523), .X(n50742) );
  inv_x1_sg U48252 ( .A(n9609), .X(n50712) );
  nand_x1_sg U48253 ( .A(n8488), .B(n9608), .X(n9607) );
  nand_x1_sg U48254 ( .A(n8548), .B(n22485), .X(n22484) );
  inv_x2_sg U48255 ( .A(n23666), .X(n45332) );
  nor_x1_sg U48256 ( .A(n23715), .B(n50700), .X(n23666) );
  nand_x1_sg U48257 ( .A(n8628), .B(n23468), .X(n23467) );
  inv_x1_sg U48258 ( .A(n22325), .X(n50755) );
  inv_x1_sg U48259 ( .A(n22755), .X(n50721) );
  nand_x1_sg U48260 ( .A(n8568), .B(n22754), .X(n22753) );
  inv_x1_sg U48261 ( .A(n23250), .X(n50751) );
  inv_x1_sg U48262 ( .A(n23713), .X(n50696) );
  nand_x1_sg U48263 ( .A(n8648), .B(n50730), .X(n23722) );
  inv_x1_sg U48264 ( .A(n23682), .X(n50732) );
  inv_x1_sg U48265 ( .A(n9657), .X(n50664) );
  nand_x1_sg U48266 ( .A(n8489), .B(n9656), .X(n9655) );
  nand_x1_sg U48267 ( .A(n8549), .B(n22479), .X(n22478) );
  inv_x2_sg U48268 ( .A(n23837), .X(n45382) );
  nor_x1_sg U48269 ( .A(n23886), .B(n50683), .X(n23837) );
  nand_x1_sg U48270 ( .A(n8629), .B(n23462), .X(n23461) );
  inv_x1_sg U48271 ( .A(n22319), .X(n50708) );
  inv_x1_sg U48272 ( .A(n22749), .X(n50673) );
  nand_x1_sg U48273 ( .A(n8569), .B(n22748), .X(n22747) );
  inv_x1_sg U48274 ( .A(n23244), .X(n50704) );
  inv_x1_sg U48275 ( .A(n23884), .X(n50651) );
  nand_x1_sg U48276 ( .A(n8630), .B(n23456), .X(n23455) );
  inv_x1_sg U48277 ( .A(n22313), .X(n50660) );
  inv_x1_sg U48278 ( .A(n22743), .X(n50626) );
  nand_x1_sg U48279 ( .A(n8570), .B(n22742), .X(n22741) );
  inv_x1_sg U48280 ( .A(n23238), .X(n50657) );
  inv_x1_sg U48281 ( .A(n9704), .X(n50617) );
  nand_x1_sg U48282 ( .A(n8490), .B(n9703), .X(n9702) );
  inv_x1_sg U48283 ( .A(n24037), .X(n50638) );
  inv_x1_sg U48284 ( .A(n24006), .X(n50641) );
  inv_x1_sg U48285 ( .A(n9752), .X(n50568) );
  nand_x1_sg U48286 ( .A(n8491), .B(n9751), .X(n9750) );
  nand_x1_sg U48287 ( .A(n8551), .B(n22467), .X(n22466) );
  inv_x2_sg U48288 ( .A(n23825), .X(n45380) );
  nor_x1_sg U48289 ( .A(n23827), .B(n50587), .X(n23825) );
  nand_x1_sg U48290 ( .A(n8631), .B(n23450), .X(n23449) );
  inv_x1_sg U48291 ( .A(n22307), .X(n50613) );
  inv_x1_sg U48292 ( .A(n22737), .X(n50577) );
  nand_x1_sg U48293 ( .A(n8571), .B(n22736), .X(n22735) );
  inv_x1_sg U48294 ( .A(n23232), .X(n50609) );
  inv_x1_sg U48295 ( .A(n24040), .X(n50588) );
  inv_x1_sg U48296 ( .A(n9800), .X(n50521) );
  nand_x1_sg U48297 ( .A(n8492), .B(n9799), .X(n9798) );
  nand_x1_sg U48298 ( .A(n8552), .B(n22461), .X(n22460) );
  inv_x2_sg U48299 ( .A(n23819), .X(n45378) );
  nor_x1_sg U48300 ( .A(n23821), .B(n50541), .X(n23819) );
  nand_x1_sg U48301 ( .A(n8632), .B(n23444), .X(n23443) );
  inv_x1_sg U48302 ( .A(n22301), .X(n50564) );
  inv_x1_sg U48303 ( .A(n22731), .X(n50530) );
  nand_x1_sg U48304 ( .A(n8572), .B(n22730), .X(n22729) );
  inv_x1_sg U48305 ( .A(n23226), .X(n50560) );
  inv_x1_sg U48306 ( .A(n24043), .X(n50542) );
  inv_x1_sg U48307 ( .A(n24266), .X(n50549) );
  inv_x1_sg U48308 ( .A(n9848), .X(n50474) );
  nand_x1_sg U48309 ( .A(n8493), .B(n9847), .X(n9846) );
  nand_x1_sg U48310 ( .A(n8553), .B(n22455), .X(n22454) );
  inv_x2_sg U48311 ( .A(n23813), .X(n45368) );
  nor_x1_sg U48312 ( .A(n23815), .B(n50493), .X(n23813) );
  nand_x1_sg U48313 ( .A(n8633), .B(n23438), .X(n23437) );
  inv_x1_sg U48314 ( .A(n22295), .X(n50517) );
  inv_x1_sg U48315 ( .A(n22725), .X(n50483) );
  nand_x1_sg U48316 ( .A(n8573), .B(n22724), .X(n22723) );
  inv_x1_sg U48317 ( .A(n23220), .X(n50513) );
  inv_x1_sg U48318 ( .A(n24046), .X(n50494) );
  inv_x1_sg U48319 ( .A(n24253), .X(n50507) );
  inv_x2_sg U48320 ( .A(n24127), .X(n44526) );
  nor_x1_sg U48321 ( .A(n24129), .B(n50497), .X(n24127) );
  inv_x1_sg U48322 ( .A(n9896), .X(n50428) );
  nand_x1_sg U48323 ( .A(n8494), .B(n9895), .X(n9894) );
  nand_x1_sg U48324 ( .A(n8554), .B(n22449), .X(n22448) );
  inv_x2_sg U48325 ( .A(n23807), .X(n45366) );
  nor_x1_sg U48326 ( .A(n23809), .B(n50447), .X(n23807) );
  nand_x1_sg U48327 ( .A(n8634), .B(n23432), .X(n23431) );
  inv_x1_sg U48328 ( .A(n22289), .X(n50470) );
  inv_x1_sg U48329 ( .A(n22719), .X(n50437) );
  nand_x1_sg U48330 ( .A(n8574), .B(n22718), .X(n22717) );
  inv_x1_sg U48331 ( .A(n23214), .X(n50466) );
  inv_x1_sg U48332 ( .A(n24049), .X(n50448) );
  inv_x1_sg U48333 ( .A(n24247), .X(n50460) );
  inv_x2_sg U48334 ( .A(n24120), .X(n44524) );
  nor_x1_sg U48335 ( .A(n24122), .B(n50451), .X(n24120) );
  inv_x1_sg U48336 ( .A(n9944), .X(n50381) );
  nand_x1_sg U48337 ( .A(n8495), .B(n9943), .X(n9942) );
  nand_x1_sg U48338 ( .A(n8555), .B(n22443), .X(n22442) );
  inv_x2_sg U48339 ( .A(n23801), .X(n45364) );
  nor_x1_sg U48340 ( .A(n23803), .B(n50401), .X(n23801) );
  nand_x1_sg U48341 ( .A(n8635), .B(n23426), .X(n23425) );
  inv_x1_sg U48342 ( .A(n22283), .X(n50424) );
  inv_x1_sg U48343 ( .A(n22713), .X(n50390) );
  nand_x1_sg U48344 ( .A(n8575), .B(n22712), .X(n22711) );
  inv_x1_sg U48345 ( .A(n23208), .X(n50420) );
  inv_x1_sg U48346 ( .A(n24052), .X(n50402) );
  inv_x1_sg U48347 ( .A(n24241), .X(n50414) );
  inv_x2_sg U48348 ( .A(n24113), .X(n44522) );
  nor_x1_sg U48349 ( .A(n24115), .B(n50405), .X(n24113) );
  nand_x1_sg U48350 ( .A(n50412), .B(n50364), .X(n24438) );
  inv_x1_sg U48351 ( .A(n24440), .X(n50412) );
  inv_x2_sg U48352 ( .A(n24351), .X(n45492) );
  nor_x1_sg U48353 ( .A(n24353), .B(n50410), .X(n24351) );
  inv_x1_sg U48354 ( .A(n23202), .X(n50373) );
  inv_x2_sg U48355 ( .A(n22959), .X(n44642) );
  nor_x1_sg U48356 ( .A(n22961), .B(n50345), .X(n22959) );
  inv_x1_sg U48357 ( .A(n22707), .X(n50343) );
  nand_x1_sg U48358 ( .A(n8576), .B(n22706), .X(n22705) );
  nand_x1_sg U48359 ( .A(n8776), .B(n40805), .X(n24436) );
  inv_x2_sg U48360 ( .A(n23795), .X(n45376) );
  nor_x1_sg U48361 ( .A(n23797), .B(n50353), .X(n23795) );
  inv_x1_sg U48362 ( .A(n9993), .X(n50334) );
  nand_x1_sg U48363 ( .A(n8496), .B(n9992), .X(n9991) );
  nand_x1_sg U48364 ( .A(n8636), .B(n23420), .X(n23419) );
  inv_x1_sg U48365 ( .A(n22277), .X(n50377) );
  inv_x1_sg U48366 ( .A(n24055), .X(n50354) );
  inv_x1_sg U48367 ( .A(n24235), .X(n50367) );
  inv_x2_sg U48368 ( .A(n24106), .X(n44628) );
  nor_x1_sg U48369 ( .A(n24108), .B(n50357), .X(n24106) );
  nand_x1_sg U48370 ( .A(n8756), .B(n24348), .X(n24347) );
  inv_x1_sg U48371 ( .A(n10041), .X(n50288) );
  nand_x1_sg U48372 ( .A(n8497), .B(n10040), .X(n10039) );
  nand_x1_sg U48373 ( .A(n8557), .B(n22431), .X(n22430) );
  inv_x2_sg U48374 ( .A(n23789), .X(n45362) );
  nor_x1_sg U48375 ( .A(n23791), .B(n50307), .X(n23789) );
  nand_x1_sg U48376 ( .A(n8637), .B(n23414), .X(n23413) );
  inv_x1_sg U48377 ( .A(n22271), .X(n50330) );
  inv_x1_sg U48378 ( .A(n22701), .X(n50297) );
  nand_x1_sg U48379 ( .A(n8577), .B(n22700), .X(n22699) );
  inv_x1_sg U48380 ( .A(n23196), .X(n50326) );
  inv_x1_sg U48381 ( .A(n24058), .X(n50308) );
  inv_x1_sg U48382 ( .A(n24229), .X(n50320) );
  inv_x2_sg U48383 ( .A(n24099), .X(n44520) );
  nor_x1_sg U48384 ( .A(n24101), .B(n50311), .X(n24099) );
  inv_x1_sg U48385 ( .A(n24429), .X(n50318) );
  inv_x2_sg U48386 ( .A(n24338), .X(n45494) );
  nor_x1_sg U48387 ( .A(n24340), .B(n50316), .X(n24338) );
  inv_x1_sg U48388 ( .A(n23190), .X(n50280) );
  inv_x2_sg U48389 ( .A(n22945), .X(n44640) );
  nor_x1_sg U48390 ( .A(n22947), .B(n50253), .X(n22945) );
  inv_x1_sg U48391 ( .A(n22695), .X(n50251) );
  nand_x1_sg U48392 ( .A(n8578), .B(n22694), .X(n22693) );
  inv_x1_sg U48393 ( .A(n10090), .X(n50242) );
  nand_x1_sg U48394 ( .A(n8498), .B(n10089), .X(n10088) );
  nand_x1_sg U48395 ( .A(n8638), .B(n23408), .X(n23407) );
  inv_x1_sg U48396 ( .A(n22265), .X(n50284) );
  inv_x1_sg U48397 ( .A(n23756), .X(n50259) );
  nand_x1_sg U48398 ( .A(n8659), .B(n23755), .X(n23754) );
  inv_x2_sg U48399 ( .A(n23783), .X(n45374) );
  nor_x1_sg U48400 ( .A(n23785), .B(n50262), .X(n23783) );
  nand_x1_sg U48401 ( .A(n8758), .B(n24335), .X(n24334) );
  inv_x1_sg U48402 ( .A(n23949), .X(n50264) );
  nand_x1_sg U48403 ( .A(n8698), .B(n23948), .X(n23947) );
  inv_x1_sg U48404 ( .A(n24223), .X(n50274) );
  inv_x2_sg U48405 ( .A(n24092), .X(n44626) );
  nor_x1_sg U48406 ( .A(n24094), .B(n50266), .X(n24092) );
  inv_x1_sg U48407 ( .A(n23184), .X(n50234) );
  inv_x2_sg U48408 ( .A(n22938), .X(n44650) );
  nor_x1_sg U48409 ( .A(n22940), .B(n50209), .X(n22938) );
  inv_x1_sg U48410 ( .A(n22689), .X(n50207) );
  nand_x1_sg U48411 ( .A(n8579), .B(n22688), .X(n22687) );
  inv_x1_sg U48412 ( .A(n10139), .X(n50198) );
  nand_x1_sg U48413 ( .A(n8499), .B(n10138), .X(n10137) );
  nand_x1_sg U48414 ( .A(n8639), .B(n23402), .X(n23401) );
  inv_x1_sg U48415 ( .A(n22259), .X(n50238) );
  inv_x2_sg U48416 ( .A(n23777), .X(n45372) );
  nor_x1_sg U48417 ( .A(n23779), .B(n50217), .X(n23777) );
  nand_x1_sg U48418 ( .A(n8759), .B(n24329), .X(n24328) );
  inv_x1_sg U48419 ( .A(n23943), .X(n50219) );
  nand_x1_sg U48420 ( .A(n8699), .B(n23942), .X(n23941) );
  inv_x1_sg U48421 ( .A(n24217), .X(n50228) );
  inv_x2_sg U48422 ( .A(n24085), .X(n44624) );
  nor_x1_sg U48423 ( .A(n24087), .B(n50221), .X(n24085) );
  inv_x1_sg U48424 ( .A(n23178), .X(n50190) );
  inv_x2_sg U48425 ( .A(n22931), .X(n44071) );
  nor_x1_sg U48426 ( .A(n22933), .B(n50163), .X(n22931) );
  inv_x1_sg U48427 ( .A(n22683), .X(n50161) );
  nand_x1_sg U48428 ( .A(n8580), .B(n22682), .X(n22681) );
  inv_x1_sg U48429 ( .A(n10186), .X(n50155) );
  nand_x1_sg U48430 ( .A(n8500), .B(n10185), .X(n10184) );
  nand_x1_sg U48431 ( .A(n8640), .B(n23396), .X(n23395) );
  inv_x1_sg U48432 ( .A(n22253), .X(n50194) );
  inv_x1_sg U48433 ( .A(n24211), .X(n50184) );
  inv_x2_sg U48434 ( .A(n24078), .X(n44518) );
  nor_x1_sg U48435 ( .A(n24080), .B(n50173), .X(n24078) );
  nand_x1_sg U48436 ( .A(n8660), .B(n23595), .X(n23594) );
  nand_x1_sg U48437 ( .A(n24410), .B(n24411), .X(n24408) );
  inv_x1_sg U48438 ( .A(n24410), .X(n50182) );
  inv_x2_sg U48439 ( .A(n24319), .X(n44246) );
  nor_x1_sg U48440 ( .A(n24321), .B(n50177), .X(n24319) );
  nand_x1_sg U48441 ( .A(n23172), .B(n50132), .X(n23171) );
  inv_x1_sg U48442 ( .A(n23173), .X(n50132) );
  nand_x2_sg U48443 ( .A(n22675), .B(n22676), .X(n22674) );
  nand_x1_sg U48444 ( .A(n22924), .B(n50131), .X(n22923) );
  inv_x1_sg U48445 ( .A(n22925), .X(n50131) );
  inv_x1_sg U48446 ( .A(n24405), .X(n50140) );
  nand_x2_sg U48447 ( .A(n23767), .B(n23768), .X(n23766) );
  nand_x1_sg U48448 ( .A(n10213), .B(n50129), .X(n22403) );
  nand_x1_sg U48449 ( .A(n22404), .B(n50151), .X(n22402) );
  inv_x1_sg U48450 ( .A(n22404), .X(n50129) );
  nand_x2_sg U48451 ( .A(n10228), .B(n10229), .X(n10227) );
  inv_x1_sg U48452 ( .A(n10227), .X(n50126) );
  nand_x1_sg U48453 ( .A(n22056), .B(n50127), .X(n22055) );
  inv_x1_sg U48454 ( .A(n22057), .X(n50127) );
  nand_x1_sg U48455 ( .A(n22247), .B(n50128), .X(n22246) );
  inv_x1_sg U48456 ( .A(n22248), .X(n50128) );
  nand_x2_sg U48457 ( .A(n24073), .B(n24074), .X(n24072) );
  nand_x1_sg U48458 ( .A(n24205), .B(n50138), .X(n24204) );
  inv_x1_sg U48459 ( .A(n24206), .X(n50138) );
  nand_x2_sg U48460 ( .A(n23929), .B(n23930), .X(n23928) );
  nand_x1_sg U48461 ( .A(n24312), .B(n50139), .X(n24311) );
  inv_x1_sg U48462 ( .A(n24313), .X(n50139) );
  nand_x2_sg U48463 ( .A(n23586), .B(n23587), .X(n23585) );
  nand_x2_sg U48464 ( .A(n25608), .B(n25609), .X(n25607) );
  inv_x1_sg U48465 ( .A(n25607), .X(n51255) );
  inv_x1_sg U48466 ( .A(n25597), .X(n43873) );
  inv_x1_sg U48467 ( .A(n10423), .X(n51273) );
  inv_x2_sg U48468 ( .A(n10411), .X(n44474) );
  nor_x1_sg U48469 ( .A(n10419), .B(n10420), .X(n10411) );
  inv_x2_sg U48470 ( .A(n10428), .X(n44368) );
  nor_x1_sg U48471 ( .A(n51269), .B(n10424), .X(n10428) );
  nand_x1_sg U48472 ( .A(n10408), .B(n10458), .X(n10456) );
  nand_x1_sg U48473 ( .A(n10475), .B(n10476), .X(n10474) );
  nand_x1_sg U48474 ( .A(n46564), .B(n10477), .X(n10476) );
  inv_x2_sg U48475 ( .A(n10467), .X(n44105) );
  nor_x1_sg U48476 ( .A(n51325), .B(n10479), .X(n10467) );
  nand_x1_sg U48477 ( .A(n10534), .B(n51349), .X(n10533) );
  inv_x1_sg U48478 ( .A(n10535), .X(n51349) );
  inv_x2_sg U48479 ( .A(n10465), .X(n45484) );
  nand_x1_sg U48480 ( .A(n44106), .B(n51314), .X(n10465) );
  nand_x4_sg U48481 ( .A(n10593), .B(n10594), .X(n10586) );
  nand_x1_sg U48482 ( .A(n51369), .B(n10595), .X(n10594) );
  nand_x1_sg U48483 ( .A(n51401), .B(n10596), .X(n10593) );
  nand_x4_sg U48484 ( .A(n10632), .B(n10633), .X(n10623) );
  nand_x1_sg U48485 ( .A(n10634), .B(n51424), .X(n10633) );
  inv_x1_sg U48486 ( .A(n10635), .X(n51424) );
  nand_x1_sg U48487 ( .A(n10683), .B(n10682), .X(n10680) );
  inv_x1_sg U48488 ( .A(n10682), .X(n51412) );
  inv_x2_sg U48489 ( .A(n10671), .X(n45402) );
  nor_x1_sg U48490 ( .A(n51430), .B(n10677), .X(n10671) );
  nand_x4_sg U48491 ( .A(n10665), .B(n51409), .X(n10631) );
  inv_x1_sg U48492 ( .A(n10666), .X(n51409) );
  inv_x1_sg U48493 ( .A(n10629), .X(n51411) );
  nand_x1_sg U48494 ( .A(n10631), .B(n10630), .X(n10628) );
  inv_x1_sg U48495 ( .A(n10623), .X(n51425) );
  nand_x4_sg U48496 ( .A(n10639), .B(n10640), .X(n10630) );
  nand_x1_sg U48497 ( .A(n51369), .B(n51401), .X(n10640) );
  inv_x1_sg U48498 ( .A(n10724), .X(n51469) );
  nand_x1_sg U48499 ( .A(n51423), .B(n10722), .X(n10721) );
  inv_x1_sg U48500 ( .A(n10723), .X(n51423) );
  inv_x1_sg U48501 ( .A(n10824), .X(n51507) );
  nand_x1_sg U48502 ( .A(n40566), .B(n10773), .X(n10770) );
  inv_x2_sg U48503 ( .A(n10761), .X(n45454) );
  nor_x1_sg U48504 ( .A(n51493), .B(n10767), .X(n10761) );
  nand_x4_sg U48505 ( .A(n10825), .B(n10826), .X(n10365) );
  nand_x1_sg U48506 ( .A(n42382), .B(n10773), .X(n10826) );
  inv_x1_sg U48507 ( .A(n10874), .X(n51444) );
  inv_x1_sg U48508 ( .A(n10926), .X(n51514) );
  nand_x2_sg U48509 ( .A(n25889), .B(n25890), .X(n25888) );
  inv_x1_sg U48510 ( .A(n25888), .X(n51531) );
  inv_x1_sg U48511 ( .A(n25878), .X(n44019) );
  nand_x1_sg U48512 ( .A(n51543), .B(n46547), .X(n11172) );
  nand_x1_sg U48513 ( .A(n11194), .B(n46540), .X(n11193) );
  inv_x2_sg U48514 ( .A(n11196), .X(n45600) );
  nand_x1_sg U48515 ( .A(n11211), .B(n11207), .X(n11212) );
  nand_x1_sg U48516 ( .A(n11251), .B(n11252), .X(n11250) );
  nand_x1_sg U48517 ( .A(n46540), .B(n11231), .X(n11252) );
  inv_x2_sg U48518 ( .A(n11243), .X(n43995) );
  nor_x1_sg U48519 ( .A(n51600), .B(n11255), .X(n11243) );
  nand_x1_sg U48520 ( .A(n46540), .B(n51589), .X(n11230) );
  nand_x1_sg U48521 ( .A(n46541), .B(n11231), .X(n11229) );
  inv_x1_sg U48522 ( .A(n11231), .X(n51589) );
  inv_x1_sg U48523 ( .A(n11222), .X(n51584) );
  inv_x1_sg U48524 ( .A(n11237), .X(n51582) );
  nand_x1_sg U48525 ( .A(n11239), .B(n11238), .X(n11236) );
  inv_x1_sg U48526 ( .A(n11215), .X(n51571) );
  inv_x2_sg U48527 ( .A(n11270), .X(n44075) );
  nor_x1_sg U48528 ( .A(n11279), .B(n11280), .X(n11270) );
  inv_x1_sg U48529 ( .A(n11308), .X(n51632) );
  inv_x2_sg U48530 ( .A(n11241), .X(n45482) );
  nand_x1_sg U48531 ( .A(n43996), .B(n41939), .X(n11241) );
  nand_x1_sg U48532 ( .A(n45551), .B(n11360), .X(n11358) );
  nand_x4_sg U48533 ( .A(n11370), .B(n11371), .X(n11363) );
  nand_x1_sg U48534 ( .A(n51640), .B(n11372), .X(n11371) );
  nand_x1_sg U48535 ( .A(n51678), .B(n11373), .X(n11370) );
  nand_x4_sg U48536 ( .A(n11411), .B(n11412), .X(n11401) );
  nand_x1_sg U48537 ( .A(n11413), .B(n11414), .X(n11412) );
  nand_x4_sg U48538 ( .A(n11445), .B(n51687), .X(n11410) );
  inv_x1_sg U48539 ( .A(n11446), .X(n51687) );
  inv_x1_sg U48540 ( .A(n11408), .X(n51689) );
  nand_x1_sg U48541 ( .A(n11410), .B(n11409), .X(n11407) );
  inv_x1_sg U48542 ( .A(n11401), .X(n51699) );
  nand_x4_sg U48543 ( .A(n11418), .B(n11419), .X(n11409) );
  nand_x1_sg U48544 ( .A(n51640), .B(n51678), .X(n11419) );
  nand_x1_sg U48545 ( .A(n51704), .B(n11503), .X(n11502) );
  inv_x1_sg U48546 ( .A(n11504), .X(n51704) );
  inv_x1_sg U48547 ( .A(n11505), .X(n51749) );
  inv_x1_sg U48548 ( .A(n11604), .X(n51787) );
  inv_x2_sg U48549 ( .A(n11601), .X(n45450) );
  nor_x1_sg U48550 ( .A(n11661), .B(n45453), .X(n11601) );
  nand_x1_sg U48551 ( .A(n40567), .B(n11552), .X(n11549) );
  inv_x2_sg U48552 ( .A(n11543), .X(n44192) );
  nor_x1_sg U48553 ( .A(n51772), .B(n11553), .X(n11543) );
  inv_x1_sg U48554 ( .A(n11654), .X(n51734) );
  nand_x1_sg U48555 ( .A(n11656), .B(n11655), .X(n11653) );
  nand_x4_sg U48556 ( .A(n11605), .B(n11606), .X(n11132) );
  nand_x1_sg U48557 ( .A(n42384), .B(n11552), .X(n11606) );
  inv_x1_sg U48558 ( .A(n11670), .X(n51800) );
  nand_x2_sg U48559 ( .A(n26169), .B(n26170), .X(n26168) );
  inv_x1_sg U48560 ( .A(n26168), .X(n51813) );
  inv_x1_sg U48561 ( .A(n26158), .X(n44031) );
  nand_x1_sg U48562 ( .A(n51819), .B(n46525), .X(n11946) );
  inv_x2_sg U48563 ( .A(n11975), .X(n45592) );
  nand_x4_sg U48564 ( .A(n11970), .B(n11971), .X(n11961) );
  nand_x1_sg U48565 ( .A(n11973), .B(n11974), .X(n11970) );
  nand_x1_sg U48566 ( .A(n11972), .B(n46517), .X(n11971) );
  nand_x1_sg U48567 ( .A(n46517), .B(n46525), .X(n11974) );
  nand_x1_sg U48568 ( .A(n12027), .B(n12028), .X(n12026) );
  nand_x1_sg U48569 ( .A(n46517), .B(n12031), .X(n12027) );
  inv_x2_sg U48570 ( .A(n12019), .X(n43993) );
  nor_x1_sg U48571 ( .A(n51881), .B(n12032), .X(n12019) );
  nand_x1_sg U48572 ( .A(n46518), .B(n12008), .X(n12006) );
  nand_x4_sg U48573 ( .A(n12009), .B(n51860), .X(n11997) );
  inv_x1_sg U48574 ( .A(n12010), .X(n51860) );
  nand_x1_sg U48575 ( .A(n12011), .B(n12012), .X(n12009) );
  nand_x4_sg U48576 ( .A(n12013), .B(n12014), .X(n12011) );
  nand_x1_sg U48577 ( .A(n51846), .B(n12015), .X(n12014) );
  nand_x1_sg U48578 ( .A(n51859), .B(n12016), .X(n12013) );
  inv_x1_sg U48579 ( .A(n12015), .X(n51859) );
  inv_x2_sg U48580 ( .A(n12049), .X(n45528) );
  nor_x1_sg U48581 ( .A(n12058), .B(n12059), .X(n12049) );
  inv_x1_sg U48582 ( .A(n12088), .X(n51913) );
  inv_x2_sg U48583 ( .A(n12017), .X(n45480) );
  nand_x1_sg U48584 ( .A(n43994), .B(n51874), .X(n12017) );
  nand_x1_sg U48585 ( .A(n45549), .B(n12140), .X(n12138) );
  nand_x4_sg U48586 ( .A(n12150), .B(n12151), .X(n12143) );
  nand_x1_sg U48587 ( .A(n51921), .B(n12152), .X(n12151) );
  nand_x1_sg U48588 ( .A(n51959), .B(n12153), .X(n12150) );
  nand_x4_sg U48589 ( .A(n12191), .B(n12192), .X(n12181) );
  nand_x1_sg U48590 ( .A(n12193), .B(n51979), .X(n12192) );
  inv_x1_sg U48591 ( .A(n12194), .X(n51979) );
  nand_x4_sg U48592 ( .A(n12198), .B(n12199), .X(n12189) );
  nand_x1_sg U48593 ( .A(n51921), .B(n51959), .X(n12199) );
  inv_x1_sg U48594 ( .A(n12190), .X(n51968) );
  nand_x4_sg U48595 ( .A(n12187), .B(n51969), .X(n12180) );
  inv_x1_sg U48596 ( .A(n12188), .X(n51969) );
  nand_x1_sg U48597 ( .A(n12190), .B(n12189), .X(n12187) );
  nand_x1_sg U48598 ( .A(n51978), .B(n12283), .X(n12282) );
  inv_x1_sg U48599 ( .A(n12284), .X(n51978) );
  inv_x1_sg U48600 ( .A(n12285), .X(n52032) );
  nand_x1_sg U48601 ( .A(n40545), .B(n11915), .X(n12384) );
  nand_x1_sg U48602 ( .A(n43302), .B(n12332), .X(n12329) );
  inv_x2_sg U48603 ( .A(n12323), .X(n44190) );
  nor_x1_sg U48604 ( .A(n52052), .B(n12333), .X(n12323) );
  inv_x1_sg U48605 ( .A(n12434), .X(n52012) );
  nand_x1_sg U48606 ( .A(n12436), .B(n12435), .X(n12433) );
  inv_x1_sg U48607 ( .A(n12450), .X(n52076) );
  nand_x2_sg U48608 ( .A(n26448), .B(n26449), .X(n26447) );
  inv_x1_sg U48609 ( .A(n26447), .X(n52089) );
  inv_x1_sg U48610 ( .A(n26437), .X(n43897) );
  nand_x1_sg U48611 ( .A(n46500), .B(n46503), .X(n12723) );
  nand_x1_sg U48612 ( .A(n52100), .B(n46503), .X(n12733) );
  nand_x1_sg U48613 ( .A(n12755), .B(n46496), .X(n12754) );
  inv_x2_sg U48614 ( .A(n12757), .X(n45598) );
  nand_x1_sg U48615 ( .A(n12772), .B(n12768), .X(n12773) );
  nand_x1_sg U48616 ( .A(n12812), .B(n12813), .X(n12811) );
  nand_x1_sg U48617 ( .A(n46496), .B(n12792), .X(n12813) );
  inv_x2_sg U48618 ( .A(n12804), .X(n43991) );
  nor_x1_sg U48619 ( .A(n52158), .B(n12816), .X(n12804) );
  nand_x1_sg U48620 ( .A(n46496), .B(n52147), .X(n12791) );
  nand_x1_sg U48621 ( .A(n12734), .B(n12792), .X(n12790) );
  inv_x1_sg U48622 ( .A(n12792), .X(n52147) );
  inv_x1_sg U48623 ( .A(n12783), .X(n52142) );
  inv_x1_sg U48624 ( .A(n12798), .X(n52140) );
  nand_x1_sg U48625 ( .A(n12800), .B(n12799), .X(n12797) );
  inv_x1_sg U48626 ( .A(n12776), .X(n52128) );
  inv_x2_sg U48627 ( .A(n12831), .X(n44282) );
  nor_x1_sg U48628 ( .A(n12840), .B(n12841), .X(n12831) );
  inv_x2_sg U48629 ( .A(n12802), .X(n45478) );
  nand_x1_sg U48630 ( .A(n43992), .B(n41938), .X(n12802) );
  nand_x1_sg U48631 ( .A(n45547), .B(n12921), .X(n12919) );
  nand_x4_sg U48632 ( .A(n12931), .B(n12932), .X(n12924) );
  nand_x1_sg U48633 ( .A(n52196), .B(n12933), .X(n12932) );
  nand_x1_sg U48634 ( .A(n52234), .B(n12934), .X(n12931) );
  nand_x4_sg U48635 ( .A(n12972), .B(n12973), .X(n12962) );
  nand_x1_sg U48636 ( .A(n12974), .B(n12975), .X(n12973) );
  nand_x4_sg U48637 ( .A(n13006), .B(n52242), .X(n12971) );
  inv_x1_sg U48638 ( .A(n13007), .X(n52242) );
  inv_x1_sg U48639 ( .A(n12969), .X(n52244) );
  nand_x1_sg U48640 ( .A(n12971), .B(n12970), .X(n12968) );
  inv_x1_sg U48641 ( .A(n12962), .X(n52255) );
  nand_x4_sg U48642 ( .A(n12979), .B(n12980), .X(n12970) );
  nand_x1_sg U48643 ( .A(n52196), .B(n52234), .X(n12980) );
  nand_x1_sg U48644 ( .A(n52260), .B(n13064), .X(n13063) );
  inv_x1_sg U48645 ( .A(n13065), .X(n52260) );
  inv_x1_sg U48646 ( .A(n13066), .X(n52307) );
  nand_x1_sg U48647 ( .A(n40547), .B(n12693), .X(n13164) );
  inv_x1_sg U48648 ( .A(n13111), .X(n52305) );
  inv_x2_sg U48649 ( .A(n13104), .X(n44188) );
  nor_x1_sg U48650 ( .A(n52329), .B(n13114), .X(n13104) );
  inv_x1_sg U48651 ( .A(n13215), .X(n52289) );
  nand_x1_sg U48652 ( .A(n13217), .B(n13216), .X(n13214) );
  nand_x4_sg U48653 ( .A(n13166), .B(n13167), .X(n12693) );
  nand_x1_sg U48654 ( .A(n44413), .B(n13112), .X(n13167) );
  nand_x1_sg U48655 ( .A(n52299), .B(n13193), .X(n13166) );
  inv_x1_sg U48656 ( .A(n13231), .X(n52354) );
  nand_x1_sg U48657 ( .A(n46582), .B(n26078), .X(n29593) );
  inv_x1_sg U48658 ( .A(n26724), .X(n52366) );
  inv_x1_sg U48659 ( .A(n26715), .X(n43885) );
  nand_x1_sg U48660 ( .A(n46478), .B(n46481), .X(n13508) );
  inv_x2_sg U48661 ( .A(n13536), .X(n45590) );
  nand_x4_sg U48662 ( .A(n13531), .B(n13532), .X(n13522) );
  nand_x1_sg U48663 ( .A(n13533), .B(n46474), .X(n13532) );
  nand_x1_sg U48664 ( .A(n13534), .B(n13535), .X(n13531) );
  nand_x1_sg U48665 ( .A(n13592), .B(n13593), .X(n13591) );
  nand_x1_sg U48666 ( .A(n46474), .B(n13596), .X(n13592) );
  inv_x2_sg U48667 ( .A(n13580), .X(n43849) );
  nor_x1_sg U48668 ( .A(n52432), .B(n13586), .X(n13580) );
  nand_x1_sg U48669 ( .A(n46475), .B(n13569), .X(n13567) );
  nand_x4_sg U48670 ( .A(n13570), .B(n52412), .X(n13558) );
  inv_x1_sg U48671 ( .A(n13571), .X(n52412) );
  nand_x1_sg U48672 ( .A(n13572), .B(n13573), .X(n13570) );
  nand_x4_sg U48673 ( .A(n13574), .B(n13575), .X(n13572) );
  nand_x1_sg U48674 ( .A(n52398), .B(n13576), .X(n13575) );
  nand_x1_sg U48675 ( .A(n52411), .B(n13577), .X(n13574) );
  inv_x1_sg U48676 ( .A(n13576), .X(n52411) );
  inv_x1_sg U48677 ( .A(n13649), .X(n52465) );
  inv_x2_sg U48678 ( .A(n13578), .X(n45476) );
  nand_x1_sg U48679 ( .A(n52426), .B(n43850), .X(n13578) );
  nand_x1_sg U48680 ( .A(n45545), .B(n13701), .X(n13699) );
  nand_x4_sg U48681 ( .A(n13711), .B(n13712), .X(n13704) );
  nand_x1_sg U48682 ( .A(n52473), .B(n13713), .X(n13712) );
  nand_x1_sg U48683 ( .A(n52511), .B(n13714), .X(n13711) );
  nand_x4_sg U48684 ( .A(n13752), .B(n13753), .X(n13742) );
  nand_x1_sg U48685 ( .A(n13754), .B(n13755), .X(n13753) );
  nand_x4_sg U48686 ( .A(n13759), .B(n13760), .X(n13750) );
  nand_x1_sg U48687 ( .A(n52473), .B(n52511), .X(n13760) );
  inv_x1_sg U48688 ( .A(n13751), .X(n52519) );
  nand_x4_sg U48689 ( .A(n13748), .B(n52520), .X(n13741) );
  inv_x1_sg U48690 ( .A(n13749), .X(n52520) );
  nand_x1_sg U48691 ( .A(n13751), .B(n13750), .X(n13748) );
  nand_x1_sg U48692 ( .A(n52536), .B(n13844), .X(n13843) );
  inv_x1_sg U48693 ( .A(n13845), .X(n52536) );
  inv_x1_sg U48694 ( .A(n13846), .X(n52582) );
  nand_x1_sg U48695 ( .A(n40549), .B(n13477), .X(n13944) );
  inv_x1_sg U48696 ( .A(n13891), .X(n52580) );
  inv_x2_sg U48697 ( .A(n13884), .X(n44186) );
  nor_x1_sg U48698 ( .A(n52604), .B(n13894), .X(n13884) );
  inv_x1_sg U48699 ( .A(n13995), .X(n52564) );
  nand_x1_sg U48700 ( .A(n13997), .B(n13996), .X(n13994) );
  nand_x4_sg U48701 ( .A(n13946), .B(n13947), .X(n13477) );
  nand_x1_sg U48702 ( .A(n44411), .B(n13892), .X(n13947) );
  nand_x1_sg U48703 ( .A(n52574), .B(n13973), .X(n13946) );
  inv_x1_sg U48704 ( .A(n14011), .X(n52629) );
  nand_x2_sg U48705 ( .A(n27005), .B(n27006), .X(n27004) );
  inv_x1_sg U48706 ( .A(n27004), .X(n52642) );
  inv_x1_sg U48707 ( .A(n26994), .X(n44027) );
  nand_x1_sg U48708 ( .A(n52648), .B(n46458), .X(n14288) );
  inv_x1_sg U48709 ( .A(n14316), .X(n52662) );
  inv_x2_sg U48710 ( .A(n14303), .X(n44472) );
  nor_x1_sg U48711 ( .A(n14311), .B(n14312), .X(n14303) );
  nand_x1_sg U48712 ( .A(n46451), .B(n14347), .X(n14345) );
  nand_x1_sg U48713 ( .A(n14367), .B(n14368), .X(n14366) );
  nand_x1_sg U48714 ( .A(n46450), .B(n14369), .X(n14368) );
  inv_x2_sg U48715 ( .A(n14359), .X(n44103) );
  nor_x1_sg U48716 ( .A(n52715), .B(n14371), .X(n14359) );
  nand_x1_sg U48717 ( .A(n14426), .B(n52739), .X(n14425) );
  inv_x1_sg U48718 ( .A(n14427), .X(n52739) );
  inv_x2_sg U48719 ( .A(n14357), .X(n45474) );
  nand_x1_sg U48720 ( .A(n44104), .B(n52703), .X(n14357) );
  nand_x1_sg U48721 ( .A(n42146), .B(n14456), .X(n14454) );
  nand_x4_sg U48722 ( .A(n14485), .B(n14486), .X(n14478) );
  nand_x1_sg U48723 ( .A(n52746), .B(n14487), .X(n14486) );
  nand_x1_sg U48724 ( .A(n52790), .B(n14488), .X(n14485) );
  nand_x1_sg U48725 ( .A(n14575), .B(n14574), .X(n14572) );
  inv_x1_sg U48726 ( .A(n14574), .X(n52801) );
  inv_x2_sg U48727 ( .A(n14563), .X(n45400) );
  nor_x1_sg U48728 ( .A(n52820), .B(n14569), .X(n14563) );
  nand_x4_sg U48729 ( .A(n14524), .B(n14525), .X(n14515) );
  nand_x1_sg U48730 ( .A(n14526), .B(n52814), .X(n14525) );
  inv_x1_sg U48731 ( .A(n14527), .X(n52814) );
  nand_x4_sg U48732 ( .A(n14531), .B(n14532), .X(n14522) );
  nand_x1_sg U48733 ( .A(n52746), .B(n52790), .X(n14532) );
  inv_x1_sg U48734 ( .A(n14523), .X(n52799) );
  nand_x4_sg U48735 ( .A(n14520), .B(n52800), .X(n14514) );
  inv_x1_sg U48736 ( .A(n14521), .X(n52800) );
  nand_x1_sg U48737 ( .A(n14523), .B(n14522), .X(n14520) );
  nand_x1_sg U48738 ( .A(n52813), .B(n14614), .X(n14613) );
  inv_x1_sg U48739 ( .A(n14615), .X(n52813) );
  inv_x1_sg U48740 ( .A(n14616), .X(n52858) );
  nand_x1_sg U48741 ( .A(n40568), .B(n14662), .X(n14659) );
  inv_x2_sg U48742 ( .A(n14653), .X(n44454) );
  nor_x1_sg U48743 ( .A(n52882), .B(n14663), .X(n14653) );
  nand_x4_sg U48744 ( .A(n14765), .B(n52834), .X(n14252) );
  inv_x1_sg U48745 ( .A(n14766), .X(n52834) );
  nand_x1_sg U48746 ( .A(n14768), .B(n14767), .X(n14765) );
  nand_x4_sg U48747 ( .A(n14717), .B(n14718), .X(n14256) );
  nand_x1_sg U48748 ( .A(n42392), .B(n14662), .X(n14718) );
  inv_x1_sg U48749 ( .A(n14782), .X(n52910) );
  nand_x2_sg U48750 ( .A(n27285), .B(n27286), .X(n27284) );
  inv_x1_sg U48751 ( .A(n27284), .X(n52923) );
  inv_x1_sg U48752 ( .A(n27274), .X(n43893) );
  nand_x1_sg U48753 ( .A(n46432), .B(n46435), .X(n15056) );
  nand_x1_sg U48754 ( .A(n52934), .B(n46435), .X(n15066) );
  nand_x1_sg U48755 ( .A(n15088), .B(n46428), .X(n15087) );
  inv_x2_sg U48756 ( .A(n15090), .X(n45596) );
  nand_x1_sg U48757 ( .A(n15105), .B(n15101), .X(n15106) );
  nand_x1_sg U48758 ( .A(n15145), .B(n15146), .X(n15144) );
  nand_x1_sg U48759 ( .A(n46428), .B(n15125), .X(n15146) );
  inv_x2_sg U48760 ( .A(n15137), .X(n43989) );
  nor_x1_sg U48761 ( .A(n52992), .B(n15149), .X(n15137) );
  nand_x1_sg U48762 ( .A(n46428), .B(n52981), .X(n15124) );
  nand_x1_sg U48763 ( .A(n15067), .B(n15125), .X(n15123) );
  inv_x1_sg U48764 ( .A(n15125), .X(n52981) );
  inv_x1_sg U48765 ( .A(n15116), .X(n52976) );
  inv_x1_sg U48766 ( .A(n15131), .X(n52974) );
  nand_x1_sg U48767 ( .A(n15133), .B(n15132), .X(n15130) );
  inv_x1_sg U48768 ( .A(n15109), .X(n52962) );
  inv_x2_sg U48769 ( .A(n15164), .X(n44280) );
  nor_x1_sg U48770 ( .A(n15173), .B(n15174), .X(n15164) );
  inv_x2_sg U48771 ( .A(n15135), .X(n45472) );
  nand_x1_sg U48772 ( .A(n43990), .B(n41937), .X(n15135) );
  nand_x1_sg U48773 ( .A(n45543), .B(n15254), .X(n15252) );
  nand_x4_sg U48774 ( .A(n15264), .B(n15265), .X(n15257) );
  nand_x1_sg U48775 ( .A(n53030), .B(n15266), .X(n15265) );
  nand_x1_sg U48776 ( .A(n53068), .B(n15267), .X(n15264) );
  nand_x4_sg U48777 ( .A(n15305), .B(n15306), .X(n15295) );
  nand_x1_sg U48778 ( .A(n15307), .B(n15308), .X(n15306) );
  nand_x4_sg U48779 ( .A(n15339), .B(n53076), .X(n15304) );
  inv_x1_sg U48780 ( .A(n15340), .X(n53076) );
  inv_x1_sg U48781 ( .A(n15302), .X(n53078) );
  nand_x1_sg U48782 ( .A(n15304), .B(n15303), .X(n15301) );
  inv_x1_sg U48783 ( .A(n15295), .X(n53089) );
  nand_x4_sg U48784 ( .A(n15312), .B(n15313), .X(n15303) );
  nand_x1_sg U48785 ( .A(n53030), .B(n53068), .X(n15313) );
  nand_x1_sg U48786 ( .A(n53094), .B(n15397), .X(n15396) );
  inv_x1_sg U48787 ( .A(n15398), .X(n53094) );
  inv_x1_sg U48788 ( .A(n15399), .X(n53141) );
  nand_x1_sg U48789 ( .A(n40553), .B(n15026), .X(n15497) );
  inv_x1_sg U48790 ( .A(n15444), .X(n53139) );
  inv_x2_sg U48791 ( .A(n15437), .X(n44184) );
  nor_x1_sg U48792 ( .A(n53163), .B(n15447), .X(n15437) );
  inv_x1_sg U48793 ( .A(n15548), .X(n53123) );
  nand_x1_sg U48794 ( .A(n15550), .B(n15549), .X(n15547) );
  nand_x4_sg U48795 ( .A(n15499), .B(n15500), .X(n15026) );
  nand_x1_sg U48796 ( .A(n44409), .B(n15445), .X(n15500) );
  nand_x1_sg U48797 ( .A(n53133), .B(n15526), .X(n15499) );
  inv_x1_sg U48798 ( .A(n15564), .X(n53188) );
  nand_x2_sg U48799 ( .A(n27564), .B(n27565), .X(n27563) );
  inv_x1_sg U48800 ( .A(n27563), .X(n53201) );
  inv_x1_sg U48801 ( .A(n27553), .X(n44023) );
  nand_x1_sg U48802 ( .A(n53207), .B(n46413), .X(n15841) );
  nand_x1_sg U48803 ( .A(n46405), .B(n46413), .X(n15869) );
  nand_x1_sg U48804 ( .A(n15922), .B(n15923), .X(n15921) );
  nand_x1_sg U48805 ( .A(n46405), .B(n15926), .X(n15922) );
  inv_x2_sg U48806 ( .A(n15914), .X(n43987) );
  nor_x1_sg U48807 ( .A(n53268), .B(n15927), .X(n15914) );
  nand_x1_sg U48808 ( .A(n15852), .B(n15903), .X(n15901) );
  nand_x4_sg U48809 ( .A(n15904), .B(n53246), .X(n15892) );
  inv_x1_sg U48810 ( .A(n15905), .X(n53246) );
  nand_x1_sg U48811 ( .A(n15906), .B(n15907), .X(n15904) );
  nand_x4_sg U48812 ( .A(n15908), .B(n15909), .X(n15906) );
  nand_x1_sg U48813 ( .A(n53232), .B(n15910), .X(n15909) );
  nand_x1_sg U48814 ( .A(n53245), .B(n15911), .X(n15908) );
  inv_x1_sg U48815 ( .A(n15910), .X(n53245) );
  inv_x2_sg U48816 ( .A(n15944), .X(n44694) );
  nor_x1_sg U48817 ( .A(n15953), .B(n15954), .X(n15944) );
  inv_x1_sg U48818 ( .A(n15983), .X(n53300) );
  inv_x2_sg U48819 ( .A(n15912), .X(n45470) );
  nand_x1_sg U48820 ( .A(n43988), .B(n53261), .X(n15912) );
  nand_x1_sg U48821 ( .A(n45541), .B(n16035), .X(n16033) );
  nand_x4_sg U48822 ( .A(n16045), .B(n16046), .X(n16038) );
  nand_x1_sg U48823 ( .A(n53308), .B(n16047), .X(n16046) );
  nand_x1_sg U48824 ( .A(n53347), .B(n16048), .X(n16045) );
  nand_x4_sg U48825 ( .A(n16086), .B(n16087), .X(n16076) );
  nand_x1_sg U48826 ( .A(n16088), .B(n53368), .X(n16087) );
  inv_x1_sg U48827 ( .A(n16089), .X(n53368) );
  nand_x4_sg U48828 ( .A(n16093), .B(n16094), .X(n16084) );
  nand_x1_sg U48829 ( .A(n53308), .B(n53347), .X(n16094) );
  inv_x1_sg U48830 ( .A(n16085), .X(n53357) );
  nand_x4_sg U48831 ( .A(n16082), .B(n53358), .X(n16075) );
  inv_x1_sg U48832 ( .A(n16083), .X(n53358) );
  nand_x1_sg U48833 ( .A(n16085), .B(n16084), .X(n16082) );
  nand_x1_sg U48834 ( .A(n53367), .B(n16178), .X(n16177) );
  inv_x1_sg U48835 ( .A(n16179), .X(n53367) );
  inv_x1_sg U48836 ( .A(n16180), .X(n53418) );
  inv_x1_sg U48837 ( .A(n16280), .X(n53457) );
  nand_x1_sg U48838 ( .A(n40569), .B(n16230), .X(n16227) );
  inv_x2_sg U48839 ( .A(n16218), .X(n44438) );
  nor_x1_sg U48840 ( .A(n53442), .B(n16224), .X(n16218) );
  nand_x4_sg U48841 ( .A(n16281), .B(n16282), .X(n15811) );
  nand_x1_sg U48842 ( .A(n42380), .B(n16230), .X(n16282) );
  inv_x1_sg U48843 ( .A(n16329), .X(n53404) );
  nand_x1_sg U48844 ( .A(n16331), .B(n16330), .X(n16328) );
  inv_x1_sg U48845 ( .A(n16384), .X(n53454) );
  nand_x2_sg U48846 ( .A(n27843), .B(n27844), .X(n27842) );
  inv_x1_sg U48847 ( .A(n27842), .X(n53481) );
  inv_x1_sg U48848 ( .A(n27832), .X(n43889) );
  nand_x1_sg U48849 ( .A(n46388), .B(n46391), .X(n16622) );
  nand_x1_sg U48850 ( .A(n53492), .B(n46391), .X(n16632) );
  nand_x1_sg U48851 ( .A(n16654), .B(n46384), .X(n16653) );
  inv_x2_sg U48852 ( .A(n16656), .X(n45594) );
  nand_x1_sg U48853 ( .A(n16671), .B(n16667), .X(n16672) );
  nand_x1_sg U48854 ( .A(n16711), .B(n16712), .X(n16710) );
  nand_x1_sg U48855 ( .A(n46384), .B(n16691), .X(n16712) );
  inv_x2_sg U48856 ( .A(n16703), .X(n43985) );
  nor_x1_sg U48857 ( .A(n53550), .B(n16715), .X(n16703) );
  nand_x1_sg U48858 ( .A(n46384), .B(n53539), .X(n16690) );
  nand_x1_sg U48859 ( .A(n16633), .B(n16691), .X(n16689) );
  inv_x1_sg U48860 ( .A(n16691), .X(n53539) );
  inv_x1_sg U48861 ( .A(n16682), .X(n53534) );
  inv_x1_sg U48862 ( .A(n16697), .X(n53532) );
  nand_x1_sg U48863 ( .A(n16699), .B(n16698), .X(n16696) );
  inv_x1_sg U48864 ( .A(n16675), .X(n53520) );
  inv_x2_sg U48865 ( .A(n16730), .X(n44278) );
  nor_x1_sg U48866 ( .A(n16739), .B(n16740), .X(n16730) );
  inv_x2_sg U48867 ( .A(n16701), .X(n45468) );
  nand_x1_sg U48868 ( .A(n43986), .B(n41936), .X(n16701) );
  nand_x1_sg U48869 ( .A(n45539), .B(n16820), .X(n16818) );
  nand_x4_sg U48870 ( .A(n16830), .B(n16831), .X(n16823) );
  nand_x1_sg U48871 ( .A(n53588), .B(n16832), .X(n16831) );
  nand_x1_sg U48872 ( .A(n53626), .B(n16833), .X(n16830) );
  nand_x4_sg U48873 ( .A(n16871), .B(n16872), .X(n16861) );
  nand_x1_sg U48874 ( .A(n16873), .B(n16874), .X(n16872) );
  nand_x4_sg U48875 ( .A(n16905), .B(n53634), .X(n16870) );
  inv_x1_sg U48876 ( .A(n16906), .X(n53634) );
  inv_x1_sg U48877 ( .A(n16868), .X(n53636) );
  nand_x1_sg U48878 ( .A(n16870), .B(n16869), .X(n16867) );
  inv_x1_sg U48879 ( .A(n16861), .X(n53647) );
  nand_x4_sg U48880 ( .A(n16878), .B(n16879), .X(n16869) );
  nand_x1_sg U48881 ( .A(n53588), .B(n53626), .X(n16879) );
  nand_x1_sg U48882 ( .A(n53652), .B(n16963), .X(n16962) );
  inv_x1_sg U48883 ( .A(n16964), .X(n53652) );
  inv_x1_sg U48884 ( .A(n16965), .X(n53699) );
  nand_x1_sg U48885 ( .A(n40556), .B(n16592), .X(n17063) );
  inv_x1_sg U48886 ( .A(n17010), .X(n53697) );
  inv_x2_sg U48887 ( .A(n17003), .X(n44182) );
  nor_x1_sg U48888 ( .A(n53721), .B(n17013), .X(n17003) );
  inv_x1_sg U48889 ( .A(n17114), .X(n53681) );
  nand_x1_sg U48890 ( .A(n17116), .B(n17115), .X(n17113) );
  nand_x4_sg U48891 ( .A(n17065), .B(n17066), .X(n16592) );
  nand_x1_sg U48892 ( .A(n44407), .B(n17011), .X(n17066) );
  nand_x1_sg U48893 ( .A(n53691), .B(n17092), .X(n17065) );
  inv_x1_sg U48894 ( .A(n17130), .X(n53746) );
  nand_x2_sg U48895 ( .A(n28124), .B(n28125), .X(n28123) );
  inv_x1_sg U48896 ( .A(n28123), .X(n53759) );
  inv_x1_sg U48897 ( .A(n28113), .X(n44015) );
  nand_x1_sg U48898 ( .A(n53765), .B(n46368), .X(n17407) );
  nand_x1_sg U48899 ( .A(n46363), .B(n46368), .X(n17416) );
  inv_x1_sg U48900 ( .A(n17438), .X(n53779) );
  inv_x2_sg U48901 ( .A(n17424), .X(n44208) );
  nor_x1_sg U48902 ( .A(n17433), .B(n17434), .X(n17424) );
  inv_x2_sg U48903 ( .A(n17443), .X(n44366) );
  nor_x1_sg U48904 ( .A(n17439), .B(n53774), .X(n17443) );
  nand_x1_sg U48905 ( .A(n46361), .B(n53817), .X(n17472) );
  nand_x1_sg U48906 ( .A(n46362), .B(n17473), .X(n17471) );
  inv_x1_sg U48907 ( .A(n17473), .X(n53817) );
  inv_x2_sg U48908 ( .A(n17461), .X(n44460) );
  nor_x1_sg U48909 ( .A(n53807), .B(n17468), .X(n17461) );
  nand_x1_sg U48910 ( .A(n17489), .B(n17490), .X(n17488) );
  nand_x1_sg U48911 ( .A(n46361), .B(n17473), .X(n17490) );
  inv_x2_sg U48912 ( .A(n17481), .X(n44384) );
  nor_x1_sg U48913 ( .A(n53829), .B(n17493), .X(n17481) );
  nand_x1_sg U48914 ( .A(n17546), .B(n53859), .X(n17545) );
  inv_x1_sg U48915 ( .A(n17547), .X(n53859) );
  inv_x2_sg U48916 ( .A(n17479), .X(n45466) );
  nand_x1_sg U48917 ( .A(n44385), .B(n41942), .X(n17479) );
  nand_x1_sg U48918 ( .A(n42144), .B(n17576), .X(n17574) );
  nand_x4_sg U48919 ( .A(n17606), .B(n17607), .X(n17599) );
  nand_x1_sg U48920 ( .A(n53866), .B(n17608), .X(n17607) );
  nand_x1_sg U48921 ( .A(n53910), .B(n17609), .X(n17606) );
  nand_x1_sg U48922 ( .A(n17696), .B(n17695), .X(n17693) );
  inv_x1_sg U48923 ( .A(n17695), .X(n53922) );
  inv_x2_sg U48924 ( .A(n17684), .X(n45398) );
  nor_x1_sg U48925 ( .A(n53940), .B(n17690), .X(n17684) );
  nand_x4_sg U48926 ( .A(n17645), .B(n17646), .X(n17636) );
  nand_x1_sg U48927 ( .A(n17647), .B(n53934), .X(n17646) );
  inv_x1_sg U48928 ( .A(n17648), .X(n53934) );
  nand_x4_sg U48929 ( .A(n17652), .B(n17653), .X(n17643) );
  nand_x1_sg U48930 ( .A(n53866), .B(n53910), .X(n17653) );
  inv_x1_sg U48931 ( .A(n17644), .X(n53920) );
  nand_x4_sg U48932 ( .A(n17641), .B(n53921), .X(n17635) );
  inv_x1_sg U48933 ( .A(n17642), .X(n53921) );
  nand_x1_sg U48934 ( .A(n17644), .B(n17643), .X(n17641) );
  nand_x1_sg U48935 ( .A(n53933), .B(n17735), .X(n17734) );
  inv_x1_sg U48936 ( .A(n17736), .X(n53933) );
  inv_x1_sg U48937 ( .A(n17737), .X(n53978) );
  nand_x1_sg U48938 ( .A(n40570), .B(n17783), .X(n17780) );
  inv_x2_sg U48939 ( .A(n17774), .X(n44452) );
  nor_x1_sg U48940 ( .A(n54002), .B(n17784), .X(n17774) );
  nand_x4_sg U48941 ( .A(n17886), .B(n53954), .X(n17371) );
  inv_x1_sg U48942 ( .A(n17887), .X(n53954) );
  nand_x1_sg U48943 ( .A(n17889), .B(n17888), .X(n17886) );
  nand_x4_sg U48944 ( .A(n17838), .B(n17839), .X(n17375) );
  nand_x1_sg U48945 ( .A(n42390), .B(n17783), .X(n17839) );
  inv_x1_sg U48946 ( .A(n17903), .X(n54030) );
  nand_x2_sg U48947 ( .A(n28403), .B(n28404), .X(n28402) );
  inv_x1_sg U48948 ( .A(n28402), .X(n54043) );
  nand_x1_sg U48949 ( .A(n28393), .B(n28394), .X(n28395) );
  nand_x1_sg U48950 ( .A(n46345), .B(n46348), .X(n18178) );
  inv_x1_sg U48951 ( .A(n18206), .X(n54065) );
  inv_x2_sg U48952 ( .A(n18191), .X(n45456) );
  nor_x1_sg U48953 ( .A(n18199), .B(n18200), .X(n18191) );
  inv_x1_sg U48954 ( .A(n18190), .X(n54072) );
  nand_x1_sg U48955 ( .A(n46338), .B(n18240), .X(n18237) );
  nand_x1_sg U48956 ( .A(n54090), .B(n18257), .X(n18256) );
  inv_x1_sg U48957 ( .A(n18259), .X(n54090) );
  inv_x2_sg U48958 ( .A(n18249), .X(n44476) );
  nor_x1_sg U48959 ( .A(n54116), .B(n18261), .X(n18249) );
  nand_x4_sg U48960 ( .A(n18286), .B(n18285), .X(n18279) );
  nand_x1_sg U48961 ( .A(n18316), .B(n54139), .X(n18315) );
  inv_x1_sg U48962 ( .A(n18317), .X(n54139) );
  nand_x1_sg U48963 ( .A(n18279), .B(n54132), .X(n18278) );
  nand_x1_sg U48964 ( .A(n42138), .B(n18346), .X(n18344) );
  nand_x4_sg U48965 ( .A(n18375), .B(n18376), .X(n18368) );
  nand_x1_sg U48966 ( .A(n54158), .B(n18377), .X(n18376) );
  nand_x1_sg U48967 ( .A(n54190), .B(n18378), .X(n18375) );
  nand_x4_sg U48968 ( .A(n18414), .B(n18415), .X(n18405) );
  nand_x1_sg U48969 ( .A(n18416), .B(n54214), .X(n18415) );
  inv_x1_sg U48970 ( .A(n18417), .X(n54214) );
  nand_x1_sg U48971 ( .A(n18465), .B(n18464), .X(n18462) );
  inv_x1_sg U48972 ( .A(n18464), .X(n54205) );
  inv_x2_sg U48973 ( .A(n18453), .X(n45396) );
  nor_x1_sg U48974 ( .A(n54222), .B(n18459), .X(n18453) );
  nand_x4_sg U48975 ( .A(n18447), .B(n54202), .X(n18413) );
  inv_x1_sg U48976 ( .A(n18448), .X(n54202) );
  inv_x1_sg U48977 ( .A(n18411), .X(n54204) );
  nand_x1_sg U48978 ( .A(n18413), .B(n18412), .X(n18410) );
  inv_x1_sg U48979 ( .A(n18405), .X(n54215) );
  nand_x4_sg U48980 ( .A(n18421), .B(n18422), .X(n18412) );
  nand_x1_sg U48981 ( .A(n54158), .B(n54190), .X(n18422) );
  nand_x1_sg U48982 ( .A(n54220), .B(n18504), .X(n18503) );
  inv_x1_sg U48983 ( .A(n18505), .X(n54220) );
  inv_x1_sg U48984 ( .A(n18506), .X(n54262) );
  inv_x1_sg U48985 ( .A(n18604), .X(n54299) );
  inv_x2_sg U48986 ( .A(n18601), .X(n45438) );
  nor_x1_sg U48987 ( .A(n18663), .B(n45441), .X(n18601) );
  nand_x1_sg U48988 ( .A(n40571), .B(n18551), .X(n18548) );
  inv_x2_sg U48989 ( .A(n18542), .X(n44180) );
  nor_x1_sg U48990 ( .A(n54284), .B(n18552), .X(n18542) );
  nand_x4_sg U48991 ( .A(n18605), .B(n18606), .X(n18146) );
  nand_x1_sg U48992 ( .A(n43300), .B(n18551), .X(n18606) );
  inv_x1_sg U48993 ( .A(n18672), .X(n54311) );
  nand_x2_sg U48994 ( .A(n28682), .B(n28683), .X(n28681) );
  inv_x1_sg U48995 ( .A(n28681), .X(n54324) );
  inv_x1_sg U48996 ( .A(n28671), .X(n44011) );
  nand_x1_sg U48997 ( .A(n54330), .B(n46321), .X(n18952) );
  nand_x1_sg U48998 ( .A(n46316), .B(n46321), .X(n18961) );
  inv_x1_sg U48999 ( .A(n18983), .X(n54344) );
  inv_x2_sg U49000 ( .A(n18969), .X(n44206) );
  nor_x1_sg U49001 ( .A(n18978), .B(n18979), .X(n18969) );
  inv_x2_sg U49002 ( .A(n18988), .X(n44364) );
  nor_x1_sg U49003 ( .A(n18984), .B(n54339), .X(n18988) );
  nand_x1_sg U49004 ( .A(n46314), .B(n54382), .X(n19017) );
  nand_x1_sg U49005 ( .A(n46315), .B(n19018), .X(n19016) );
  inv_x1_sg U49006 ( .A(n19018), .X(n54382) );
  inv_x2_sg U49007 ( .A(n19006), .X(n44458) );
  nor_x1_sg U49008 ( .A(n54372), .B(n19013), .X(n19006) );
  nand_x1_sg U49009 ( .A(n19034), .B(n19035), .X(n19033) );
  nand_x1_sg U49010 ( .A(n46314), .B(n19018), .X(n19035) );
  inv_x2_sg U49011 ( .A(n19026), .X(n44382) );
  nor_x1_sg U49012 ( .A(n54394), .B(n19038), .X(n19026) );
  nand_x1_sg U49013 ( .A(n19091), .B(n54424), .X(n19090) );
  inv_x1_sg U49014 ( .A(n19092), .X(n54424) );
  inv_x2_sg U49015 ( .A(n19024), .X(n45464) );
  nand_x1_sg U49016 ( .A(n44383), .B(n41941), .X(n19024) );
  nand_x1_sg U49017 ( .A(n42142), .B(n19121), .X(n19119) );
  nand_x4_sg U49018 ( .A(n19151), .B(n19152), .X(n19144) );
  nand_x1_sg U49019 ( .A(n54431), .B(n19153), .X(n19152) );
  nand_x1_sg U49020 ( .A(n54475), .B(n19154), .X(n19151) );
  nand_x1_sg U49021 ( .A(n19241), .B(n19240), .X(n19238) );
  inv_x1_sg U49022 ( .A(n19240), .X(n54487) );
  inv_x2_sg U49023 ( .A(n19229), .X(n45394) );
  nor_x1_sg U49024 ( .A(n54505), .B(n19235), .X(n19229) );
  nand_x4_sg U49025 ( .A(n19190), .B(n19191), .X(n19181) );
  nand_x1_sg U49026 ( .A(n19192), .B(n54499), .X(n19191) );
  inv_x1_sg U49027 ( .A(n19193), .X(n54499) );
  nand_x4_sg U49028 ( .A(n19197), .B(n19198), .X(n19188) );
  nand_x1_sg U49029 ( .A(n54431), .B(n54475), .X(n19198) );
  inv_x1_sg U49030 ( .A(n19189), .X(n54485) );
  nand_x4_sg U49031 ( .A(n19186), .B(n54486), .X(n19180) );
  inv_x1_sg U49032 ( .A(n19187), .X(n54486) );
  nand_x1_sg U49033 ( .A(n19189), .B(n19188), .X(n19186) );
  nand_x1_sg U49034 ( .A(n54498), .B(n19280), .X(n19279) );
  inv_x1_sg U49035 ( .A(n19281), .X(n54498) );
  inv_x1_sg U49036 ( .A(n19282), .X(n54543) );
  nand_x1_sg U49037 ( .A(n40572), .B(n19328), .X(n19325) );
  inv_x2_sg U49038 ( .A(n19319), .X(n44450) );
  nor_x1_sg U49039 ( .A(n54567), .B(n19329), .X(n19319) );
  nand_x4_sg U49040 ( .A(n19431), .B(n54519), .X(n18916) );
  inv_x1_sg U49041 ( .A(n19432), .X(n54519) );
  nand_x1_sg U49042 ( .A(n19434), .B(n19433), .X(n19431) );
  nand_x4_sg U49043 ( .A(n19383), .B(n19384), .X(n18920) );
  nand_x1_sg U49044 ( .A(n42388), .B(n19328), .X(n19384) );
  inv_x1_sg U49045 ( .A(n19448), .X(n54595) );
  nand_x2_sg U49046 ( .A(n28960), .B(n28961), .X(n28959) );
  inv_x1_sg U49047 ( .A(n28959), .X(n54608) );
  inv_x1_sg U49048 ( .A(n28949), .X(n43877) );
  nand_x1_sg U49049 ( .A(n54614), .B(n46301), .X(n19723) );
  inv_x1_sg U49050 ( .A(n19750), .X(n54627) );
  inv_x2_sg U49051 ( .A(n19738), .X(n44470) );
  nor_x1_sg U49052 ( .A(n19746), .B(n19747), .X(n19738) );
  nand_x1_sg U49053 ( .A(n19735), .B(n19785), .X(n19783) );
  nand_x1_sg U49054 ( .A(n19802), .B(n19803), .X(n19801) );
  nand_x1_sg U49055 ( .A(n46294), .B(n19804), .X(n19803) );
  inv_x2_sg U49056 ( .A(n19794), .X(n43983) );
  nor_x1_sg U49057 ( .A(n54679), .B(n19806), .X(n19794) );
  nand_x1_sg U49058 ( .A(n19861), .B(n54703), .X(n19860) );
  inv_x1_sg U49059 ( .A(n19862), .X(n54703) );
  inv_x2_sg U49060 ( .A(n19792), .X(n45462) );
  nand_x1_sg U49061 ( .A(n43984), .B(n54668), .X(n19792) );
  nand_x4_sg U49062 ( .A(n19920), .B(n19921), .X(n19913) );
  nand_x1_sg U49063 ( .A(n54723), .B(n19922), .X(n19921) );
  nand_x1_sg U49064 ( .A(n54757), .B(n19923), .X(n19920) );
  nand_x4_sg U49065 ( .A(n19959), .B(n19960), .X(n19950) );
  nand_x1_sg U49066 ( .A(n19961), .B(n54783), .X(n19960) );
  inv_x1_sg U49067 ( .A(n19962), .X(n54783) );
  nand_x1_sg U49068 ( .A(n20010), .B(n20009), .X(n20007) );
  inv_x1_sg U49069 ( .A(n20009), .X(n54773) );
  inv_x2_sg U49070 ( .A(n19998), .X(n45392) );
  nor_x1_sg U49071 ( .A(n54789), .B(n20004), .X(n19998) );
  nand_x4_sg U49072 ( .A(n19992), .B(n54770), .X(n19958) );
  inv_x1_sg U49073 ( .A(n19993), .X(n54770) );
  inv_x1_sg U49074 ( .A(n19956), .X(n54772) );
  nand_x1_sg U49075 ( .A(n19958), .B(n19957), .X(n19955) );
  inv_x1_sg U49076 ( .A(n19950), .X(n54784) );
  nand_x4_sg U49077 ( .A(n19966), .B(n19967), .X(n19957) );
  nand_x1_sg U49078 ( .A(n54723), .B(n54757), .X(n19967) );
  nand_x1_sg U49079 ( .A(n54782), .B(n20049), .X(n20048) );
  inv_x1_sg U49080 ( .A(n20050), .X(n54782) );
  inv_x1_sg U49081 ( .A(n20051), .X(n54829) );
  inv_x1_sg U49082 ( .A(n20150), .X(n54867) );
  inv_x2_sg U49083 ( .A(n20147), .X(n45430) );
  nor_x1_sg U49084 ( .A(n20208), .B(n45433), .X(n20147) );
  nand_x1_sg U49085 ( .A(n40573), .B(n20096), .X(n20093) );
  inv_x2_sg U49086 ( .A(n20087), .X(n44178) );
  nor_x1_sg U49087 ( .A(n54852), .B(n20097), .X(n20087) );
  nand_x4_sg U49088 ( .A(n20151), .B(n20152), .X(n19691) );
  nand_x1_sg U49089 ( .A(n43298), .B(n20096), .X(n20152) );
  inv_x1_sg U49090 ( .A(n20217), .X(n54879) );
  nand_x2_sg U49091 ( .A(n29243), .B(n29244), .X(n29242) );
  inv_x1_sg U49092 ( .A(n29242), .X(n54892) );
  inv_x1_sg U49093 ( .A(n29232), .X(n44007) );
  nand_x1_sg U49094 ( .A(n54898), .B(n46276), .X(n20496) );
  nand_x1_sg U49095 ( .A(n46271), .B(n46276), .X(n20505) );
  inv_x1_sg U49096 ( .A(n20527), .X(n54912) );
  inv_x2_sg U49097 ( .A(n20513), .X(n44204) );
  nor_x1_sg U49098 ( .A(n20522), .B(n20523), .X(n20513) );
  inv_x2_sg U49099 ( .A(n20532), .X(n44362) );
  nor_x1_sg U49100 ( .A(n20528), .B(n54907), .X(n20532) );
  nand_x1_sg U49101 ( .A(n46269), .B(n54950), .X(n20561) );
  nand_x1_sg U49102 ( .A(n46270), .B(n20562), .X(n20560) );
  inv_x1_sg U49103 ( .A(n20562), .X(n54950) );
  inv_x2_sg U49104 ( .A(n20550), .X(n44456) );
  nor_x1_sg U49105 ( .A(n54940), .B(n20557), .X(n20550) );
  nand_x1_sg U49106 ( .A(n20578), .B(n20579), .X(n20577) );
  nand_x1_sg U49107 ( .A(n46269), .B(n20562), .X(n20579) );
  inv_x2_sg U49108 ( .A(n20570), .X(n44380) );
  nor_x1_sg U49109 ( .A(n54962), .B(n20582), .X(n20570) );
  nand_x1_sg U49110 ( .A(n20635), .B(n54992), .X(n20634) );
  inv_x1_sg U49111 ( .A(n20636), .X(n54992) );
  inv_x2_sg U49112 ( .A(n20568), .X(n45460) );
  nand_x1_sg U49113 ( .A(n44381), .B(n41940), .X(n20568) );
  nand_x1_sg U49114 ( .A(n42140), .B(n20665), .X(n20663) );
  nand_x4_sg U49115 ( .A(n20695), .B(n20696), .X(n20688) );
  nand_x1_sg U49116 ( .A(n54999), .B(n20697), .X(n20696) );
  nand_x1_sg U49117 ( .A(n55043), .B(n20698), .X(n20695) );
  nand_x1_sg U49118 ( .A(n20785), .B(n20784), .X(n20782) );
  inv_x1_sg U49119 ( .A(n20784), .X(n55055) );
  inv_x2_sg U49120 ( .A(n20773), .X(n45390) );
  nor_x1_sg U49121 ( .A(n55073), .B(n20779), .X(n20773) );
  nand_x4_sg U49122 ( .A(n20734), .B(n20735), .X(n20725) );
  nand_x1_sg U49123 ( .A(n20736), .B(n55067), .X(n20735) );
  inv_x1_sg U49124 ( .A(n20737), .X(n55067) );
  nand_x4_sg U49125 ( .A(n20741), .B(n20742), .X(n20732) );
  nand_x1_sg U49126 ( .A(n54999), .B(n55043), .X(n20742) );
  inv_x1_sg U49127 ( .A(n20733), .X(n55053) );
  nand_x4_sg U49128 ( .A(n20730), .B(n55054), .X(n20724) );
  inv_x1_sg U49129 ( .A(n20731), .X(n55054) );
  nand_x1_sg U49130 ( .A(n20733), .B(n20732), .X(n20730) );
  nand_x1_sg U49131 ( .A(n55066), .B(n20824), .X(n20823) );
  inv_x1_sg U49132 ( .A(n20825), .X(n55066) );
  inv_x1_sg U49133 ( .A(n20826), .X(n55111) );
  nand_x1_sg U49134 ( .A(n40574), .B(n20872), .X(n20869) );
  inv_x2_sg U49135 ( .A(n20863), .X(n44448) );
  nor_x1_sg U49136 ( .A(n55135), .B(n20873), .X(n20863) );
  nand_x4_sg U49137 ( .A(n20975), .B(n55087), .X(n20460) );
  inv_x1_sg U49138 ( .A(n20976), .X(n55087) );
  nand_x1_sg U49139 ( .A(n20978), .B(n20977), .X(n20975) );
  nand_x4_sg U49140 ( .A(n20927), .B(n20928), .X(n20464) );
  nand_x1_sg U49141 ( .A(n42386), .B(n20872), .X(n20928) );
  inv_x1_sg U49142 ( .A(n20992), .X(n55163) );
  nand_x2_sg U49143 ( .A(n29521), .B(n29522), .X(n29520) );
  inv_x1_sg U49144 ( .A(n29520), .X(n55176) );
  inv_x1_sg U49145 ( .A(n29510), .X(n43881) );
  nand_x1_sg U49146 ( .A(n55182), .B(n46256), .X(n21268) );
  inv_x1_sg U49147 ( .A(n21295), .X(n55195) );
  inv_x2_sg U49148 ( .A(n21283), .X(n44468) );
  nor_x1_sg U49149 ( .A(n21291), .B(n21292), .X(n21283) );
  nand_x1_sg U49150 ( .A(n21280), .B(n21330), .X(n21328) );
  nand_x1_sg U49151 ( .A(n21347), .B(n21348), .X(n21346) );
  nand_x1_sg U49152 ( .A(n46249), .B(n21349), .X(n21348) );
  inv_x2_sg U49153 ( .A(n21339), .X(n43981) );
  nor_x1_sg U49154 ( .A(n55247), .B(n21351), .X(n21339) );
  nand_x1_sg U49155 ( .A(n21406), .B(n55271), .X(n21405) );
  inv_x1_sg U49156 ( .A(n21407), .X(n55271) );
  inv_x2_sg U49157 ( .A(n21337), .X(n45458) );
  nand_x1_sg U49158 ( .A(n43982), .B(n55236), .X(n21337) );
  nand_x4_sg U49159 ( .A(n21465), .B(n21466), .X(n21458) );
  nand_x1_sg U49160 ( .A(n55291), .B(n21467), .X(n21466) );
  nand_x1_sg U49161 ( .A(n55325), .B(n21468), .X(n21465) );
  nand_x4_sg U49162 ( .A(n21504), .B(n21505), .X(n21495) );
  nand_x1_sg U49163 ( .A(n21506), .B(n55351), .X(n21505) );
  inv_x1_sg U49164 ( .A(n21507), .X(n55351) );
  nand_x1_sg U49165 ( .A(n21555), .B(n21554), .X(n21552) );
  inv_x1_sg U49166 ( .A(n21554), .X(n55341) );
  inv_x2_sg U49167 ( .A(n21543), .X(n45388) );
  nor_x1_sg U49168 ( .A(n55357), .B(n21549), .X(n21543) );
  nand_x4_sg U49169 ( .A(n21537), .B(n55338), .X(n21503) );
  inv_x1_sg U49170 ( .A(n21538), .X(n55338) );
  inv_x1_sg U49171 ( .A(n21501), .X(n55340) );
  nand_x1_sg U49172 ( .A(n21503), .B(n21502), .X(n21500) );
  inv_x1_sg U49173 ( .A(n21495), .X(n55352) );
  nand_x4_sg U49174 ( .A(n21511), .B(n21512), .X(n21502) );
  nand_x1_sg U49175 ( .A(n55291), .B(n55325), .X(n21512) );
  nand_x1_sg U49176 ( .A(n55350), .B(n21594), .X(n21593) );
  inv_x1_sg U49177 ( .A(n21595), .X(n55350) );
  inv_x1_sg U49178 ( .A(n21596), .X(n55397) );
  inv_x1_sg U49179 ( .A(n21695), .X(n55435) );
  inv_x2_sg U49180 ( .A(n21692), .X(n45422) );
  nor_x1_sg U49181 ( .A(n21753), .B(n45425), .X(n21692) );
  nand_x1_sg U49182 ( .A(n40575), .B(n21641), .X(n21638) );
  inv_x2_sg U49183 ( .A(n21632), .X(n44176) );
  nor_x1_sg U49184 ( .A(n55420), .B(n21642), .X(n21632) );
  nand_x4_sg U49185 ( .A(n21696), .B(n21697), .X(n21236) );
  nand_x1_sg U49186 ( .A(n43296), .B(n21641), .X(n21697) );
  inv_x1_sg U49187 ( .A(n21762), .X(n55447) );
  inv_x1_sg U49188 ( .A(n29663), .X(n50089) );
  nand_x1_sg U49189 ( .A(n8183), .B(n29662), .X(n29661) );
  nand_x1_sg U49190 ( .A(n8243), .B(n30281), .X(n30280) );
  nand_x1_sg U49191 ( .A(n8323), .B(n30253), .X(n30252) );
  inv_x1_sg U49192 ( .A(n29649), .X(n50082) );
  nand_x1_sg U49193 ( .A(n8223), .B(n29648), .X(n29647) );
  inv_x1_sg U49194 ( .A(n30274), .X(n50078) );
  nand_x1_sg U49195 ( .A(n8263), .B(n30273), .X(n30272) );
  inv_x1_sg U49196 ( .A(n30260), .X(n50072) );
  nand_x1_sg U49197 ( .A(n8303), .B(n30259), .X(n30258) );
  nand_x1_sg U49198 ( .A(n30203), .B(n40741), .X(n30202) );
  nand_x1_sg U49199 ( .A(n8463), .B(n40806), .X(n30205) );
  nand_x1_sg U49200 ( .A(out_L1[19]), .B(n40807), .X(n30206) );
  inv_x1_sg U49201 ( .A(n30216), .X(n50055) );
  nand_x1_sg U49202 ( .A(n8423), .B(n30215), .X(n30214) );
  inv_x2_sg U49203 ( .A(n30183), .X(n45360) );
  nor_x1_sg U49204 ( .A(n30236), .B(n50064), .X(n30183) );
  nand_x1_sg U49205 ( .A(n8343), .B(n30245), .X(n30244) );
  inv_x1_sg U49206 ( .A(n30223), .X(n50059) );
  nand_x1_sg U49207 ( .A(n8403), .B(n30222), .X(n30221) );
  nor_x1_sg U49208 ( .A(n29628), .B(n30195), .X(n30194) );
  inv_x1_sg U49209 ( .A(n30231), .X(n50061) );
  nand_x1_sg U49210 ( .A(n8383), .B(n30230), .X(n30229) );
  inv_x1_sg U49211 ( .A(n24522), .X(n50042) );
  nand_x1_sg U49212 ( .A(n8184), .B(n24521), .X(n24520) );
  nand_x1_sg U49213 ( .A(n8244), .B(n29849), .X(n29848) );
  nand_x1_sg U49214 ( .A(n8324), .B(n30257), .X(n30517) );
  inv_x1_sg U49215 ( .A(n29851), .X(n50037) );
  nand_x1_sg U49216 ( .A(n8224), .B(n29653), .X(n29850) );
  inv_x1_sg U49217 ( .A(n30535), .X(n50049) );
  nand_x1_sg U49218 ( .A(n8264), .B(n30278), .X(n30534) );
  inv_x1_sg U49219 ( .A(n30523), .X(n50030) );
  nand_x1_sg U49220 ( .A(n8304), .B(n30264), .X(n30522) );
  inv_x2_sg U49221 ( .A(n30473), .X(n44732) );
  inv_x2_sg U49222 ( .A(n30513), .X(n44736) );
  inv_x2_sg U49223 ( .A(n30469), .X(n44622) );
  nor_x1_sg U49224 ( .A(n30479), .B(n50008), .X(n30469) );
  inv_x1_sg U49225 ( .A(n30500), .X(n50018) );
  nand_x1_sg U49226 ( .A(n8384), .B(n30235), .X(n30499) );
  inv_x1_sg U49227 ( .A(n24571), .X(n49993) );
  nand_x1_sg U49228 ( .A(n8185), .B(n24570), .X(n24569) );
  nand_x1_sg U49229 ( .A(n8245), .B(n30015), .X(n30014) );
  inv_x1_sg U49230 ( .A(n30439), .X(n50001) );
  nand_x1_sg U49231 ( .A(n8265), .B(n30438), .X(n30437) );
  inv_x1_sg U49232 ( .A(n30780), .X(n49985) );
  nand_x1_sg U49233 ( .A(n8305), .B(n30527), .X(n30779) );
  nand_x1_sg U49234 ( .A(n8325), .B(n30521), .X(n30774) );
  nand_x1_sg U49235 ( .A(n8346), .B(n30771), .X(n30770) );
  inv_x2_sg U49236 ( .A(n30711), .X(n45358) );
  nor_x1_sg U49237 ( .A(n30760), .B(n49977), .X(n30711) );
  inv_x1_sg U49238 ( .A(n30755), .X(n49974) );
  nand_x1_sg U49239 ( .A(n8385), .B(n30504), .X(n30754) );
  inv_x1_sg U49240 ( .A(n24620), .X(n49948) );
  nand_x1_sg U49241 ( .A(n8186), .B(n24619), .X(n24618) );
  nand_x1_sg U49242 ( .A(n8246), .B(n30162), .X(n30161) );
  inv_x2_sg U49243 ( .A(n30937), .X(n45330) );
  nor_x1_sg U49244 ( .A(n30986), .B(n49933), .X(n30937) );
  inv_x1_sg U49245 ( .A(n30433), .X(n49957) );
  nand_x1_sg U49246 ( .A(n8266), .B(n30432), .X(n30431) );
  inv_x1_sg U49247 ( .A(n31004), .X(n49961) );
  nand_x1_sg U49248 ( .A(n8306), .B(n30784), .X(n31003) );
  nand_x1_sg U49249 ( .A(n8326), .B(n30778), .X(n30998) );
  inv_x1_sg U49250 ( .A(n30002), .X(n49989) );
  inv_x2_sg U49251 ( .A(n30994), .X(n44292) );
  inv_x1_sg U49252 ( .A(n30953), .X(n49963) );
  inv_x1_sg U49253 ( .A(n30981), .X(n49930) );
  nand_x1_sg U49254 ( .A(n8386), .B(n30759), .X(n30980) );
  inv_x1_sg U49255 ( .A(n24669), .X(n49900) );
  nand_x1_sg U49256 ( .A(n8187), .B(n24668), .X(n24667) );
  nand_x1_sg U49257 ( .A(n8247), .B(n30156), .X(n30155) );
  inv_x1_sg U49258 ( .A(n30427), .X(n49909) );
  nand_x1_sg U49259 ( .A(n8267), .B(n30426), .X(n30425) );
  inv_x1_sg U49260 ( .A(n30926), .X(n49913) );
  nand_x1_sg U49261 ( .A(n8307), .B(n30925), .X(n30924) );
  nand_x1_sg U49262 ( .A(n8327), .B(n31002), .X(n31205) );
  inv_x1_sg U49263 ( .A(n29996), .X(n49944) );
  nand_x1_sg U49264 ( .A(n8348), .B(n31202), .X(n31201) );
  inv_x2_sg U49265 ( .A(n31142), .X(n45356) );
  nor_x1_sg U49266 ( .A(n31191), .B(n49887), .X(n31142) );
  inv_x1_sg U49267 ( .A(n31186), .X(n49884) );
  nand_x1_sg U49268 ( .A(n8387), .B(n30985), .X(n31185) );
  inv_x1_sg U49269 ( .A(n24717), .X(n49853) );
  nand_x1_sg U49270 ( .A(n8188), .B(n24716), .X(n24715) );
  nand_x1_sg U49271 ( .A(n8248), .B(n30150), .X(n30149) );
  inv_x2_sg U49272 ( .A(n31332), .X(n45328) );
  nor_x1_sg U49273 ( .A(n31381), .B(n49841), .X(n31332) );
  nand_x1_sg U49274 ( .A(n8328), .B(n31134), .X(n31133) );
  inv_x1_sg U49275 ( .A(n29990), .X(n49896) );
  inv_x1_sg U49276 ( .A(n30421), .X(n49862) );
  nand_x1_sg U49277 ( .A(n8268), .B(n30420), .X(n30419) );
  inv_x1_sg U49278 ( .A(n30916), .X(n49892) );
  inv_x2_sg U49279 ( .A(n31389), .X(n44290) );
  inv_x1_sg U49280 ( .A(n31348), .X(n49873) );
  inv_x1_sg U49281 ( .A(n31376), .X(n49838) );
  nand_x1_sg U49282 ( .A(n8388), .B(n31190), .X(n31375) );
  inv_x1_sg U49283 ( .A(n24765), .X(n49805) );
  nand_x1_sg U49284 ( .A(n8189), .B(n24764), .X(n24763) );
  nand_x1_sg U49285 ( .A(n8249), .B(n30144), .X(n30143) );
  nand_x1_sg U49286 ( .A(n8329), .B(n31128), .X(n31127) );
  inv_x1_sg U49287 ( .A(n29984), .X(n49849) );
  inv_x1_sg U49288 ( .A(n30415), .X(n49814) );
  nand_x1_sg U49289 ( .A(n8269), .B(n30414), .X(n30413) );
  inv_x1_sg U49290 ( .A(n30910), .X(n49845) );
  nand_x1_sg U49291 ( .A(n8350), .B(n31394), .X(n31393) );
  inv_x2_sg U49292 ( .A(n31503), .X(n45354) );
  nor_x1_sg U49293 ( .A(n31552), .B(n49824), .X(n31503) );
  inv_x1_sg U49294 ( .A(n31547), .X(n49793) );
  nand_x1_sg U49295 ( .A(n8389), .B(n31380), .X(n31546) );
  nand_x1_sg U49296 ( .A(n8330), .B(n31122), .X(n31121) );
  inv_x1_sg U49297 ( .A(n29978), .X(n49801) );
  inv_x1_sg U49298 ( .A(n30409), .X(n49767) );
  nand_x1_sg U49299 ( .A(n8270), .B(n30408), .X(n30407) );
  inv_x1_sg U49300 ( .A(n30904), .X(n49798) );
  inv_x1_sg U49301 ( .A(n24812), .X(n49758) );
  nand_x1_sg U49302 ( .A(n8190), .B(n24811), .X(n24810) );
  inv_x1_sg U49303 ( .A(n31672), .X(n49782) );
  inv_x1_sg U49304 ( .A(n31700), .X(n49780) );
  nand_x1_sg U49305 ( .A(n8390), .B(n31551), .X(n31699) );
  inv_x1_sg U49306 ( .A(n24860), .X(n49709) );
  nand_x1_sg U49307 ( .A(n8191), .B(n24859), .X(n24858) );
  nand_x1_sg U49308 ( .A(n8251), .B(n30132), .X(n30131) );
  nand_x1_sg U49309 ( .A(n8331), .B(n31116), .X(n31115) );
  inv_x1_sg U49310 ( .A(n29972), .X(n49754) );
  inv_x1_sg U49311 ( .A(n30403), .X(n49718) );
  nand_x1_sg U49312 ( .A(n8271), .B(n30402), .X(n30401) );
  inv_x1_sg U49313 ( .A(n30898), .X(n49750) );
  inv_x2_sg U49314 ( .A(n31491), .X(n45352) );
  nor_x1_sg U49315 ( .A(n31493), .B(n49728), .X(n31491) );
  inv_x1_sg U49316 ( .A(n31657), .X(n49730) );
  nand_x1_sg U49317 ( .A(n8391), .B(n31656), .X(n31655) );
  inv_x1_sg U49318 ( .A(n24908), .X(n49662) );
  nand_x1_sg U49319 ( .A(n8192), .B(n24907), .X(n24906) );
  nand_x1_sg U49320 ( .A(n8252), .B(n30126), .X(n30125) );
  nand_x1_sg U49321 ( .A(n8332), .B(n31110), .X(n31109) );
  inv_x1_sg U49322 ( .A(n29966), .X(n49705) );
  inv_x1_sg U49323 ( .A(n30397), .X(n49671) );
  nand_x1_sg U49324 ( .A(n8272), .B(n30396), .X(n30395) );
  inv_x1_sg U49325 ( .A(n30892), .X(n49701) );
  inv_x2_sg U49326 ( .A(n31485), .X(n45350) );
  nor_x1_sg U49327 ( .A(n31487), .B(n49682), .X(n31485) );
  inv_x1_sg U49328 ( .A(n31932), .X(n49690) );
  inv_x1_sg U49329 ( .A(n31651), .X(n49684) );
  nand_x1_sg U49330 ( .A(n8392), .B(n31650), .X(n31649) );
  inv_x1_sg U49331 ( .A(n24956), .X(n49615) );
  nand_x1_sg U49332 ( .A(n8193), .B(n24955), .X(n24954) );
  nand_x1_sg U49333 ( .A(n8253), .B(n30120), .X(n30119) );
  nand_x1_sg U49334 ( .A(n8333), .B(n31104), .X(n31103) );
  inv_x1_sg U49335 ( .A(n29960), .X(n49658) );
  inv_x1_sg U49336 ( .A(n30391), .X(n49624) );
  nand_x1_sg U49337 ( .A(n8273), .B(n30390), .X(n30389) );
  inv_x1_sg U49338 ( .A(n30886), .X(n49654) );
  inv_x2_sg U49339 ( .A(n31479), .X(n45348) );
  nor_x1_sg U49340 ( .A(n31481), .B(n49634), .X(n31479) );
  inv_x1_sg U49341 ( .A(n31919), .X(n49648) );
  inv_x2_sg U49342 ( .A(n31793), .X(n44516) );
  nor_x1_sg U49343 ( .A(n31795), .B(n49638), .X(n31793) );
  inv_x1_sg U49344 ( .A(n31645), .X(n49636) );
  nand_x1_sg U49345 ( .A(n8393), .B(n31644), .X(n31643) );
  inv_x1_sg U49346 ( .A(n25004), .X(n49569) );
  nand_x1_sg U49347 ( .A(n8194), .B(n25003), .X(n25002) );
  nand_x1_sg U49348 ( .A(n8254), .B(n30114), .X(n30113) );
  nand_x1_sg U49349 ( .A(n8334), .B(n31098), .X(n31097) );
  inv_x1_sg U49350 ( .A(n29954), .X(n49611) );
  inv_x1_sg U49351 ( .A(n30385), .X(n49578) );
  nand_x1_sg U49352 ( .A(n8274), .B(n30384), .X(n30383) );
  inv_x1_sg U49353 ( .A(n30880), .X(n49607) );
  inv_x2_sg U49354 ( .A(n31473), .X(n45346) );
  nor_x1_sg U49355 ( .A(n31475), .B(n49588), .X(n31473) );
  inv_x1_sg U49356 ( .A(n31913), .X(n49601) );
  inv_x2_sg U49357 ( .A(n31786), .X(n44514) );
  nor_x1_sg U49358 ( .A(n31788), .B(n49592), .X(n31786) );
  inv_x1_sg U49359 ( .A(n31639), .X(n49590) );
  nand_x1_sg U49360 ( .A(n8394), .B(n31638), .X(n31637) );
  inv_x1_sg U49361 ( .A(n25052), .X(n49522) );
  nand_x1_sg U49362 ( .A(n8195), .B(n25051), .X(n25050) );
  nand_x1_sg U49363 ( .A(n8255), .B(n30108), .X(n30107) );
  nand_x1_sg U49364 ( .A(n8335), .B(n31092), .X(n31091) );
  inv_x1_sg U49365 ( .A(n29948), .X(n49565) );
  inv_x1_sg U49366 ( .A(n30379), .X(n49531) );
  nand_x1_sg U49367 ( .A(n8275), .B(n30378), .X(n30377) );
  inv_x1_sg U49368 ( .A(n30874), .X(n49561) );
  inv_x2_sg U49369 ( .A(n31467), .X(n45344) );
  nor_x1_sg U49370 ( .A(n31469), .B(n49542), .X(n31467) );
  inv_x1_sg U49371 ( .A(n31907), .X(n49555) );
  inv_x2_sg U49372 ( .A(n31779), .X(n44512) );
  nor_x1_sg U49373 ( .A(n31781), .B(n49546), .X(n31779) );
  nand_x1_sg U49374 ( .A(n49553), .B(n49505), .X(n32104) );
  inv_x1_sg U49375 ( .A(n32106), .X(n49553) );
  inv_x2_sg U49376 ( .A(n32017), .X(n45490) );
  nor_x1_sg U49377 ( .A(n32019), .B(n49551), .X(n32017) );
  inv_x1_sg U49378 ( .A(n31633), .X(n49544) );
  nand_x1_sg U49379 ( .A(n8395), .B(n31632), .X(n31631) );
  inv_x1_sg U49380 ( .A(n30868), .X(n49514) );
  inv_x2_sg U49381 ( .A(n30625), .X(n44636) );
  nor_x1_sg U49382 ( .A(n30627), .B(n49486), .X(n30625) );
  inv_x1_sg U49383 ( .A(n30373), .X(n49484) );
  nand_x1_sg U49384 ( .A(n8276), .B(n30372), .X(n30371) );
  nand_x1_sg U49385 ( .A(n8476), .B(n40808), .X(n32102) );
  inv_x1_sg U49386 ( .A(n25101), .X(n49475) );
  nand_x1_sg U49387 ( .A(n8196), .B(n25100), .X(n25099) );
  nand_x1_sg U49388 ( .A(n8336), .B(n31086), .X(n31085) );
  inv_x1_sg U49389 ( .A(n29942), .X(n49518) );
  inv_x2_sg U49390 ( .A(n31461), .X(n45342) );
  nor_x1_sg U49391 ( .A(n31463), .B(n49494), .X(n31461) );
  inv_x1_sg U49392 ( .A(n31901), .X(n49508) );
  inv_x2_sg U49393 ( .A(n31772), .X(n44510) );
  nor_x1_sg U49394 ( .A(n31774), .B(n49498), .X(n31772) );
  nand_x1_sg U49395 ( .A(n8456), .B(n32014), .X(n32013) );
  inv_x1_sg U49396 ( .A(n31627), .X(n49496) );
  nand_x1_sg U49397 ( .A(n8396), .B(n31626), .X(n31625) );
  inv_x1_sg U49398 ( .A(n25149), .X(n49429) );
  nand_x1_sg U49399 ( .A(n8197), .B(n25148), .X(n25147) );
  nand_x1_sg U49400 ( .A(n8257), .B(n30096), .X(n30095) );
  nand_x1_sg U49401 ( .A(n8337), .B(n31080), .X(n31079) );
  inv_x1_sg U49402 ( .A(n29936), .X(n49471) );
  inv_x1_sg U49403 ( .A(n30367), .X(n49438) );
  nand_x1_sg U49404 ( .A(n8277), .B(n30366), .X(n30365) );
  inv_x1_sg U49405 ( .A(n30862), .X(n49467) );
  inv_x2_sg U49406 ( .A(n31455), .X(n45340) );
  nor_x1_sg U49407 ( .A(n31457), .B(n49448), .X(n31455) );
  inv_x1_sg U49408 ( .A(n31895), .X(n49461) );
  inv_x2_sg U49409 ( .A(n31765), .X(n44508) );
  nor_x1_sg U49410 ( .A(n31767), .B(n49452), .X(n31765) );
  inv_x1_sg U49411 ( .A(n32095), .X(n49459) );
  inv_x2_sg U49412 ( .A(n32004), .X(n45488) );
  nor_x1_sg U49413 ( .A(n32006), .B(n49457), .X(n32004) );
  inv_x1_sg U49414 ( .A(n31621), .X(n49450) );
  nand_x1_sg U49415 ( .A(n8397), .B(n31620), .X(n31619) );
  inv_x1_sg U49416 ( .A(n30856), .X(n49421) );
  inv_x2_sg U49417 ( .A(n30611), .X(n44634) );
  nor_x1_sg U49418 ( .A(n30613), .B(n49394), .X(n30611) );
  inv_x1_sg U49419 ( .A(n30361), .X(n49392) );
  nand_x1_sg U49420 ( .A(n8278), .B(n30360), .X(n30359) );
  inv_x1_sg U49421 ( .A(n25198), .X(n49383) );
  nand_x1_sg U49422 ( .A(n8198), .B(n25197), .X(n25196) );
  nand_x1_sg U49423 ( .A(n8338), .B(n31074), .X(n31073) );
  inv_x1_sg U49424 ( .A(n29930), .X(n49425) );
  inv_x1_sg U49425 ( .A(n31422), .X(n49400) );
  nand_x1_sg U49426 ( .A(n8359), .B(n31421), .X(n31420) );
  inv_x2_sg U49427 ( .A(n31449), .X(n45338) );
  nor_x1_sg U49428 ( .A(n31451), .B(n49403), .X(n31449) );
  nand_x1_sg U49429 ( .A(n8458), .B(n32001), .X(n32000) );
  inv_x1_sg U49430 ( .A(n31889), .X(n49415) );
  inv_x2_sg U49431 ( .A(n31758), .X(n44506) );
  nor_x1_sg U49432 ( .A(n31760), .B(n49407), .X(n31758) );
  inv_x1_sg U49433 ( .A(n31615), .X(n49405) );
  nand_x1_sg U49434 ( .A(n8398), .B(n31614), .X(n31613) );
  inv_x1_sg U49435 ( .A(n30850), .X(n49375) );
  inv_x2_sg U49436 ( .A(n30604), .X(n44648) );
  nor_x1_sg U49437 ( .A(n30606), .B(n49350), .X(n30604) );
  inv_x1_sg U49438 ( .A(n30355), .X(n49348) );
  nand_x1_sg U49439 ( .A(n8279), .B(n30354), .X(n30353) );
  inv_x1_sg U49440 ( .A(n25247), .X(n49339) );
  nand_x1_sg U49441 ( .A(n8199), .B(n25246), .X(n25245) );
  nand_x1_sg U49442 ( .A(n8339), .B(n31068), .X(n31067) );
  inv_x1_sg U49443 ( .A(n29924), .X(n49379) );
  inv_x2_sg U49444 ( .A(n31443), .X(n45336) );
  nor_x1_sg U49445 ( .A(n31445), .B(n49358), .X(n31443) );
  nand_x1_sg U49446 ( .A(n8459), .B(n31995), .X(n31994) );
  inv_x1_sg U49447 ( .A(n31883), .X(n49369) );
  inv_x2_sg U49448 ( .A(n31751), .X(n44504) );
  nor_x1_sg U49449 ( .A(n31753), .B(n49362), .X(n31751) );
  inv_x1_sg U49450 ( .A(n31609), .X(n49360) );
  nand_x1_sg U49451 ( .A(n8399), .B(n31608), .X(n31607) );
  inv_x1_sg U49452 ( .A(n30844), .X(n49331) );
  inv_x2_sg U49453 ( .A(n30597), .X(n44067) );
  nor_x1_sg U49454 ( .A(n30599), .B(n49304), .X(n30597) );
  inv_x1_sg U49455 ( .A(n30349), .X(n49302) );
  nand_x1_sg U49456 ( .A(n8280), .B(n30348), .X(n30347) );
  inv_x1_sg U49457 ( .A(n25294), .X(n49296) );
  nand_x1_sg U49458 ( .A(n8200), .B(n25293), .X(n25292) );
  nand_x1_sg U49459 ( .A(n8340), .B(n31062), .X(n31061) );
  inv_x1_sg U49460 ( .A(n29918), .X(n49335) );
  nand_x1_sg U49461 ( .A(n8380), .B(n31441), .X(n31440) );
  inv_x1_sg U49462 ( .A(n31877), .X(n49325) );
  inv_x2_sg U49463 ( .A(n31744), .X(n44620) );
  nor_x1_sg U49464 ( .A(n31746), .B(n49314), .X(n31744) );
  nand_x1_sg U49465 ( .A(n32076), .B(n32077), .X(n32074) );
  inv_x1_sg U49466 ( .A(n32076), .X(n49323) );
  inv_x2_sg U49467 ( .A(n31985), .X(n44244) );
  nor_x1_sg U49468 ( .A(n31987), .B(n49318), .X(n31985) );
  inv_x1_sg U49469 ( .A(n31603), .X(n49312) );
  nand_x1_sg U49470 ( .A(n8400), .B(n31602), .X(n31601) );
  nand_x1_sg U49471 ( .A(n30838), .B(n49273), .X(n30837) );
  inv_x1_sg U49472 ( .A(n30839), .X(n49273) );
  nand_x2_sg U49473 ( .A(n30341), .B(n30342), .X(n30340) );
  nand_x1_sg U49474 ( .A(n30590), .B(n49272), .X(n30589) );
  inv_x1_sg U49475 ( .A(n30591), .X(n49272) );
  inv_x1_sg U49476 ( .A(n32071), .X(n49281) );
  nand_x1_sg U49477 ( .A(n31871), .B(n49279), .X(n31870) );
  inv_x1_sg U49478 ( .A(n31872), .X(n49279) );
  nand_x1_sg U49479 ( .A(n25321), .B(n49270), .X(n30068) );
  nand_x1_sg U49480 ( .A(n30069), .B(n49292), .X(n30067) );
  inv_x1_sg U49481 ( .A(n30069), .X(n49270) );
  nand_x2_sg U49482 ( .A(n25336), .B(n25337), .X(n25335) );
  nand_x1_sg U49483 ( .A(n29721), .B(n49268), .X(n29720) );
  inv_x1_sg U49484 ( .A(n29722), .X(n49268) );
  inv_x1_sg U49485 ( .A(n25335), .X(n49267) );
  nand_x1_sg U49486 ( .A(n25308), .B(n49274), .X(n31052) );
  nand_x1_sg U49487 ( .A(n31053), .B(n49288), .X(n31051) );
  inv_x1_sg U49488 ( .A(n31053), .X(n49274) );
  nand_x1_sg U49489 ( .A(n29912), .B(n49269), .X(n29911) );
  inv_x1_sg U49490 ( .A(n29913), .X(n49269) );
  nand_x2_sg U49491 ( .A(n31433), .B(n31434), .X(n31432) );
  nand_x1_sg U49492 ( .A(n31978), .B(n49280), .X(n31977) );
  inv_x1_sg U49493 ( .A(n31979), .X(n49280) );
  nand_x2_sg U49494 ( .A(n31595), .B(n31596), .X(n31594) );
  nand_x1_sg U49495 ( .A(n31737), .B(n49278), .X(n31736) );
  inv_x1_sg U49496 ( .A(n31738), .X(n49278) );
  nand_x1_sg U49497 ( .A(n51279), .B(n25582), .X(n25579) );
  inv_x1_sg U49498 ( .A(n25570), .X(n51305) );
  nand_x1_sg U49499 ( .A(n51303), .B(n51318), .X(n25562) );
  nand_x1_sg U49500 ( .A(n25563), .B(n25564), .X(n25561) );
  nand_x4_sg U49501 ( .A(n25566), .B(n25642), .X(n25557) );
  nand_x1_sg U49502 ( .A(n25565), .B(n25564), .X(n25642) );
  nand_x2_sg U49503 ( .A(n45121), .B(n51375), .X(n25549) );
  nand_x2_sg U49504 ( .A(n45123), .B(n51351), .X(n25553) );
  inv_x1_sg U49505 ( .A(n25540), .X(n51395) );
  nand_x1_sg U49506 ( .A(n25542), .B(n25541), .X(n25539) );
  nand_x2_sg U49507 ( .A(n45183), .B(n51416), .X(n25537) );
  nand_x2_sg U49508 ( .A(n45119), .B(n51394), .X(n25543) );
  nand_x4_sg U49509 ( .A(n25550), .B(n25639), .X(n25541) );
  nand_x1_sg U49510 ( .A(n25547), .B(n25549), .X(n25639) );
  nand_x2_sg U49511 ( .A(n45117), .B(n51433), .X(n25531) );
  nand_x4_sg U49512 ( .A(n25538), .B(n25637), .X(n25529) );
  nand_x1_sg U49513 ( .A(n25535), .B(n25537), .X(n25637) );
  nand_x2_sg U49514 ( .A(n45115), .B(n51456), .X(n25525) );
  nor_x1_sg U49515 ( .A(n51559), .B(n25860), .X(n11199) );
  nand_x1_sg U49516 ( .A(n51585), .B(n51597), .X(n25843) );
  nand_x1_sg U49517 ( .A(n25844), .B(n25845), .X(n25842) );
  nand_x2_sg U49518 ( .A(n45159), .B(n51613), .X(n25840) );
  nand_x2_sg U49519 ( .A(n45113), .B(n51596), .X(n25846) );
  nand_x1_sg U49520 ( .A(n25850), .B(n50992), .X(n25922) );
  nand_x1_sg U49521 ( .A(n46029), .B(n51573), .X(n25923) );
  inv_x1_sg U49522 ( .A(n25924), .X(n51573) );
  nand_x2_sg U49523 ( .A(n45109), .B(n51648), .X(n25828) );
  nand_x2_sg U49524 ( .A(n45111), .B(n51628), .X(n25834) );
  nand_x4_sg U49525 ( .A(n25841), .B(n25920), .X(n25832) );
  nand_x1_sg U49526 ( .A(n25838), .B(n25840), .X(n25920) );
  nand_x4_sg U49527 ( .A(n25829), .B(n25918), .X(n25820) );
  nand_x1_sg U49528 ( .A(n25826), .B(n25828), .X(n25918) );
  nand_x2_sg U49529 ( .A(n45147), .B(n51691), .X(n25816) );
  nand_x4_sg U49530 ( .A(n25823), .B(n25917), .X(n25814) );
  nand_x1_sg U49531 ( .A(n25820), .B(n25822), .X(n25917) );
  nand_x2_sg U49532 ( .A(n45105), .B(n51715), .X(n25810) );
  nand_x2_sg U49533 ( .A(n45103), .B(n51736), .X(n25804) );
  nand_x1_sg U49534 ( .A(n25903), .B(n25902), .X(n25904) );
  nand_x1_sg U49535 ( .A(n51838), .B(n26143), .X(n26140) );
  inv_x1_sg U49536 ( .A(n26131), .X(n51866) );
  nand_x1_sg U49537 ( .A(n51864), .B(n51878), .X(n26123) );
  nand_x1_sg U49538 ( .A(n26124), .B(n26125), .X(n26122) );
  nand_x2_sg U49539 ( .A(n45173), .B(n51894), .X(n26120) );
  nand_x2_sg U49540 ( .A(n45097), .B(n51877), .X(n26126) );
  inv_x1_sg U49541 ( .A(n26204), .X(n51863) );
  nand_x2_sg U49542 ( .A(n45093), .B(n51929), .X(n26108) );
  nand_x2_sg U49543 ( .A(n45095), .B(n51909), .X(n26114) );
  nand_x4_sg U49544 ( .A(n26121), .B(n26200), .X(n26112) );
  nand_x1_sg U49545 ( .A(n26118), .B(n26120), .X(n26200) );
  nand_x4_sg U49546 ( .A(n26109), .B(n26198), .X(n26100) );
  nand_x1_sg U49547 ( .A(n26106), .B(n26108), .X(n26198) );
  nand_x2_sg U49548 ( .A(n45089), .B(n51993), .X(n26090) );
  nand_x2_sg U49549 ( .A(n45153), .B(n51972), .X(n26096) );
  nand_x4_sg U49550 ( .A(n26103), .B(n26197), .X(n26094) );
  nand_x1_sg U49551 ( .A(n26100), .B(n26102), .X(n26197) );
  nand_x2_sg U49552 ( .A(n45087), .B(n52015), .X(n26084) );
  nand_x4_sg U49553 ( .A(n26091), .B(n26195), .X(n26082) );
  nand_x1_sg U49554 ( .A(n26088), .B(n26090), .X(n26195) );
  nand_x1_sg U49555 ( .A(n26183), .B(n26182), .X(n26184) );
  nor_x1_sg U49556 ( .A(n52116), .B(n26419), .X(n12760) );
  nand_x1_sg U49557 ( .A(n52143), .B(n52155), .X(n26402) );
  nand_x1_sg U49558 ( .A(n26403), .B(n26404), .X(n26401) );
  nand_x2_sg U49559 ( .A(n45169), .B(n52171), .X(n26399) );
  nand_x2_sg U49560 ( .A(n45081), .B(n52154), .X(n26405) );
  nand_x1_sg U49561 ( .A(n45217), .B(n52130), .X(n26482) );
  nand_x1_sg U49562 ( .A(n26409), .B(n51030), .X(n26481) );
  inv_x1_sg U49563 ( .A(n26483), .X(n52130) );
  nand_x2_sg U49564 ( .A(n45143), .B(n52204), .X(n26387) );
  nand_x2_sg U49565 ( .A(n45079), .B(n52185), .X(n26393) );
  nand_x4_sg U49566 ( .A(n26400), .B(n26479), .X(n26391) );
  nand_x1_sg U49567 ( .A(n26397), .B(n26399), .X(n26479) );
  nand_x2_sg U49568 ( .A(n45179), .B(n52247), .X(n26375) );
  nand_x2_sg U49569 ( .A(n45077), .B(n52225), .X(n26381) );
  nand_x4_sg U49570 ( .A(n26388), .B(n26477), .X(n26379) );
  nand_x1_sg U49571 ( .A(n26385), .B(n26387), .X(n26477) );
  nand_x4_sg U49572 ( .A(n26376), .B(n26475), .X(n26367) );
  nand_x1_sg U49573 ( .A(n26373), .B(n26375), .X(n26475) );
  nand_x2_sg U49574 ( .A(n45073), .B(n52291), .X(n26363) );
  nand_x4_sg U49575 ( .A(n26370), .B(n26474), .X(n26361) );
  nand_x1_sg U49576 ( .A(n26367), .B(n26369), .X(n26474) );
  nand_x1_sg U49577 ( .A(n26462), .B(n26461), .X(n26463) );
  nand_x1_sg U49578 ( .A(n52390), .B(n26700), .X(n26697) );
  inv_x1_sg U49579 ( .A(n26688), .X(n52418) );
  nand_x1_sg U49580 ( .A(n52416), .B(n52429), .X(n26680) );
  nand_x1_sg U49581 ( .A(n26681), .B(n26682), .X(n26679) );
  nand_x4_sg U49582 ( .A(n26684), .B(n26758), .X(n26675) );
  nand_x1_sg U49583 ( .A(n26683), .B(n26682), .X(n26758) );
  nand_x2_sg U49584 ( .A(n45137), .B(n52481), .X(n26665) );
  nand_x2_sg U49585 ( .A(n45065), .B(n52461), .X(n26671) );
  nand_x4_sg U49586 ( .A(n26678), .B(n26757), .X(n26669) );
  nand_x1_sg U49587 ( .A(n26675), .B(n26677), .X(n26757) );
  nand_x2_sg U49588 ( .A(n45163), .B(n52523), .X(n26653) );
  nand_x2_sg U49589 ( .A(n45063), .B(n52502), .X(n26659) );
  nand_x4_sg U49590 ( .A(n26666), .B(n26755), .X(n26657) );
  nand_x1_sg U49591 ( .A(n26663), .B(n26665), .X(n26755) );
  nand_x4_sg U49592 ( .A(n26654), .B(n26753), .X(n26645) );
  nand_x1_sg U49593 ( .A(n26651), .B(n26653), .X(n26753) );
  nand_x2_sg U49594 ( .A(n45059), .B(n52566), .X(n26641) );
  nand_x4_sg U49595 ( .A(n26648), .B(n26752), .X(n26639) );
  nand_x1_sg U49596 ( .A(n26645), .B(n26647), .X(n26752) );
  nand_x1_sg U49597 ( .A(n26740), .B(n26739), .X(n26741) );
  nand_x1_sg U49598 ( .A(n52669), .B(n26979), .X(n26976) );
  inv_x1_sg U49599 ( .A(n26967), .X(n52694) );
  nand_x2_sg U49600 ( .A(n26962), .B(n26963), .X(n26960) );
  inv_x1_sg U49601 ( .A(n26961), .X(n52692) );
  nand_x2_sg U49602 ( .A(n45199), .B(n52722), .X(n26956) );
  nand_x2_sg U49603 ( .A(n45053), .B(n52705), .X(n26962) );
  nand_x1_sg U49604 ( .A(n44320), .B(n51069), .X(n27038) );
  nand_x2_sg U49605 ( .A(n45049), .B(n52761), .X(n26944) );
  nand_x2_sg U49606 ( .A(n45051), .B(n52740), .X(n26950) );
  nand_x4_sg U49607 ( .A(n26957), .B(n27036), .X(n26948) );
  nand_x1_sg U49608 ( .A(n26954), .B(n26956), .X(n27036) );
  nand_x2_sg U49609 ( .A(n45047), .B(n52804), .X(n26932) );
  nand_x2_sg U49610 ( .A(n45185), .B(n52781), .X(n26938) );
  nand_x4_sg U49611 ( .A(n26945), .B(n27034), .X(n26936) );
  nand_x1_sg U49612 ( .A(n26942), .B(n26944), .X(n27034) );
  nand_x2_sg U49613 ( .A(n45129), .B(n52822), .X(n26926) );
  nand_x4_sg U49614 ( .A(n26933), .B(n27032), .X(n26924) );
  nand_x1_sg U49615 ( .A(n26930), .B(n26932), .X(n27032) );
  nand_x2_sg U49616 ( .A(n45045), .B(n52846), .X(n26920) );
  nand_x1_sg U49617 ( .A(n27019), .B(n27018), .X(n27020) );
  nor_x1_sg U49618 ( .A(n52950), .B(n27256), .X(n15093) );
  nand_x1_sg U49619 ( .A(n52977), .B(n52989), .X(n27239) );
  nand_x1_sg U49620 ( .A(n27240), .B(n27241), .X(n27238) );
  nand_x2_sg U49621 ( .A(n45167), .B(n53005), .X(n27236) );
  nand_x2_sg U49622 ( .A(n45039), .B(n52988), .X(n27242) );
  nand_x1_sg U49623 ( .A(n45215), .B(n52964), .X(n27319) );
  nand_x1_sg U49624 ( .A(n27246), .B(n51088), .X(n27318) );
  inv_x1_sg U49625 ( .A(n27320), .X(n52964) );
  nand_x2_sg U49626 ( .A(n45141), .B(n53038), .X(n27224) );
  nand_x2_sg U49627 ( .A(n45037), .B(n53019), .X(n27230) );
  nand_x4_sg U49628 ( .A(n27237), .B(n27316), .X(n27228) );
  nand_x1_sg U49629 ( .A(n27234), .B(n27236), .X(n27316) );
  nand_x2_sg U49630 ( .A(n45177), .B(n53081), .X(n27212) );
  nand_x2_sg U49631 ( .A(n45035), .B(n53059), .X(n27218) );
  nand_x4_sg U49632 ( .A(n27225), .B(n27314), .X(n27216) );
  nand_x1_sg U49633 ( .A(n27222), .B(n27224), .X(n27314) );
  nand_x4_sg U49634 ( .A(n27213), .B(n27312), .X(n27204) );
  nand_x1_sg U49635 ( .A(n27210), .B(n27212), .X(n27312) );
  nand_x2_sg U49636 ( .A(n45031), .B(n53125), .X(n27200) );
  nand_x4_sg U49637 ( .A(n27207), .B(n27311), .X(n27198) );
  nand_x1_sg U49638 ( .A(n27204), .B(n27206), .X(n27311) );
  nand_x1_sg U49639 ( .A(n27299), .B(n27298), .X(n27300) );
  nand_x1_sg U49640 ( .A(n53226), .B(n27538), .X(n27535) );
  inv_x1_sg U49641 ( .A(n27526), .X(n53252) );
  nand_x1_sg U49642 ( .A(n53250), .B(n53265), .X(n27518) );
  nand_x1_sg U49643 ( .A(n27519), .B(n27520), .X(n27517) );
  nand_x4_sg U49644 ( .A(n27522), .B(n27596), .X(n27513) );
  nand_x1_sg U49645 ( .A(n27521), .B(n27520), .X(n27596) );
  nand_x2_sg U49646 ( .A(n45021), .B(n53317), .X(n27503) );
  nand_x2_sg U49647 ( .A(n45023), .B(n53296), .X(n27509) );
  nand_x4_sg U49648 ( .A(n27516), .B(n27595), .X(n27507) );
  nand_x1_sg U49649 ( .A(n27513), .B(n27515), .X(n27595) );
  nand_x4_sg U49650 ( .A(n27504), .B(n27593), .X(n27495) );
  nand_x1_sg U49651 ( .A(n27501), .B(n27503), .X(n27593) );
  nand_x2_sg U49652 ( .A(n45161), .B(n53361), .X(n27491) );
  nand_x4_sg U49653 ( .A(n27498), .B(n27592), .X(n27489) );
  nand_x1_sg U49654 ( .A(n27495), .B(n27497), .X(n27592) );
  nand_x2_sg U49655 ( .A(n45017), .B(n53382), .X(n27485) );
  nand_x2_sg U49656 ( .A(n45015), .B(n53406), .X(n27479) );
  nand_x1_sg U49657 ( .A(n27578), .B(n27577), .X(n27579) );
  nor_x1_sg U49658 ( .A(n53508), .B(n27814), .X(n16659) );
  nand_x1_sg U49659 ( .A(n53535), .B(n53547), .X(n27797) );
  nand_x1_sg U49660 ( .A(n27798), .B(n27799), .X(n27796) );
  nand_x2_sg U49661 ( .A(n45165), .B(n53563), .X(n27794) );
  nand_x2_sg U49662 ( .A(n45009), .B(n53546), .X(n27800) );
  nand_x1_sg U49663 ( .A(n45213), .B(n53522), .X(n27877) );
  nand_x1_sg U49664 ( .A(n27804), .B(n51126), .X(n27876) );
  inv_x1_sg U49665 ( .A(n27878), .X(n53522) );
  nand_x2_sg U49666 ( .A(n45139), .B(n53596), .X(n27782) );
  nand_x2_sg U49667 ( .A(n45007), .B(n53577), .X(n27788) );
  nand_x4_sg U49668 ( .A(n27795), .B(n27874), .X(n27786) );
  nand_x1_sg U49669 ( .A(n27792), .B(n27794), .X(n27874) );
  nand_x2_sg U49670 ( .A(n45175), .B(n53639), .X(n27770) );
  nand_x2_sg U49671 ( .A(n45005), .B(n53617), .X(n27776) );
  nand_x4_sg U49672 ( .A(n27783), .B(n27872), .X(n27774) );
  nand_x1_sg U49673 ( .A(n27780), .B(n27782), .X(n27872) );
  nand_x4_sg U49674 ( .A(n27771), .B(n27870), .X(n27762) );
  nand_x1_sg U49675 ( .A(n27768), .B(n27770), .X(n27870) );
  nand_x2_sg U49676 ( .A(n45001), .B(n53683), .X(n27758) );
  nand_x4_sg U49677 ( .A(n27765), .B(n27869), .X(n27756) );
  nand_x1_sg U49678 ( .A(n27762), .B(n27764), .X(n27869) );
  nand_x1_sg U49679 ( .A(n27857), .B(n27856), .X(n27858) );
  inv_x2_sg U49680 ( .A(n17436), .X(n44003) );
  nor_x1_sg U49681 ( .A(n53787), .B(n28095), .X(n17436) );
  inv_x1_sg U49682 ( .A(n28094), .X(n53800) );
  inv_x1_sg U49683 ( .A(n28165), .X(n53776) );
  nand_x2_sg U49684 ( .A(n28081), .B(n28082), .X(n28079) );
  inv_x1_sg U49685 ( .A(n28080), .X(n53811) );
  nand_x2_sg U49686 ( .A(n45197), .B(n53842), .X(n28075) );
  nand_x2_sg U49687 ( .A(n44995), .B(n53825), .X(n28081) );
  nand_x1_sg U49688 ( .A(n28085), .B(n51145), .X(n28157) );
  nand_x1_sg U49689 ( .A(n45981), .B(n53799), .X(n28158) );
  inv_x1_sg U49690 ( .A(n28159), .X(n53799) );
  nand_x2_sg U49691 ( .A(n44991), .B(n53881), .X(n28063) );
  nand_x2_sg U49692 ( .A(n44993), .B(n53860), .X(n28069) );
  nand_x4_sg U49693 ( .A(n28076), .B(n28155), .X(n28067) );
  nand_x1_sg U49694 ( .A(n28073), .B(n28075), .X(n28155) );
  nand_x2_sg U49695 ( .A(n44989), .B(n53924), .X(n28051) );
  nand_x2_sg U49696 ( .A(n45191), .B(n53901), .X(n28057) );
  nand_x4_sg U49697 ( .A(n28064), .B(n28153), .X(n28055) );
  nand_x1_sg U49698 ( .A(n28061), .B(n28063), .X(n28153) );
  nand_x2_sg U49699 ( .A(n45135), .B(n53942), .X(n28045) );
  nand_x4_sg U49700 ( .A(n28052), .B(n28151), .X(n28043) );
  nand_x1_sg U49701 ( .A(n28049), .B(n28051), .X(n28151) );
  nand_x2_sg U49702 ( .A(n44987), .B(n53966), .X(n28039) );
  nand_x1_sg U49703 ( .A(n28138), .B(n28137), .X(n28139) );
  nand_x1_sg U49704 ( .A(n54069), .B(n54058), .X(n28375) );
  nand_x1_sg U49705 ( .A(n28376), .B(n28377), .X(n28374) );
  nand_x1_sg U49706 ( .A(n54094), .B(n54108), .X(n28357) );
  nand_x1_sg U49707 ( .A(n28358), .B(n28359), .X(n28356) );
  nand_x4_sg U49708 ( .A(n28361), .B(n28435), .X(n28352) );
  nand_x1_sg U49709 ( .A(n28360), .B(n28359), .X(n28435) );
  nand_x2_sg U49710 ( .A(n44977), .B(n54163), .X(n28344) );
  nand_x2_sg U49711 ( .A(n44979), .B(n54140), .X(n28348) );
  nand_x2_sg U49712 ( .A(n44973), .B(n54207), .X(n28332) );
  nand_x2_sg U49713 ( .A(n44975), .B(n54182), .X(n28338) );
  nand_x4_sg U49714 ( .A(n28345), .B(n28432), .X(n28336) );
  nand_x1_sg U49715 ( .A(n28342), .B(n28344), .X(n28432) );
  nand_x2_sg U49716 ( .A(n44971), .B(n54227), .X(n28326) );
  nand_x4_sg U49717 ( .A(n28333), .B(n28430), .X(n28324) );
  nand_x1_sg U49718 ( .A(n28330), .B(n28332), .X(n28430) );
  nand_x2_sg U49719 ( .A(n44969), .B(n54248), .X(n28320) );
  nand_x1_sg U49720 ( .A(n28417), .B(n28416), .X(n28418) );
  inv_x2_sg U49721 ( .A(n18981), .X(n44001) );
  nor_x1_sg U49722 ( .A(n54352), .B(n28653), .X(n18981) );
  inv_x1_sg U49723 ( .A(n28652), .X(n54365) );
  inv_x1_sg U49724 ( .A(n28723), .X(n54341) );
  nand_x2_sg U49725 ( .A(n28639), .B(n28640), .X(n28637) );
  inv_x1_sg U49726 ( .A(n28638), .X(n54376) );
  nand_x2_sg U49727 ( .A(n45195), .B(n54407), .X(n28633) );
  nand_x2_sg U49728 ( .A(n44963), .B(n54390), .X(n28639) );
  nand_x1_sg U49729 ( .A(n28643), .B(n51182), .X(n28715) );
  nand_x1_sg U49730 ( .A(n45979), .B(n54364), .X(n28716) );
  inv_x1_sg U49731 ( .A(n28717), .X(n54364) );
  nand_x2_sg U49732 ( .A(n44959), .B(n54446), .X(n28621) );
  nand_x2_sg U49733 ( .A(n44961), .B(n54425), .X(n28627) );
  nand_x4_sg U49734 ( .A(n28634), .B(n28713), .X(n28625) );
  nand_x1_sg U49735 ( .A(n28631), .B(n28633), .X(n28713) );
  nand_x2_sg U49736 ( .A(n44957), .B(n54489), .X(n28609) );
  nand_x2_sg U49737 ( .A(n45189), .B(n54466), .X(n28615) );
  nand_x4_sg U49738 ( .A(n28622), .B(n28711), .X(n28613) );
  nand_x1_sg U49739 ( .A(n28619), .B(n28621), .X(n28711) );
  nand_x2_sg U49740 ( .A(n45133), .B(n54507), .X(n28603) );
  nand_x4_sg U49741 ( .A(n28610), .B(n28709), .X(n28601) );
  nand_x1_sg U49742 ( .A(n28607), .B(n28609), .X(n28709) );
  nand_x2_sg U49743 ( .A(n44955), .B(n54531), .X(n28597) );
  nand_x1_sg U49744 ( .A(n28696), .B(n28695), .X(n28697) );
  nand_x1_sg U49745 ( .A(n54633), .B(n28934), .X(n28931) );
  inv_x1_sg U49746 ( .A(n28922), .X(n54659) );
  nand_x1_sg U49747 ( .A(n54657), .B(n54672), .X(n28914) );
  nand_x1_sg U49748 ( .A(n28915), .B(n28916), .X(n28913) );
  nand_x2_sg U49749 ( .A(n44949), .B(n54671), .X(n28917) );
  inv_x1_sg U49750 ( .A(n28995), .X(n54656) );
  nand_x2_sg U49751 ( .A(n44945), .B(n54729), .X(n28901) );
  nand_x2_sg U49752 ( .A(n44947), .B(n54705), .X(n28905) );
  nand_x2_sg U49753 ( .A(n45151), .B(n54774), .X(n28889) );
  nand_x2_sg U49754 ( .A(n44943), .B(n54749), .X(n28895) );
  nand_x4_sg U49755 ( .A(n28902), .B(n28989), .X(n28893) );
  nand_x1_sg U49756 ( .A(n28899), .B(n28901), .X(n28989) );
  nand_x2_sg U49757 ( .A(n45157), .B(n54792), .X(n28883) );
  nand_x4_sg U49758 ( .A(n28890), .B(n28987), .X(n28881) );
  nand_x1_sg U49759 ( .A(n28887), .B(n28889), .X(n28987) );
  nand_x2_sg U49760 ( .A(n44941), .B(n54816), .X(n28877) );
  nand_x1_sg U49761 ( .A(n28974), .B(n28973), .X(n28975) );
  inv_x2_sg U49762 ( .A(n20525), .X(n43999) );
  nor_x1_sg U49763 ( .A(n54920), .B(n29214), .X(n20525) );
  inv_x1_sg U49764 ( .A(n29213), .X(n54933) );
  inv_x1_sg U49765 ( .A(n29284), .X(n54909) );
  nand_x2_sg U49766 ( .A(n29200), .B(n29201), .X(n29198) );
  inv_x1_sg U49767 ( .A(n29199), .X(n54944) );
  nand_x2_sg U49768 ( .A(n45193), .B(n54975), .X(n29194) );
  nand_x2_sg U49769 ( .A(n44935), .B(n54958), .X(n29200) );
  nand_x1_sg U49770 ( .A(n29204), .B(n51220), .X(n29276) );
  nand_x1_sg U49771 ( .A(n45977), .B(n54932), .X(n29277) );
  inv_x1_sg U49772 ( .A(n29278), .X(n54932) );
  nand_x2_sg U49773 ( .A(n44931), .B(n55014), .X(n29182) );
  nand_x2_sg U49774 ( .A(n44933), .B(n54993), .X(n29188) );
  nand_x4_sg U49775 ( .A(n29195), .B(n29274), .X(n29186) );
  nand_x1_sg U49776 ( .A(n29192), .B(n29194), .X(n29274) );
  nand_x2_sg U49777 ( .A(n44929), .B(n55057), .X(n29170) );
  nand_x2_sg U49778 ( .A(n45187), .B(n55034), .X(n29176) );
  nand_x4_sg U49779 ( .A(n29183), .B(n29272), .X(n29174) );
  nand_x1_sg U49780 ( .A(n29180), .B(n29182), .X(n29272) );
  nand_x2_sg U49781 ( .A(n45131), .B(n55075), .X(n29164) );
  nand_x4_sg U49782 ( .A(n29171), .B(n29270), .X(n29162) );
  nand_x1_sg U49783 ( .A(n29168), .B(n29170), .X(n29270) );
  nand_x2_sg U49784 ( .A(n44927), .B(n55099), .X(n29158) );
  nand_x1_sg U49785 ( .A(n29257), .B(n29256), .X(n29258) );
  nand_x1_sg U49786 ( .A(n55201), .B(n29495), .X(n29492) );
  inv_x1_sg U49787 ( .A(n29487), .X(n55214) );
  nand_x1_sg U49788 ( .A(n29488), .B(n29489), .X(n29486) );
  inv_x1_sg U49789 ( .A(n29483), .X(n55227) );
  nand_x1_sg U49790 ( .A(n55225), .B(n55240), .X(n29475) );
  nand_x1_sg U49791 ( .A(n29476), .B(n29477), .X(n29474) );
  nand_x4_sg U49792 ( .A(n29479), .B(n29553), .X(n29470) );
  nand_x1_sg U49793 ( .A(n29478), .B(n29477), .X(n29553) );
  nand_x4_sg U49794 ( .A(n29467), .B(n29551), .X(n29460) );
  nand_x1_sg U49795 ( .A(n29464), .B(n29466), .X(n29551) );
  nand_x4_sg U49796 ( .A(n29463), .B(n29550), .X(n29454) );
  nand_x1_sg U49797 ( .A(n29460), .B(n29462), .X(n29550) );
  nand_x4_sg U49798 ( .A(n29457), .B(n29549), .X(n29448) );
  nand_x1_sg U49799 ( .A(n29454), .B(n29456), .X(n29549) );
  nand_x2_sg U49800 ( .A(n45155), .B(n55360), .X(n29444) );
  nand_x4_sg U49801 ( .A(n29451), .B(n29548), .X(n29442) );
  nand_x1_sg U49802 ( .A(n29448), .B(n29450), .X(n29548) );
  nand_x2_sg U49803 ( .A(n44913), .B(n55384), .X(n29438) );
  nand_x1_sg U49804 ( .A(n29535), .B(n29534), .X(n29536) );
  inv_x1_sg U49805 ( .A(n21973), .X(n50966) );
  nand_x4_sg U49806 ( .A(n22501), .B(n50962), .X(n21958) );
  inv_x1_sg U49807 ( .A(n22502), .X(n50962) );
  nand_x1_sg U49808 ( .A(n22503), .B(n21959), .X(n22501) );
  nand_x4_sg U49809 ( .A(n50957), .B(n22516), .X(n21968) );
  inv_x1_sg U49810 ( .A(n22518), .X(n50957) );
  nand_x1_sg U49811 ( .A(n21940), .B(n45371), .X(n22516) );
  inv_x2_sg U49812 ( .A(n22514), .X(n44099) );
  nor_x1_sg U49813 ( .A(n22577), .B(n50951), .X(n22514) );
  inv_x2_sg U49814 ( .A(n22528), .X(n44748) );
  inv_x1_sg U49815 ( .A(n9409), .X(n50946) );
  inv_x1_sg U49816 ( .A(n9459), .X(n50899) );
  inv_x1_sg U49817 ( .A(n23089), .X(n50833) );
  nand_x1_sg U49818 ( .A(n8685), .B(n22838), .X(n23088) );
  inv_x1_sg U49819 ( .A(n9508), .X(n50850) );
  inv_x1_sg U49820 ( .A(n23272), .X(n50837) );
  inv_x1_sg U49821 ( .A(n23315), .X(n50789) );
  nand_x1_sg U49822 ( .A(n8686), .B(n23093), .X(n23314) );
  inv_x1_sg U49823 ( .A(n9557), .X(n50805) );
  inv_x1_sg U49824 ( .A(n23520), .X(n50743) );
  nand_x1_sg U49825 ( .A(n8687), .B(n23319), .X(n23519) );
  inv_x1_sg U49826 ( .A(n9605), .X(n50757) );
  inv_x1_sg U49827 ( .A(n23667), .X(n50747) );
  inv_x1_sg U49828 ( .A(n23710), .X(n50697) );
  nand_x1_sg U49829 ( .A(n8688), .B(n23524), .X(n23709) );
  inv_x1_sg U49830 ( .A(n9653), .X(n50710) );
  inv_x1_sg U49831 ( .A(n23881), .X(n50652) );
  nand_x1_sg U49832 ( .A(n8689), .B(n23714), .X(n23880) );
  inv_x1_sg U49833 ( .A(n9700), .X(n50662) );
  inv_x1_sg U49834 ( .A(n24034), .X(n50639) );
  nand_x1_sg U49835 ( .A(n8690), .B(n23885), .X(n24033) );
  inv_x1_sg U49836 ( .A(n9748), .X(n50615) );
  inv_x1_sg U49837 ( .A(n23991), .X(n50589) );
  nand_x1_sg U49838 ( .A(n8691), .B(n23990), .X(n23989) );
  inv_x1_sg U49839 ( .A(n9796), .X(n50566) );
  inv_x1_sg U49840 ( .A(n23985), .X(n50543) );
  nand_x1_sg U49841 ( .A(n8692), .B(n23984), .X(n23983) );
  inv_x1_sg U49842 ( .A(n9844), .X(n50519) );
  inv_x1_sg U49843 ( .A(n23979), .X(n50495) );
  nand_x1_sg U49844 ( .A(n8693), .B(n23978), .X(n23977) );
  inv_x1_sg U49845 ( .A(n9892), .X(n50472) );
  inv_x1_sg U49846 ( .A(n23973), .X(n50449) );
  nand_x1_sg U49847 ( .A(n8694), .B(n23972), .X(n23971) );
  inv_x1_sg U49848 ( .A(n9940), .X(n50426) );
  inv_x1_sg U49849 ( .A(n23967), .X(n50403) );
  nand_x1_sg U49850 ( .A(n8695), .B(n23966), .X(n23965) );
  inv_x1_sg U49851 ( .A(n9989), .X(n50379) );
  inv_x1_sg U49852 ( .A(n23961), .X(n50355) );
  nand_x1_sg U49853 ( .A(n8696), .B(n23960), .X(n23959) );
  inv_x1_sg U49854 ( .A(n10037), .X(n50332) );
  inv_x1_sg U49855 ( .A(n23955), .X(n50309) );
  nand_x1_sg U49856 ( .A(n8697), .B(n23954), .X(n23953) );
  inv_x1_sg U49857 ( .A(n10086), .X(n50286) );
  inv_x1_sg U49858 ( .A(n10135), .X(n50240) );
  inv_x2_sg U49859 ( .A(n23597), .X(n44372) );
  nor_x1_sg U49860 ( .A(n23599), .B(n23600), .X(n23597) );
  inv_x1_sg U49861 ( .A(n10182), .X(n50196) );
  inv_x1_sg U49862 ( .A(n23937), .X(n50171) );
  nand_x1_sg U49863 ( .A(n8700), .B(n23936), .X(n23935) );
  inv_x1_sg U49864 ( .A(n22674), .X(n50130) );
  nand_x4_sg U49865 ( .A(n23764), .B(n23765), .X(n10220) );
  nand_x1_sg U49866 ( .A(n10200), .B(n50135), .X(n23765) );
  nand_x1_sg U49867 ( .A(n23766), .B(n50145), .X(n23764) );
  inv_x1_sg U49868 ( .A(n23766), .X(n50135) );
  nand_x1_sg U49869 ( .A(n10226), .B(n50126), .X(n10225) );
  nand_x1_sg U49870 ( .A(n24071), .B(n50137), .X(n24070) );
  inv_x1_sg U49871 ( .A(n24072), .X(n50137) );
  inv_x1_sg U49872 ( .A(n23928), .X(n50136) );
  inv_x1_sg U49873 ( .A(n23585), .X(n50134) );
  inv_x1_sg U49874 ( .A(n10273), .X(n50109) );
  inv_x2_sg U49875 ( .A(n10290), .X(n43871) );
  nor_x1_sg U49876 ( .A(n43874), .B(n25598), .X(n10290) );
  nand_x1_sg U49877 ( .A(n10394), .B(n46572), .X(n10393) );
  inv_x1_sg U49878 ( .A(n10410), .X(n51282) );
  nand_x2_sg U49879 ( .A(n51310), .B(n10444), .X(n10431) );
  inv_x1_sg U49880 ( .A(n10445), .X(n51310) );
  nand_x1_sg U49881 ( .A(n10409), .B(n10415), .X(n10417) );
  inv_x1_sg U49882 ( .A(n10466), .X(n51326) );
  nand_x4_sg U49883 ( .A(n10452), .B(n10444), .X(n10450) );
  inv_x1_sg U49884 ( .A(n10431), .X(n51311) );
  nand_x1_sg U49885 ( .A(n51294), .B(n51289), .X(n10437) );
  inv_x1_sg U49886 ( .A(n10527), .X(n51362) );
  nand_x1_sg U49887 ( .A(n10525), .B(n10526), .X(n10524) );
  inv_x1_sg U49888 ( .A(n10556), .X(n51386) );
  nand_x1_sg U49889 ( .A(n10586), .B(n10587), .X(n10584) );
  inv_x1_sg U49890 ( .A(n10586), .X(n51402) );
  nand_x1_sg U49891 ( .A(n51388), .B(n10586), .X(n10592) );
  inv_x1_sg U49892 ( .A(n10621), .X(n51427) );
  nand_x1_sg U49893 ( .A(n10622), .B(n10623), .X(n10620) );
  inv_x1_sg U49894 ( .A(n10377), .X(n51426) );
  nand_x4_sg U49895 ( .A(n10626), .B(n10627), .X(n10377) );
  nand_x1_sg U49896 ( .A(n51410), .B(n10630), .X(n10626) );
  nand_x1_sg U49897 ( .A(n51425), .B(n10622), .X(n10627) );
  inv_x1_sg U49898 ( .A(n10631), .X(n51410) );
  inv_x1_sg U49899 ( .A(n10717), .X(n51471) );
  inv_x1_sg U49900 ( .A(n10822), .X(n51508) );
  nand_x4_sg U49901 ( .A(n10718), .B(n10719), .X(n10717) );
  nand_x1_sg U49902 ( .A(n51470), .B(n51451), .X(n10719) );
  nand_x1_sg U49903 ( .A(n10361), .B(n42093), .X(n10359) );
  inv_x1_sg U49904 ( .A(n10886), .X(n51520) );
  nand_x1_sg U49905 ( .A(n51509), .B(n10371), .X(n10370) );
  inv_x2_sg U49906 ( .A(n11058), .X(n44017) );
  nor_x1_sg U49907 ( .A(n44020), .B(n25879), .X(n11058) );
  nand_x4_sg U49908 ( .A(n11158), .B(n11159), .X(n11061) );
  nand_x1_sg U49909 ( .A(n11161), .B(n11162), .X(n11158) );
  nand_x1_sg U49910 ( .A(n11160), .B(n51537), .X(n11159) );
  nand_x1_sg U49911 ( .A(n51537), .B(n46547), .X(n11162) );
  nand_x1_sg U49912 ( .A(n11170), .B(n51543), .X(n11169) );
  nand_x1_sg U49913 ( .A(n51537), .B(n11061), .X(n11157) );
  inv_x2_sg U49914 ( .A(n11179), .X(n44675) );
  nor_x1_sg U49915 ( .A(n11181), .B(n11182), .X(n11179) );
  inv_x2_sg U49916 ( .A(n11189), .X(n43842) );
  nand_x1_sg U49917 ( .A(n11184), .B(n11183), .X(n11189) );
  nand_x4_sg U49918 ( .A(n46536), .B(n46551), .X(n11207) );
  inv_x1_sg U49919 ( .A(n11242), .X(n51601) );
  nand_x4_sg U49920 ( .A(n11227), .B(n11228), .X(n11225) );
  nand_x1_sg U49921 ( .A(n51570), .B(n11233), .X(n11227) );
  nand_x1_sg U49922 ( .A(n51584), .B(n11221), .X(n11228) );
  inv_x1_sg U49923 ( .A(n11234), .X(n51570) );
  nand_x1_sg U49924 ( .A(n51576), .B(n11211), .X(n11210) );
  inv_x1_sg U49925 ( .A(n11304), .X(n51633) );
  nand_x1_sg U49926 ( .A(n11302), .B(n11303), .X(n11301) );
  inv_x2_sg U49927 ( .A(n11307), .X(n44708) );
  nor_x1_sg U49928 ( .A(n51654), .B(n11326), .X(n11307) );
  inv_x1_sg U49929 ( .A(n11327), .X(n51653) );
  nand_x1_sg U49930 ( .A(n51679), .B(n51660), .X(n11362) );
  nand_x1_sg U49931 ( .A(n11363), .B(n11364), .X(n11361) );
  inv_x1_sg U49932 ( .A(n11363), .X(n51679) );
  inv_x1_sg U49933 ( .A(n11399), .X(n51700) );
  nand_x1_sg U49934 ( .A(n11400), .B(n11401), .X(n11398) );
  inv_x1_sg U49935 ( .A(n11451), .X(n51722) );
  nand_x1_sg U49936 ( .A(n51688), .B(n11409), .X(n11405) );
  nand_x1_sg U49937 ( .A(n51699), .B(n11400), .X(n11406) );
  inv_x1_sg U49938 ( .A(n11410), .X(n51688) );
  inv_x1_sg U49939 ( .A(n11498), .X(n51751) );
  nand_x4_sg U49940 ( .A(n11499), .B(n11500), .X(n11498) );
  nand_x1_sg U49941 ( .A(n51750), .B(n51730), .X(n11500) );
  nand_x1_sg U49942 ( .A(n11128), .B(n42091), .X(n11126) );
  inv_x2_sg U49943 ( .A(n11841), .X(n44029) );
  nor_x1_sg U49944 ( .A(n44032), .B(n26159), .X(n11841) );
  nand_x1_sg U49945 ( .A(n11944), .B(n51819), .X(n11943) );
  inv_x2_sg U49946 ( .A(n11955), .X(n44326) );
  nor_x1_sg U49947 ( .A(n11959), .B(n11960), .X(n11955) );
  inv_x2_sg U49948 ( .A(n11967), .X(n43937) );
  nand_x1_sg U49949 ( .A(n11962), .B(n11961), .X(n11967) );
  inv_x2_sg U49950 ( .A(n11966), .X(n44202) );
  nor_x1_sg U49951 ( .A(n51856), .B(n11978), .X(n11966) );
  inv_x1_sg U49952 ( .A(n12018), .X(n51882) );
  nand_x4_sg U49953 ( .A(n12004), .B(n12005), .X(n12002) );
  nand_x1_sg U49954 ( .A(n51850), .B(n12011), .X(n12004) );
  nand_x1_sg U49955 ( .A(n11997), .B(n11999), .X(n12005) );
  inv_x1_sg U49956 ( .A(n12012), .X(n51850) );
  nand_x1_sg U49957 ( .A(n51855), .B(n51849), .X(n11989) );
  inv_x1_sg U49958 ( .A(n12084), .X(n51914) );
  nand_x1_sg U49959 ( .A(n12082), .B(n12083), .X(n12081) );
  inv_x2_sg U49960 ( .A(n12087), .X(n44706) );
  nor_x1_sg U49961 ( .A(n51935), .B(n12106), .X(n12087) );
  inv_x1_sg U49962 ( .A(n12107), .X(n51934) );
  nand_x1_sg U49963 ( .A(n51960), .B(n51941), .X(n12142) );
  nand_x1_sg U49964 ( .A(n12143), .B(n12144), .X(n12141) );
  inv_x1_sg U49965 ( .A(n12143), .X(n51960) );
  inv_x1_sg U49966 ( .A(n12179), .X(n51981) );
  nand_x1_sg U49967 ( .A(n12180), .B(n12181), .X(n12178) );
  inv_x1_sg U49968 ( .A(n12231), .X(n52000) );
  nand_x1_sg U49969 ( .A(n51980), .B(n12180), .X(n12186) );
  nand_x1_sg U49970 ( .A(n51968), .B(n12189), .X(n12185) );
  inv_x1_sg U49971 ( .A(n12181), .X(n51980) );
  inv_x1_sg U49972 ( .A(n12278), .X(n52034) );
  nand_x4_sg U49973 ( .A(n12279), .B(n12280), .X(n12278) );
  nand_x1_sg U49974 ( .A(n52033), .B(n52008), .X(n12280) );
  nand_x1_sg U49975 ( .A(n11911), .B(n42079), .X(n11909) );
  inv_x2_sg U49976 ( .A(n12619), .X(n43895) );
  nor_x1_sg U49977 ( .A(n43898), .B(n26438), .X(n12619) );
  nand_x1_sg U49978 ( .A(n12721), .B(n46500), .X(n12720) );
  nand_x1_sg U49979 ( .A(n12731), .B(n52100), .X(n12730) );
  nand_x1_sg U49980 ( .A(n46500), .B(n12622), .X(n12718) );
  inv_x2_sg U49981 ( .A(n12740), .X(n44673) );
  nor_x1_sg U49982 ( .A(n12742), .B(n12743), .X(n12740) );
  inv_x2_sg U49983 ( .A(n12750), .X(n43840) );
  nand_x1_sg U49984 ( .A(n12745), .B(n12744), .X(n12750) );
  nand_x4_sg U49985 ( .A(n52133), .B(n46507), .X(n12768) );
  inv_x1_sg U49986 ( .A(n12803), .X(n52159) );
  nand_x4_sg U49987 ( .A(n12788), .B(n12789), .X(n12786) );
  nand_x1_sg U49988 ( .A(n52127), .B(n12794), .X(n12788) );
  nand_x1_sg U49989 ( .A(n52142), .B(n12782), .X(n12789) );
  inv_x1_sg U49990 ( .A(n12795), .X(n52127) );
  nand_x1_sg U49991 ( .A(n52134), .B(n12772), .X(n12771) );
  inv_x1_sg U49992 ( .A(n12865), .X(n52189) );
  nand_x1_sg U49993 ( .A(n12863), .B(n12864), .X(n12862) );
  inv_x2_sg U49994 ( .A(n12868), .X(n44704) );
  nor_x1_sg U49995 ( .A(n52210), .B(n12887), .X(n12868) );
  inv_x1_sg U49996 ( .A(n12888), .X(n52209) );
  nand_x1_sg U49997 ( .A(n52235), .B(n52216), .X(n12923) );
  nand_x1_sg U49998 ( .A(n12924), .B(n12925), .X(n12922) );
  inv_x1_sg U49999 ( .A(n12924), .X(n52235) );
  inv_x1_sg U50000 ( .A(n12960), .X(n52256) );
  nand_x1_sg U50001 ( .A(n12961), .B(n12962), .X(n12959) );
  inv_x1_sg U50002 ( .A(n13012), .X(n52276) );
  nand_x1_sg U50003 ( .A(n52243), .B(n12970), .X(n12966) );
  nand_x1_sg U50004 ( .A(n52255), .B(n12961), .X(n12967) );
  inv_x1_sg U50005 ( .A(n12971), .X(n52243) );
  inv_x1_sg U50006 ( .A(n13059), .X(n52309) );
  nand_x4_sg U50007 ( .A(n13060), .B(n13061), .X(n13059) );
  nand_x1_sg U50008 ( .A(n52308), .B(n52286), .X(n13061) );
  nand_x1_sg U50009 ( .A(n12689), .B(n42077), .X(n12687) );
  nand_x1_sg U50010 ( .A(n26724), .B(n26725), .X(n26722) );
  inv_x2_sg U50011 ( .A(n13403), .X(n43883) );
  nor_x1_sg U50012 ( .A(n43886), .B(n26716), .X(n13403) );
  nand_x1_sg U50013 ( .A(n13506), .B(n46478), .X(n13505) );
  inv_x2_sg U50014 ( .A(n13516), .X(n44324) );
  nor_x1_sg U50015 ( .A(n13520), .B(n13521), .X(n13516) );
  inv_x2_sg U50016 ( .A(n13528), .X(n43935) );
  nand_x1_sg U50017 ( .A(n13523), .B(n13522), .X(n13528) );
  inv_x2_sg U50018 ( .A(n13527), .X(n44200) );
  nor_x1_sg U50019 ( .A(n52408), .B(n13539), .X(n13527) );
  nand_x1_sg U50020 ( .A(n52407), .B(n52401), .X(n13550) );
  inv_x1_sg U50021 ( .A(n13579), .X(n52433) );
  nand_x4_sg U50022 ( .A(n13565), .B(n13566), .X(n13563) );
  nand_x1_sg U50023 ( .A(n52402), .B(n13572), .X(n13565) );
  nand_x1_sg U50024 ( .A(n13558), .B(n13560), .X(n13566) );
  inv_x1_sg U50025 ( .A(n13573), .X(n52402) );
  inv_x1_sg U50026 ( .A(n13645), .X(n52466) );
  nand_x1_sg U50027 ( .A(n13643), .B(n13644), .X(n13642) );
  inv_x2_sg U50028 ( .A(n13648), .X(n44702) );
  nor_x1_sg U50029 ( .A(n52487), .B(n13667), .X(n13648) );
  inv_x1_sg U50030 ( .A(n13668), .X(n52486) );
  nand_x1_sg U50031 ( .A(n52512), .B(n52493), .X(n13703) );
  nand_x1_sg U50032 ( .A(n13704), .B(n13705), .X(n13702) );
  inv_x1_sg U50033 ( .A(n13704), .X(n52512) );
  inv_x1_sg U50034 ( .A(n13740), .X(n52532) );
  nand_x1_sg U50035 ( .A(n13741), .B(n13742), .X(n13739) );
  inv_x1_sg U50036 ( .A(n13792), .X(n52551) );
  nand_x1_sg U50037 ( .A(n52531), .B(n13741), .X(n13747) );
  nand_x1_sg U50038 ( .A(n52519), .B(n13750), .X(n13746) );
  inv_x1_sg U50039 ( .A(n13742), .X(n52531) );
  inv_x1_sg U50040 ( .A(n13839), .X(n52584) );
  nand_x4_sg U50041 ( .A(n13840), .B(n13841), .X(n13839) );
  nand_x1_sg U50042 ( .A(n52583), .B(n52561), .X(n13841) );
  nand_x1_sg U50043 ( .A(n13473), .B(n40550), .X(n13471) );
  nor_x1_sg U50044 ( .A(n44028), .B(n26995), .X(n14182) );
  nand_x1_sg U50045 ( .A(n14286), .B(n52648), .X(n14285) );
  inv_x1_sg U50046 ( .A(n14302), .X(n52672) );
  inv_x2_sg U50047 ( .A(n14308), .X(n44198) );
  nor_x1_sg U50048 ( .A(n52685), .B(n14318), .X(n14308) );
  nand_x2_sg U50049 ( .A(n52699), .B(n14336), .X(n14323) );
  inv_x1_sg U50050 ( .A(n14337), .X(n52699) );
  nand_x1_sg U50051 ( .A(n14301), .B(n14307), .X(n14309) );
  inv_x1_sg U50052 ( .A(n14358), .X(n52716) );
  nand_x4_sg U50053 ( .A(n14344), .B(n14336), .X(n14342) );
  inv_x1_sg U50054 ( .A(n14323), .X(n52700) );
  nand_x1_sg U50055 ( .A(n52684), .B(n52679), .X(n14329) );
  inv_x1_sg U50056 ( .A(n14419), .X(n52752) );
  nand_x1_sg U50057 ( .A(n14417), .B(n14418), .X(n14416) );
  inv_x1_sg U50058 ( .A(n14448), .X(n52773) );
  nand_x1_sg U50059 ( .A(n14478), .B(n14479), .X(n14476) );
  inv_x1_sg U50060 ( .A(n14478), .X(n52791) );
  nand_x1_sg U50061 ( .A(n52776), .B(n14478), .X(n14484) );
  inv_x1_sg U50062 ( .A(n14513), .X(n52817) );
  nand_x1_sg U50063 ( .A(n14514), .B(n14515), .X(n14512) );
  inv_x1_sg U50064 ( .A(n14269), .X(n52816) );
  nand_x4_sg U50065 ( .A(n14518), .B(n14519), .X(n14269) );
  nand_x1_sg U50066 ( .A(n52815), .B(n14514), .X(n14519) );
  nand_x1_sg U50067 ( .A(n52799), .B(n14522), .X(n14518) );
  inv_x1_sg U50068 ( .A(n14515), .X(n52815) );
  inv_x1_sg U50069 ( .A(n14609), .X(n52860) );
  nand_x4_sg U50070 ( .A(n14610), .B(n14611), .X(n14609) );
  nand_x1_sg U50071 ( .A(n52859), .B(n52842), .X(n14611) );
  nand_x1_sg U50072 ( .A(n14252), .B(n42089), .X(n14250) );
  inv_x2_sg U50073 ( .A(n14258), .X(n43950) );
  nor_x1_sg U50074 ( .A(n14240), .B(n14261), .X(n14258) );
  inv_x2_sg U50075 ( .A(n14952), .X(n43891) );
  nor_x1_sg U50076 ( .A(n43894), .B(n27275), .X(n14952) );
  nand_x1_sg U50077 ( .A(n15054), .B(n46432), .X(n15053) );
  nand_x1_sg U50078 ( .A(n15064), .B(n52934), .X(n15063) );
  nand_x1_sg U50079 ( .A(n46432), .B(n14955), .X(n15051) );
  inv_x2_sg U50080 ( .A(n15073), .X(n44671) );
  nor_x1_sg U50081 ( .A(n15075), .B(n15076), .X(n15073) );
  inv_x2_sg U50082 ( .A(n15083), .X(n43838) );
  nand_x1_sg U50083 ( .A(n15078), .B(n15077), .X(n15083) );
  nand_x4_sg U50084 ( .A(n52967), .B(n46439), .X(n15101) );
  inv_x1_sg U50085 ( .A(n15136), .X(n52993) );
  nand_x4_sg U50086 ( .A(n15121), .B(n15122), .X(n15119) );
  nand_x1_sg U50087 ( .A(n52961), .B(n15127), .X(n15121) );
  nand_x1_sg U50088 ( .A(n52976), .B(n15115), .X(n15122) );
  inv_x1_sg U50089 ( .A(n15128), .X(n52961) );
  nand_x1_sg U50090 ( .A(n52968), .B(n15105), .X(n15104) );
  inv_x1_sg U50091 ( .A(n15198), .X(n53023) );
  nand_x1_sg U50092 ( .A(n15196), .B(n15197), .X(n15195) );
  inv_x2_sg U50093 ( .A(n15201), .X(n44700) );
  nor_x1_sg U50094 ( .A(n53044), .B(n15220), .X(n15201) );
  inv_x1_sg U50095 ( .A(n15221), .X(n53043) );
  nand_x1_sg U50096 ( .A(n53069), .B(n53050), .X(n15256) );
  nand_x1_sg U50097 ( .A(n15257), .B(n15258), .X(n15255) );
  inv_x1_sg U50098 ( .A(n15257), .X(n53069) );
  inv_x1_sg U50099 ( .A(n15293), .X(n53090) );
  nand_x1_sg U50100 ( .A(n15294), .B(n15295), .X(n15292) );
  inv_x1_sg U50101 ( .A(n15345), .X(n53110) );
  nand_x1_sg U50102 ( .A(n53077), .B(n15303), .X(n15299) );
  nand_x1_sg U50103 ( .A(n53089), .B(n15294), .X(n15300) );
  inv_x1_sg U50104 ( .A(n15304), .X(n53077) );
  inv_x1_sg U50105 ( .A(n15392), .X(n53143) );
  nand_x4_sg U50106 ( .A(n15393), .B(n15394), .X(n15392) );
  nand_x1_sg U50107 ( .A(n53142), .B(n53120), .X(n15394) );
  nand_x1_sg U50108 ( .A(n15022), .B(n42073), .X(n15020) );
  nor_x1_sg U50109 ( .A(n44024), .B(n27554), .X(n15736) );
  nand_x1_sg U50110 ( .A(n15839), .B(n53207), .X(n15838) );
  inv_x2_sg U50111 ( .A(n15861), .X(n44196) );
  nor_x1_sg U50112 ( .A(n53242), .B(n15873), .X(n15861) );
  inv_x1_sg U50113 ( .A(n15913), .X(n53269) );
  nand_x4_sg U50114 ( .A(n15899), .B(n15900), .X(n15897) );
  nand_x1_sg U50115 ( .A(n53236), .B(n15906), .X(n15899) );
  nand_x1_sg U50116 ( .A(n15892), .B(n15894), .X(n15900) );
  inv_x1_sg U50117 ( .A(n15907), .X(n53236) );
  nand_x1_sg U50118 ( .A(n53241), .B(n53235), .X(n15884) );
  inv_x1_sg U50119 ( .A(n15979), .X(n53301) );
  nand_x1_sg U50120 ( .A(n15977), .B(n15978), .X(n15976) );
  inv_x2_sg U50121 ( .A(n15982), .X(n44698) );
  nor_x1_sg U50122 ( .A(n53323), .B(n16001), .X(n15982) );
  inv_x1_sg U50123 ( .A(n16002), .X(n53322) );
  nand_x1_sg U50124 ( .A(n53348), .B(n53329), .X(n16037) );
  nand_x1_sg U50125 ( .A(n16038), .B(n16039), .X(n16036) );
  inv_x1_sg U50126 ( .A(n16038), .X(n53348) );
  inv_x1_sg U50127 ( .A(n16074), .X(n53370) );
  nand_x1_sg U50128 ( .A(n16075), .B(n16076), .X(n16073) );
  inv_x1_sg U50129 ( .A(n16126), .X(n53389) );
  nand_x1_sg U50130 ( .A(n53369), .B(n16075), .X(n16081) );
  nand_x1_sg U50131 ( .A(n53357), .B(n16084), .X(n16080) );
  inv_x1_sg U50132 ( .A(n16076), .X(n53369) );
  inv_x1_sg U50133 ( .A(n16173), .X(n53420) );
  inv_x1_sg U50134 ( .A(n16278), .X(n53458) );
  nand_x4_sg U50135 ( .A(n16174), .B(n16175), .X(n16173) );
  nand_x1_sg U50136 ( .A(n53419), .B(n53399), .X(n16175) );
  nand_x1_sg U50137 ( .A(n15807), .B(n42087), .X(n15805) );
  inv_x1_sg U50138 ( .A(n16341), .X(n53469) );
  nand_x1_sg U50139 ( .A(n53459), .B(n15817), .X(n15816) );
  inv_x2_sg U50140 ( .A(n16518), .X(n43887) );
  nor_x1_sg U50141 ( .A(n43890), .B(n27833), .X(n16518) );
  nand_x1_sg U50142 ( .A(n16620), .B(n46388), .X(n16619) );
  nand_x1_sg U50143 ( .A(n16630), .B(n53492), .X(n16629) );
  nand_x1_sg U50144 ( .A(n46388), .B(n16521), .X(n16617) );
  inv_x2_sg U50145 ( .A(n16639), .X(n44669) );
  nor_x1_sg U50146 ( .A(n16641), .B(n16642), .X(n16639) );
  inv_x2_sg U50147 ( .A(n16649), .X(n43836) );
  nand_x1_sg U50148 ( .A(n16644), .B(n16643), .X(n16649) );
  nand_x4_sg U50149 ( .A(n53525), .B(n46395), .X(n16667) );
  inv_x1_sg U50150 ( .A(n16702), .X(n53551) );
  nand_x4_sg U50151 ( .A(n16687), .B(n16688), .X(n16685) );
  nand_x1_sg U50152 ( .A(n53519), .B(n16693), .X(n16687) );
  nand_x1_sg U50153 ( .A(n53534), .B(n16681), .X(n16688) );
  inv_x1_sg U50154 ( .A(n16694), .X(n53519) );
  nand_x1_sg U50155 ( .A(n53526), .B(n16671), .X(n16670) );
  inv_x1_sg U50156 ( .A(n16764), .X(n53581) );
  nand_x1_sg U50157 ( .A(n16762), .B(n16763), .X(n16761) );
  inv_x2_sg U50158 ( .A(n16767), .X(n44696) );
  nor_x1_sg U50159 ( .A(n53602), .B(n16786), .X(n16767) );
  inv_x1_sg U50160 ( .A(n16787), .X(n53601) );
  nand_x1_sg U50161 ( .A(n53627), .B(n53608), .X(n16822) );
  nand_x1_sg U50162 ( .A(n16823), .B(n16824), .X(n16821) );
  inv_x1_sg U50163 ( .A(n16823), .X(n53627) );
  inv_x1_sg U50164 ( .A(n16859), .X(n53648) );
  nand_x1_sg U50165 ( .A(n16860), .B(n16861), .X(n16858) );
  inv_x1_sg U50166 ( .A(n16911), .X(n53668) );
  nand_x1_sg U50167 ( .A(n53635), .B(n16869), .X(n16865) );
  nand_x1_sg U50168 ( .A(n53647), .B(n16860), .X(n16866) );
  inv_x1_sg U50169 ( .A(n16870), .X(n53635) );
  inv_x1_sg U50170 ( .A(n16958), .X(n53701) );
  nand_x4_sg U50171 ( .A(n16959), .B(n16960), .X(n16958) );
  nand_x1_sg U50172 ( .A(n53700), .B(n53678), .X(n16960) );
  nand_x1_sg U50173 ( .A(n16588), .B(n42069), .X(n16586) );
  inv_x2_sg U50174 ( .A(n17301), .X(n44013) );
  nor_x1_sg U50175 ( .A(n44016), .B(n28114), .X(n17301) );
  nand_x1_sg U50176 ( .A(n17405), .B(n53765), .X(n17404) );
  nand_x1_sg U50177 ( .A(n17414), .B(n46363), .X(n17413) );
  nand_x2_sg U50178 ( .A(n17422), .B(n53791), .X(n17419) );
  inv_x1_sg U50179 ( .A(n17423), .X(n53791) );
  nand_x2_sg U50180 ( .A(n53783), .B(n53793), .X(n17399) );
  inv_x1_sg U50181 ( .A(n17419), .X(n53793) );
  inv_x2_sg U50182 ( .A(n17446), .X(n53819) );
  nor_x1_sg U50183 ( .A(n17459), .B(n53818), .X(n17446) );
  nand_x1_sg U50184 ( .A(n17422), .B(n17428), .X(n17430) );
  inv_x1_sg U50185 ( .A(n17480), .X(n53830) );
  nand_x4_sg U50186 ( .A(n17467), .B(n17460), .X(n17465) );
  inv_x1_sg U50187 ( .A(n53819), .X(n44156) );
  nand_x1_sg U50188 ( .A(n53803), .B(n53798), .X(n17452) );
  inv_x1_sg U50189 ( .A(n17539), .X(n53872) );
  nand_x1_sg U50190 ( .A(n17537), .B(n17538), .X(n17536) );
  inv_x1_sg U50191 ( .A(n17568), .X(n53893) );
  nand_x1_sg U50192 ( .A(n17599), .B(n17600), .X(n17597) );
  inv_x1_sg U50193 ( .A(n17599), .X(n53911) );
  nand_x1_sg U50194 ( .A(n53896), .B(n17599), .X(n17605) );
  inv_x1_sg U50195 ( .A(n17634), .X(n53937) );
  nand_x1_sg U50196 ( .A(n17635), .B(n17636), .X(n17633) );
  inv_x1_sg U50197 ( .A(n17388), .X(n53936) );
  nand_x4_sg U50198 ( .A(n17639), .B(n17640), .X(n17388) );
  nand_x1_sg U50199 ( .A(n53935), .B(n17635), .X(n17640) );
  nand_x1_sg U50200 ( .A(n53920), .B(n17643), .X(n17639) );
  inv_x1_sg U50201 ( .A(n17636), .X(n53935) );
  inv_x1_sg U50202 ( .A(n17730), .X(n53980) );
  nand_x4_sg U50203 ( .A(n17731), .B(n17732), .X(n17730) );
  nand_x1_sg U50204 ( .A(n53979), .B(n53962), .X(n17732) );
  nand_x1_sg U50205 ( .A(n17371), .B(n42085), .X(n17369) );
  inv_x2_sg U50206 ( .A(n17377), .X(n43948) );
  nor_x1_sg U50207 ( .A(n17359), .B(n17380), .X(n17377) );
  inv_x2_sg U50208 ( .A(n18073), .X(n43857) );
  nor_x1_sg U50209 ( .A(n54049), .B(n28392), .X(n18073) );
  nand_x1_sg U50210 ( .A(n18176), .B(n46345), .X(n18175) );
  inv_x2_sg U50211 ( .A(n18196), .X(n44194) );
  nor_x1_sg U50212 ( .A(n54086), .B(n18207), .X(n18196) );
  nand_x2_sg U50213 ( .A(n54100), .B(n18225), .X(n18212) );
  inv_x1_sg U50214 ( .A(n18226), .X(n54100) );
  nand_x1_sg U50215 ( .A(n18189), .B(n18195), .X(n18197) );
  inv_x1_sg U50216 ( .A(n18248), .X(n54117) );
  inv_x1_sg U50217 ( .A(n18212), .X(n54101) );
  nand_x1_sg U50218 ( .A(n54085), .B(n54079), .X(n18218) );
  nor_x1_sg U50219 ( .A(n18252), .B(n54121), .X(n18251) );
  inv_x1_sg U50220 ( .A(n18309), .X(n54151) );
  nand_x1_sg U50221 ( .A(n18307), .B(n18308), .X(n18306) );
  nand_x1_sg U50222 ( .A(n54118), .B(n18231), .X(n18167) );
  inv_x1_sg U50223 ( .A(n18338), .X(n54174) );
  nand_x1_sg U50224 ( .A(n18368), .B(n18369), .X(n18366) );
  inv_x1_sg U50225 ( .A(n18368), .X(n54191) );
  nand_x1_sg U50226 ( .A(n54176), .B(n18368), .X(n18374) );
  inv_x1_sg U50227 ( .A(n18403), .X(n54217) );
  nand_x1_sg U50228 ( .A(n18404), .B(n18405), .X(n18402) );
  inv_x1_sg U50229 ( .A(n18159), .X(n54216) );
  nand_x4_sg U50230 ( .A(n18408), .B(n18409), .X(n18159) );
  nand_x1_sg U50231 ( .A(n54203), .B(n18412), .X(n18408) );
  nand_x1_sg U50232 ( .A(n54215), .B(n18404), .X(n18409) );
  inv_x1_sg U50233 ( .A(n18413), .X(n54203) );
  inv_x1_sg U50234 ( .A(n18499), .X(n54264) );
  nand_x4_sg U50235 ( .A(n18500), .B(n18501), .X(n18499) );
  nand_x1_sg U50236 ( .A(n54263), .B(n54244), .X(n18501) );
  nand_x1_sg U50237 ( .A(n54239), .B(n40558), .X(n18141) );
  inv_x2_sg U50238 ( .A(n18846), .X(n44009) );
  nor_x1_sg U50239 ( .A(n44012), .B(n28672), .X(n18846) );
  nand_x1_sg U50240 ( .A(n18950), .B(n54330), .X(n18949) );
  nand_x1_sg U50241 ( .A(n18959), .B(n46316), .X(n18958) );
  nand_x2_sg U50242 ( .A(n18967), .B(n54356), .X(n18964) );
  inv_x1_sg U50243 ( .A(n18968), .X(n54356) );
  nand_x2_sg U50244 ( .A(n54348), .B(n54358), .X(n18944) );
  inv_x1_sg U50245 ( .A(n18964), .X(n54358) );
  inv_x2_sg U50246 ( .A(n18991), .X(n54384) );
  nor_x1_sg U50247 ( .A(n19004), .B(n54383), .X(n18991) );
  nand_x1_sg U50248 ( .A(n18967), .B(n18973), .X(n18975) );
  inv_x1_sg U50249 ( .A(n19025), .X(n54395) );
  nand_x4_sg U50250 ( .A(n19012), .B(n19005), .X(n19010) );
  inv_x1_sg U50251 ( .A(n54384), .X(n44155) );
  nand_x1_sg U50252 ( .A(n54368), .B(n54363), .X(n18997) );
  inv_x1_sg U50253 ( .A(n19084), .X(n54437) );
  nand_x1_sg U50254 ( .A(n19082), .B(n19083), .X(n19081) );
  inv_x1_sg U50255 ( .A(n19113), .X(n54458) );
  nand_x1_sg U50256 ( .A(n19144), .B(n19145), .X(n19142) );
  inv_x1_sg U50257 ( .A(n19144), .X(n54476) );
  nand_x1_sg U50258 ( .A(n54461), .B(n19144), .X(n19150) );
  inv_x1_sg U50259 ( .A(n19179), .X(n54502) );
  nand_x1_sg U50260 ( .A(n19180), .B(n19181), .X(n19178) );
  inv_x1_sg U50261 ( .A(n18933), .X(n54501) );
  nand_x4_sg U50262 ( .A(n19184), .B(n19185), .X(n18933) );
  nand_x1_sg U50263 ( .A(n54500), .B(n19180), .X(n19185) );
  nand_x1_sg U50264 ( .A(n54485), .B(n19188), .X(n19184) );
  inv_x1_sg U50265 ( .A(n19181), .X(n54500) );
  inv_x1_sg U50266 ( .A(n19275), .X(n54545) );
  nand_x4_sg U50267 ( .A(n19276), .B(n19277), .X(n19275) );
  nand_x1_sg U50268 ( .A(n54544), .B(n54527), .X(n19277) );
  nand_x1_sg U50269 ( .A(n18916), .B(n42083), .X(n18914) );
  inv_x2_sg U50270 ( .A(n18922), .X(n43946) );
  nor_x1_sg U50271 ( .A(n18904), .B(n18925), .X(n18922) );
  inv_x2_sg U50272 ( .A(n19618), .X(n43875) );
  nor_x1_sg U50273 ( .A(n43878), .B(n28950), .X(n19618) );
  nand_x1_sg U50274 ( .A(n19721), .B(n54614), .X(n19720) );
  inv_x1_sg U50275 ( .A(n19737), .X(n54636) );
  nand_x2_sg U50276 ( .A(n54664), .B(n19771), .X(n19758) );
  inv_x1_sg U50277 ( .A(n19772), .X(n54664) );
  nand_x1_sg U50278 ( .A(n19736), .B(n19742), .X(n19744) );
  inv_x1_sg U50279 ( .A(n19793), .X(n54680) );
  nand_x4_sg U50280 ( .A(n19779), .B(n19771), .X(n19777) );
  inv_x1_sg U50281 ( .A(n19758), .X(n54665) );
  nand_x1_sg U50282 ( .A(n54648), .B(n54643), .X(n19764) );
  inv_x1_sg U50283 ( .A(n19854), .X(n54716) );
  nand_x1_sg U50284 ( .A(n19852), .B(n19853), .X(n19851) );
  inv_x1_sg U50285 ( .A(n19883), .X(n54740) );
  nand_x1_sg U50286 ( .A(n19913), .B(n19914), .X(n19911) );
  inv_x1_sg U50287 ( .A(n19913), .X(n54758) );
  nand_x1_sg U50288 ( .A(n54743), .B(n19913), .X(n19919) );
  inv_x1_sg U50289 ( .A(n19948), .X(n54786) );
  nand_x1_sg U50290 ( .A(n19949), .B(n19950), .X(n19947) );
  inv_x1_sg U50291 ( .A(n19704), .X(n54785) );
  nand_x4_sg U50292 ( .A(n19953), .B(n19954), .X(n19704) );
  nand_x1_sg U50293 ( .A(n54771), .B(n19957), .X(n19953) );
  nand_x1_sg U50294 ( .A(n54784), .B(n19949), .X(n19954) );
  inv_x1_sg U50295 ( .A(n19958), .X(n54771) );
  inv_x1_sg U50296 ( .A(n20044), .X(n54831) );
  nand_x4_sg U50297 ( .A(n20045), .B(n20046), .X(n20044) );
  nand_x1_sg U50298 ( .A(n54830), .B(n54812), .X(n20046) );
  nand_x1_sg U50299 ( .A(n54804), .B(n42097), .X(n19686) );
  inv_x2_sg U50300 ( .A(n20390), .X(n44005) );
  nor_x1_sg U50301 ( .A(n44008), .B(n29233), .X(n20390) );
  nand_x1_sg U50302 ( .A(n20494), .B(n54898), .X(n20493) );
  nand_x1_sg U50303 ( .A(n20503), .B(n46271), .X(n20502) );
  nand_x2_sg U50304 ( .A(n20511), .B(n54924), .X(n20508) );
  inv_x1_sg U50305 ( .A(n20512), .X(n54924) );
  nand_x2_sg U50306 ( .A(n54916), .B(n54926), .X(n20488) );
  inv_x1_sg U50307 ( .A(n20508), .X(n54926) );
  inv_x2_sg U50308 ( .A(n20535), .X(n54952) );
  nor_x1_sg U50309 ( .A(n20548), .B(n54951), .X(n20535) );
  nand_x1_sg U50310 ( .A(n20511), .B(n20517), .X(n20519) );
  inv_x1_sg U50311 ( .A(n20569), .X(n54963) );
  nand_x4_sg U50312 ( .A(n20556), .B(n20549), .X(n20554) );
  inv_x1_sg U50313 ( .A(n54952), .X(n44154) );
  nand_x1_sg U50314 ( .A(n54936), .B(n54931), .X(n20541) );
  inv_x1_sg U50315 ( .A(n20628), .X(n55005) );
  nand_x1_sg U50316 ( .A(n20626), .B(n20627), .X(n20625) );
  inv_x1_sg U50317 ( .A(n20657), .X(n55026) );
  nand_x1_sg U50318 ( .A(n20688), .B(n20689), .X(n20686) );
  inv_x1_sg U50319 ( .A(n20688), .X(n55044) );
  nand_x1_sg U50320 ( .A(n55029), .B(n20688), .X(n20694) );
  inv_x1_sg U50321 ( .A(n20723), .X(n55070) );
  nand_x1_sg U50322 ( .A(n20724), .B(n20725), .X(n20722) );
  inv_x1_sg U50323 ( .A(n20477), .X(n55069) );
  nand_x4_sg U50324 ( .A(n20728), .B(n20729), .X(n20477) );
  nand_x1_sg U50325 ( .A(n55068), .B(n20724), .X(n20729) );
  nand_x1_sg U50326 ( .A(n55053), .B(n20732), .X(n20728) );
  inv_x1_sg U50327 ( .A(n20725), .X(n55068) );
  inv_x1_sg U50328 ( .A(n20819), .X(n55113) );
  nand_x4_sg U50329 ( .A(n20820), .B(n20821), .X(n20819) );
  nand_x1_sg U50330 ( .A(n55112), .B(n55095), .X(n20821) );
  nand_x1_sg U50331 ( .A(n20460), .B(n42081), .X(n20458) );
  inv_x2_sg U50332 ( .A(n20466), .X(n43944) );
  nor_x1_sg U50333 ( .A(n20448), .B(n20469), .X(n20466) );
  inv_x2_sg U50334 ( .A(n21163), .X(n43879) );
  nor_x1_sg U50335 ( .A(n43882), .B(n29511), .X(n21163) );
  nand_x1_sg U50336 ( .A(n21266), .B(n55182), .X(n21265) );
  inv_x1_sg U50337 ( .A(n21282), .X(n55204) );
  nand_x2_sg U50338 ( .A(n55232), .B(n21316), .X(n21303) );
  inv_x1_sg U50339 ( .A(n21317), .X(n55232) );
  nand_x1_sg U50340 ( .A(n21281), .B(n21287), .X(n21289) );
  inv_x1_sg U50341 ( .A(n21338), .X(n55248) );
  nand_x4_sg U50342 ( .A(n21324), .B(n21316), .X(n21322) );
  inv_x1_sg U50343 ( .A(n21303), .X(n55233) );
  nand_x1_sg U50344 ( .A(n55216), .B(n55211), .X(n21309) );
  inv_x1_sg U50345 ( .A(n21399), .X(n55284) );
  nand_x1_sg U50346 ( .A(n21397), .B(n21398), .X(n21396) );
  inv_x1_sg U50347 ( .A(n21428), .X(n55308) );
  nand_x1_sg U50348 ( .A(n21458), .B(n21459), .X(n21456) );
  inv_x1_sg U50349 ( .A(n21458), .X(n55326) );
  nand_x1_sg U50350 ( .A(n55311), .B(n21458), .X(n21464) );
  inv_x1_sg U50351 ( .A(n21493), .X(n55354) );
  nand_x1_sg U50352 ( .A(n21494), .B(n21495), .X(n21492) );
  inv_x1_sg U50353 ( .A(n21249), .X(n55353) );
  nand_x4_sg U50354 ( .A(n21498), .B(n21499), .X(n21249) );
  nand_x1_sg U50355 ( .A(n55339), .B(n21502), .X(n21498) );
  nand_x1_sg U50356 ( .A(n55352), .B(n21494), .X(n21499) );
  inv_x1_sg U50357 ( .A(n21503), .X(n55339) );
  inv_x1_sg U50358 ( .A(n21589), .X(n55399) );
  nand_x4_sg U50359 ( .A(n21590), .B(n21591), .X(n21589) );
  nand_x1_sg U50360 ( .A(n55398), .B(n55380), .X(n21591) );
  nand_x1_sg U50361 ( .A(n55372), .B(n42095), .X(n21231) );
  inv_x1_sg U50362 ( .A(n29638), .X(n50107) );
  nand_x4_sg U50363 ( .A(n30167), .B(n50103), .X(n29615) );
  inv_x1_sg U50364 ( .A(n30168), .X(n50103) );
  nand_x1_sg U50365 ( .A(n30169), .B(n29618), .X(n30167) );
  nand_x4_sg U50366 ( .A(n50098), .B(n30182), .X(n29631) );
  inv_x1_sg U50367 ( .A(n30184), .X(n50098) );
  nand_x1_sg U50368 ( .A(n29592), .B(n45361), .X(n30182) );
  inv_x2_sg U50369 ( .A(n30180), .X(n44097) );
  nor_x1_sg U50370 ( .A(n30243), .B(n50092), .X(n30180) );
  inv_x2_sg U50371 ( .A(n30194), .X(n44746) );
  inv_x1_sg U50372 ( .A(n24518), .X(n50087) );
  inv_x1_sg U50373 ( .A(n24567), .X(n50040) );
  inv_x1_sg U50374 ( .A(n24616), .X(n49991) );
  inv_x1_sg U50375 ( .A(n30938), .X(n49978) );
  nand_x1_sg U50376 ( .A(n8346), .B(n49936), .X(n30993) );
  inv_x1_sg U50377 ( .A(n24665), .X(n49946) );
  inv_x1_sg U50378 ( .A(n24713), .X(n49898) );
  inv_x1_sg U50379 ( .A(n31333), .X(n49888) );
  nand_x1_sg U50380 ( .A(n8348), .B(n49871), .X(n31388) );
  inv_x1_sg U50381 ( .A(n24761), .X(n49851) );
  inv_x1_sg U50382 ( .A(n24808), .X(n49803) );
  inv_x1_sg U50383 ( .A(n24856), .X(n49756) );
  inv_x1_sg U50384 ( .A(n24904), .X(n49707) );
  inv_x1_sg U50385 ( .A(n24952), .X(n49660) );
  inv_x1_sg U50386 ( .A(n25000), .X(n49613) );
  inv_x1_sg U50387 ( .A(n25048), .X(n49567) );
  inv_x1_sg U50388 ( .A(n25097), .X(n49520) );
  inv_x1_sg U50389 ( .A(n25145), .X(n49473) );
  inv_x1_sg U50390 ( .A(n25194), .X(n49427) );
  inv_x1_sg U50391 ( .A(n25243), .X(n49381) );
  inv_x2_sg U50392 ( .A(n31263), .X(n44370) );
  nor_x1_sg U50393 ( .A(n31265), .B(n31266), .X(n31263) );
  inv_x1_sg U50394 ( .A(n25290), .X(n49337) );
  nand_x1_sg U50395 ( .A(n8360), .B(n31261), .X(n31260) );
  inv_x1_sg U50396 ( .A(n30340), .X(n49271) );
  nand_x1_sg U50397 ( .A(n25334), .B(n49267), .X(n25333) );
  nand_x2_sg U50398 ( .A(n31252), .B(n31253), .X(n31251) );
  nand_x4_sg U50399 ( .A(n31430), .B(n31431), .X(n25328) );
  nand_x1_sg U50400 ( .A(n25307), .B(n49276), .X(n31431) );
  nand_x1_sg U50401 ( .A(n31432), .B(n49286), .X(n31430) );
  inv_x1_sg U50402 ( .A(n31432), .X(n49276) );
  inv_x1_sg U50403 ( .A(n31594), .X(n49277) );
  inv_x1_sg U50404 ( .A(n25379), .X(n49250) );
  nand_x4_sg U50405 ( .A(n11039), .B(n51352), .X(n25459) );
  inv_x1_sg U50406 ( .A(n11038), .X(n51352) );
  nand_x4_sg U50407 ( .A(n25554), .B(n25640), .X(n25547) );
  nand_x1_sg U50408 ( .A(n25551), .B(n25553), .X(n25640) );
  nand_x4_sg U50409 ( .A(n25544), .B(n25638), .X(n25535) );
  nand_x1_sg U50410 ( .A(n25541), .B(n25543), .X(n25638) );
  nand_x4_sg U50411 ( .A(n25532), .B(n25636), .X(n25523) );
  nand_x1_sg U50412 ( .A(n25529), .B(n25531), .X(n25636) );
  nand_x1_sg U50413 ( .A(n25622), .B(n25621), .X(n25623) );
  nand_x4_sg U50414 ( .A(n25526), .B(n25635), .X(n25616) );
  nand_x1_sg U50415 ( .A(n25523), .B(n25525), .X(n25635) );
  nand_x4_sg U50416 ( .A(n25847), .B(n25921), .X(n25838) );
  nand_x1_sg U50417 ( .A(n25846), .B(n25845), .X(n25921) );
  nand_x4_sg U50418 ( .A(n25835), .B(n25919), .X(n25826) );
  nand_x1_sg U50419 ( .A(n25832), .B(n25834), .X(n25919) );
  nand_x4_sg U50420 ( .A(n25817), .B(n25916), .X(n25808) );
  nand_x1_sg U50421 ( .A(n25814), .B(n25816), .X(n25916) );
  nand_x4_sg U50422 ( .A(n25811), .B(n25915), .X(n25802) );
  nand_x1_sg U50423 ( .A(n25808), .B(n25810), .X(n25915) );
  nand_x4_sg U50424 ( .A(n25805), .B(n25914), .X(n25897) );
  nand_x1_sg U50425 ( .A(n25802), .B(n25804), .X(n25914) );
  inv_x2_sg U50426 ( .A(n25674), .X(n44165) );
  nor_x1_sg U50427 ( .A(n51806), .B(n25901), .X(n25674) );
  nand_x4_sg U50428 ( .A(n11829), .B(n51779), .X(n25783) );
  inv_x1_sg U50429 ( .A(n11828), .X(n51779) );
  nand_x4_sg U50430 ( .A(n26127), .B(n26201), .X(n26118) );
  nand_x1_sg U50431 ( .A(n26126), .B(n26125), .X(n26201) );
  nand_x4_sg U50432 ( .A(n26115), .B(n26199), .X(n26106) );
  nand_x1_sg U50433 ( .A(n26112), .B(n26114), .X(n26199) );
  inv_x4_sg U50434 ( .A(n12295), .X(n51952) );
  nand_x4_sg U50435 ( .A(n26097), .B(n26196), .X(n26088) );
  nand_x1_sg U50436 ( .A(n26094), .B(n26096), .X(n26196) );
  nand_x4_sg U50437 ( .A(n26085), .B(n26194), .X(n26177) );
  nand_x1_sg U50438 ( .A(n26082), .B(n26084), .X(n26194) );
  inv_x2_sg U50439 ( .A(n25952), .X(n44167) );
  nor_x1_sg U50440 ( .A(n52082), .B(n26181), .X(n25952) );
  nand_x4_sg U50441 ( .A(n12608), .B(n52059), .X(n26062) );
  inv_x1_sg U50442 ( .A(n12607), .X(n52059) );
  nand_x4_sg U50443 ( .A(n26406), .B(n26480), .X(n26397) );
  nand_x1_sg U50444 ( .A(n26405), .B(n26404), .X(n26480) );
  nand_x4_sg U50445 ( .A(n26394), .B(n26478), .X(n26385) );
  nand_x1_sg U50446 ( .A(n26391), .B(n26393), .X(n26478) );
  inv_x4_sg U50447 ( .A(n13076), .X(n52227) );
  nand_x4_sg U50448 ( .A(n26382), .B(n26476), .X(n26373) );
  nand_x1_sg U50449 ( .A(n26379), .B(n26381), .X(n26476) );
  nand_x4_sg U50450 ( .A(n26364), .B(n26473), .X(n26456) );
  nand_x1_sg U50451 ( .A(n26361), .B(n26363), .X(n26473) );
  inv_x2_sg U50452 ( .A(n26233), .X(n43791) );
  nor_x1_sg U50453 ( .A(n52360), .B(n26460), .X(n26233) );
  nand_x4_sg U50454 ( .A(n13390), .B(n52336), .X(n26343) );
  inv_x1_sg U50455 ( .A(n13389), .X(n52336) );
  nand_x4_sg U50456 ( .A(n26672), .B(n26756), .X(n26663) );
  nand_x1_sg U50457 ( .A(n26669), .B(n26671), .X(n26756) );
  inv_x4_sg U50458 ( .A(n13856), .X(n52504) );
  nand_x4_sg U50459 ( .A(n26660), .B(n26754), .X(n26651) );
  nand_x1_sg U50460 ( .A(n26657), .B(n26659), .X(n26754) );
  nand_x4_sg U50461 ( .A(n26642), .B(n26751), .X(n26734) );
  nand_x1_sg U50462 ( .A(n26639), .B(n26641), .X(n26751) );
  inv_x2_sg U50463 ( .A(n26512), .X(n43808) );
  nor_x1_sg U50464 ( .A(n52635), .B(n26738), .X(n26512) );
  nand_x4_sg U50465 ( .A(n14170), .B(n52611), .X(n26622) );
  inv_x1_sg U50466 ( .A(n14169), .X(n52611) );
  inv_x1_sg U50467 ( .A(n26960), .X(n52706) );
  nand_x4_sg U50468 ( .A(n26963), .B(n27037), .X(n26954) );
  nand_x1_sg U50469 ( .A(n26962), .B(n26961), .X(n27037) );
  nand_x4_sg U50470 ( .A(n26951), .B(n27035), .X(n26942) );
  nand_x1_sg U50471 ( .A(n26948), .B(n26950), .X(n27035) );
  nand_x4_sg U50472 ( .A(n26939), .B(n27033), .X(n26930) );
  nand_x1_sg U50473 ( .A(n26936), .B(n26938), .X(n27033) );
  nand_x4_sg U50474 ( .A(n26927), .B(n27031), .X(n26918) );
  nand_x1_sg U50475 ( .A(n26924), .B(n26926), .X(n27031) );
  nand_x4_sg U50476 ( .A(n26921), .B(n27030), .X(n27013) );
  nand_x1_sg U50477 ( .A(n26918), .B(n26920), .X(n27030) );
  inv_x2_sg U50478 ( .A(n26790), .X(n43785) );
  nor_x1_sg U50479 ( .A(n52916), .B(n27017), .X(n26790) );
  nand_x4_sg U50480 ( .A(n14941), .B(n52889), .X(n26899) );
  inv_x1_sg U50481 ( .A(n14940), .X(n52889) );
  nand_x4_sg U50482 ( .A(n27243), .B(n27317), .X(n27234) );
  nand_x1_sg U50483 ( .A(n27242), .B(n27241), .X(n27317) );
  nand_x4_sg U50484 ( .A(n27231), .B(n27315), .X(n27222) );
  nand_x1_sg U50485 ( .A(n27228), .B(n27230), .X(n27315) );
  inv_x4_sg U50486 ( .A(n15409), .X(n53061) );
  nand_x4_sg U50487 ( .A(n27219), .B(n27313), .X(n27210) );
  nand_x1_sg U50488 ( .A(n27216), .B(n27218), .X(n27313) );
  nand_x4_sg U50489 ( .A(n27201), .B(n27310), .X(n27293) );
  nand_x1_sg U50490 ( .A(n27198), .B(n27200), .X(n27310) );
  inv_x2_sg U50491 ( .A(n27069), .X(n43789) );
  nor_x1_sg U50492 ( .A(n53194), .B(n27297), .X(n27069) );
  nand_x4_sg U50493 ( .A(n15723), .B(n53170), .X(n27179) );
  inv_x1_sg U50494 ( .A(n15722), .X(n53170) );
  nand_x4_sg U50495 ( .A(n27510), .B(n27594), .X(n27501) );
  nand_x1_sg U50496 ( .A(n27507), .B(n27509), .X(n27594) );
  nand_x4_sg U50497 ( .A(n27492), .B(n27591), .X(n27483) );
  nand_x1_sg U50498 ( .A(n27489), .B(n27491), .X(n27591) );
  nand_x4_sg U50499 ( .A(n27486), .B(n27590), .X(n27477) );
  nand_x1_sg U50500 ( .A(n27483), .B(n27485), .X(n27590) );
  nand_x4_sg U50501 ( .A(n27480), .B(n27589), .X(n27572) );
  nand_x1_sg U50502 ( .A(n27477), .B(n27479), .X(n27589) );
  inv_x2_sg U50503 ( .A(n27349), .X(n44163) );
  nor_x1_sg U50504 ( .A(n53474), .B(n27576), .X(n27349) );
  nand_x4_sg U50505 ( .A(n16506), .B(n53448), .X(n27458) );
  inv_x1_sg U50506 ( .A(n16505), .X(n53448) );
  nand_x4_sg U50507 ( .A(n27801), .B(n27875), .X(n27792) );
  nand_x1_sg U50508 ( .A(n27800), .B(n27799), .X(n27875) );
  nand_x4_sg U50509 ( .A(n27789), .B(n27873), .X(n27780) );
  nand_x1_sg U50510 ( .A(n27786), .B(n27788), .X(n27873) );
  inv_x4_sg U50511 ( .A(n16975), .X(n53619) );
  nand_x4_sg U50512 ( .A(n27777), .B(n27871), .X(n27768) );
  nand_x1_sg U50513 ( .A(n27774), .B(n27776), .X(n27871) );
  nand_x4_sg U50514 ( .A(n27759), .B(n27868), .X(n27851) );
  nand_x1_sg U50515 ( .A(n27756), .B(n27758), .X(n27868) );
  inv_x2_sg U50516 ( .A(n27629), .X(n43853) );
  nor_x1_sg U50517 ( .A(n53752), .B(n27855), .X(n27629) );
  nand_x4_sg U50518 ( .A(n17289), .B(n53728), .X(n27739) );
  inv_x1_sg U50519 ( .A(n17288), .X(n53728) );
  inv_x1_sg U50520 ( .A(n28079), .X(n53826) );
  nand_x4_sg U50521 ( .A(n28082), .B(n28156), .X(n28073) );
  nand_x1_sg U50522 ( .A(n28081), .B(n28080), .X(n28156) );
  nand_x4_sg U50523 ( .A(n28070), .B(n28154), .X(n28061) );
  nand_x1_sg U50524 ( .A(n28067), .B(n28069), .X(n28154) );
  nand_x4_sg U50525 ( .A(n28058), .B(n28152), .X(n28049) );
  nand_x1_sg U50526 ( .A(n28055), .B(n28057), .X(n28152) );
  nand_x4_sg U50527 ( .A(n28046), .B(n28150), .X(n28037) );
  nand_x1_sg U50528 ( .A(n28043), .B(n28045), .X(n28150) );
  nand_x4_sg U50529 ( .A(n28040), .B(n28149), .X(n28132) );
  nand_x1_sg U50530 ( .A(n28037), .B(n28039), .X(n28149) );
  inv_x2_sg U50531 ( .A(n27909), .X(n43766) );
  nor_x1_sg U50532 ( .A(n54036), .B(n28136), .X(n27909) );
  nand_x4_sg U50533 ( .A(n18062), .B(n54009), .X(n28018) );
  inv_x1_sg U50534 ( .A(n18061), .X(n54009) );
  nand_x4_sg U50535 ( .A(n18826), .B(n54141), .X(n28252) );
  inv_x1_sg U50536 ( .A(n18825), .X(n54141) );
  nand_x4_sg U50537 ( .A(n28349), .B(n28433), .X(n28342) );
  nand_x1_sg U50538 ( .A(n28346), .B(n28348), .X(n28433) );
  nand_x4_sg U50539 ( .A(n28339), .B(n28431), .X(n28330) );
  nand_x1_sg U50540 ( .A(n28336), .B(n28338), .X(n28431) );
  nand_x4_sg U50541 ( .A(n28327), .B(n28429), .X(n28318) );
  nand_x1_sg U50542 ( .A(n28324), .B(n28326), .X(n28429) );
  nand_x4_sg U50543 ( .A(n28321), .B(n28428), .X(n28411) );
  nand_x1_sg U50544 ( .A(n28318), .B(n28320), .X(n28428) );
  inv_x2_sg U50545 ( .A(n28188), .X(n43806) );
  nor_x1_sg U50546 ( .A(n54317), .B(n28415), .X(n28188) );
  nand_x4_sg U50547 ( .A(n18834), .B(n54291), .X(n28298) );
  inv_x1_sg U50548 ( .A(n18833), .X(n54291) );
  inv_x1_sg U50549 ( .A(n28637), .X(n54391) );
  nand_x4_sg U50550 ( .A(n28640), .B(n28714), .X(n28631) );
  nand_x1_sg U50551 ( .A(n28639), .B(n28638), .X(n28714) );
  nand_x4_sg U50552 ( .A(n28628), .B(n28712), .X(n28619) );
  nand_x1_sg U50553 ( .A(n28625), .B(n28627), .X(n28712) );
  nand_x4_sg U50554 ( .A(n28616), .B(n28710), .X(n28607) );
  nand_x1_sg U50555 ( .A(n28613), .B(n28615), .X(n28710) );
  nand_x4_sg U50556 ( .A(n28604), .B(n28708), .X(n28595) );
  nand_x1_sg U50557 ( .A(n28601), .B(n28603), .X(n28708) );
  nand_x4_sg U50558 ( .A(n28598), .B(n28707), .X(n28690) );
  nand_x1_sg U50559 ( .A(n28595), .B(n28597), .X(n28707) );
  inv_x2_sg U50560 ( .A(n28467), .X(n44161) );
  nor_x1_sg U50561 ( .A(n54601), .B(n28694), .X(n28467) );
  nand_x4_sg U50562 ( .A(n19607), .B(n54574), .X(n28576) );
  inv_x1_sg U50563 ( .A(n19606), .X(n54574) );
  nand_x4_sg U50564 ( .A(n28918), .B(n28992), .X(n28909) );
  nand_x1_sg U50565 ( .A(n28917), .B(n28916), .X(n28992) );
  nand_x4_sg U50566 ( .A(n20371), .B(n54706), .X(n28810) );
  inv_x1_sg U50567 ( .A(n20370), .X(n54706) );
  nand_x4_sg U50568 ( .A(n28906), .B(n28990), .X(n28899) );
  nand_x1_sg U50569 ( .A(n28903), .B(n28905), .X(n28990) );
  nand_x4_sg U50570 ( .A(n28896), .B(n28988), .X(n28887) );
  nand_x1_sg U50571 ( .A(n28893), .B(n28895), .X(n28988) );
  nand_x4_sg U50572 ( .A(n28884), .B(n28986), .X(n28875) );
  nand_x1_sg U50573 ( .A(n28881), .B(n28883), .X(n28986) );
  nand_x4_sg U50574 ( .A(n28878), .B(n28985), .X(n28968) );
  nand_x1_sg U50575 ( .A(n28875), .B(n28877), .X(n28985) );
  inv_x2_sg U50576 ( .A(n28746), .X(n43851) );
  nor_x1_sg U50577 ( .A(n54885), .B(n28972), .X(n28746) );
  nand_x4_sg U50578 ( .A(n20379), .B(n54859), .X(n28856) );
  inv_x1_sg U50579 ( .A(n20378), .X(n54859) );
  inv_x1_sg U50580 ( .A(n29198), .X(n54959) );
  nand_x4_sg U50581 ( .A(n29201), .B(n29275), .X(n29192) );
  nand_x1_sg U50582 ( .A(n29200), .B(n29199), .X(n29275) );
  nand_x4_sg U50583 ( .A(n29189), .B(n29273), .X(n29180) );
  nand_x1_sg U50584 ( .A(n29186), .B(n29188), .X(n29273) );
  nand_x4_sg U50585 ( .A(n29177), .B(n29271), .X(n29168) );
  nand_x1_sg U50586 ( .A(n29174), .B(n29176), .X(n29271) );
  nand_x4_sg U50587 ( .A(n29165), .B(n29269), .X(n29156) );
  nand_x1_sg U50588 ( .A(n29162), .B(n29164), .X(n29269) );
  nand_x4_sg U50589 ( .A(n29159), .B(n29268), .X(n29251) );
  nand_x1_sg U50590 ( .A(n29156), .B(n29158), .X(n29268) );
  inv_x2_sg U50591 ( .A(n29026), .X(n43787) );
  nor_x1_sg U50592 ( .A(n55169), .B(n29255), .X(n29026) );
  nand_x4_sg U50593 ( .A(n21151), .B(n55142), .X(n29135) );
  inv_x1_sg U50594 ( .A(n21150), .X(n55142) );
  nand_x4_sg U50595 ( .A(n21916), .B(n55274), .X(n29371) );
  inv_x1_sg U50596 ( .A(n21915), .X(n55274) );
  nand_x4_sg U50597 ( .A(n29445), .B(n29547), .X(n29436) );
  nand_x1_sg U50598 ( .A(n29442), .B(n29444), .X(n29547) );
  nand_x4_sg U50599 ( .A(n29439), .B(n29546), .X(n29529) );
  nand_x1_sg U50600 ( .A(n29436), .B(n29438), .X(n29546) );
  inv_x2_sg U50601 ( .A(n29307), .X(n44159) );
  nor_x1_sg U50602 ( .A(n55453), .B(n29533), .X(n29307) );
  nand_x4_sg U50603 ( .A(n21924), .B(n55427), .X(n29417) );
  inv_x1_sg U50604 ( .A(n21923), .X(n55427) );
  nand_x1_sg U50605 ( .A(n46600), .B(n21968), .X(n21967) );
  nand_x4_sg U50606 ( .A(n50958), .B(n22513), .X(n21941) );
  inv_x1_sg U50607 ( .A(n22515), .X(n50958) );
  nand_x1_sg U50608 ( .A(n21968), .B(n44100), .X(n22513) );
  nand_x1_sg U50609 ( .A(n46607), .B(n9388), .X(n9387) );
  nand_x1_sg U50610 ( .A(n46600), .B(n9454), .X(n9453) );
  nand_x1_sg U50611 ( .A(n50866), .B(n46608), .X(n9450) );
  nand_x1_sg U50612 ( .A(n46600), .B(n9503), .X(n9502) );
  nand_x1_sg U50613 ( .A(n50823), .B(n46608), .X(n9499) );
  nand_x1_sg U50614 ( .A(n46600), .B(n9552), .X(n9551) );
  nand_x1_sg U50615 ( .A(n50779), .B(n46608), .X(n9548) );
  nand_x1_sg U50616 ( .A(n46600), .B(n9600), .X(n9599) );
  nand_x1_sg U50617 ( .A(n50733), .B(n46608), .X(n9596) );
  nand_x1_sg U50618 ( .A(n46600), .B(n9648), .X(n9647) );
  nand_x1_sg U50619 ( .A(n50687), .B(n46608), .X(n9644) );
  nand_x1_sg U50620 ( .A(n50642), .B(n46608), .X(n9692) );
  nand_x1_sg U50621 ( .A(n46600), .B(n9743), .X(n9742) );
  nand_x1_sg U50622 ( .A(n50596), .B(n46608), .X(n9739) );
  nand_x1_sg U50623 ( .A(n46600), .B(n9791), .X(n9790) );
  nand_x1_sg U50624 ( .A(n50550), .B(n46608), .X(n9787) );
  nand_x1_sg U50625 ( .A(n46600), .B(n9839), .X(n9838) );
  nand_x1_sg U50626 ( .A(n50505), .B(n46608), .X(n9835) );
  nand_x1_sg U50627 ( .A(n46600), .B(n9887), .X(n9886) );
  nand_x1_sg U50628 ( .A(n50459), .B(n46608), .X(n9883) );
  nand_x1_sg U50629 ( .A(n46600), .B(n9935), .X(n9934) );
  nand_x1_sg U50630 ( .A(n46600), .B(n9984), .X(n9983) );
  nand_x1_sg U50631 ( .A(n46600), .B(n10032), .X(n10031) );
  nand_x1_sg U50632 ( .A(n46600), .B(n10081), .X(n10080) );
  nand_x1_sg U50633 ( .A(n46600), .B(n10130), .X(n10129) );
  nor_x1_sg U50634 ( .A(n10211), .B(n10212), .X(n10209) );
  nand_x1_sg U50635 ( .A(n46600), .B(n10220), .X(n10219) );
  nand_x1_sg U50636 ( .A(n46600), .B(n50116), .X(n10275) );
  inv_x1_sg U50637 ( .A(n10276), .X(n50116) );
  inv_x1_sg U50638 ( .A(n10251), .X(n55466) );
  inv_x1_sg U50639 ( .A(n10259), .X(n55463) );
  nand_x1_sg U50640 ( .A(n46598), .B(n50112), .X(n10271) );
  nand_x1_sg U50641 ( .A(n50109), .B(n46608), .X(n10270) );
  inv_x1_sg U50642 ( .A(n10272), .X(n50112) );
  nand_x2_sg U50643 ( .A(n10291), .B(n10292), .X(n10289) );
  inv_x2_sg U50644 ( .A(n10297), .X(n44139) );
  nor_x1_sg U50645 ( .A(n10398), .B(n51274), .X(n10297) );
  inv_x2_sg U50646 ( .A(n10296), .X(n43772) );
  nor_x1_sg U50647 ( .A(n51262), .B(n10391), .X(n10296) );
  nand_x2_sg U50648 ( .A(n42605), .B(n10413), .X(n10304) );
  nand_x1_sg U50649 ( .A(n10414), .B(n10415), .X(n10413) );
  inv_x1_sg U50650 ( .A(n10304), .X(n51296) );
  nand_x2_sg U50651 ( .A(n10386), .B(n10429), .X(n10308) );
  nand_x1_sg U50652 ( .A(n10430), .B(n10431), .X(n10429) );
  inv_x1_sg U50653 ( .A(n10308), .X(n51312) );
  nand_x1_sg U50654 ( .A(n51313), .B(n51327), .X(n10449) );
  inv_x1_sg U50655 ( .A(n10450), .X(n51313) );
  inv_x2_sg U50656 ( .A(n10328), .X(n51404) );
  nor_x1_sg U50657 ( .A(n51403), .B(n10557), .X(n10328) );
  inv_x1_sg U50658 ( .A(n51404), .X(n44356) );
  nand_x1_sg U50659 ( .A(n51440), .B(n10377), .X(n10624) );
  inv_x1_sg U50660 ( .A(n10376), .X(n51440) );
  nand_x1_sg U50661 ( .A(n51495), .B(n10717), .X(n10714) );
  inv_x1_sg U50662 ( .A(n10716), .X(n51495) );
  inv_x1_sg U50663 ( .A(n10371), .X(n51497) );
  inv_x1_sg U50664 ( .A(n10367), .X(n51521) );
  nand_x1_sg U50665 ( .A(n10369), .B(n10368), .X(n10366) );
  nand_x2_sg U50666 ( .A(n11059), .B(n51544), .X(n11057) );
  inv_x1_sg U50667 ( .A(n11060), .X(n51544) );
  inv_x1_sg U50668 ( .A(n11167), .X(n51553) );
  inv_x2_sg U50669 ( .A(n11064), .X(n44684) );
  nor_x1_sg U50670 ( .A(n11062), .B(n51546), .X(n11064) );
  nand_x2_sg U50671 ( .A(n42617), .B(n11185), .X(n11072) );
  nand_x1_sg U50672 ( .A(n11186), .B(n11187), .X(n11185) );
  inv_x1_sg U50673 ( .A(n11072), .X(n51578) );
  nand_x2_sg U50674 ( .A(n11153), .B(n11203), .X(n11076) );
  inv_x1_sg U50675 ( .A(n11076), .X(n51592) );
  nand_x1_sg U50676 ( .A(n51593), .B(n51602), .X(n11224) );
  inv_x1_sg U50677 ( .A(n11225), .X(n51593) );
  inv_x2_sg U50678 ( .A(n11096), .X(n51681) );
  nor_x1_sg U50679 ( .A(n51680), .B(n11330), .X(n11096) );
  inv_x1_sg U50680 ( .A(n51681), .X(n44355) );
  nand_x1_sg U50681 ( .A(n43276), .B(n11498), .X(n11495) );
  inv_x1_sg U50682 ( .A(n11136), .X(n51802) );
  nand_x2_sg U50683 ( .A(n11842), .B(n11843), .X(n11840) );
  inv_x2_sg U50684 ( .A(n11847), .X(n43754) );
  nor_x1_sg U50685 ( .A(n51821), .B(n11941), .X(n11847) );
  nand_x2_sg U50686 ( .A(n11937), .B(n11963), .X(n11855) );
  nand_x1_sg U50687 ( .A(n11964), .B(n11965), .X(n11963) );
  nand_x1_sg U50688 ( .A(n51836), .B(n51842), .X(n11938) );
  inv_x1_sg U50689 ( .A(n11855), .X(n51857) );
  nand_x2_sg U50690 ( .A(n11936), .B(n11981), .X(n11859) );
  inv_x1_sg U50691 ( .A(n11859), .X(n51872) );
  nand_x1_sg U50692 ( .A(n51873), .B(n51883), .X(n12001) );
  inv_x1_sg U50693 ( .A(n12002), .X(n51873) );
  inv_x2_sg U50694 ( .A(n11879), .X(n51962) );
  nor_x1_sg U50695 ( .A(n51961), .B(n12110), .X(n11879) );
  inv_x1_sg U50696 ( .A(n51962), .X(n44354) );
  nand_x1_sg U50697 ( .A(n42378), .B(n12278), .X(n12275) );
  inv_x1_sg U50698 ( .A(n11919), .X(n52078) );
  nand_x2_sg U50699 ( .A(n12620), .B(n52101), .X(n12618) );
  inv_x1_sg U50700 ( .A(n12621), .X(n52101) );
  inv_x1_sg U50701 ( .A(n12728), .X(n52110) );
  inv_x2_sg U50702 ( .A(n12625), .X(n44682) );
  nor_x1_sg U50703 ( .A(n12623), .B(n52103), .X(n12625) );
  nand_x2_sg U50704 ( .A(n42615), .B(n12746), .X(n12633) );
  nand_x1_sg U50705 ( .A(n12747), .B(n12748), .X(n12746) );
  inv_x1_sg U50706 ( .A(n12633), .X(n52136) );
  nand_x2_sg U50707 ( .A(n12714), .B(n12764), .X(n12637) );
  inv_x1_sg U50708 ( .A(n12637), .X(n52150) );
  nand_x1_sg U50709 ( .A(n52151), .B(n52160), .X(n12785) );
  inv_x1_sg U50710 ( .A(n12786), .X(n52151) );
  inv_x2_sg U50711 ( .A(n12657), .X(n52237) );
  nor_x1_sg U50712 ( .A(n52236), .B(n12891), .X(n12657) );
  inv_x1_sg U50713 ( .A(n52237), .X(n44353) );
  nand_x1_sg U50714 ( .A(n43274), .B(n13059), .X(n13056) );
  inv_x1_sg U50715 ( .A(n12697), .X(n52356) );
  nand_x2_sg U50716 ( .A(n13404), .B(n13405), .X(n13402) );
  inv_x2_sg U50717 ( .A(n13409), .X(n43799) );
  nor_x1_sg U50718 ( .A(n52373), .B(n13503), .X(n13409) );
  nand_x2_sg U50719 ( .A(n13499), .B(n13524), .X(n13417) );
  nand_x1_sg U50720 ( .A(n13525), .B(n13526), .X(n13524) );
  nand_x1_sg U50721 ( .A(n52388), .B(n52394), .X(n13500) );
  inv_x1_sg U50722 ( .A(n13417), .X(n52409) );
  nand_x2_sg U50723 ( .A(n13498), .B(n13542), .X(n13421) );
  inv_x1_sg U50724 ( .A(n13421), .X(n52424) );
  nand_x1_sg U50725 ( .A(n52425), .B(n52434), .X(n13562) );
  nand_x1_sg U50726 ( .A(n13564), .B(n13563), .X(n13561) );
  inv_x1_sg U50727 ( .A(n13563), .X(n52425) );
  inv_x2_sg U50728 ( .A(n13441), .X(n52514) );
  nor_x1_sg U50729 ( .A(n52513), .B(n13671), .X(n13441) );
  inv_x1_sg U50730 ( .A(n52514), .X(n44352) );
  nand_x1_sg U50731 ( .A(n43272), .B(n13839), .X(n13836) );
  inv_x1_sg U50732 ( .A(n13481), .X(n52631) );
  nand_x2_sg U50733 ( .A(n14183), .B(n14184), .X(n14181) );
  inv_x2_sg U50734 ( .A(n14188), .X(n43801) );
  nor_x1_sg U50735 ( .A(n52650), .B(n14283), .X(n14188) );
  inv_x2_sg U50736 ( .A(n14189), .X(n44404) );
  nor_x1_sg U50737 ( .A(n14290), .B(n52663), .X(n14189) );
  nand_x2_sg U50738 ( .A(n14279), .B(n14305), .X(n14196) );
  nand_x1_sg U50739 ( .A(n14306), .B(n14307), .X(n14305) );
  inv_x1_sg U50740 ( .A(n14196), .X(n52686) );
  nand_x2_sg U50741 ( .A(n14278), .B(n14321), .X(n14200) );
  nand_x1_sg U50742 ( .A(n14322), .B(n14323), .X(n14321) );
  inv_x1_sg U50743 ( .A(n14200), .X(n52701) );
  nand_x1_sg U50744 ( .A(n52702), .B(n52717), .X(n14341) );
  inv_x1_sg U50745 ( .A(n14342), .X(n52702) );
  inv_x2_sg U50746 ( .A(n14220), .X(n52793) );
  nor_x1_sg U50747 ( .A(n52792), .B(n14449), .X(n14220) );
  inv_x1_sg U50748 ( .A(n52793), .X(n44351) );
  nand_x1_sg U50749 ( .A(n52829), .B(n14269), .X(n14516) );
  inv_x1_sg U50750 ( .A(n14268), .X(n52829) );
  nand_x1_sg U50751 ( .A(n43294), .B(n14609), .X(n14606) );
  inv_x2_sg U50752 ( .A(n14241), .X(n44692) );
  nor_x1_sg U50753 ( .A(n14655), .B(n14656), .X(n14241) );
  inv_x1_sg U50754 ( .A(n14260), .X(n52912) );
  nand_x1_sg U50755 ( .A(n46576), .B(n15726), .X(n15725) );
  nand_x2_sg U50756 ( .A(n14953), .B(n52935), .X(n14951) );
  inv_x1_sg U50757 ( .A(n14954), .X(n52935) );
  inv_x1_sg U50758 ( .A(n15061), .X(n52944) );
  inv_x2_sg U50759 ( .A(n14958), .X(n44680) );
  nor_x1_sg U50760 ( .A(n14956), .B(n52937), .X(n14958) );
  nand_x2_sg U50761 ( .A(n42613), .B(n15079), .X(n14966) );
  nand_x1_sg U50762 ( .A(n15080), .B(n15081), .X(n15079) );
  inv_x1_sg U50763 ( .A(n14966), .X(n52970) );
  nand_x2_sg U50764 ( .A(n15047), .B(n15097), .X(n14970) );
  inv_x1_sg U50765 ( .A(n14970), .X(n52984) );
  nand_x1_sg U50766 ( .A(n52985), .B(n52994), .X(n15118) );
  inv_x1_sg U50767 ( .A(n15119), .X(n52985) );
  inv_x2_sg U50768 ( .A(n14990), .X(n53071) );
  nor_x1_sg U50769 ( .A(n53070), .B(n15224), .X(n14990) );
  inv_x1_sg U50770 ( .A(n53071), .X(n44350) );
  nand_x1_sg U50771 ( .A(n43270), .B(n15392), .X(n15389) );
  inv_x1_sg U50772 ( .A(n15030), .X(n53190) );
  nand_x2_sg U50773 ( .A(n15737), .B(n15738), .X(n15735) );
  inv_x2_sg U50774 ( .A(n15742), .X(n43770) );
  nor_x1_sg U50775 ( .A(n53209), .B(n15836), .X(n15742) );
  nand_x2_sg U50776 ( .A(n15832), .B(n15858), .X(n15750) );
  nand_x1_sg U50777 ( .A(n15859), .B(n15860), .X(n15858) );
  nand_x1_sg U50778 ( .A(n53224), .B(n43140), .X(n15833) );
  inv_x1_sg U50779 ( .A(n15750), .X(n53243) );
  nand_x2_sg U50780 ( .A(n15831), .B(n15876), .X(n15754) );
  inv_x1_sg U50781 ( .A(n15754), .X(n53259) );
  nand_x1_sg U50782 ( .A(n53260), .B(n53270), .X(n15896) );
  inv_x1_sg U50783 ( .A(n15897), .X(n53260) );
  inv_x2_sg U50784 ( .A(n15774), .X(n53350) );
  nor_x1_sg U50785 ( .A(n53349), .B(n16005), .X(n15774) );
  inv_x1_sg U50786 ( .A(n53350), .X(n44349) );
  nand_x1_sg U50787 ( .A(n43266), .B(n16173), .X(n16170) );
  inv_x1_sg U50788 ( .A(n15817), .X(n53445) );
  inv_x1_sg U50789 ( .A(n15813), .X(n53470) );
  nand_x1_sg U50790 ( .A(n15815), .B(n15814), .X(n15812) );
  nand_x2_sg U50791 ( .A(n16519), .B(n53493), .X(n16517) );
  inv_x1_sg U50792 ( .A(n16520), .X(n53493) );
  inv_x1_sg U50793 ( .A(n16627), .X(n53502) );
  inv_x2_sg U50794 ( .A(n16524), .X(n44678) );
  nor_x1_sg U50795 ( .A(n16522), .B(n53495), .X(n16524) );
  nand_x2_sg U50796 ( .A(n42611), .B(n16645), .X(n16532) );
  nand_x1_sg U50797 ( .A(n16646), .B(n16647), .X(n16645) );
  inv_x1_sg U50798 ( .A(n16532), .X(n53528) );
  nand_x2_sg U50799 ( .A(n16613), .B(n16663), .X(n16536) );
  inv_x1_sg U50800 ( .A(n16536), .X(n53542) );
  nand_x1_sg U50801 ( .A(n53543), .B(n53552), .X(n16684) );
  inv_x1_sg U50802 ( .A(n16685), .X(n53543) );
  inv_x2_sg U50803 ( .A(n16556), .X(n53629) );
  nor_x1_sg U50804 ( .A(n53628), .B(n16790), .X(n16556) );
  inv_x1_sg U50805 ( .A(n53629), .X(n44348) );
  nand_x1_sg U50806 ( .A(n43268), .B(n16958), .X(n16955) );
  inv_x1_sg U50807 ( .A(n16596), .X(n53748) );
  nand_x2_sg U50808 ( .A(n17302), .B(n17303), .X(n17300) );
  inv_x1_sg U50809 ( .A(n17411), .X(n53780) );
  nand_x2_sg U50810 ( .A(n42624), .B(n17426), .X(n17315) );
  nand_x1_sg U50811 ( .A(n17427), .B(n17428), .X(n17426) );
  inv_x2_sg U50812 ( .A(n17316), .X(n53795) );
  nand_x1_sg U50813 ( .A(n53794), .B(n17399), .X(n17316) );
  inv_x1_sg U50814 ( .A(n53795), .X(n45420) );
  inv_x1_sg U50815 ( .A(n17315), .X(n53805) );
  nand_x2_sg U50816 ( .A(n17397), .B(n17444), .X(n17319) );
  nand_x1_sg U50817 ( .A(n17445), .B(n53819), .X(n17444) );
  inv_x1_sg U50818 ( .A(n17319), .X(n53820) );
  nand_x1_sg U50819 ( .A(n53821), .B(n53831), .X(n17464) );
  inv_x1_sg U50820 ( .A(n17465), .X(n53821) );
  inv_x2_sg U50821 ( .A(n17339), .X(n53913) );
  nor_x1_sg U50822 ( .A(n53912), .B(n17569), .X(n17339) );
  inv_x1_sg U50823 ( .A(n53913), .X(n44347) );
  nand_x1_sg U50824 ( .A(n53949), .B(n17388), .X(n17637) );
  inv_x1_sg U50825 ( .A(n17387), .X(n53949) );
  nand_x1_sg U50826 ( .A(n43292), .B(n17730), .X(n17727) );
  inv_x2_sg U50827 ( .A(n17360), .X(n44690) );
  nor_x1_sg U50828 ( .A(n17776), .B(n17777), .X(n17360) );
  inv_x1_sg U50829 ( .A(n17379), .X(n54032) );
  nand_x2_sg U50830 ( .A(n18074), .B(n18075), .X(n18072) );
  inv_x2_sg U50831 ( .A(n18080), .X(n44402) );
  nor_x1_sg U50832 ( .A(n18179), .B(n54060), .X(n18080) );
  inv_x2_sg U50833 ( .A(n18079), .X(n43972) );
  nor_x1_sg U50834 ( .A(n54051), .B(n18173), .X(n18079) );
  inv_x2_sg U50835 ( .A(n18084), .X(n43997) );
  nor_x1_sg U50836 ( .A(n18185), .B(n18186), .X(n18084) );
  nand_x2_sg U50837 ( .A(n18169), .B(n18193), .X(n18087) );
  nand_x1_sg U50838 ( .A(n18194), .B(n18195), .X(n18193) );
  inv_x1_sg U50839 ( .A(n18087), .X(n54087) );
  nand_x2_sg U50840 ( .A(n18168), .B(n18210), .X(n18091) );
  nand_x1_sg U50841 ( .A(n18211), .B(n18212), .X(n18210) );
  inv_x1_sg U50842 ( .A(n18091), .X(n54102) );
  inv_x1_sg U50843 ( .A(n18231), .X(n54103) );
  inv_x2_sg U50844 ( .A(n18251), .X(n44720) );
  inv_x2_sg U50845 ( .A(n18111), .X(n54193) );
  nor_x1_sg U50846 ( .A(n54192), .B(n18339), .X(n18111) );
  inv_x1_sg U50847 ( .A(n54193), .X(n44346) );
  nand_x1_sg U50848 ( .A(n54234), .B(n18159), .X(n18406) );
  inv_x1_sg U50849 ( .A(n18158), .X(n54234) );
  nand_x1_sg U50850 ( .A(n42376), .B(n18499), .X(n18496) );
  inv_x1_sg U50851 ( .A(n18150), .X(n54313) );
  nand_x2_sg U50852 ( .A(n18847), .B(n18848), .X(n18845) );
  inv_x1_sg U50853 ( .A(n18956), .X(n54345) );
  nand_x2_sg U50854 ( .A(n42622), .B(n18971), .X(n18860) );
  nand_x1_sg U50855 ( .A(n18972), .B(n18973), .X(n18971) );
  inv_x2_sg U50856 ( .A(n18861), .X(n54360) );
  nand_x1_sg U50857 ( .A(n54359), .B(n18944), .X(n18861) );
  inv_x1_sg U50858 ( .A(n54360), .X(n45419) );
  inv_x1_sg U50859 ( .A(n18860), .X(n54370) );
  nand_x2_sg U50860 ( .A(n18942), .B(n18989), .X(n18864) );
  nand_x1_sg U50861 ( .A(n18990), .B(n54384), .X(n18989) );
  inv_x1_sg U50862 ( .A(n18864), .X(n54385) );
  nand_x1_sg U50863 ( .A(n54386), .B(n54396), .X(n19009) );
  inv_x1_sg U50864 ( .A(n19010), .X(n54386) );
  inv_x2_sg U50865 ( .A(n18884), .X(n54478) );
  nor_x1_sg U50866 ( .A(n54477), .B(n19114), .X(n18884) );
  inv_x1_sg U50867 ( .A(n54478), .X(n44345) );
  nand_x1_sg U50868 ( .A(n54514), .B(n18933), .X(n19182) );
  inv_x1_sg U50869 ( .A(n18932), .X(n54514) );
  nand_x1_sg U50870 ( .A(n43290), .B(n19275), .X(n19272) );
  inv_x2_sg U50871 ( .A(n18905), .X(n44688) );
  nor_x1_sg U50872 ( .A(n19321), .B(n19322), .X(n18905) );
  inv_x1_sg U50873 ( .A(n18924), .X(n54597) );
  nand_x2_sg U50874 ( .A(n19619), .B(n19620), .X(n19617) );
  nand_x2_sg U50875 ( .A(n42609), .B(n19740), .X(n19632) );
  nand_x1_sg U50876 ( .A(n19741), .B(n19742), .X(n19740) );
  inv_x1_sg U50877 ( .A(n19632), .X(n54650) );
  nand_x2_sg U50878 ( .A(n19713), .B(n19756), .X(n19636) );
  nand_x1_sg U50879 ( .A(n19757), .B(n19758), .X(n19756) );
  inv_x1_sg U50880 ( .A(n19636), .X(n54666) );
  nand_x1_sg U50881 ( .A(n54667), .B(n54681), .X(n19776) );
  inv_x1_sg U50882 ( .A(n19777), .X(n54667) );
  inv_x2_sg U50883 ( .A(n19656), .X(n54760) );
  nor_x1_sg U50884 ( .A(n54759), .B(n19884), .X(n19656) );
  inv_x1_sg U50885 ( .A(n54760), .X(n44344) );
  nand_x1_sg U50886 ( .A(n54799), .B(n19704), .X(n19951) );
  inv_x1_sg U50887 ( .A(n19703), .X(n54799) );
  nand_x1_sg U50888 ( .A(n42374), .B(n20044), .X(n20041) );
  inv_x1_sg U50889 ( .A(n19695), .X(n54881) );
  nand_x2_sg U50890 ( .A(n20391), .B(n20392), .X(n20389) );
  inv_x1_sg U50891 ( .A(n20500), .X(n54913) );
  nand_x2_sg U50892 ( .A(n42620), .B(n20515), .X(n20404) );
  nand_x1_sg U50893 ( .A(n20516), .B(n20517), .X(n20515) );
  inv_x2_sg U50894 ( .A(n20405), .X(n54928) );
  nand_x1_sg U50895 ( .A(n54927), .B(n20488), .X(n20405) );
  inv_x1_sg U50896 ( .A(n54928), .X(n45418) );
  inv_x1_sg U50897 ( .A(n20404), .X(n54938) );
  nand_x2_sg U50898 ( .A(n20486), .B(n20533), .X(n20408) );
  nand_x1_sg U50899 ( .A(n20534), .B(n54952), .X(n20533) );
  inv_x1_sg U50900 ( .A(n20408), .X(n54953) );
  nand_x1_sg U50901 ( .A(n54954), .B(n54964), .X(n20553) );
  inv_x1_sg U50902 ( .A(n20554), .X(n54954) );
  inv_x2_sg U50903 ( .A(n20428), .X(n55046) );
  nor_x1_sg U50904 ( .A(n55045), .B(n20658), .X(n20428) );
  inv_x1_sg U50905 ( .A(n55046), .X(n44343) );
  nand_x1_sg U50906 ( .A(n55082), .B(n20477), .X(n20726) );
  inv_x1_sg U50907 ( .A(n20476), .X(n55082) );
  nand_x1_sg U50908 ( .A(n43288), .B(n20819), .X(n20816) );
  inv_x2_sg U50909 ( .A(n20449), .X(n44686) );
  nor_x1_sg U50910 ( .A(n20865), .B(n20866), .X(n20449) );
  inv_x1_sg U50911 ( .A(n20468), .X(n55165) );
  nand_x2_sg U50912 ( .A(n21164), .B(n21165), .X(n21162) );
  inv_x2_sg U50913 ( .A(n21170), .X(n44137) );
  nor_x1_sg U50914 ( .A(n21270), .B(n55196), .X(n21170) );
  nand_x2_sg U50915 ( .A(n42607), .B(n21285), .X(n21177) );
  nand_x1_sg U50916 ( .A(n21286), .B(n21287), .X(n21285) );
  inv_x1_sg U50917 ( .A(n21177), .X(n55218) );
  nand_x2_sg U50918 ( .A(n21258), .B(n21301), .X(n21181) );
  nand_x1_sg U50919 ( .A(n21302), .B(n21303), .X(n21301) );
  inv_x1_sg U50920 ( .A(n21181), .X(n55234) );
  nand_x1_sg U50921 ( .A(n55235), .B(n55249), .X(n21321) );
  inv_x1_sg U50922 ( .A(n21322), .X(n55235) );
  inv_x2_sg U50923 ( .A(n21201), .X(n55328) );
  nor_x1_sg U50924 ( .A(n55327), .B(n21429), .X(n21201) );
  inv_x1_sg U50925 ( .A(n55328), .X(n44342) );
  nand_x1_sg U50926 ( .A(n55367), .B(n21249), .X(n21496) );
  inv_x1_sg U50927 ( .A(n21248), .X(n55367) );
  nand_x1_sg U50928 ( .A(n42372), .B(n21589), .X(n21586) );
  inv_x1_sg U50929 ( .A(n21240), .X(n55449) );
  nand_x1_sg U50930 ( .A(n9403), .B(n29631), .X(n29630) );
  nand_x4_sg U50931 ( .A(n50099), .B(n30179), .X(n29594) );
  inv_x1_sg U50932 ( .A(n30181), .X(n50099) );
  nand_x1_sg U50933 ( .A(n29631), .B(n44098), .X(n30179) );
  nand_x1_sg U50934 ( .A(n46600), .B(n24562), .X(n24561) );
  nand_x1_sg U50935 ( .A(n50007), .B(n46608), .X(n24558) );
  nand_x1_sg U50936 ( .A(n46600), .B(n24611), .X(n24610) );
  nand_x1_sg U50937 ( .A(n49964), .B(n46608), .X(n24607) );
  nand_x1_sg U50938 ( .A(n46600), .B(n24660), .X(n24659) );
  nand_x1_sg U50939 ( .A(n49920), .B(n46608), .X(n24656) );
  nand_x1_sg U50940 ( .A(n46600), .B(n24708), .X(n24707) );
  nand_x1_sg U50941 ( .A(n49874), .B(n46608), .X(n24704) );
  nand_x1_sg U50942 ( .A(n46600), .B(n24756), .X(n24755) );
  nand_x1_sg U50943 ( .A(n49828), .B(n46608), .X(n24752) );
  nand_x1_sg U50944 ( .A(n49783), .B(n46608), .X(n24800) );
  nand_x1_sg U50945 ( .A(n46600), .B(n24851), .X(n24850) );
  nand_x1_sg U50946 ( .A(n49737), .B(n46608), .X(n24847) );
  nand_x1_sg U50947 ( .A(n46600), .B(n24899), .X(n24898) );
  nand_x1_sg U50948 ( .A(n49691), .B(n46608), .X(n24895) );
  nand_x1_sg U50949 ( .A(n46600), .B(n24947), .X(n24946) );
  nand_x1_sg U50950 ( .A(n49646), .B(n46608), .X(n24943) );
  nand_x1_sg U50951 ( .A(n46600), .B(n24995), .X(n24994) );
  nand_x1_sg U50952 ( .A(n49600), .B(n46608), .X(n24991) );
  nand_x1_sg U50953 ( .A(n46600), .B(n25043), .X(n25042) );
  nand_x1_sg U50954 ( .A(n46600), .B(n25092), .X(n25091) );
  nand_x1_sg U50955 ( .A(n46600), .B(n25140), .X(n25139) );
  nand_x1_sg U50956 ( .A(n46600), .B(n25189), .X(n25188) );
  nand_x1_sg U50957 ( .A(n46600), .B(n25238), .X(n25237) );
  nor_x1_sg U50958 ( .A(n25319), .B(n25320), .X(n25317) );
  nand_x1_sg U50959 ( .A(n46600), .B(n25328), .X(n25327) );
  inv_x1_sg U50960 ( .A(n31251), .X(n49275) );
  nand_x1_sg U50961 ( .A(n49257), .B(n46600), .X(n25381) );
  inv_x1_sg U50962 ( .A(n25382), .X(n49257) );
  inv_x1_sg U50963 ( .A(n25366), .X(n55464) );
  inv_x1_sg U50964 ( .A(n25359), .X(n55467) );
  nand_x1_sg U50965 ( .A(n49253), .B(n9399), .X(n25377) );
  nand_x1_sg U50966 ( .A(n49250), .B(n46610), .X(n25376) );
  inv_x1_sg U50967 ( .A(n25378), .X(n49253) );
  nand_x1_sg U50968 ( .A(n10490), .B(n46231), .X(n25438) );
  nand_x1_sg U50969 ( .A(n46232), .B(n25437), .X(n25436) );
  nand_x1_sg U50970 ( .A(n46231), .B(n46559), .X(n25445) );
  inv_x1_sg U50971 ( .A(n25443), .X(n51526) );
  nand_x1_sg U50972 ( .A(n46231), .B(n25459), .X(n25460) );
  nand_x1_sg U50973 ( .A(n51374), .B(n25458), .X(n25457) );
  inv_x1_sg U50974 ( .A(n25459), .X(n51374) );
  nand_x1_sg U50975 ( .A(n46231), .B(n46555), .X(n25474) );
  nand_x1_sg U50976 ( .A(n46554), .B(n25473), .X(n25472) );
  nand_x1_sg U50977 ( .A(n46231), .B(n10843), .X(n25488) );
  inv_x2_sg U50978 ( .A(n25395), .X(n44157) );
  nor_x1_sg U50979 ( .A(n51524), .B(n25620), .X(n25395) );
  inv_x2_sg U50980 ( .A(n25632), .X(n44248) );
  nor_x1_sg U50981 ( .A(n25664), .B(n25665), .X(n25632) );
  nand_x4_sg U50982 ( .A(n11045), .B(n51500), .X(n25505) );
  inv_x1_sg U50983 ( .A(n11044), .X(n51500) );
  nand_x1_sg U50984 ( .A(n46201), .B(n46229), .X(n25717) );
  nand_x1_sg U50985 ( .A(n46230), .B(n25716), .X(n25715) );
  nand_x1_sg U50986 ( .A(n46229), .B(n11290), .X(n25724) );
  inv_x1_sg U50987 ( .A(n25722), .X(n51808) );
  nand_x1_sg U50988 ( .A(n46229), .B(n11394), .X(n25738) );
  nand_x1_sg U50989 ( .A(n51630), .B(n25737), .X(n25736) );
  nand_x1_sg U50990 ( .A(n46229), .B(n11515), .X(n25752) );
  nor_x2_sg U50991 ( .A(n25763), .B(n51738), .X(n25770) );
  nand_x1_sg U50992 ( .A(n12043), .B(n46227), .X(n25995) );
  nand_x1_sg U50993 ( .A(n46228), .B(n25994), .X(n25993) );
  nand_x1_sg U50994 ( .A(n46227), .B(n12070), .X(n26002) );
  inv_x1_sg U50995 ( .A(n26000), .X(n52084) );
  nand_x1_sg U50996 ( .A(n46227), .B(n12174), .X(n26016) );
  nand_x1_sg U50997 ( .A(n51911), .B(n26015), .X(n26014) );
  nand_x1_sg U50998 ( .A(n46227), .B(n12295), .X(n26030) );
  inv_x1_sg U50999 ( .A(n42515), .X(n52016) );
  nand_x1_sg U51000 ( .A(n43745), .B(n46225), .X(n26276) );
  nand_x1_sg U51001 ( .A(n46226), .B(n26275), .X(n26274) );
  nand_x1_sg U51002 ( .A(n46225), .B(n12851), .X(n26283) );
  inv_x1_sg U51003 ( .A(n26281), .X(n52362) );
  nand_x1_sg U51004 ( .A(n46225), .B(n12955), .X(n26297) );
  nand_x1_sg U51005 ( .A(n52187), .B(n26296), .X(n26295) );
  nand_x1_sg U51006 ( .A(n46225), .B(n13076), .X(n26311) );
  nand_x1_sg U51007 ( .A(n46225), .B(n13184), .X(n26325) );
  inv_x1_sg U51008 ( .A(n42513), .X(n52292) );
  nand_x1_sg U51009 ( .A(n46469), .B(n46223), .X(n26555) );
  nand_x1_sg U51010 ( .A(n46224), .B(n26554), .X(n26553) );
  nand_x1_sg U51011 ( .A(n46223), .B(n13631), .X(n26562) );
  inv_x1_sg U51012 ( .A(n26560), .X(n52637) );
  nand_x1_sg U51013 ( .A(n46223), .B(n13735), .X(n26576) );
  nand_x1_sg U51014 ( .A(n52463), .B(n26575), .X(n26574) );
  nand_x1_sg U51015 ( .A(n46223), .B(n13856), .X(n26590) );
  nand_x1_sg U51016 ( .A(n46223), .B(n13964), .X(n26604) );
  inv_x1_sg U51017 ( .A(n42511), .X(n52567) );
  nand_x1_sg U51018 ( .A(n46445), .B(n46221), .X(n26833) );
  nand_x1_sg U51019 ( .A(n46222), .B(n26832), .X(n26831) );
  nand_x1_sg U51020 ( .A(n46221), .B(n14411), .X(n26840) );
  inv_x1_sg U51021 ( .A(n26838), .X(n52918) );
  nand_x1_sg U51022 ( .A(n46221), .B(n14507), .X(n26854) );
  nand_x1_sg U51023 ( .A(n46221), .B(n14627), .X(n26868) );
  nand_x1_sg U51024 ( .A(n46221), .B(n14735), .X(n26882) );
  nand_x1_sg U51025 ( .A(n43746), .B(n46219), .X(n27112) );
  nand_x1_sg U51026 ( .A(n46220), .B(n27111), .X(n27110) );
  nand_x1_sg U51027 ( .A(n46219), .B(n15184), .X(n27119) );
  inv_x1_sg U51028 ( .A(n27117), .X(n53196) );
  nand_x1_sg U51029 ( .A(n46219), .B(n15288), .X(n27133) );
  nand_x1_sg U51030 ( .A(n53021), .B(n27132), .X(n27131) );
  nand_x1_sg U51031 ( .A(n46219), .B(n15409), .X(n27147) );
  nand_x1_sg U51032 ( .A(n46219), .B(n15517), .X(n27161) );
  inv_x1_sg U51033 ( .A(n42509), .X(n53126) );
  nand_x1_sg U51034 ( .A(n15938), .B(n46217), .X(n27392) );
  nand_x1_sg U51035 ( .A(n46218), .B(n27391), .X(n27390) );
  nand_x1_sg U51036 ( .A(n46217), .B(n15965), .X(n27399) );
  inv_x1_sg U51037 ( .A(n27397), .X(n53476) );
  nand_x1_sg U51038 ( .A(n46217), .B(n16069), .X(n27413) );
  nand_x1_sg U51039 ( .A(n46217), .B(n16190), .X(n27427) );
  nor_x2_sg U51040 ( .A(n27438), .B(n53408), .X(n27445) );
  nand_x1_sg U51041 ( .A(n43747), .B(n46215), .X(n27672) );
  nand_x1_sg U51042 ( .A(n46216), .B(n27671), .X(n27670) );
  nand_x1_sg U51043 ( .A(n46215), .B(n16750), .X(n27679) );
  inv_x1_sg U51044 ( .A(n27677), .X(n53754) );
  nand_x1_sg U51045 ( .A(n46215), .B(n16854), .X(n27693) );
  nand_x1_sg U51046 ( .A(n53579), .B(n27692), .X(n27691) );
  nand_x1_sg U51047 ( .A(n46215), .B(n16975), .X(n27707) );
  nand_x1_sg U51048 ( .A(n46215), .B(n17083), .X(n27721) );
  inv_x1_sg U51049 ( .A(n42507), .X(n53684) );
  nand_x1_sg U51050 ( .A(n53814), .B(n46213), .X(n27952) );
  nand_x1_sg U51051 ( .A(n46214), .B(n27951), .X(n27950) );
  nand_x1_sg U51052 ( .A(n46213), .B(n17524), .X(n27959) );
  inv_x1_sg U51053 ( .A(n27957), .X(n54038) );
  nand_x1_sg U51054 ( .A(n46213), .B(n17628), .X(n27973) );
  nand_x1_sg U51055 ( .A(n46213), .B(n17748), .X(n27987) );
  nand_x1_sg U51056 ( .A(n46213), .B(n17856), .X(n28001) );
  nand_x1_sg U51057 ( .A(n54097), .B(n46211), .X(n28231) );
  nand_x1_sg U51058 ( .A(n46212), .B(n28230), .X(n28229) );
  nand_x1_sg U51059 ( .A(n46211), .B(n18301), .X(n28238) );
  inv_x1_sg U51060 ( .A(n28236), .X(n54319) );
  nand_x1_sg U51061 ( .A(n46211), .B(n28252), .X(n28253) );
  nand_x1_sg U51062 ( .A(n54162), .B(n28251), .X(n28250) );
  inv_x1_sg U51063 ( .A(n28252), .X(n54162) );
  nand_x1_sg U51064 ( .A(n46211), .B(n18574), .X(n28267) );
  nand_x1_sg U51065 ( .A(n46211), .B(n18623), .X(n28281) );
  nand_x1_sg U51066 ( .A(n54379), .B(n46209), .X(n28510) );
  nand_x1_sg U51067 ( .A(n46210), .B(n28509), .X(n28508) );
  nand_x1_sg U51068 ( .A(n46209), .B(n19069), .X(n28517) );
  inv_x1_sg U51069 ( .A(n28515), .X(n54603) );
  nand_x1_sg U51070 ( .A(n46209), .B(n19173), .X(n28531) );
  nand_x1_sg U51071 ( .A(n46209), .B(n19293), .X(n28545) );
  nand_x1_sg U51072 ( .A(n46209), .B(n19401), .X(n28559) );
  nand_x1_sg U51073 ( .A(n19817), .B(n46207), .X(n28789) );
  nand_x1_sg U51074 ( .A(n46208), .B(n28788), .X(n28787) );
  nand_x1_sg U51075 ( .A(n46207), .B(n46287), .X(n28796) );
  inv_x1_sg U51076 ( .A(n28794), .X(n54887) );
  nand_x1_sg U51077 ( .A(n46207), .B(n28810), .X(n28811) );
  nand_x1_sg U51078 ( .A(n54728), .B(n28809), .X(n28808) );
  inv_x1_sg U51079 ( .A(n28810), .X(n54728) );
  nand_x1_sg U51080 ( .A(n46207), .B(n20229), .X(n28825) );
  nand_x1_sg U51081 ( .A(n46207), .B(n20169), .X(n28839) );
  nand_x1_sg U51082 ( .A(n54947), .B(n46205), .X(n29069) );
  nand_x1_sg U51083 ( .A(n46206), .B(n29068), .X(n29067) );
  nand_x1_sg U51084 ( .A(n46205), .B(n20613), .X(n29076) );
  inv_x1_sg U51085 ( .A(n29074), .X(n55171) );
  nand_x1_sg U51086 ( .A(n46205), .B(n20717), .X(n29090) );
  nand_x1_sg U51087 ( .A(n46205), .B(n20837), .X(n29104) );
  nand_x1_sg U51088 ( .A(n46205), .B(n20945), .X(n29118) );
  nand_x1_sg U51089 ( .A(n21362), .B(n46203), .X(n29350) );
  nand_x1_sg U51090 ( .A(n46204), .B(n29349), .X(n29348) );
  nand_x1_sg U51091 ( .A(n46203), .B(n46242), .X(n29357) );
  inv_x1_sg U51092 ( .A(n29355), .X(n55455) );
  nand_x1_sg U51093 ( .A(n46203), .B(n29371), .X(n29372) );
  nand_x1_sg U51094 ( .A(n55296), .B(n29370), .X(n29369) );
  inv_x1_sg U51095 ( .A(n29371), .X(n55296) );
  nand_x1_sg U51096 ( .A(n46203), .B(n21774), .X(n29386) );
  nand_x1_sg U51097 ( .A(n46203), .B(n21714), .X(n29400) );
  inv_x2_sg U51098 ( .A(n9049), .X(n43952) );
  nor_x1_sg U51099 ( .A(n40870), .B(n10285), .X(n9049) );
  nor_x1_sg U51100 ( .A(n10283), .B(n51261), .X(n10284) );
  nand_x1_sg U51101 ( .A(n10289), .B(n43872), .X(n10287) );
  inv_x1_sg U51102 ( .A(n10289), .X(n51268) );
  inv_x1_sg U51103 ( .A(n10299), .X(n51285) );
  nand_x1_sg U51104 ( .A(n51286), .B(n10304), .X(n10303) );
  inv_x1_sg U51105 ( .A(n10305), .X(n51286) );
  nand_x1_sg U51106 ( .A(n51297), .B(n10308), .X(n10307) );
  inv_x1_sg U51107 ( .A(n10309), .X(n51297) );
  inv_x1_sg U51108 ( .A(n10311), .X(n51328) );
  inv_x1_sg U51109 ( .A(n10319), .X(n51364) );
  nand_x1_sg U51110 ( .A(n10327), .B(n51404), .X(n10326) );
  inv_x1_sg U51111 ( .A(n10336), .X(n51441) );
  inv_x2_sg U51112 ( .A(n9043), .X(n44400) );
  nor_x1_sg U51113 ( .A(n10339), .B(n51473), .X(n9043) );
  inv_x1_sg U51114 ( .A(n10344), .X(n51496) );
  inv_x1_sg U51115 ( .A(n10348), .X(n51510) );
  inv_x1_sg U51116 ( .A(n10352), .X(n51522) );
  nand_x1_sg U51117 ( .A(n11057), .B(n44018), .X(n11055) );
  nand_x1_sg U51118 ( .A(n51537), .B(n51545), .X(n11056) );
  inv_x1_sg U51119 ( .A(n11057), .X(n51545) );
  inv_x1_sg U51120 ( .A(n11066), .X(n51554) );
  nand_x1_sg U51121 ( .A(n51566), .B(n11072), .X(n11071) );
  inv_x1_sg U51122 ( .A(n11073), .X(n51566) );
  nand_x1_sg U51123 ( .A(n51579), .B(n11076), .X(n11075) );
  inv_x1_sg U51124 ( .A(n11077), .X(n51579) );
  inv_x1_sg U51125 ( .A(n11079), .X(n51603) );
  inv_x1_sg U51126 ( .A(n11087), .X(n51635) );
  nand_x1_sg U51127 ( .A(n11095), .B(n51681), .X(n11094) );
  inv_x2_sg U51128 ( .A(n8878), .X(n44135) );
  nor_x1_sg U51129 ( .A(n11103), .B(n51724), .X(n8878) );
  inv_x2_sg U51130 ( .A(n8864), .X(n44133) );
  nor_x1_sg U51131 ( .A(n11107), .B(n51753), .X(n8864) );
  inv_x1_sg U51132 ( .A(n11112), .X(n51774) );
  inv_x1_sg U51133 ( .A(n11116), .X(n51790) );
  inv_x1_sg U51134 ( .A(n11119), .X(n51803) );
  inv_x2_sg U51135 ( .A(n8108), .X(n44174) );
  nor_x1_sg U51136 ( .A(n11831), .B(n12609), .X(n8108) );
  inv_x2_sg U51137 ( .A(n8902), .X(n44095) );
  nor_x1_sg U51138 ( .A(n11835), .B(n11836), .X(n8902) );
  nand_x1_sg U51139 ( .A(n11840), .B(n44030), .X(n11838) );
  nand_x1_sg U51140 ( .A(n51819), .B(n51829), .X(n11839) );
  inv_x1_sg U51141 ( .A(n11840), .X(n51829) );
  inv_x1_sg U51142 ( .A(n11850), .X(n51843) );
  nand_x1_sg U51143 ( .A(n51844), .B(n11855), .X(n11854) );
  inv_x1_sg U51144 ( .A(n11856), .X(n51844) );
  nand_x1_sg U51145 ( .A(n51858), .B(n11859), .X(n11858) );
  inv_x1_sg U51146 ( .A(n11860), .X(n51858) );
  inv_x1_sg U51147 ( .A(n11862), .X(n51884) );
  inv_x1_sg U51148 ( .A(n11870), .X(n51916) );
  nand_x1_sg U51149 ( .A(n11878), .B(n51962), .X(n11877) );
  inv_x2_sg U51150 ( .A(n8935), .X(n44131) );
  nor_x1_sg U51151 ( .A(n11886), .B(n52002), .X(n8935) );
  inv_x2_sg U51152 ( .A(n8927), .X(n44129) );
  nor_x1_sg U51153 ( .A(n11890), .B(n52036), .X(n8927) );
  inv_x1_sg U51154 ( .A(n11895), .X(n52054) );
  inv_x1_sg U51155 ( .A(n11902), .X(n52079) );
  nand_x1_sg U51156 ( .A(n46500), .B(n52102), .X(n12617) );
  nand_x1_sg U51157 ( .A(n12618), .B(n43896), .X(n12616) );
  inv_x1_sg U51158 ( .A(n12618), .X(n52102) );
  inv_x1_sg U51159 ( .A(n12627), .X(n52111) );
  nand_x1_sg U51160 ( .A(n52123), .B(n12633), .X(n12632) );
  inv_x1_sg U51161 ( .A(n12634), .X(n52123) );
  nand_x1_sg U51162 ( .A(n52137), .B(n12637), .X(n12636) );
  inv_x1_sg U51163 ( .A(n12638), .X(n52137) );
  inv_x1_sg U51164 ( .A(n12640), .X(n52161) );
  inv_x1_sg U51165 ( .A(n12648), .X(n52191) );
  nand_x1_sg U51166 ( .A(n12656), .B(n52237), .X(n12655) );
  inv_x2_sg U51167 ( .A(n8840), .X(n44127) );
  nor_x1_sg U51168 ( .A(n12664), .B(n52278), .X(n8840) );
  inv_x2_sg U51169 ( .A(n8826), .X(n44125) );
  nor_x1_sg U51170 ( .A(n12668), .B(n52311), .X(n8826) );
  inv_x1_sg U51171 ( .A(n12673), .X(n52331) );
  inv_x1_sg U51172 ( .A(n12677), .X(n52346) );
  inv_x1_sg U51173 ( .A(n12680), .X(n52357) );
  inv_x2_sg U51174 ( .A(n8793), .X(n44093) );
  nor_x1_sg U51175 ( .A(n13397), .B(n13398), .X(n8793) );
  nand_x1_sg U51176 ( .A(n46478), .B(n52381), .X(n13401) );
  nand_x1_sg U51177 ( .A(n13402), .B(n43884), .X(n13400) );
  inv_x1_sg U51178 ( .A(n13402), .X(n52381) );
  inv_x1_sg U51179 ( .A(n13412), .X(n52395) );
  nand_x1_sg U51180 ( .A(n52396), .B(n13417), .X(n13416) );
  inv_x1_sg U51181 ( .A(n13418), .X(n52396) );
  nand_x1_sg U51182 ( .A(n52410), .B(n13421), .X(n13420) );
  inv_x1_sg U51183 ( .A(n13422), .X(n52410) );
  inv_x1_sg U51184 ( .A(n13424), .X(n52435) );
  inv_x1_sg U51185 ( .A(n13432), .X(n52468) );
  nand_x1_sg U51186 ( .A(n13440), .B(n52514), .X(n13439) );
  inv_x2_sg U51187 ( .A(n8795), .X(n44123) );
  nor_x1_sg U51188 ( .A(n13448), .B(n52553), .X(n8795) );
  inv_x2_sg U51189 ( .A(n8791), .X(n44121) );
  nor_x1_sg U51190 ( .A(n13452), .B(n52586), .X(n8791) );
  inv_x1_sg U51191 ( .A(n13457), .X(n52606) );
  inv_x1_sg U51192 ( .A(n13461), .X(n52621) );
  inv_x1_sg U51193 ( .A(n13464), .X(n52632) );
  inv_x2_sg U51194 ( .A(n9004), .X(n44091) );
  nor_x1_sg U51195 ( .A(n14176), .B(n14177), .X(n9004) );
  nand_x1_sg U51196 ( .A(n14181), .B(n46456), .X(n14179) );
  nand_x1_sg U51197 ( .A(n52648), .B(n52657), .X(n14180) );
  inv_x1_sg U51198 ( .A(n14181), .X(n52657) );
  inv_x1_sg U51199 ( .A(n14191), .X(n52675) );
  nand_x1_sg U51200 ( .A(n52676), .B(n14196), .X(n14195) );
  inv_x1_sg U51201 ( .A(n14197), .X(n52676) );
  nand_x1_sg U51202 ( .A(n52687), .B(n14200), .X(n14199) );
  inv_x1_sg U51203 ( .A(n14201), .X(n52687) );
  inv_x1_sg U51204 ( .A(n14203), .X(n52718) );
  inv_x1_sg U51205 ( .A(n14211), .X(n52754) );
  nand_x1_sg U51206 ( .A(n14219), .B(n52793), .X(n14218) );
  inv_x1_sg U51207 ( .A(n14228), .X(n52830) );
  inv_x2_sg U51208 ( .A(n8942), .X(n44398) );
  nor_x1_sg U51209 ( .A(n14231), .B(n52862), .X(n8942) );
  inv_x1_sg U51210 ( .A(n14236), .X(n52884) );
  inv_x1_sg U51211 ( .A(n14240), .X(n52900) );
  inv_x1_sg U51212 ( .A(n14243), .X(n52913) );
  inv_x2_sg U51213 ( .A(n8074), .X(n44172) );
  nor_x1_sg U51214 ( .A(n14942), .B(n15724), .X(n8074) );
  nand_x1_sg U51215 ( .A(n46432), .B(n52936), .X(n14950) );
  nand_x1_sg U51216 ( .A(n14951), .B(n43892), .X(n14949) );
  inv_x1_sg U51217 ( .A(n14951), .X(n52936) );
  inv_x1_sg U51218 ( .A(n14960), .X(n52945) );
  nand_x1_sg U51219 ( .A(n52957), .B(n14966), .X(n14965) );
  inv_x1_sg U51220 ( .A(n14967), .X(n52957) );
  nand_x1_sg U51221 ( .A(n52971), .B(n14970), .X(n14969) );
  inv_x1_sg U51222 ( .A(n14971), .X(n52971) );
  inv_x1_sg U51223 ( .A(n14973), .X(n52995) );
  inv_x1_sg U51224 ( .A(n14981), .X(n53025) );
  nand_x1_sg U51225 ( .A(n14989), .B(n53071), .X(n14988) );
  inv_x2_sg U51226 ( .A(n8979), .X(n44119) );
  nor_x1_sg U51227 ( .A(n14997), .B(n53112), .X(n8979) );
  inv_x2_sg U51228 ( .A(n8965), .X(n44117) );
  nor_x1_sg U51229 ( .A(n15001), .B(n53145), .X(n8965) );
  inv_x1_sg U51230 ( .A(n15006), .X(n53165) );
  inv_x1_sg U51231 ( .A(n15010), .X(n53180) );
  inv_x1_sg U51232 ( .A(n15013), .X(n53191) );
  inv_x2_sg U51233 ( .A(n9338), .X(n44089) );
  nor_x1_sg U51234 ( .A(n15730), .B(n15731), .X(n9338) );
  nand_x1_sg U51235 ( .A(n15735), .B(n46411), .X(n15733) );
  nand_x1_sg U51236 ( .A(n53207), .B(n53217), .X(n15734) );
  inv_x1_sg U51237 ( .A(n15735), .X(n53217) );
  inv_x1_sg U51238 ( .A(n15745), .X(n53229) );
  nand_x1_sg U51239 ( .A(n53230), .B(n15750), .X(n15749) );
  inv_x1_sg U51240 ( .A(n15751), .X(n53230) );
  nand_x1_sg U51241 ( .A(n53244), .B(n15754), .X(n15753) );
  inv_x1_sg U51242 ( .A(n15755), .X(n53244) );
  inv_x1_sg U51243 ( .A(n15757), .X(n53271) );
  inv_x1_sg U51244 ( .A(n15765), .X(n53303) );
  nand_x1_sg U51245 ( .A(n15773), .B(n53350), .X(n15772) );
  inv_x2_sg U51246 ( .A(n9328), .X(n44115) );
  nor_x1_sg U51247 ( .A(n15781), .B(n53391), .X(n9328) );
  inv_x2_sg U51248 ( .A(n9318), .X(n44113) );
  nor_x1_sg U51249 ( .A(n15785), .B(n53422), .X(n9318) );
  inv_x1_sg U51250 ( .A(n15790), .X(n53444) );
  inv_x1_sg U51251 ( .A(n15794), .X(n53460) );
  inv_x1_sg U51252 ( .A(n15798), .X(n53471) );
  nand_x1_sg U51253 ( .A(n46388), .B(n53494), .X(n16516) );
  nand_x1_sg U51254 ( .A(n16517), .B(n43888), .X(n16515) );
  inv_x1_sg U51255 ( .A(n16517), .X(n53494) );
  inv_x1_sg U51256 ( .A(n16526), .X(n53503) );
  nand_x1_sg U51257 ( .A(n53515), .B(n16532), .X(n16531) );
  inv_x1_sg U51258 ( .A(n16533), .X(n53515) );
  nand_x1_sg U51259 ( .A(n53529), .B(n16536), .X(n16535) );
  inv_x1_sg U51260 ( .A(n16537), .X(n53529) );
  inv_x1_sg U51261 ( .A(n16539), .X(n53553) );
  inv_x1_sg U51262 ( .A(n16547), .X(n53583) );
  nand_x1_sg U51263 ( .A(n16555), .B(n53629), .X(n16554) );
  inv_x2_sg U51264 ( .A(n9296), .X(n44111) );
  nor_x1_sg U51265 ( .A(n16563), .B(n53670), .X(n9296) );
  inv_x2_sg U51266 ( .A(n9282), .X(n44109) );
  nor_x1_sg U51267 ( .A(n16567), .B(n53703), .X(n9282) );
  inv_x1_sg U51268 ( .A(n16572), .X(n53723) );
  inv_x1_sg U51269 ( .A(n16576), .X(n53738) );
  inv_x1_sg U51270 ( .A(n16579), .X(n53749) );
  nand_x1_sg U51271 ( .A(n17300), .B(n44014), .X(n17298) );
  nand_x1_sg U51272 ( .A(n53765), .B(n53773), .X(n17299) );
  inv_x1_sg U51273 ( .A(n17300), .X(n53773) );
  inv_x1_sg U51274 ( .A(n17309), .X(n53781) );
  nand_x1_sg U51275 ( .A(n53795), .B(n17315), .X(n17314) );
  nand_x1_sg U51276 ( .A(n53806), .B(n17319), .X(n17318) );
  inv_x1_sg U51277 ( .A(n17320), .X(n53806) );
  inv_x1_sg U51278 ( .A(n17322), .X(n53832) );
  inv_x1_sg U51279 ( .A(n17330), .X(n53874) );
  nand_x1_sg U51280 ( .A(n17338), .B(n53913), .X(n17337) );
  inv_x1_sg U51281 ( .A(n17347), .X(n53950) );
  inv_x2_sg U51282 ( .A(n9244), .X(n44396) );
  nor_x1_sg U51283 ( .A(n17350), .B(n53982), .X(n9244) );
  inv_x1_sg U51284 ( .A(n17355), .X(n54004) );
  inv_x1_sg U51285 ( .A(n17359), .X(n54020) );
  inv_x1_sg U51286 ( .A(n17362), .X(n54033) );
  inv_x2_sg U51287 ( .A(n8034), .X(n44428) );
  nor_x1_sg U51288 ( .A(n18063), .B(n18835), .X(n8034) );
  inv_x2_sg U51289 ( .A(n9056), .X(n44087) );
  nor_x1_sg U51290 ( .A(n18067), .B(n18068), .X(n9056) );
  nand_x1_sg U51291 ( .A(n46345), .B(n54055), .X(n18071) );
  nand_x1_sg U51292 ( .A(n18072), .B(n46346), .X(n18070) );
  inv_x1_sg U51293 ( .A(n18072), .X(n54055) );
  inv_x1_sg U51294 ( .A(n18082), .X(n54075) );
  nand_x1_sg U51295 ( .A(n54076), .B(n18087), .X(n18086) );
  inv_x1_sg U51296 ( .A(n18088), .X(n54076) );
  nand_x1_sg U51297 ( .A(n54088), .B(n18091), .X(n18090) );
  inv_x1_sg U51298 ( .A(n18092), .X(n54088) );
  inv_x1_sg U51299 ( .A(n18094), .X(n54119) );
  inv_x2_sg U51300 ( .A(n9052), .X(n44107) );
  nor_x1_sg U51301 ( .A(n18097), .B(n54135), .X(n9052) );
  inv_x1_sg U51302 ( .A(n18102), .X(n54153) );
  nand_x1_sg U51303 ( .A(n18110), .B(n54193), .X(n18109) );
  inv_x1_sg U51304 ( .A(n18119), .X(n54235) );
  inv_x2_sg U51305 ( .A(n9059), .X(n44394) );
  nor_x1_sg U51306 ( .A(n18122), .B(n54266), .X(n9059) );
  inv_x1_sg U51307 ( .A(n18127), .X(n54286) );
  inv_x1_sg U51308 ( .A(n18134), .X(n54314) );
  nand_x1_sg U51309 ( .A(n18845), .B(n44010), .X(n18843) );
  nand_x1_sg U51310 ( .A(n54330), .B(n54338), .X(n18844) );
  inv_x1_sg U51311 ( .A(n18845), .X(n54338) );
  inv_x1_sg U51312 ( .A(n18854), .X(n54346) );
  nand_x1_sg U51313 ( .A(n54360), .B(n18860), .X(n18859) );
  nand_x1_sg U51314 ( .A(n54371), .B(n18864), .X(n18863) );
  inv_x1_sg U51315 ( .A(n18865), .X(n54371) );
  inv_x1_sg U51316 ( .A(n18867), .X(n54397) );
  inv_x1_sg U51317 ( .A(n18875), .X(n54439) );
  nand_x1_sg U51318 ( .A(n18883), .B(n54478), .X(n18882) );
  inv_x1_sg U51319 ( .A(n18892), .X(n54515) );
  inv_x2_sg U51320 ( .A(n9206), .X(n44392) );
  nor_x1_sg U51321 ( .A(n18895), .B(n54547), .X(n9206) );
  inv_x1_sg U51322 ( .A(n18900), .X(n54569) );
  inv_x1_sg U51323 ( .A(n18904), .X(n54585) );
  inv_x1_sg U51324 ( .A(n18907), .X(n54598) );
  inv_x2_sg U51325 ( .A(n7978), .X(n43855) );
  nor_x1_sg U51326 ( .A(n19608), .B(n20380), .X(n7978) );
  inv_x2_sg U51327 ( .A(n9168), .X(n44085) );
  nor_x1_sg U51328 ( .A(n19612), .B(n19613), .X(n9168) );
  nand_x1_sg U51329 ( .A(n19617), .B(n43876), .X(n19615) );
  nand_x1_sg U51330 ( .A(n54614), .B(n54622), .X(n19616) );
  inv_x1_sg U51331 ( .A(n19617), .X(n54622) );
  inv_x1_sg U51332 ( .A(n19627), .X(n54639) );
  nand_x1_sg U51333 ( .A(n54640), .B(n19632), .X(n19631) );
  inv_x1_sg U51334 ( .A(n19633), .X(n54640) );
  nand_x1_sg U51335 ( .A(n54651), .B(n19636), .X(n19635) );
  inv_x1_sg U51336 ( .A(n19637), .X(n54651) );
  inv_x1_sg U51337 ( .A(n19639), .X(n54682) );
  inv_x1_sg U51338 ( .A(n19647), .X(n54718) );
  nand_x1_sg U51339 ( .A(n19655), .B(n54760), .X(n19654) );
  inv_x1_sg U51340 ( .A(n19664), .X(n54800) );
  inv_x2_sg U51341 ( .A(n9185), .X(n44390) );
  nor_x1_sg U51342 ( .A(n19667), .B(n54833), .X(n9185) );
  inv_x1_sg U51343 ( .A(n19672), .X(n54854) );
  inv_x1_sg U51344 ( .A(n19679), .X(n54882) );
  inv_x2_sg U51345 ( .A(n7988), .X(n44170) );
  nor_x1_sg U51346 ( .A(n19608), .B(n21152), .X(n7988) );
  nand_x1_sg U51347 ( .A(n20389), .B(n44006), .X(n20387) );
  nand_x1_sg U51348 ( .A(n54898), .B(n54906), .X(n20388) );
  inv_x1_sg U51349 ( .A(n20389), .X(n54906) );
  inv_x1_sg U51350 ( .A(n20398), .X(n54914) );
  nand_x1_sg U51351 ( .A(n54928), .B(n20404), .X(n20403) );
  nand_x1_sg U51352 ( .A(n54939), .B(n20408), .X(n20407) );
  inv_x1_sg U51353 ( .A(n20409), .X(n54939) );
  inv_x1_sg U51354 ( .A(n20411), .X(n54965) );
  inv_x1_sg U51355 ( .A(n20419), .X(n55007) );
  nand_x1_sg U51356 ( .A(n20427), .B(n55046), .X(n20426) );
  inv_x1_sg U51357 ( .A(n20436), .X(n55083) );
  inv_x2_sg U51358 ( .A(n9130), .X(n44388) );
  nor_x1_sg U51359 ( .A(n20439), .B(n55115), .X(n9130) );
  inv_x1_sg U51360 ( .A(n20444), .X(n55137) );
  inv_x1_sg U51361 ( .A(n20448), .X(n55153) );
  inv_x1_sg U51362 ( .A(n20451), .X(n55166) );
  inv_x2_sg U51363 ( .A(n9092), .X(n44083) );
  nor_x1_sg U51364 ( .A(n21157), .B(n21158), .X(n9092) );
  nand_x1_sg U51365 ( .A(n21162), .B(n43880), .X(n21160) );
  nand_x1_sg U51366 ( .A(n55182), .B(n55190), .X(n21161) );
  inv_x1_sg U51367 ( .A(n21162), .X(n55190) );
  inv_x1_sg U51368 ( .A(n21172), .X(n55207) );
  nand_x1_sg U51369 ( .A(n55208), .B(n21177), .X(n21176) );
  inv_x1_sg U51370 ( .A(n21178), .X(n55208) );
  nand_x1_sg U51371 ( .A(n55219), .B(n21181), .X(n21180) );
  inv_x1_sg U51372 ( .A(n21182), .X(n55219) );
  inv_x1_sg U51373 ( .A(n21184), .X(n55250) );
  inv_x1_sg U51374 ( .A(n21192), .X(n55286) );
  nand_x1_sg U51375 ( .A(n21200), .B(n55328), .X(n21199) );
  inv_x1_sg U51376 ( .A(n21209), .X(n55368) );
  inv_x2_sg U51377 ( .A(n9125), .X(n44386) );
  nor_x1_sg U51378 ( .A(n21212), .B(n55401), .X(n9125) );
  inv_x1_sg U51379 ( .A(n21217), .X(n55422) );
  inv_x1_sg U51380 ( .A(n21224), .X(n55450) );
  inv_x2_sg U51381 ( .A(n25432), .X(n44500) );
  nor_x1_sg U51382 ( .A(n25433), .B(n25434), .X(n25432) );
  inv_x2_sg U51383 ( .A(n25439), .X(n44242) );
  nor_x1_sg U51384 ( .A(n25440), .B(n25441), .X(n25439) );
  inv_x2_sg U51385 ( .A(n25453), .X(n44063) );
  nor_x1_sg U51386 ( .A(n25454), .B(n25455), .X(n25453) );
  inv_x2_sg U51387 ( .A(n25468), .X(n43933) );
  nor_x1_sg U51388 ( .A(n25469), .B(n25470), .X(n25468) );
  inv_x2_sg U51389 ( .A(n25482), .X(n43834) );
  nor_x1_sg U51390 ( .A(n25483), .B(n25484), .X(n25482) );
  nand_x1_sg U51391 ( .A(n29627), .B(n26358), .X(n32137) );
  inv_x2_sg U51392 ( .A(n25711), .X(n44061) );
  nor_x1_sg U51393 ( .A(n25712), .B(n25713), .X(n25711) );
  inv_x2_sg U51394 ( .A(n25718), .X(n44498) );
  nor_x1_sg U51395 ( .A(n25719), .B(n25720), .X(n25718) );
  inv_x2_sg U51396 ( .A(n25732), .X(n43931) );
  nor_x1_sg U51397 ( .A(n25733), .B(n25734), .X(n25732) );
  inv_x2_sg U51398 ( .A(n25746), .X(n44059) );
  nor_x1_sg U51399 ( .A(n25747), .B(n25748), .X(n25746) );
  nand_x1_sg U51400 ( .A(n46229), .B(n11623), .X(n25766) );
  inv_x2_sg U51401 ( .A(n25989), .X(n44496) );
  nor_x1_sg U51402 ( .A(n25990), .B(n25991), .X(n25989) );
  inv_x2_sg U51403 ( .A(n25996), .X(n44240) );
  nor_x1_sg U51404 ( .A(n25997), .B(n25998), .X(n25996) );
  inv_x2_sg U51405 ( .A(n26010), .X(n43929) );
  nor_x1_sg U51406 ( .A(n26011), .B(n26012), .X(n26010) );
  inv_x2_sg U51407 ( .A(n26024), .X(n43832) );
  nor_x1_sg U51408 ( .A(n26025), .B(n26026), .X(n26024) );
  nand_x1_sg U51409 ( .A(n46227), .B(n12404), .X(n26044) );
  inv_x2_sg U51410 ( .A(n26270), .X(n44057) );
  nor_x1_sg U51411 ( .A(n26271), .B(n26272), .X(n26270) );
  inv_x2_sg U51412 ( .A(n26277), .X(n44494) );
  nor_x1_sg U51413 ( .A(n26278), .B(n26279), .X(n26277) );
  inv_x2_sg U51414 ( .A(n26291), .X(n44238) );
  nor_x1_sg U51415 ( .A(n26292), .B(n26293), .X(n26291) );
  inv_x2_sg U51416 ( .A(n26305), .X(n43830) );
  nor_x1_sg U51417 ( .A(n26306), .B(n26307), .X(n26305) );
  inv_x2_sg U51418 ( .A(n26319), .X(n43927) );
  nor_x1_sg U51419 ( .A(n26320), .B(n26321), .X(n26319) );
  inv_x2_sg U51420 ( .A(n26549), .X(n44055) );
  nor_x1_sg U51421 ( .A(n26550), .B(n26551), .X(n26549) );
  inv_x2_sg U51422 ( .A(n26556), .X(n44492) );
  nor_x1_sg U51423 ( .A(n26557), .B(n26558), .X(n26556) );
  inv_x2_sg U51424 ( .A(n26570), .X(n43925) );
  nor_x1_sg U51425 ( .A(n26571), .B(n26572), .X(n26570) );
  inv_x2_sg U51426 ( .A(n26584), .X(n43923) );
  nor_x1_sg U51427 ( .A(n26585), .B(n26586), .X(n26584) );
  inv_x2_sg U51428 ( .A(n26598), .X(n44236) );
  nor_x1_sg U51429 ( .A(n26599), .B(n26600), .X(n26598) );
  inv_x2_sg U51430 ( .A(n26827), .X(n43921) );
  nor_x1_sg U51431 ( .A(n26828), .B(n26829), .X(n26827) );
  inv_x2_sg U51432 ( .A(n26834), .X(n44234) );
  nor_x1_sg U51433 ( .A(n26835), .B(n26836), .X(n26834) );
  inv_x2_sg U51434 ( .A(n26848), .X(n44053) );
  nor_x1_sg U51435 ( .A(n26849), .B(n26850), .X(n26848) );
  inv_x2_sg U51436 ( .A(n26862), .X(n43919) );
  nor_x1_sg U51437 ( .A(n26863), .B(n26864), .X(n26862) );
  inv_x2_sg U51438 ( .A(n26876), .X(n43828) );
  nor_x1_sg U51439 ( .A(n26877), .B(n26878), .X(n26876) );
  inv_x2_sg U51440 ( .A(n27106), .X(n44051) );
  nor_x1_sg U51441 ( .A(n27107), .B(n27108), .X(n27106) );
  inv_x2_sg U51442 ( .A(n27113), .X(n44490) );
  nor_x1_sg U51443 ( .A(n27114), .B(n27115), .X(n27113) );
  inv_x2_sg U51444 ( .A(n27127), .X(n44232) );
  nor_x1_sg U51445 ( .A(n27128), .B(n27129), .X(n27127) );
  inv_x2_sg U51446 ( .A(n27141), .X(n43826) );
  nor_x1_sg U51447 ( .A(n27142), .B(n27143), .X(n27141) );
  inv_x2_sg U51448 ( .A(n27155), .X(n43917) );
  nor_x1_sg U51449 ( .A(n27156), .B(n27157), .X(n27155) );
  nand_x1_sg U51450 ( .A(n46584), .B(n26358), .X(n27620) );
  inv_x2_sg U51451 ( .A(n27386), .X(n44488) );
  nor_x1_sg U51452 ( .A(n27387), .B(n27388), .X(n27386) );
  inv_x2_sg U51453 ( .A(n27393), .X(n45486) );
  nor_x1_sg U51454 ( .A(n27394), .B(n27395), .X(n27393) );
  inv_x2_sg U51455 ( .A(n27407), .X(n43915) );
  nor_x1_sg U51456 ( .A(n27408), .B(n27409), .X(n27407) );
  inv_x2_sg U51457 ( .A(n27421), .X(n43824) );
  nor_x1_sg U51458 ( .A(n27422), .B(n27423), .X(n27421) );
  nand_x1_sg U51459 ( .A(n46217), .B(n16299), .X(n27441) );
  nand_x1_sg U51460 ( .A(n27900), .B(n26358), .X(n27899) );
  inv_x2_sg U51461 ( .A(n27666), .X(n44049) );
  nor_x1_sg U51462 ( .A(n27667), .B(n27668), .X(n27666) );
  inv_x2_sg U51463 ( .A(n27673), .X(n44486) );
  nor_x1_sg U51464 ( .A(n27674), .B(n27675), .X(n27673) );
  inv_x2_sg U51465 ( .A(n27687), .X(n44230) );
  nor_x1_sg U51466 ( .A(n27688), .B(n27689), .X(n27687) );
  inv_x2_sg U51467 ( .A(n27701), .X(n43795) );
  nor_x1_sg U51468 ( .A(n27702), .B(n27703), .X(n27701) );
  inv_x2_sg U51469 ( .A(n27715), .X(n43768) );
  nor_x1_sg U51470 ( .A(n27716), .B(n27717), .X(n27715) );
  inv_x2_sg U51471 ( .A(n27946), .X(n44047) );
  nor_x1_sg U51472 ( .A(n27947), .B(n27948), .X(n27946) );
  inv_x2_sg U51473 ( .A(n27953), .X(n44228) );
  nor_x1_sg U51474 ( .A(n27954), .B(n27955), .X(n27953) );
  inv_x2_sg U51475 ( .A(n27967), .X(n43913) );
  nor_x1_sg U51476 ( .A(n27968), .B(n27969), .X(n27967) );
  inv_x2_sg U51477 ( .A(n27981), .X(n43822) );
  nor_x1_sg U51478 ( .A(n27982), .B(n27983), .X(n27981) );
  inv_x2_sg U51479 ( .A(n27995), .X(n43793) );
  nor_x1_sg U51480 ( .A(n27996), .B(n27997), .X(n27995) );
  inv_x2_sg U51481 ( .A(n28225), .X(n43911) );
  nor_x1_sg U51482 ( .A(n28226), .B(n28227), .X(n28225) );
  inv_x2_sg U51483 ( .A(n28232), .X(n44484) );
  nor_x1_sg U51484 ( .A(n28233), .B(n28234), .X(n28232) );
  inv_x2_sg U51485 ( .A(n28246), .X(n44482) );
  nor_x1_sg U51486 ( .A(n28247), .B(n28248), .X(n28246) );
  inv_x2_sg U51487 ( .A(n28261), .X(n43909) );
  nor_x1_sg U51488 ( .A(n28262), .B(n28263), .X(n28261) );
  inv_x2_sg U51489 ( .A(n28275), .X(n44226) );
  nor_x1_sg U51490 ( .A(n28276), .B(n28277), .X(n28275) );
  inv_x2_sg U51491 ( .A(n28504), .X(n44045) );
  nor_x1_sg U51492 ( .A(n28505), .B(n28506), .X(n28504) );
  inv_x2_sg U51493 ( .A(n28511), .X(n43907) );
  nor_x1_sg U51494 ( .A(n28512), .B(n28513), .X(n28511) );
  inv_x2_sg U51495 ( .A(n28525), .X(n43820) );
  nor_x1_sg U51496 ( .A(n28526), .B(n28527), .X(n28525) );
  inv_x2_sg U51497 ( .A(n28539), .X(n43818) );
  nor_x1_sg U51498 ( .A(n28540), .B(n28541), .X(n28539) );
  inv_x2_sg U51499 ( .A(n28553), .X(n43905) );
  nor_x1_sg U51500 ( .A(n28554), .B(n28555), .X(n28553) );
  inv_x2_sg U51501 ( .A(n28783), .X(n44480) );
  nor_x1_sg U51502 ( .A(n28784), .B(n28785), .X(n28783) );
  inv_x2_sg U51503 ( .A(n28790), .X(n44224) );
  nor_x1_sg U51504 ( .A(n28791), .B(n28792), .X(n28790) );
  inv_x2_sg U51505 ( .A(n28804), .X(n44222) );
  nor_x1_sg U51506 ( .A(n28805), .B(n28806), .X(n28804) );
  inv_x2_sg U51507 ( .A(n28819), .X(n44220) );
  nor_x1_sg U51508 ( .A(n28820), .B(n28821), .X(n28819) );
  inv_x2_sg U51509 ( .A(n28833), .X(n44043) );
  nor_x1_sg U51510 ( .A(n28834), .B(n28835), .X(n28833) );
  inv_x2_sg U51511 ( .A(n29063), .X(n44041) );
  nor_x1_sg U51512 ( .A(n29064), .B(n29065), .X(n29063) );
  inv_x2_sg U51513 ( .A(n29070), .X(n44218) );
  nor_x1_sg U51514 ( .A(n29071), .B(n29072), .X(n29070) );
  inv_x2_sg U51515 ( .A(n29084), .X(n43903) );
  nor_x1_sg U51516 ( .A(n29085), .B(n29086), .X(n29084) );
  inv_x2_sg U51517 ( .A(n29098), .X(n43901) );
  nor_x1_sg U51518 ( .A(n29099), .B(n29100), .X(n29098) );
  inv_x2_sg U51519 ( .A(n29112), .X(n43816) );
  nor_x1_sg U51520 ( .A(n29113), .B(n29114), .X(n29112) );
  inv_x2_sg U51521 ( .A(n29344), .X(n44478) );
  nor_x1_sg U51522 ( .A(n29345), .B(n29346), .X(n29344) );
  inv_x2_sg U51523 ( .A(n29351), .X(n44216) );
  nor_x1_sg U51524 ( .A(n29352), .B(n29353), .X(n29351) );
  inv_x2_sg U51525 ( .A(n29365), .X(n44039) );
  nor_x1_sg U51526 ( .A(n29366), .B(n29367), .X(n29365) );
  inv_x2_sg U51527 ( .A(n29380), .X(n43899) );
  nor_x1_sg U51528 ( .A(n29381), .B(n29382), .X(n29380) );
  inv_x2_sg U51529 ( .A(n29394), .X(n43814) );
  nor_x1_sg U51530 ( .A(n29395), .B(n29396), .X(n29394) );
  nand_x1_sg U51531 ( .A(n39291), .B(n39292), .X(out[0]) );
  nand_x1_sg U51532 ( .A(out_L2[0]), .B(n46670), .X(n39291) );
  nand_x1_sg U51533 ( .A(out_L1[0]), .B(n46672), .X(n39292) );
  nand_x1_sg U51534 ( .A(n39269), .B(n39270), .X(out[1]) );
  nand_x1_sg U51535 ( .A(out_L2[1]), .B(n46671), .X(n39269) );
  nand_x1_sg U51536 ( .A(out_L1[1]), .B(n46672), .X(n39270) );
  nand_x1_sg U51537 ( .A(n39267), .B(n39268), .X(out[2]) );
  nand_x1_sg U51538 ( .A(out_L2[2]), .B(n46665), .X(n39267) );
  nand_x1_sg U51539 ( .A(out_L1[2]), .B(n46672), .X(n39268) );
  nand_x1_sg U51540 ( .A(n39265), .B(n39266), .X(out[3]) );
  nand_x1_sg U51541 ( .A(out_L2[3]), .B(n46665), .X(n39265) );
  nand_x1_sg U51542 ( .A(out_L1[3]), .B(n46672), .X(n39266) );
  nand_x1_sg U51543 ( .A(n39263), .B(n39264), .X(out[4]) );
  nand_x1_sg U51544 ( .A(out_L2[4]), .B(n46664), .X(n39263) );
  nand_x1_sg U51545 ( .A(out_L1[4]), .B(n46672), .X(n39264) );
  nand_x1_sg U51546 ( .A(n39261), .B(n39262), .X(out[5]) );
  nand_x1_sg U51547 ( .A(out_L2[5]), .B(n46664), .X(n39261) );
  nand_x1_sg U51548 ( .A(out_L1[5]), .B(n46672), .X(n39262) );
  nand_x1_sg U51549 ( .A(n39259), .B(n39260), .X(out[6]) );
  nand_x1_sg U51550 ( .A(out_L2[6]), .B(n46662), .X(n39259) );
  nand_x1_sg U51551 ( .A(out_L1[6]), .B(n46672), .X(n39260) );
  nand_x1_sg U51552 ( .A(n39257), .B(n39258), .X(out[7]) );
  nand_x1_sg U51553 ( .A(out_L2[7]), .B(n46661), .X(n39257) );
  nand_x1_sg U51554 ( .A(out_L1[7]), .B(n46672), .X(n39258) );
  nand_x1_sg U51555 ( .A(n39255), .B(n39256), .X(out[8]) );
  nand_x1_sg U51556 ( .A(out_L2[8]), .B(n46663), .X(n39255) );
  nand_x1_sg U51557 ( .A(out_L1[8]), .B(n46672), .X(n39256) );
  nand_x1_sg U51558 ( .A(n39253), .B(n39254), .X(out[9]) );
  nand_x1_sg U51559 ( .A(out_L2[9]), .B(n46663), .X(n39253) );
  nand_x1_sg U51560 ( .A(n46672), .B(out_L1[9]), .X(n39254) );
  nand_x1_sg U51561 ( .A(n39289), .B(n39290), .X(out[10]) );
  nand_x1_sg U51562 ( .A(out_L2[10]), .B(n46670), .X(n39289) );
  nand_x1_sg U51563 ( .A(out_L1[10]), .B(n46672), .X(n39290) );
  nand_x1_sg U51564 ( .A(n39287), .B(n39288), .X(out[11]) );
  nand_x1_sg U51565 ( .A(out_L2[11]), .B(n46669), .X(n39287) );
  nand_x1_sg U51566 ( .A(out_L1[11]), .B(n46672), .X(n39288) );
  nand_x1_sg U51567 ( .A(n39285), .B(n39286), .X(out[12]) );
  nand_x1_sg U51568 ( .A(out_L2[12]), .B(n46669), .X(n39285) );
  nand_x1_sg U51569 ( .A(out_L1[12]), .B(n46672), .X(n39286) );
  nand_x1_sg U51570 ( .A(n39283), .B(n39284), .X(out[13]) );
  nand_x1_sg U51571 ( .A(out_L2[13]), .B(n46668), .X(n39283) );
  nand_x1_sg U51572 ( .A(out_L1[13]), .B(n46672), .X(n39284) );
  nand_x1_sg U51573 ( .A(n39281), .B(n39282), .X(out[14]) );
  nand_x1_sg U51574 ( .A(out_L2[14]), .B(n46668), .X(n39281) );
  nand_x1_sg U51575 ( .A(out_L1[14]), .B(n46672), .X(n39282) );
  nand_x1_sg U51576 ( .A(n39279), .B(n39280), .X(out[15]) );
  nand_x1_sg U51577 ( .A(out_L2[15]), .B(n46667), .X(n39279) );
  nand_x1_sg U51578 ( .A(out_L1[15]), .B(n46672), .X(n39280) );
  nand_x1_sg U51579 ( .A(n39277), .B(n39278), .X(out[16]) );
  nand_x1_sg U51580 ( .A(out_L2[16]), .B(n46667), .X(n39277) );
  nand_x1_sg U51581 ( .A(out_L1[16]), .B(n46672), .X(n39278) );
  nand_x1_sg U51582 ( .A(n39275), .B(n39276), .X(out[17]) );
  nand_x1_sg U51583 ( .A(out_L2[17]), .B(n46666), .X(n39275) );
  nand_x1_sg U51584 ( .A(out_L1[17]), .B(n46672), .X(n39276) );
  nand_x1_sg U51585 ( .A(n39273), .B(n39274), .X(out[18]) );
  nand_x1_sg U51586 ( .A(out_L2[18]), .B(n46666), .X(n39273) );
  nand_x1_sg U51587 ( .A(out_L1[18]), .B(n46672), .X(n39274) );
  nand_x1_sg U51588 ( .A(n39271), .B(n39272), .X(out[19]) );
  nand_x1_sg U51589 ( .A(out_L2[19]), .B(n46673), .X(n39271) );
  nand_x1_sg U51590 ( .A(out_L1[19]), .B(n46672), .X(n39272) );
  nand_x1_sg U51591 ( .A(n9012), .B(n21930), .X(\L2_0/n2903 ) );
  nand_x1_sg U51592 ( .A(n21931), .B(n55490), .X(n21930) );
  inv_x1_sg U51593 ( .A(n21929), .X(n55490) );
  nand_x1_sg U51594 ( .A(n9012), .B(n9358), .X(\L2_0/n4219 ) );
  nand_x1_sg U51595 ( .A(n9359), .B(n55471), .X(n9358) );
  inv_x1_sg U51596 ( .A(n9357), .X(n55471) );
  nand_x1_sg U51597 ( .A(n9012), .B(n9419), .X(\L2_0/n4215 ) );
  nand_x1_sg U51598 ( .A(n9420), .B(n55472), .X(n9419) );
  inv_x1_sg U51599 ( .A(n9418), .X(n55472) );
  nand_x1_sg U51600 ( .A(n9012), .B(n9468), .X(\L2_0/n4211 ) );
  nand_x1_sg U51601 ( .A(n9469), .B(n55473), .X(n9468) );
  inv_x1_sg U51602 ( .A(n9467), .X(n55473) );
  nand_x1_sg U51603 ( .A(n9012), .B(n9517), .X(\L2_0/n4207 ) );
  nand_x1_sg U51604 ( .A(n9518), .B(n55474), .X(n9517) );
  inv_x1_sg U51605 ( .A(n9516), .X(n55474) );
  nand_x1_sg U51606 ( .A(n9012), .B(n9566), .X(\L2_0/n4203 ) );
  nand_x1_sg U51607 ( .A(n9567), .B(n55475), .X(n9566) );
  inv_x1_sg U51608 ( .A(n9565), .X(n55475) );
  nand_x1_sg U51609 ( .A(n9012), .B(n9614), .X(\L2_0/n4199 ) );
  nand_x1_sg U51610 ( .A(n9615), .B(n55476), .X(n9614) );
  inv_x1_sg U51611 ( .A(n9613), .X(n55476) );
  nand_x1_sg U51612 ( .A(n9012), .B(n9662), .X(\L2_0/n4195 ) );
  nand_x1_sg U51613 ( .A(n9663), .B(n55477), .X(n9662) );
  inv_x1_sg U51614 ( .A(n9661), .X(n55477) );
  nand_x1_sg U51615 ( .A(n9012), .B(n9709), .X(\L2_0/n4191 ) );
  nand_x1_sg U51616 ( .A(n9710), .B(n55478), .X(n9709) );
  inv_x1_sg U51617 ( .A(n9708), .X(n55478) );
  nand_x1_sg U51618 ( .A(n9012), .B(n9757), .X(\L2_0/n4187 ) );
  nand_x1_sg U51619 ( .A(n9758), .B(n55479), .X(n9757) );
  inv_x1_sg U51620 ( .A(n9756), .X(n55479) );
  nand_x1_sg U51621 ( .A(n9012), .B(n9805), .X(\L2_0/n4183 ) );
  nand_x1_sg U51622 ( .A(n9806), .B(n55480), .X(n9805) );
  inv_x1_sg U51623 ( .A(n9804), .X(n55480) );
  nand_x1_sg U51624 ( .A(n9012), .B(n9853), .X(\L2_0/n4179 ) );
  nand_x1_sg U51625 ( .A(n9854), .B(n55481), .X(n9853) );
  inv_x1_sg U51626 ( .A(n9852), .X(n55481) );
  nand_x1_sg U51627 ( .A(n9012), .B(n9901), .X(\L2_0/n4175 ) );
  nand_x1_sg U51628 ( .A(n9902), .B(n55482), .X(n9901) );
  inv_x1_sg U51629 ( .A(n9900), .X(n55482) );
  nand_x1_sg U51630 ( .A(n9012), .B(n9949), .X(\L2_0/n4171 ) );
  nand_x1_sg U51631 ( .A(n9950), .B(n55483), .X(n9949) );
  inv_x1_sg U51632 ( .A(n9948), .X(n55483) );
  nand_x1_sg U51633 ( .A(n9012), .B(n9998), .X(\L2_0/n4167 ) );
  nand_x1_sg U51634 ( .A(n9999), .B(n55484), .X(n9998) );
  inv_x1_sg U51635 ( .A(n9997), .X(n55484) );
  nand_x1_sg U51636 ( .A(n9012), .B(n10046), .X(\L2_0/n4163 ) );
  nand_x1_sg U51637 ( .A(n10047), .B(n55485), .X(n10046) );
  inv_x1_sg U51638 ( .A(n10045), .X(n55485) );
  nand_x1_sg U51639 ( .A(n9012), .B(n10095), .X(\L2_0/n4159 ) );
  nand_x1_sg U51640 ( .A(n10096), .B(n55486), .X(n10095) );
  inv_x1_sg U51641 ( .A(n10094), .X(n55486) );
  nand_x1_sg U51642 ( .A(n9012), .B(n10144), .X(\L2_0/n4155 ) );
  nand_x1_sg U51643 ( .A(n10145), .B(n55487), .X(n10144) );
  inv_x1_sg U51644 ( .A(n10143), .X(n55487) );
  nand_x1_sg U51645 ( .A(n9012), .B(n10191), .X(\L2_0/n4151 ) );
  nand_x1_sg U51646 ( .A(n10192), .B(n55488), .X(n10191) );
  inv_x1_sg U51647 ( .A(n10190), .X(n55488) );
  nand_x1_sg U51648 ( .A(n9012), .B(n10234), .X(\L2_0/n4147 ) );
  nand_x1_sg U51649 ( .A(n10235), .B(n55489), .X(n10234) );
  inv_x1_sg U51650 ( .A(n10233), .X(n55489) );
  nand_x1_sg U51651 ( .A(n9012), .B(n9037), .X(n8054) );
  nand_x1_sg U51652 ( .A(n46573), .B(n8050), .X(n9037) );
  nand_x1_sg U51653 ( .A(n9012), .B(n9035), .X(n8055) );
  nand_x1_sg U51654 ( .A(n9036), .B(n46578), .X(n9035) );
  nand_x1_sg U51655 ( .A(n9012), .B(n9048), .X(n8047) );
  nand_x1_sg U51656 ( .A(n9012), .B(n9044), .X(n8049) );
  nand_x1_sg U51657 ( .A(n9045), .B(n46577), .X(n9044) );
  nand_x1_sg U51658 ( .A(n9012), .B(n9033), .X(n8056) );
  nand_x1_sg U51659 ( .A(n9034), .B(n46577), .X(n9033) );
  nand_x1_sg U51660 ( .A(n9012), .B(n9031), .X(n8057) );
  nand_x1_sg U51661 ( .A(n9032), .B(n8050), .X(n9031) );
  nand_x1_sg U51662 ( .A(n9012), .B(n9029), .X(n8058) );
  nand_x1_sg U51663 ( .A(n9030), .B(n46578), .X(n9029) );
  nand_x1_sg U51664 ( .A(n9012), .B(n9046), .X(n8048) );
  nand_x1_sg U51665 ( .A(n9047), .B(n46578), .X(n9046) );
  nand_x1_sg U51666 ( .A(n9012), .B(n9027), .X(n8059) );
  nand_x1_sg U51667 ( .A(n9028), .B(n46577), .X(n9027) );
  nand_x1_sg U51668 ( .A(n9012), .B(n9025), .X(n8060) );
  nand_x1_sg U51669 ( .A(n9012), .B(n9040), .X(n8052) );
  nand_x1_sg U51670 ( .A(n9041), .B(n46578), .X(n9040) );
  nand_x1_sg U51671 ( .A(n9012), .B(n9038), .X(n8053) );
  nand_x1_sg U51672 ( .A(n9012), .B(n9023), .X(n8061) );
  nand_x1_sg U51673 ( .A(n9024), .B(n46578), .X(n9023) );
  nand_x1_sg U51674 ( .A(n9012), .B(n9021), .X(n8062) );
  nand_x1_sg U51675 ( .A(n9012), .B(n9019), .X(n8063) );
  nand_x1_sg U51676 ( .A(n9020), .B(n8050), .X(n9019) );
  nand_x1_sg U51677 ( .A(n9012), .B(n9042), .X(n8051) );
  nand_x1_sg U51678 ( .A(n9012), .B(n9017), .X(n8064) );
  nand_x1_sg U51679 ( .A(n9018), .B(n46578), .X(n9017) );
  nand_x1_sg U51680 ( .A(n9012), .B(n9015), .X(n8065) );
  nand_x1_sg U51681 ( .A(n46577), .B(n9016), .X(n9015) );
  nand_x1_sg U51682 ( .A(n9012), .B(n9013), .X(n8066) );
  nand_x1_sg U51683 ( .A(n9014), .B(n8050), .X(n9013) );
  nand_x1_sg U51684 ( .A(n8860), .B(n8887), .X(n8131) );
  nand_x1_sg U51685 ( .A(n46550), .B(n46553), .X(n8887) );
  nand_x1_sg U51686 ( .A(n8860), .B(n8892), .X(n8128) );
  nand_x1_sg U51687 ( .A(n46553), .B(n8893), .X(n8892) );
  nand_x1_sg U51688 ( .A(n8860), .B(n8888), .X(n8130) );
  nand_x1_sg U51689 ( .A(n8860), .B(n8896), .X(n8126) );
  nand_x1_sg U51690 ( .A(n46553), .B(n8897), .X(n8896) );
  nand_x1_sg U51691 ( .A(n8860), .B(n8861), .X(n8144) );
  nand_x1_sg U51692 ( .A(n46553), .B(n8862), .X(n8861) );
  nand_x1_sg U51693 ( .A(n8860), .B(n8873), .X(n8138) );
  nand_x1_sg U51694 ( .A(n46553), .B(n8874), .X(n8873) );
  nand_x1_sg U51695 ( .A(n8860), .B(n8885), .X(n8132) );
  nand_x1_sg U51696 ( .A(n46553), .B(n8886), .X(n8885) );
  nand_x1_sg U51697 ( .A(n8860), .B(n8869), .X(n8140) );
  nand_x1_sg U51698 ( .A(n46553), .B(n8870), .X(n8869) );
  nand_x1_sg U51699 ( .A(n8860), .B(n8871), .X(n8139) );
  nand_x1_sg U51700 ( .A(n46553), .B(n8872), .X(n8871) );
  nand_x1_sg U51701 ( .A(n8860), .B(n8890), .X(n8129) );
  nand_x1_sg U51702 ( .A(n8860), .B(n8875), .X(n8137) );
  nand_x1_sg U51703 ( .A(n46553), .B(n8876), .X(n8875) );
  nand_x1_sg U51704 ( .A(n8860), .B(n8879), .X(n8135) );
  nand_x1_sg U51705 ( .A(n8860), .B(n8865), .X(n8142) );
  nand_x1_sg U51706 ( .A(n46553), .B(n8866), .X(n8865) );
  nand_x1_sg U51707 ( .A(n8860), .B(n8883), .X(n8133) );
  nand_x1_sg U51708 ( .A(n8860), .B(n8877), .X(n8136) );
  nand_x1_sg U51709 ( .A(n8860), .B(n8863), .X(n8143) );
  nand_x1_sg U51710 ( .A(n8860), .B(n8867), .X(n8141) );
  nand_x1_sg U51711 ( .A(n46553), .B(n8868), .X(n8867) );
  nand_x1_sg U51712 ( .A(n8860), .B(n8881), .X(n8134) );
  nand_x1_sg U51713 ( .A(n46553), .B(n8882), .X(n8881) );
  nand_x1_sg U51714 ( .A(n8860), .B(n8894), .X(n8127) );
  nand_x1_sg U51715 ( .A(n46553), .B(n8895), .X(n8894) );
  nand_x1_sg U51716 ( .A(n8898), .B(n8903), .X(n8123) );
  nand_x1_sg U51717 ( .A(n46528), .B(n46531), .X(n8903) );
  nand_x1_sg U51718 ( .A(n8898), .B(n8918), .X(n8115) );
  nand_x1_sg U51719 ( .A(n46531), .B(n8919), .X(n8918) );
  nand_x1_sg U51720 ( .A(n8898), .B(n8901), .X(n8124) );
  nand_x1_sg U51721 ( .A(n8898), .B(n8930), .X(n8109) );
  nand_x1_sg U51722 ( .A(n46531), .B(n8931), .X(n8930) );
  nand_x1_sg U51723 ( .A(n8898), .B(n8914), .X(n8117) );
  nand_x1_sg U51724 ( .A(n46531), .B(n41366), .X(n8914) );
  nand_x1_sg U51725 ( .A(n8898), .B(n8908), .X(n8120) );
  nand_x1_sg U51726 ( .A(n46531), .B(n8909), .X(n8908) );
  nand_x1_sg U51727 ( .A(n8898), .B(n8932), .X(n8107) );
  nand_x1_sg U51728 ( .A(n46531), .B(n8933), .X(n8932) );
  nand_x1_sg U51729 ( .A(n8898), .B(n8922), .X(n8113) );
  nand_x1_sg U51730 ( .A(n44175), .B(n8923), .X(n8922) );
  nand_x1_sg U51731 ( .A(n8898), .B(n8906), .X(n8121) );
  nand_x1_sg U51732 ( .A(n46531), .B(n8907), .X(n8906) );
  nand_x1_sg U51733 ( .A(n8898), .B(n8924), .X(n8112) );
  nand_x1_sg U51734 ( .A(n8898), .B(n8912), .X(n8118) );
  nand_x1_sg U51735 ( .A(n46531), .B(n8913), .X(n8912) );
  nand_x1_sg U51736 ( .A(n8898), .B(n8916), .X(n8116) );
  nand_x1_sg U51737 ( .A(n8898), .B(n8904), .X(n8122) );
  nand_x1_sg U51738 ( .A(n46531), .B(n8905), .X(n8904) );
  nand_x1_sg U51739 ( .A(n8898), .B(n8920), .X(n8114) );
  nand_x1_sg U51740 ( .A(n8898), .B(n8934), .X(n8106) );
  nand_x1_sg U51741 ( .A(n8898), .B(n8926), .X(n8111) );
  nand_x1_sg U51742 ( .A(n8898), .B(n8910), .X(n8119) );
  nand_x1_sg U51743 ( .A(n46531), .B(n8911), .X(n8910) );
  nand_x1_sg U51744 ( .A(n8898), .B(n8899), .X(n8125) );
  nand_x1_sg U51745 ( .A(n46531), .B(n8900), .X(n8899) );
  nand_x1_sg U51746 ( .A(n8898), .B(n8928), .X(n8110) );
  nand_x1_sg U51747 ( .A(n46531), .B(n8929), .X(n8928) );
  nand_x1_sg U51748 ( .A(n8822), .B(n8849), .X(n8150) );
  nand_x1_sg U51749 ( .A(n46508), .B(n46510), .X(n8849) );
  nand_x1_sg U51750 ( .A(n8822), .B(n8852), .X(n8148) );
  nand_x1_sg U51751 ( .A(n46510), .B(n8853), .X(n8852) );
  nand_x1_sg U51752 ( .A(n8822), .B(n8843), .X(n8153) );
  nand_x1_sg U51753 ( .A(n8822), .B(n8845), .X(n8152) );
  nand_x1_sg U51754 ( .A(n55787), .B(n8846), .X(n8845) );
  nand_x1_sg U51755 ( .A(n8822), .B(n8823), .X(n8163) );
  nand_x1_sg U51756 ( .A(n46510), .B(n8824), .X(n8823) );
  nand_x1_sg U51757 ( .A(n8822), .B(n8835), .X(n8157) );
  nand_x1_sg U51758 ( .A(n46510), .B(n8836), .X(n8835) );
  nand_x1_sg U51759 ( .A(n8822), .B(n8856), .X(n8146) );
  nand_x1_sg U51760 ( .A(n46510), .B(n8857), .X(n8856) );
  nand_x1_sg U51761 ( .A(n8822), .B(n8831), .X(n8159) );
  nand_x1_sg U51762 ( .A(n46510), .B(n8832), .X(n8831) );
  nand_x1_sg U51763 ( .A(n8822), .B(n8833), .X(n8158) );
  nand_x1_sg U51764 ( .A(n46510), .B(n8834), .X(n8833) );
  nand_x1_sg U51765 ( .A(n8822), .B(n8854), .X(n8147) );
  nand_x1_sg U51766 ( .A(n8822), .B(n8837), .X(n8156) );
  nand_x1_sg U51767 ( .A(n46510), .B(n8838), .X(n8837) );
  nand_x1_sg U51768 ( .A(n8822), .B(n8841), .X(n8154) );
  nand_x1_sg U51769 ( .A(n8822), .B(n8827), .X(n8161) );
  nand_x1_sg U51770 ( .A(n46510), .B(n8828), .X(n8827) );
  nand_x1_sg U51771 ( .A(n8822), .B(n8850), .X(n8149) );
  nand_x1_sg U51772 ( .A(n8822), .B(n8839), .X(n8155) );
  nand_x1_sg U51773 ( .A(n8822), .B(n8825), .X(n8162) );
  nand_x1_sg U51774 ( .A(n8822), .B(n8829), .X(n8160) );
  nand_x1_sg U51775 ( .A(n46510), .B(n8830), .X(n8829) );
  nand_x1_sg U51776 ( .A(n8822), .B(n8847), .X(n8151) );
  nand_x1_sg U51777 ( .A(n46510), .B(n8848), .X(n8847) );
  nand_x1_sg U51778 ( .A(n8822), .B(n8858), .X(n8145) );
  nand_x1_sg U51779 ( .A(n46510), .B(n8859), .X(n8858) );
  nand_x1_sg U51780 ( .A(n8783), .B(n8784), .X(n8182) );
  nand_x1_sg U51781 ( .A(n46487), .B(n46485), .X(n8784) );
  nand_x1_sg U51782 ( .A(n8783), .B(n8808), .X(n8170) );
  nand_x1_sg U51783 ( .A(n46487), .B(n8809), .X(n8808) );
  nand_x1_sg U51784 ( .A(n8783), .B(n8792), .X(n8178) );
  nand_x1_sg U51785 ( .A(n8783), .B(n8804), .X(n8172) );
  nand_x1_sg U51786 ( .A(n46487), .B(n8805), .X(n8804) );
  nand_x1_sg U51787 ( .A(n8783), .B(n8814), .X(n8167) );
  nand_x1_sg U51788 ( .A(n46487), .B(n41364), .X(n8814) );
  nand_x1_sg U51789 ( .A(n8783), .B(n8788), .X(n8180) );
  nand_x1_sg U51790 ( .A(n55788), .B(n8789), .X(n8788) );
  nand_x1_sg U51791 ( .A(n8783), .B(n8818), .X(n8165) );
  nand_x1_sg U51792 ( .A(n46487), .B(n8819), .X(n8818) );
  nand_x1_sg U51793 ( .A(n8783), .B(n8800), .X(n8174) );
  nand_x1_sg U51794 ( .A(n46487), .B(n8801), .X(n8800) );
  nand_x1_sg U51795 ( .A(n8783), .B(n8786), .X(n8181) );
  nand_x1_sg U51796 ( .A(n46487), .B(n8787), .X(n8786) );
  nand_x1_sg U51797 ( .A(n8783), .B(n8816), .X(n8166) );
  nand_x1_sg U51798 ( .A(n8783), .B(n8802), .X(n8173) );
  nand_x1_sg U51799 ( .A(n46487), .B(n41362), .X(n8802) );
  nand_x1_sg U51800 ( .A(n8783), .B(n8796), .X(n8176) );
  nand_x1_sg U51801 ( .A(n8783), .B(n8806), .X(n8171) );
  nand_x1_sg U51802 ( .A(n46487), .B(n8807), .X(n8806) );
  nand_x1_sg U51803 ( .A(n8783), .B(n8810), .X(n8169) );
  nand_x1_sg U51804 ( .A(n8783), .B(n8794), .X(n8177) );
  nand_x1_sg U51805 ( .A(n8783), .B(n8790), .X(n8179) );
  nand_x1_sg U51806 ( .A(n8783), .B(n8812), .X(n8168) );
  nand_x1_sg U51807 ( .A(n46487), .B(n8813), .X(n8812) );
  nand_x1_sg U51808 ( .A(n8783), .B(n8798), .X(n8175) );
  nand_x1_sg U51809 ( .A(n46487), .B(n8799), .X(n8798) );
  nand_x1_sg U51810 ( .A(n8783), .B(n8820), .X(n8164) );
  nand_x1_sg U51811 ( .A(n46487), .B(n8821), .X(n8820) );
  nand_x1_sg U51812 ( .A(n8936), .B(n9005), .X(n8070) );
  nand_x1_sg U51813 ( .A(n46463), .B(n46465), .X(n9005) );
  nand_x1_sg U51814 ( .A(n8936), .B(n9006), .X(n8069) );
  nand_x1_sg U51815 ( .A(n46465), .B(n9007), .X(n9006) );
  nand_x1_sg U51816 ( .A(n8936), .B(n9003), .X(n8071) );
  nand_x1_sg U51817 ( .A(n8936), .B(n9010), .X(n8067) );
  nand_x1_sg U51818 ( .A(n46465), .B(n9011), .X(n9010) );
  nand_x1_sg U51819 ( .A(n8936), .B(n8939), .X(n8104) );
  nand_x1_sg U51820 ( .A(n46465), .B(n8940), .X(n8939) );
  nand_x1_sg U51821 ( .A(n8936), .B(n8949), .X(n8099) );
  nand_x1_sg U51822 ( .A(n46465), .B(n8950), .X(n8949) );
  nand_x1_sg U51823 ( .A(n8936), .B(n8959), .X(n8094) );
  nand_x1_sg U51824 ( .A(n55793), .B(n8960), .X(n8959) );
  nand_x1_sg U51825 ( .A(n8936), .B(n8937), .X(n8105) );
  nand_x1_sg U51826 ( .A(n46465), .B(n8938), .X(n8937) );
  nand_x1_sg U51827 ( .A(n8936), .B(n8947), .X(n8100) );
  nand_x1_sg U51828 ( .A(n46465), .B(n8948), .X(n8947) );
  nand_x1_sg U51829 ( .A(n8936), .B(n8957), .X(n8095) );
  nand_x1_sg U51830 ( .A(n8936), .B(n8951), .X(n8098) );
  nand_x1_sg U51831 ( .A(n46465), .B(n8952), .X(n8951) );
  nand_x1_sg U51832 ( .A(n8936), .B(n8955), .X(n8096) );
  nand_x1_sg U51833 ( .A(n8936), .B(n8943), .X(n8102) );
  nand_x1_sg U51834 ( .A(n46465), .B(n8944), .X(n8943) );
  nand_x1_sg U51835 ( .A(n8936), .B(n8999), .X(n8073) );
  nand_x1_sg U51836 ( .A(n8936), .B(n8953), .X(n8097) );
  nand_x1_sg U51837 ( .A(n46465), .B(n8954), .X(n8953) );
  nand_x1_sg U51838 ( .A(n8936), .B(n8941), .X(n8103) );
  nand_x1_sg U51839 ( .A(n8936), .B(n8945), .X(n8101) );
  nand_x1_sg U51840 ( .A(n46465), .B(n8946), .X(n8945) );
  nand_x1_sg U51841 ( .A(n8936), .B(n9001), .X(n8072) );
  nand_x1_sg U51842 ( .A(n46465), .B(n9002), .X(n9001) );
  nand_x1_sg U51843 ( .A(n8936), .B(n9008), .X(n8068) );
  nand_x1_sg U51844 ( .A(n46465), .B(n9009), .X(n9008) );
  nand_x1_sg U51845 ( .A(n8961), .B(n8986), .X(n8081) );
  nand_x1_sg U51846 ( .A(n46440), .B(n44173), .X(n8986) );
  nand_x1_sg U51847 ( .A(n8961), .B(n8995), .X(n8076) );
  nand_x1_sg U51848 ( .A(n46442), .B(n8996), .X(n8995) );
  nand_x1_sg U51849 ( .A(n8961), .B(n8982), .X(n8083) );
  nand_x1_sg U51850 ( .A(n8961), .B(n8987), .X(n8080) );
  nand_x1_sg U51851 ( .A(n46442), .B(n8988), .X(n8987) );
  nand_x1_sg U51852 ( .A(n8961), .B(n8962), .X(n8093) );
  nand_x1_sg U51853 ( .A(n46442), .B(n8963), .X(n8962) );
  nand_x1_sg U51854 ( .A(n8961), .B(n8974), .X(n8087) );
  nand_x1_sg U51855 ( .A(n8961), .B(n8989), .X(n8079) );
  nand_x1_sg U51856 ( .A(n46442), .B(n8990), .X(n8989) );
  nand_x1_sg U51857 ( .A(n8961), .B(n8970), .X(n8089) );
  nand_x1_sg U51858 ( .A(n46442), .B(n8971), .X(n8970) );
  nand_x1_sg U51859 ( .A(n8961), .B(n8972), .X(n8088) );
  nand_x1_sg U51860 ( .A(n46442), .B(n8973), .X(n8972) );
  nand_x1_sg U51861 ( .A(n8961), .B(n8984), .X(n8082) );
  nand_x1_sg U51862 ( .A(n8961), .B(n8976), .X(n8086) );
  nand_x1_sg U51863 ( .A(n46442), .B(n8977), .X(n8976) );
  nand_x1_sg U51864 ( .A(n8961), .B(n8980), .X(n8084) );
  nand_x1_sg U51865 ( .A(n8961), .B(n8966), .X(n8091) );
  nand_x1_sg U51866 ( .A(n46442), .B(n8967), .X(n8966) );
  nand_x1_sg U51867 ( .A(n8961), .B(n8993), .X(n8077) );
  nand_x1_sg U51868 ( .A(n8961), .B(n8978), .X(n8085) );
  nand_x1_sg U51869 ( .A(n8961), .B(n8964), .X(n8092) );
  nand_x1_sg U51870 ( .A(n8961), .B(n8968), .X(n8090) );
  nand_x1_sg U51871 ( .A(n46442), .B(n8969), .X(n8968) );
  nand_x1_sg U51872 ( .A(n8961), .B(n8991), .X(n8078) );
  nand_x1_sg U51873 ( .A(n46442), .B(n8992), .X(n8991) );
  nand_x1_sg U51874 ( .A(n8961), .B(n8997), .X(n8075) );
  nand_x1_sg U51875 ( .A(n46442), .B(n8998), .X(n8997) );
  nand_x1_sg U51876 ( .A(n9316), .B(n9339), .X(n7899) );
  nand_x1_sg U51877 ( .A(n46416), .B(n55792), .X(n9339) );
  nand_x1_sg U51878 ( .A(n9316), .B(n9342), .X(n7897) );
  nand_x1_sg U51879 ( .A(n46419), .B(n9343), .X(n9342) );
  nand_x1_sg U51880 ( .A(n9316), .B(n9337), .X(n7900) );
  nand_x1_sg U51881 ( .A(n9316), .B(n9325), .X(n7906) );
  nand_x1_sg U51882 ( .A(n46419), .B(n9326), .X(n9325) );
  nand_x1_sg U51883 ( .A(n9316), .B(n9352), .X(n7892) );
  nand_x1_sg U51884 ( .A(n46419), .B(n41360), .X(n9352) );
  nand_x1_sg U51885 ( .A(n9316), .B(n9333), .X(n7902) );
  nand_x1_sg U51886 ( .A(n46419), .B(n9334), .X(n9333) );
  nand_x1_sg U51887 ( .A(n9316), .B(n9321), .X(n7908) );
  nand_x1_sg U51888 ( .A(n46419), .B(n9322), .X(n9321) );
  nand_x1_sg U51889 ( .A(n9316), .B(n9346), .X(n7895) );
  nand_x1_sg U51890 ( .A(n46419), .B(n9347), .X(n9346) );
  nand_x1_sg U51891 ( .A(n9316), .B(n9331), .X(n7903) );
  nand_x1_sg U51892 ( .A(n46419), .B(n9332), .X(n9331) );
  nand_x1_sg U51893 ( .A(n9316), .B(n9319), .X(n7909) );
  nand_x1_sg U51894 ( .A(n9316), .B(n9350), .X(n7893) );
  nand_x1_sg U51895 ( .A(n46419), .B(n9351), .X(n9350) );
  nand_x1_sg U51896 ( .A(n9316), .B(n9340), .X(n7898) );
  nand_x1_sg U51897 ( .A(n9316), .B(n9329), .X(n7904) );
  nand_x1_sg U51898 ( .A(n46419), .B(n9330), .X(n9329) );
  nand_x1_sg U51899 ( .A(n9316), .B(n9344), .X(n7896) );
  nand_x1_sg U51900 ( .A(n9316), .B(n9327), .X(n7905) );
  nand_x1_sg U51901 ( .A(n9316), .B(n9317), .X(n7910) );
  nand_x1_sg U51902 ( .A(n9316), .B(n9348), .X(n7894) );
  nand_x1_sg U51903 ( .A(n46419), .B(n9349), .X(n9348) );
  nand_x1_sg U51904 ( .A(n9316), .B(n9335), .X(n7901) );
  nand_x1_sg U51905 ( .A(n46419), .B(n9336), .X(n9335) );
  nand_x1_sg U51906 ( .A(n9316), .B(n9323), .X(n7907) );
  nand_x1_sg U51907 ( .A(n46419), .B(n9324), .X(n9323) );
  nand_x1_sg U51908 ( .A(n9278), .B(n9303), .X(n7917) );
  nand_x1_sg U51909 ( .A(n46394), .B(n46398), .X(n9303) );
  nand_x1_sg U51910 ( .A(n9278), .B(n9306), .X(n7915) );
  nand_x1_sg U51911 ( .A(n55791), .B(n9307), .X(n9306) );
  nand_x1_sg U51912 ( .A(n9278), .B(n9301), .X(n7918) );
  nand_x1_sg U51913 ( .A(n9278), .B(n9312), .X(n7912) );
  nand_x1_sg U51914 ( .A(n46398), .B(n9313), .X(n9312) );
  nand_x1_sg U51915 ( .A(n9278), .B(n9279), .X(n7929) );
  nand_x1_sg U51916 ( .A(n46398), .B(n9280), .X(n9279) );
  nand_x1_sg U51917 ( .A(n9278), .B(n9291), .X(n7923) );
  nand_x1_sg U51918 ( .A(n9278), .B(n9310), .X(n7913) );
  nand_x1_sg U51919 ( .A(n46398), .B(n9311), .X(n9310) );
  nand_x1_sg U51920 ( .A(n9278), .B(n9287), .X(n7925) );
  nand_x1_sg U51921 ( .A(n46398), .B(n9288), .X(n9287) );
  nand_x1_sg U51922 ( .A(n9278), .B(n9289), .X(n7924) );
  nand_x1_sg U51923 ( .A(n46398), .B(n9290), .X(n9289) );
  nand_x1_sg U51924 ( .A(n9278), .B(n9308), .X(n7914) );
  nand_x1_sg U51925 ( .A(n9278), .B(n9293), .X(n7922) );
  nand_x1_sg U51926 ( .A(n46398), .B(n9294), .X(n9293) );
  nand_x1_sg U51927 ( .A(n9278), .B(n9297), .X(n7920) );
  nand_x1_sg U51928 ( .A(n9278), .B(n9283), .X(n7927) );
  nand_x1_sg U51929 ( .A(n46398), .B(n9284), .X(n9283) );
  nand_x1_sg U51930 ( .A(n9278), .B(n9304), .X(n7916) );
  nand_x1_sg U51931 ( .A(n9278), .B(n9295), .X(n7921) );
  nand_x1_sg U51932 ( .A(n9278), .B(n9281), .X(n7928) );
  nand_x1_sg U51933 ( .A(n9278), .B(n9285), .X(n7926) );
  nand_x1_sg U51934 ( .A(n46398), .B(n9286), .X(n9285) );
  nand_x1_sg U51935 ( .A(n9278), .B(n9299), .X(n7919) );
  nand_x1_sg U51936 ( .A(n46398), .B(n9300), .X(n9299) );
  nand_x1_sg U51937 ( .A(n9278), .B(n9314), .X(n7911) );
  nand_x1_sg U51938 ( .A(n46398), .B(n9315), .X(n9314) );
  nand_x1_sg U51939 ( .A(n9240), .B(n9265), .X(n7936) );
  nand_x1_sg U51940 ( .A(n46371), .B(n46375), .X(n9265) );
  nand_x1_sg U51941 ( .A(n9240), .B(n9268), .X(n7934) );
  nand_x1_sg U51942 ( .A(n55789), .B(n9269), .X(n9268) );
  nand_x1_sg U51943 ( .A(n9240), .B(n9263), .X(n7937) );
  nand_x1_sg U51944 ( .A(n9240), .B(n9276), .X(n7930) );
  nand_x1_sg U51945 ( .A(n46375), .B(n9277), .X(n9276) );
  nand_x1_sg U51946 ( .A(n9240), .B(n9241), .X(n7948) );
  nand_x1_sg U51947 ( .A(n46375), .B(n9242), .X(n9241) );
  nand_x1_sg U51948 ( .A(n9240), .B(n9253), .X(n7942) );
  nand_x1_sg U51949 ( .A(n46375), .B(n9254), .X(n9253) );
  nand_x1_sg U51950 ( .A(n9240), .B(n9272), .X(n7932) );
  nand_x1_sg U51951 ( .A(n46375), .B(n9273), .X(n9272) );
  nand_x1_sg U51952 ( .A(n9240), .B(n9249), .X(n7944) );
  nand_x1_sg U51953 ( .A(n46375), .B(n9250), .X(n9249) );
  nand_x1_sg U51954 ( .A(n9240), .B(n9251), .X(n7943) );
  nand_x1_sg U51955 ( .A(n46375), .B(n9252), .X(n9251) );
  nand_x1_sg U51956 ( .A(n9240), .B(n9270), .X(n7933) );
  nand_x1_sg U51957 ( .A(n9240), .B(n9255), .X(n7941) );
  nand_x1_sg U51958 ( .A(n46375), .B(n9256), .X(n9255) );
  nand_x1_sg U51959 ( .A(n9240), .B(n9259), .X(n7939) );
  nand_x1_sg U51960 ( .A(n9240), .B(n9245), .X(n7946) );
  nand_x1_sg U51961 ( .A(n46375), .B(n9246), .X(n9245) );
  nand_x1_sg U51962 ( .A(n9240), .B(n9266), .X(n7935) );
  nand_x1_sg U51963 ( .A(n9240), .B(n9257), .X(n7940) );
  nand_x1_sg U51964 ( .A(n46375), .B(n9258), .X(n9257) );
  nand_x1_sg U51965 ( .A(n9240), .B(n9243), .X(n7947) );
  nand_x1_sg U51966 ( .A(n9240), .B(n9247), .X(n7945) );
  nand_x1_sg U51967 ( .A(n46375), .B(n9248), .X(n9247) );
  nand_x1_sg U51968 ( .A(n9240), .B(n9261), .X(n7938) );
  nand_x1_sg U51969 ( .A(n46375), .B(n9262), .X(n9261) );
  nand_x1_sg U51970 ( .A(n9240), .B(n9274), .X(n7931) );
  nand_x1_sg U51971 ( .A(n46375), .B(n9275), .X(n9274) );
  nand_x1_sg U51972 ( .A(n9050), .B(n9057), .X(n8043) );
  nand_x1_sg U51973 ( .A(n46351), .B(n44429), .X(n9057) );
  nand_x1_sg U51974 ( .A(n9050), .B(n9076), .X(n8032) );
  nand_x1_sg U51975 ( .A(n46355), .B(n9077), .X(n9076) );
  nand_x1_sg U51976 ( .A(n9050), .B(n9055), .X(n8044) );
  nand_x1_sg U51977 ( .A(n9050), .B(n9070), .X(n8036) );
  nand_x1_sg U51978 ( .A(n46355), .B(n9071), .X(n9070) );
  nand_x1_sg U51979 ( .A(n9050), .B(n9082), .X(n8029) );
  nand_x1_sg U51980 ( .A(n9050), .B(n9062), .X(n8040) );
  nand_x1_sg U51981 ( .A(n46355), .B(n9063), .X(n9062) );
  nand_x1_sg U51982 ( .A(n9050), .B(n9084), .X(n8028) );
  nand_x1_sg U51983 ( .A(n46355), .B(n9085), .X(n9084) );
  nand_x1_sg U51984 ( .A(n9050), .B(n9068), .X(n8037) );
  nand_x1_sg U51985 ( .A(n46355), .B(n9069), .X(n9068) );
  nand_x1_sg U51986 ( .A(n9050), .B(n9060), .X(n8041) );
  nand_x1_sg U51987 ( .A(n46355), .B(n9061), .X(n9060) );
  nand_x1_sg U51988 ( .A(n9050), .B(n9051), .X(n8046) );
  nand_x1_sg U51989 ( .A(n9050), .B(n9074), .X(n8033) );
  nand_x1_sg U51990 ( .A(n46355), .B(n9075), .X(n9074) );
  nand_x1_sg U51991 ( .A(n9050), .B(n9066), .X(n8038) );
  nand_x1_sg U51992 ( .A(n9050), .B(n9072), .X(n8035) );
  nand_x1_sg U51993 ( .A(n46355), .B(n9073), .X(n9072) );
  nand_x1_sg U51994 ( .A(n9050), .B(n9078), .X(n8031) );
  nand_x1_sg U51995 ( .A(n9050), .B(n9064), .X(n8039) );
  nand_x1_sg U51996 ( .A(n46355), .B(n9065), .X(n9064) );
  nand_x1_sg U51997 ( .A(n9050), .B(n9058), .X(n8042) );
  nand_x1_sg U51998 ( .A(n9050), .B(n9080), .X(n8030) );
  nand_x1_sg U51999 ( .A(n46355), .B(n9081), .X(n9080) );
  nand_x1_sg U52000 ( .A(n9050), .B(n9053), .X(n8045) );
  nand_x1_sg U52001 ( .A(n46355), .B(n9054), .X(n9053) );
  nand_x1_sg U52002 ( .A(n9050), .B(n9086), .X(n8027) );
  nand_x1_sg U52003 ( .A(n46355), .B(n9087), .X(n9086) );
  nand_x1_sg U52004 ( .A(n9202), .B(n9227), .X(n7955) );
  nand_x1_sg U52005 ( .A(n46324), .B(n46327), .X(n9227) );
  nand_x1_sg U52006 ( .A(n9202), .B(n9230), .X(n7953) );
  nand_x1_sg U52007 ( .A(n46327), .B(n9231), .X(n9230) );
  nand_x1_sg U52008 ( .A(n9202), .B(n9225), .X(n7956) );
  nand_x1_sg U52009 ( .A(n9202), .B(n9238), .X(n7949) );
  nand_x1_sg U52010 ( .A(n46327), .B(n9239), .X(n9238) );
  nand_x1_sg U52011 ( .A(n9202), .B(n9203), .X(n7967) );
  nand_x1_sg U52012 ( .A(n46327), .B(n9204), .X(n9203) );
  nand_x1_sg U52013 ( .A(n9202), .B(n9215), .X(n7961) );
  nand_x1_sg U52014 ( .A(n46327), .B(n9216), .X(n9215) );
  nand_x1_sg U52015 ( .A(n9202), .B(n9234), .X(n7951) );
  nand_x1_sg U52016 ( .A(n46327), .B(n9235), .X(n9234) );
  nand_x1_sg U52017 ( .A(n9202), .B(n9211), .X(n7963) );
  nand_x1_sg U52018 ( .A(n46327), .B(n9212), .X(n9211) );
  nand_x1_sg U52019 ( .A(n9202), .B(n9213), .X(n7962) );
  nand_x1_sg U52020 ( .A(n46327), .B(n9214), .X(n9213) );
  nand_x1_sg U52021 ( .A(n9202), .B(n9232), .X(n7952) );
  nand_x1_sg U52022 ( .A(n9202), .B(n9217), .X(n7960) );
  nand_x1_sg U52023 ( .A(n46327), .B(n9218), .X(n9217) );
  nand_x1_sg U52024 ( .A(n9202), .B(n9221), .X(n7958) );
  nand_x1_sg U52025 ( .A(n9202), .B(n9207), .X(n7965) );
  nand_x1_sg U52026 ( .A(n46327), .B(n9208), .X(n9207) );
  nand_x1_sg U52027 ( .A(n9202), .B(n9228), .X(n7954) );
  nand_x1_sg U52028 ( .A(n9202), .B(n9219), .X(n7959) );
  nand_x1_sg U52029 ( .A(n46327), .B(n9220), .X(n9219) );
  nand_x1_sg U52030 ( .A(n9202), .B(n9205), .X(n7966) );
  nand_x1_sg U52031 ( .A(n9202), .B(n9209), .X(n7964) );
  nand_x1_sg U52032 ( .A(n46327), .B(n9210), .X(n9209) );
  nand_x1_sg U52033 ( .A(n9202), .B(n9223), .X(n7957) );
  nand_x1_sg U52034 ( .A(n46327), .B(n9224), .X(n9223) );
  nand_x1_sg U52035 ( .A(n9202), .B(n9236), .X(n7950) );
  nand_x1_sg U52036 ( .A(n46327), .B(n9237), .X(n9236) );
  nand_x1_sg U52037 ( .A(n9164), .B(n9169), .X(n7985) );
  nand_x1_sg U52038 ( .A(n46306), .B(n46308), .X(n9169) );
  nand_x1_sg U52039 ( .A(n9164), .B(n9190), .X(n7973) );
  nand_x1_sg U52040 ( .A(n46308), .B(n9191), .X(n9190) );
  nand_x1_sg U52041 ( .A(n9164), .B(n9167), .X(n7986) );
  nand_x1_sg U52042 ( .A(n9164), .B(n9180), .X(n7979) );
  nand_x1_sg U52043 ( .A(n46308), .B(n9181), .X(n9180) );
  nand_x1_sg U52044 ( .A(n9164), .B(n9196), .X(n7970) );
  nand_x1_sg U52045 ( .A(n9164), .B(n9194), .X(n7971) );
  nand_x1_sg U52046 ( .A(n43856), .B(n9195), .X(n9194) );
  nand_x1_sg U52047 ( .A(n9164), .B(n9176), .X(n7981) );
  nand_x1_sg U52048 ( .A(n46308), .B(n9177), .X(n9176) );
  nand_x1_sg U52049 ( .A(n9164), .B(n9172), .X(n7983) );
  nand_x1_sg U52050 ( .A(n46308), .B(n9173), .X(n9172) );
  nand_x1_sg U52051 ( .A(n9164), .B(n9192), .X(n7972) );
  nand_x1_sg U52052 ( .A(n46308), .B(n9193), .X(n9192) );
  nand_x1_sg U52053 ( .A(n9164), .B(n9174), .X(n7982) );
  nand_x1_sg U52054 ( .A(n9164), .B(n9182), .X(n7977) );
  nand_x1_sg U52055 ( .A(n46308), .B(n9183), .X(n9182) );
  nand_x1_sg U52056 ( .A(n9164), .B(n9200), .X(n7968) );
  nand_x1_sg U52057 ( .A(n9164), .B(n9186), .X(n7975) );
  nand_x1_sg U52058 ( .A(n46308), .B(n9187), .X(n9186) );
  nand_x1_sg U52059 ( .A(n9164), .B(n9188), .X(n7974) );
  nand_x1_sg U52060 ( .A(n9164), .B(n9198), .X(n7969) );
  nand_x1_sg U52061 ( .A(n46308), .B(n9199), .X(n9198) );
  nand_x1_sg U52062 ( .A(n9164), .B(n9184), .X(n7976) );
  nand_x1_sg U52063 ( .A(n9164), .B(n9170), .X(n7984) );
  nand_x1_sg U52064 ( .A(n46308), .B(n9171), .X(n9170) );
  nand_x1_sg U52065 ( .A(n9164), .B(n9165), .X(n7987) );
  nand_x1_sg U52066 ( .A(n46308), .B(n9166), .X(n9165) );
  nand_x1_sg U52067 ( .A(n9164), .B(n9178), .X(n7980) );
  nand_x1_sg U52068 ( .A(n46308), .B(n9179), .X(n9178) );
  nand_x1_sg U52069 ( .A(n9126), .B(n9151), .X(n7995) );
  nand_x1_sg U52070 ( .A(n46279), .B(n44171), .X(n9151) );
  nand_x1_sg U52071 ( .A(n9126), .B(n9154), .X(n7993) );
  nand_x1_sg U52072 ( .A(n46283), .B(n9155), .X(n9154) );
  nand_x1_sg U52073 ( .A(n9126), .B(n9149), .X(n7996) );
  nand_x1_sg U52074 ( .A(n9126), .B(n9162), .X(n7989) );
  nand_x1_sg U52075 ( .A(n46283), .B(n9163), .X(n9162) );
  nand_x1_sg U52076 ( .A(n9126), .B(n9127), .X(n8007) );
  nand_x1_sg U52077 ( .A(n46283), .B(n9128), .X(n9127) );
  nand_x1_sg U52078 ( .A(n9126), .B(n9139), .X(n8001) );
  nand_x1_sg U52079 ( .A(n9126), .B(n9158), .X(n7991) );
  nand_x1_sg U52080 ( .A(n46283), .B(n9159), .X(n9158) );
  nand_x1_sg U52081 ( .A(n9126), .B(n9135), .X(n8003) );
  nand_x1_sg U52082 ( .A(n46283), .B(n9136), .X(n9135) );
  nand_x1_sg U52083 ( .A(n9126), .B(n9137), .X(n8002) );
  nand_x1_sg U52084 ( .A(n46283), .B(n9138), .X(n9137) );
  nand_x1_sg U52085 ( .A(n9126), .B(n9156), .X(n7992) );
  nand_x1_sg U52086 ( .A(n9126), .B(n9141), .X(n8000) );
  nand_x1_sg U52087 ( .A(n46283), .B(n9142), .X(n9141) );
  nand_x1_sg U52088 ( .A(n9126), .B(n9145), .X(n7998) );
  nand_x1_sg U52089 ( .A(n9126), .B(n9131), .X(n8005) );
  nand_x1_sg U52090 ( .A(n46283), .B(n9132), .X(n9131) );
  nand_x1_sg U52091 ( .A(n9126), .B(n9152), .X(n7994) );
  nand_x1_sg U52092 ( .A(n9126), .B(n9143), .X(n7999) );
  nand_x1_sg U52093 ( .A(n46283), .B(n9144), .X(n9143) );
  nand_x1_sg U52094 ( .A(n9126), .B(n9129), .X(n8006) );
  nand_x1_sg U52095 ( .A(n9126), .B(n9133), .X(n8004) );
  nand_x1_sg U52096 ( .A(n46283), .B(n9134), .X(n9133) );
  nand_x1_sg U52097 ( .A(n9126), .B(n9147), .X(n7997) );
  nand_x1_sg U52098 ( .A(n46283), .B(n9148), .X(n9147) );
  nand_x1_sg U52099 ( .A(n9126), .B(n9160), .X(n7990) );
  nand_x1_sg U52100 ( .A(n46283), .B(n9161), .X(n9160) );
  nand_x1_sg U52101 ( .A(n9088), .B(n9093), .X(n8024) );
  nand_x1_sg U52102 ( .A(n46261), .B(n55790), .X(n9093) );
  nand_x1_sg U52103 ( .A(n9088), .B(n9102), .X(n8019) );
  nand_x1_sg U52104 ( .A(n46263), .B(n9103), .X(n9102) );
  nand_x1_sg U52105 ( .A(n9088), .B(n9091), .X(n8025) );
  nand_x1_sg U52106 ( .A(n9088), .B(n9100), .X(n8020) );
  nand_x1_sg U52107 ( .A(n46263), .B(n9101), .X(n9100) );
  nand_x1_sg U52108 ( .A(n9088), .B(n9118), .X(n8011) );
  nand_x1_sg U52109 ( .A(n46263), .B(n9119), .X(n9118) );
  nand_x1_sg U52110 ( .A(n9088), .B(n9096), .X(n8022) );
  nand_x1_sg U52111 ( .A(n46263), .B(n9097), .X(n9096) );
  nand_x1_sg U52112 ( .A(n9088), .B(n9122), .X(n8009) );
  nand_x1_sg U52113 ( .A(n46263), .B(n9123), .X(n9122) );
  nand_x1_sg U52114 ( .A(n9088), .B(n9106), .X(n8017) );
  nand_x1_sg U52115 ( .A(n46263), .B(n9107), .X(n9106) );
  nand_x1_sg U52116 ( .A(n9088), .B(n9094), .X(n8023) );
  nand_x1_sg U52117 ( .A(n46263), .B(n9095), .X(n9094) );
  nand_x1_sg U52118 ( .A(n9088), .B(n9120), .X(n8010) );
  nand_x1_sg U52119 ( .A(n9088), .B(n9116), .X(n8012) );
  nand_x1_sg U52120 ( .A(n46263), .B(n9117), .X(n9116) );
  nand_x1_sg U52121 ( .A(n9088), .B(n9110), .X(n8015) );
  nand_x1_sg U52122 ( .A(n9088), .B(n9112), .X(n8014) );
  nand_x1_sg U52123 ( .A(n46263), .B(n9113), .X(n9112) );
  nand_x1_sg U52124 ( .A(n9088), .B(n9104), .X(n8018) );
  nand_x1_sg U52125 ( .A(n9088), .B(n9108), .X(n8016) );
  nand_x1_sg U52126 ( .A(n46263), .B(n9109), .X(n9108) );
  nand_x1_sg U52127 ( .A(n9088), .B(n9124), .X(n8008) );
  nand_x1_sg U52128 ( .A(n9088), .B(n9114), .X(n8013) );
  nand_x1_sg U52129 ( .A(n46263), .B(n9115), .X(n9114) );
  nand_x1_sg U52130 ( .A(n9088), .B(n9089), .X(n8026) );
  nand_x1_sg U52131 ( .A(n46263), .B(n9090), .X(n9089) );
  nand_x1_sg U52132 ( .A(n9088), .B(n9098), .X(n8021) );
  nand_x1_sg U52133 ( .A(n46263), .B(n9099), .X(n9098) );
  nand_x1_sg U52134 ( .A(n46237), .B(n29580), .X(\L1_0/n3506 ) );
  nand_x1_sg U52135 ( .A(n29581), .B(n55510), .X(n29580) );
  inv_x1_sg U52136 ( .A(n29579), .X(n55510) );
  nand_x1_sg U52137 ( .A(n46237), .B(n24477), .X(\L1_0/n4822 ) );
  nand_x1_sg U52138 ( .A(n24478), .B(n55491), .X(n24477) );
  inv_x1_sg U52139 ( .A(n24475), .X(n55491) );
  nand_x1_sg U52140 ( .A(n24476), .B(n24527), .X(\L1_0/n4818 ) );
  nand_x1_sg U52141 ( .A(n24528), .B(n55492), .X(n24527) );
  inv_x1_sg U52142 ( .A(n24526), .X(n55492) );
  nand_x1_sg U52143 ( .A(n46238), .B(n24576), .X(\L1_0/n4814 ) );
  nand_x1_sg U52144 ( .A(n24577), .B(n55493), .X(n24576) );
  inv_x1_sg U52145 ( .A(n24575), .X(n55493) );
  nand_x1_sg U52146 ( .A(n46237), .B(n24625), .X(\L1_0/n4810 ) );
  nand_x1_sg U52147 ( .A(n24626), .B(n55494), .X(n24625) );
  inv_x1_sg U52148 ( .A(n24624), .X(n55494) );
  nand_x1_sg U52149 ( .A(n24476), .B(n24674), .X(\L1_0/n4806 ) );
  nand_x1_sg U52150 ( .A(n24675), .B(n55495), .X(n24674) );
  inv_x1_sg U52151 ( .A(n24673), .X(n55495) );
  nand_x1_sg U52152 ( .A(n46238), .B(n24722), .X(\L1_0/n4802 ) );
  nand_x1_sg U52153 ( .A(n24723), .B(n55496), .X(n24722) );
  inv_x1_sg U52154 ( .A(n24721), .X(n55496) );
  nand_x1_sg U52155 ( .A(n46237), .B(n24770), .X(\L1_0/n4798 ) );
  nand_x1_sg U52156 ( .A(n24771), .B(n55497), .X(n24770) );
  inv_x1_sg U52157 ( .A(n24769), .X(n55497) );
  nand_x1_sg U52158 ( .A(n24476), .B(n24817), .X(\L1_0/n4794 ) );
  nand_x1_sg U52159 ( .A(n24818), .B(n55498), .X(n24817) );
  inv_x1_sg U52160 ( .A(n24816), .X(n55498) );
  nand_x1_sg U52161 ( .A(n46238), .B(n24865), .X(\L1_0/n4790 ) );
  nand_x1_sg U52162 ( .A(n24866), .B(n55499), .X(n24865) );
  inv_x1_sg U52163 ( .A(n24864), .X(n55499) );
  nand_x1_sg U52164 ( .A(n46237), .B(n24913), .X(\L1_0/n4786 ) );
  nand_x1_sg U52165 ( .A(n24914), .B(n55500), .X(n24913) );
  inv_x1_sg U52166 ( .A(n24912), .X(n55500) );
  nand_x1_sg U52167 ( .A(n24476), .B(n24961), .X(\L1_0/n4782 ) );
  nand_x1_sg U52168 ( .A(n24962), .B(n55501), .X(n24961) );
  inv_x1_sg U52169 ( .A(n24960), .X(n55501) );
  nand_x1_sg U52170 ( .A(n46238), .B(n25009), .X(\L1_0/n4778 ) );
  nand_x1_sg U52171 ( .A(n25010), .B(n55502), .X(n25009) );
  inv_x1_sg U52172 ( .A(n25008), .X(n55502) );
  nand_x1_sg U52173 ( .A(n46237), .B(n25057), .X(\L1_0/n4774 ) );
  nand_x1_sg U52174 ( .A(n25058), .B(n55503), .X(n25057) );
  inv_x1_sg U52175 ( .A(n25056), .X(n55503) );
  nand_x1_sg U52176 ( .A(n24476), .B(n25106), .X(\L1_0/n4770 ) );
  nand_x1_sg U52177 ( .A(n25107), .B(n55504), .X(n25106) );
  inv_x1_sg U52178 ( .A(n25105), .X(n55504) );
  nand_x1_sg U52179 ( .A(n46238), .B(n25154), .X(\L1_0/n4766 ) );
  nand_x1_sg U52180 ( .A(n25155), .B(n55505), .X(n25154) );
  inv_x1_sg U52181 ( .A(n25153), .X(n55505) );
  nand_x1_sg U52182 ( .A(n46237), .B(n25203), .X(\L1_0/n4762 ) );
  nand_x1_sg U52183 ( .A(n25204), .B(n55506), .X(n25203) );
  inv_x1_sg U52184 ( .A(n25202), .X(n55506) );
  nand_x1_sg U52185 ( .A(n24476), .B(n25252), .X(\L1_0/n4758 ) );
  nand_x1_sg U52186 ( .A(n25253), .B(n55507), .X(n25252) );
  inv_x1_sg U52187 ( .A(n25251), .X(n55507) );
  nand_x1_sg U52188 ( .A(n46238), .B(n25299), .X(\L1_0/n4754 ) );
  nand_x1_sg U52189 ( .A(n25300), .B(n55508), .X(n25299) );
  inv_x1_sg U52190 ( .A(n25298), .X(n55508) );
  nand_x1_sg U52191 ( .A(n46237), .B(n25342), .X(\L1_0/n4750 ) );
  nand_x1_sg U52192 ( .A(n25343), .B(n55509), .X(n25342) );
  inv_x1_sg U52193 ( .A(n25341), .X(n55509) );
  nand_x1_sg U52194 ( .A(n24476), .B(n25387), .X(\L1_0/n4746 ) );
  nand_x1_sg U52195 ( .A(n46573), .B(n25388), .X(n25387) );
  nand_x1_sg U52196 ( .A(n46238), .B(n25517), .X(\L1_0/n4670 ) );
  nand_x1_sg U52197 ( .A(n25518), .B(n25388), .X(n25517) );
  nand_x1_sg U52198 ( .A(n39304), .B(n39305), .X(n2002) );
  nand_x1_sg U52199 ( .A(model), .B(n46626), .X(n39304) );
  nand_x1_sg U52200 ( .A(n46648), .B(n46672), .X(n39305) );
  nand_x1_sg U52201 ( .A(n39308), .B(n39309), .X(n2001) );
  nand_x1_sg U52202 ( .A(\yHat[0][0] ), .B(n46632), .X(n39308) );
  nand_x1_sg U52203 ( .A(n39310), .B(n39311), .X(n2000) );
  nand_x1_sg U52204 ( .A(\yHat[0][1] ), .B(n46626), .X(n39310) );
  nand_x1_sg U52205 ( .A(n39312), .B(n39313), .X(n1999) );
  nand_x1_sg U52206 ( .A(\yHat[0][2] ), .B(n46635), .X(n39312) );
  nand_x1_sg U52207 ( .A(n39314), .B(n39315), .X(n1998) );
  nand_x1_sg U52208 ( .A(\yHat[0][3] ), .B(n46634), .X(n39314) );
  nand_x1_sg U52209 ( .A(n39316), .B(n39317), .X(n1997) );
  nand_x1_sg U52210 ( .A(\yHat[0][4] ), .B(n46631), .X(n39316) );
  nand_x1_sg U52211 ( .A(n39318), .B(n39319), .X(n1996) );
  nand_x1_sg U52212 ( .A(\yHat[0][5] ), .B(n40524), .X(n39318) );
  nand_x1_sg U52213 ( .A(n39320), .B(n39321), .X(n1995) );
  nand_x1_sg U52214 ( .A(\yHat[0][6] ), .B(n46635), .X(n39320) );
  nand_x1_sg U52215 ( .A(n39322), .B(n39323), .X(n1994) );
  nand_x1_sg U52216 ( .A(\yHat[0][7] ), .B(n46634), .X(n39322) );
  nand_x1_sg U52217 ( .A(n39324), .B(n39325), .X(n1993) );
  nand_x1_sg U52218 ( .A(\yHat[0][8] ), .B(n40523), .X(n39324) );
  nand_x1_sg U52219 ( .A(n39326), .B(n39327), .X(n1992) );
  nand_x1_sg U52220 ( .A(\yHat[0][9] ), .B(n46626), .X(n39326) );
  nand_x1_sg U52221 ( .A(n39328), .B(n39329), .X(n1991) );
  nand_x1_sg U52222 ( .A(\yHat[0][10] ), .B(n46626), .X(n39328) );
  nand_x1_sg U52223 ( .A(n39330), .B(n39331), .X(n1990) );
  nand_x1_sg U52224 ( .A(\yHat[0][11] ), .B(n46632), .X(n39330) );
  nand_x1_sg U52225 ( .A(n39332), .B(n39333), .X(n1989) );
  nand_x1_sg U52226 ( .A(\yHat[0][12] ), .B(n46634), .X(n39332) );
  nand_x1_sg U52227 ( .A(n39334), .B(n39335), .X(n1988) );
  nand_x1_sg U52228 ( .A(\yHat[0][13] ), .B(n40524), .X(n39334) );
  nand_x1_sg U52229 ( .A(n39336), .B(n39337), .X(n1987) );
  nand_x1_sg U52230 ( .A(\yHat[0][14] ), .B(n46626), .X(n39336) );
  nand_x1_sg U52231 ( .A(n39338), .B(n39339), .X(n1986) );
  nand_x1_sg U52232 ( .A(\yHat[0][15] ), .B(n46632), .X(n39338) );
  nand_x1_sg U52233 ( .A(n39340), .B(n39341), .X(n1985) );
  nand_x1_sg U52234 ( .A(\yHat[0][16] ), .B(n40521), .X(n39340) );
  nand_x1_sg U52235 ( .A(n39342), .B(n39343), .X(n1984) );
  nand_x1_sg U52236 ( .A(\yHat[0][17] ), .B(n46626), .X(n39342) );
  nand_x1_sg U52237 ( .A(n39344), .B(n39345), .X(n1983) );
  nand_x1_sg U52238 ( .A(\yHat[0][18] ), .B(n46635), .X(n39344) );
  nand_x1_sg U52239 ( .A(n39346), .B(n39347), .X(n1982) );
  nand_x1_sg U52240 ( .A(\yHat[0][19] ), .B(n46634), .X(n39346) );
  nand_x1_sg U52241 ( .A(n39348), .B(n39349), .X(n1981) );
  nand_x1_sg U52242 ( .A(\yHat[1][0] ), .B(n40523), .X(n39348) );
  nand_x1_sg U52243 ( .A(n39350), .B(n39351), .X(n1980) );
  nand_x1_sg U52244 ( .A(\yHat[1][1] ), .B(n46626), .X(n39350) );
  nand_x1_sg U52245 ( .A(n39352), .B(n39353), .X(n1979) );
  nand_x1_sg U52246 ( .A(\yHat[1][2] ), .B(n46634), .X(n39352) );
  nand_x1_sg U52247 ( .A(n39354), .B(n39355), .X(n1978) );
  nand_x1_sg U52248 ( .A(\yHat[1][3] ), .B(n46632), .X(n39354) );
  nand_x1_sg U52249 ( .A(n39356), .B(n39357), .X(n1977) );
  nand_x1_sg U52250 ( .A(\yHat[1][4] ), .B(n46631), .X(n39356) );
  nand_x1_sg U52251 ( .A(n39358), .B(n39359), .X(n1976) );
  nand_x1_sg U52252 ( .A(\yHat[1][5] ), .B(n46632), .X(n39358) );
  nand_x1_sg U52253 ( .A(n39360), .B(n39361), .X(n1975) );
  nand_x1_sg U52254 ( .A(\yHat[1][6] ), .B(n40524), .X(n39360) );
  nand_x1_sg U52255 ( .A(n39362), .B(n39363), .X(n1974) );
  nand_x1_sg U52256 ( .A(\yHat[1][7] ), .B(n46635), .X(n39362) );
  nand_x1_sg U52257 ( .A(n39364), .B(n39365), .X(n1973) );
  nand_x1_sg U52258 ( .A(\yHat[1][8] ), .B(n40520), .X(n39364) );
  nand_x1_sg U52259 ( .A(n39366), .B(n39367), .X(n1972) );
  nand_x1_sg U52260 ( .A(\yHat[1][9] ), .B(n40523), .X(n39366) );
  nand_x1_sg U52261 ( .A(n39368), .B(n39369), .X(n1971) );
  nand_x1_sg U52262 ( .A(\yHat[1][10] ), .B(n46634), .X(n39368) );
  nand_x1_sg U52263 ( .A(n39370), .B(n39371), .X(n1970) );
  nand_x1_sg U52264 ( .A(\yHat[1][11] ), .B(n46635), .X(n39370) );
  nand_x1_sg U52265 ( .A(n39372), .B(n39373), .X(n1969) );
  nand_x1_sg U52266 ( .A(\yHat[1][12] ), .B(n46634), .X(n39372) );
  nand_x1_sg U52267 ( .A(n39374), .B(n39375), .X(n1968) );
  nand_x1_sg U52268 ( .A(\yHat[1][13] ), .B(n46635), .X(n39374) );
  nand_x1_sg U52269 ( .A(n39376), .B(n39377), .X(n1967) );
  nand_x1_sg U52270 ( .A(\yHat[1][14] ), .B(n46634), .X(n39376) );
  nand_x1_sg U52271 ( .A(n39378), .B(n39379), .X(n1966) );
  nand_x1_sg U52272 ( .A(\yHat[1][15] ), .B(n40524), .X(n39378) );
  nand_x1_sg U52273 ( .A(n39380), .B(n39381), .X(n1965) );
  nand_x1_sg U52274 ( .A(\yHat[1][16] ), .B(n46631), .X(n39380) );
  nand_x1_sg U52275 ( .A(n39382), .B(n39383), .X(n1964) );
  nand_x1_sg U52276 ( .A(\yHat[1][17] ), .B(n46634), .X(n39382) );
  nand_x1_sg U52277 ( .A(n39384), .B(n39385), .X(n1963) );
  nand_x1_sg U52278 ( .A(\yHat[1][18] ), .B(n46635), .X(n39384) );
  nand_x1_sg U52279 ( .A(n39386), .B(n39387), .X(n1962) );
  nand_x1_sg U52280 ( .A(\yHat[1][19] ), .B(n46626), .X(n39386) );
  nand_x1_sg U52281 ( .A(n39388), .B(n39389), .X(n1961) );
  nand_x1_sg U52282 ( .A(\yHat[2][0] ), .B(n46634), .X(n39388) );
  nand_x1_sg U52283 ( .A(n39390), .B(n39391), .X(n1960) );
  nand_x1_sg U52284 ( .A(\yHat[2][1] ), .B(n46634), .X(n39390) );
  nand_x1_sg U52285 ( .A(n39392), .B(n39393), .X(n1959) );
  nand_x1_sg U52286 ( .A(\yHat[2][2] ), .B(n40521), .X(n39392) );
  nand_x1_sg U52287 ( .A(n39394), .B(n39395), .X(n1958) );
  nand_x1_sg U52288 ( .A(\yHat[2][3] ), .B(n46631), .X(n39394) );
  nand_x1_sg U52289 ( .A(n39396), .B(n39397), .X(n1957) );
  nand_x1_sg U52290 ( .A(\yHat[2][4] ), .B(n46631), .X(n39396) );
  nand_x1_sg U52291 ( .A(n39398), .B(n39399), .X(n1956) );
  nand_x1_sg U52292 ( .A(\yHat[2][5] ), .B(n40521), .X(n39398) );
  nand_x1_sg U52293 ( .A(n39400), .B(n39401), .X(n1955) );
  nand_x1_sg U52294 ( .A(\yHat[2][6] ), .B(n46634), .X(n39400) );
  nand_x1_sg U52295 ( .A(n39402), .B(n39403), .X(n1954) );
  nand_x1_sg U52296 ( .A(\yHat[2][7] ), .B(n46635), .X(n39402) );
  nand_x1_sg U52297 ( .A(n39404), .B(n39405), .X(n1953) );
  nand_x1_sg U52298 ( .A(\yHat[2][8] ), .B(n46632), .X(n39404) );
  nand_x1_sg U52299 ( .A(n39406), .B(n39407), .X(n1952) );
  nand_x1_sg U52300 ( .A(\yHat[2][9] ), .B(n40523), .X(n39406) );
  nand_x1_sg U52301 ( .A(n39408), .B(n39409), .X(n1951) );
  nand_x1_sg U52302 ( .A(\yHat[2][10] ), .B(n46632), .X(n39408) );
  nand_x1_sg U52303 ( .A(n39410), .B(n39411), .X(n1950) );
  nand_x1_sg U52304 ( .A(\yHat[2][11] ), .B(n46626), .X(n39410) );
  nand_x1_sg U52305 ( .A(n39412), .B(n39413), .X(n1949) );
  nand_x1_sg U52306 ( .A(\yHat[2][12] ), .B(n46626), .X(n39412) );
  nand_x1_sg U52307 ( .A(n39414), .B(n39415), .X(n1948) );
  nand_x1_sg U52308 ( .A(\yHat[2][13] ), .B(n46632), .X(n39414) );
  nand_x1_sg U52309 ( .A(n39416), .B(n39417), .X(n1947) );
  nand_x1_sg U52310 ( .A(\yHat[2][14] ), .B(n40523), .X(n39416) );
  nand_x1_sg U52311 ( .A(n39418), .B(n39419), .X(n1946) );
  nand_x1_sg U52312 ( .A(\yHat[2][15] ), .B(n40523), .X(n39418) );
  nand_x1_sg U52313 ( .A(n39420), .B(n39421), .X(n1945) );
  nand_x1_sg U52314 ( .A(\yHat[2][16] ), .B(n46631), .X(n39420) );
  nand_x1_sg U52315 ( .A(n39422), .B(n39423), .X(n1944) );
  nand_x1_sg U52316 ( .A(\yHat[2][17] ), .B(n46635), .X(n39422) );
  nand_x1_sg U52317 ( .A(n39424), .B(n39425), .X(n1943) );
  nand_x1_sg U52318 ( .A(\yHat[2][18] ), .B(n46634), .X(n39424) );
  nand_x1_sg U52319 ( .A(n39426), .B(n39427), .X(n1942) );
  nand_x1_sg U52320 ( .A(\yHat[2][19] ), .B(n46635), .X(n39426) );
  nand_x1_sg U52321 ( .A(n39428), .B(n39429), .X(n1941) );
  nand_x1_sg U52322 ( .A(\yHat[3][0] ), .B(n46626), .X(n39428) );
  nand_x1_sg U52323 ( .A(n39430), .B(n39431), .X(n1940) );
  nand_x1_sg U52324 ( .A(\yHat[3][1] ), .B(n46635), .X(n39430) );
  nand_x1_sg U52325 ( .A(n39432), .B(n39433), .X(n1939) );
  nand_x1_sg U52326 ( .A(\yHat[3][2] ), .B(n46635), .X(n39432) );
  nand_x1_sg U52327 ( .A(n39434), .B(n39435), .X(n1938) );
  nand_x1_sg U52328 ( .A(\yHat[3][3] ), .B(n40524), .X(n39434) );
  nand_x1_sg U52329 ( .A(n39436), .B(n39437), .X(n1937) );
  nand_x1_sg U52330 ( .A(\yHat[3][4] ), .B(n40524), .X(n39436) );
  nand_x1_sg U52331 ( .A(n39438), .B(n39439), .X(n1936) );
  nand_x1_sg U52332 ( .A(\yHat[3][5] ), .B(n46632), .X(n39438) );
  nand_x1_sg U52333 ( .A(n39440), .B(n39441), .X(n1935) );
  nand_x1_sg U52334 ( .A(\yHat[3][6] ), .B(n46635), .X(n39440) );
  nand_x1_sg U52335 ( .A(n39442), .B(n39443), .X(n1934) );
  nand_x1_sg U52336 ( .A(\yHat[3][7] ), .B(n46626), .X(n39442) );
  nand_x1_sg U52337 ( .A(n39444), .B(n39445), .X(n1933) );
  nand_x1_sg U52338 ( .A(\yHat[3][8] ), .B(n46634), .X(n39444) );
  nand_x1_sg U52339 ( .A(n39446), .B(n39447), .X(n1932) );
  nand_x1_sg U52340 ( .A(\yHat[3][9] ), .B(n40524), .X(n39446) );
  nand_x1_sg U52341 ( .A(n39448), .B(n39449), .X(n1931) );
  nand_x1_sg U52342 ( .A(\yHat[3][10] ), .B(n46632), .X(n39448) );
  nand_x1_sg U52343 ( .A(n39450), .B(n39451), .X(n1930) );
  nand_x1_sg U52344 ( .A(\yHat[3][11] ), .B(n46635), .X(n39450) );
  nand_x1_sg U52345 ( .A(n39452), .B(n39453), .X(n1929) );
  nand_x1_sg U52346 ( .A(\yHat[3][12] ), .B(n40520), .X(n39452) );
  nand_x1_sg U52347 ( .A(n39454), .B(n39455), .X(n1928) );
  nand_x1_sg U52348 ( .A(\yHat[3][13] ), .B(n46631), .X(n39454) );
  nand_x1_sg U52349 ( .A(n39456), .B(n39457), .X(n1927) );
  nand_x1_sg U52350 ( .A(\yHat[3][14] ), .B(n46634), .X(n39456) );
  nand_x1_sg U52351 ( .A(n39458), .B(n39459), .X(n1926) );
  nand_x1_sg U52352 ( .A(\yHat[3][15] ), .B(n46635), .X(n39458) );
  nand_x1_sg U52353 ( .A(n39460), .B(n39461), .X(n1925) );
  nand_x1_sg U52354 ( .A(\yHat[3][16] ), .B(n40523), .X(n39460) );
  nand_x1_sg U52355 ( .A(n39462), .B(n39463), .X(n1924) );
  nand_x1_sg U52356 ( .A(\yHat[3][17] ), .B(n46626), .X(n39462) );
  nand_x1_sg U52357 ( .A(n39464), .B(n39465), .X(n1923) );
  nand_x1_sg U52358 ( .A(\yHat[3][18] ), .B(n46632), .X(n39464) );
  nand_x1_sg U52359 ( .A(n39466), .B(n39467), .X(n1922) );
  nand_x1_sg U52360 ( .A(\yHat[3][19] ), .B(n40521), .X(n39466) );
  nand_x1_sg U52361 ( .A(n39468), .B(n39469), .X(n1921) );
  nand_x1_sg U52362 ( .A(\yHat[4][0] ), .B(n46634), .X(n39468) );
  nand_x1_sg U52363 ( .A(n39470), .B(n39471), .X(n1920) );
  nand_x1_sg U52364 ( .A(\yHat[4][1] ), .B(n40521), .X(n39470) );
  nand_x1_sg U52365 ( .A(n39472), .B(n39473), .X(n1919) );
  nand_x1_sg U52366 ( .A(\yHat[4][2] ), .B(n46631), .X(n39472) );
  nand_x1_sg U52367 ( .A(n39474), .B(n39475), .X(n1918) );
  nand_x1_sg U52368 ( .A(\yHat[4][3] ), .B(n46626), .X(n39474) );
  nand_x1_sg U52369 ( .A(n39476), .B(n39477), .X(n1917) );
  nand_x1_sg U52370 ( .A(\yHat[4][4] ), .B(n46632), .X(n39476) );
  nand_x1_sg U52371 ( .A(n39478), .B(n39479), .X(n1916) );
  nand_x1_sg U52372 ( .A(\yHat[4][5] ), .B(n40520), .X(n39478) );
  nand_x1_sg U52373 ( .A(n39480), .B(n39481), .X(n1915) );
  nand_x1_sg U52374 ( .A(\yHat[4][6] ), .B(n46635), .X(n39480) );
  nand_x1_sg U52375 ( .A(n39482), .B(n39483), .X(n1914) );
  nand_x1_sg U52376 ( .A(\yHat[4][7] ), .B(n40524), .X(n39482) );
  nand_x1_sg U52377 ( .A(n39484), .B(n39485), .X(n1913) );
  nand_x1_sg U52378 ( .A(\yHat[4][8] ), .B(n46631), .X(n39484) );
  nand_x1_sg U52379 ( .A(n39486), .B(n39487), .X(n1912) );
  nand_x1_sg U52380 ( .A(\yHat[4][9] ), .B(n46631), .X(n39486) );
  nand_x1_sg U52381 ( .A(n39488), .B(n39489), .X(n1911) );
  nand_x1_sg U52382 ( .A(\yHat[4][10] ), .B(n46634), .X(n39488) );
  nand_x1_sg U52383 ( .A(n39490), .B(n39491), .X(n1910) );
  nand_x1_sg U52384 ( .A(\yHat[4][11] ), .B(n46635), .X(n39490) );
  nand_x1_sg U52385 ( .A(n39492), .B(n39493), .X(n1909) );
  nand_x1_sg U52386 ( .A(\yHat[4][12] ), .B(n40523), .X(n39492) );
  nand_x1_sg U52387 ( .A(n39494), .B(n39495), .X(n1908) );
  nand_x1_sg U52388 ( .A(\yHat[4][13] ), .B(n46626), .X(n39494) );
  nand_x1_sg U52389 ( .A(n39496), .B(n39497), .X(n1907) );
  nand_x1_sg U52390 ( .A(\yHat[4][14] ), .B(n46632), .X(n39496) );
  nand_x1_sg U52391 ( .A(n39498), .B(n39499), .X(n1906) );
  nand_x1_sg U52392 ( .A(\yHat[4][15] ), .B(n46634), .X(n39498) );
  nand_x1_sg U52393 ( .A(n39500), .B(n39501), .X(n1905) );
  nand_x1_sg U52394 ( .A(\yHat[4][16] ), .B(n40520), .X(n39500) );
  nand_x1_sg U52395 ( .A(n39502), .B(n39503), .X(n1904) );
  nand_x1_sg U52396 ( .A(\yHat[4][17] ), .B(n46631), .X(n39502) );
  nand_x1_sg U52397 ( .A(n39504), .B(n39505), .X(n1903) );
  nand_x1_sg U52398 ( .A(\yHat[4][18] ), .B(n46634), .X(n39504) );
  nand_x1_sg U52399 ( .A(n39506), .B(n39507), .X(n1902) );
  nand_x1_sg U52400 ( .A(\yHat[4][19] ), .B(n40523), .X(n39506) );
  nand_x1_sg U52401 ( .A(n39508), .B(n39509), .X(n1901) );
  nand_x1_sg U52402 ( .A(\yHat[5][0] ), .B(n46631), .X(n39508) );
  nand_x1_sg U52403 ( .A(n39510), .B(n39511), .X(n1900) );
  nand_x1_sg U52404 ( .A(\yHat[5][1] ), .B(n46631), .X(n39510) );
  nand_x1_sg U52405 ( .A(n39512), .B(n39513), .X(n1899) );
  nand_x1_sg U52406 ( .A(\yHat[5][2] ), .B(n40520), .X(n39512) );
  nand_x1_sg U52407 ( .A(n39514), .B(n39515), .X(n1898) );
  nand_x1_sg U52408 ( .A(\yHat[5][3] ), .B(n40521), .X(n39514) );
  nand_x1_sg U52409 ( .A(n39516), .B(n39517), .X(n1897) );
  nand_x1_sg U52410 ( .A(\yHat[5][4] ), .B(n46631), .X(n39516) );
  nand_x1_sg U52411 ( .A(n39518), .B(n39519), .X(n1896) );
  nand_x1_sg U52412 ( .A(\yHat[5][5] ), .B(n46635), .X(n39518) );
  nand_x1_sg U52413 ( .A(n39520), .B(n39521), .X(n1895) );
  nand_x1_sg U52414 ( .A(\yHat[5][6] ), .B(n46634), .X(n39520) );
  nand_x1_sg U52415 ( .A(n39522), .B(n39523), .X(n1894) );
  nand_x1_sg U52416 ( .A(\yHat[5][7] ), .B(n40524), .X(n39522) );
  nand_x1_sg U52417 ( .A(n39524), .B(n39525), .X(n1893) );
  nand_x1_sg U52418 ( .A(\yHat[5][8] ), .B(n40521), .X(n39524) );
  nand_x1_sg U52419 ( .A(n39526), .B(n39527), .X(n1892) );
  nand_x1_sg U52420 ( .A(\yHat[5][9] ), .B(n46631), .X(n39526) );
  nand_x1_sg U52421 ( .A(n39528), .B(n39529), .X(n1891) );
  nand_x1_sg U52422 ( .A(\yHat[5][10] ), .B(n46626), .X(n39528) );
  nand_x1_sg U52423 ( .A(n39530), .B(n39531), .X(n1890) );
  nand_x1_sg U52424 ( .A(\yHat[5][11] ), .B(n46632), .X(n39530) );
  nand_x1_sg U52425 ( .A(n39532), .B(n39533), .X(n1889) );
  nand_x1_sg U52426 ( .A(\yHat[5][12] ), .B(n40524), .X(n39532) );
  nand_x1_sg U52427 ( .A(n39534), .B(n39535), .X(n1888) );
  nand_x1_sg U52428 ( .A(\yHat[5][13] ), .B(n46635), .X(n39534) );
  nand_x1_sg U52429 ( .A(n39536), .B(n39537), .X(n1887) );
  nand_x1_sg U52430 ( .A(\yHat[5][14] ), .B(n46634), .X(n39536) );
  nand_x1_sg U52431 ( .A(n39538), .B(n39539), .X(n1886) );
  nand_x1_sg U52432 ( .A(\yHat[5][15] ), .B(n46632), .X(n39538) );
  nand_x1_sg U52433 ( .A(n39540), .B(n39541), .X(n1885) );
  nand_x1_sg U52434 ( .A(\yHat[5][16] ), .B(n46631), .X(n39540) );
  nand_x1_sg U52435 ( .A(n39542), .B(n39543), .X(n1884) );
  nand_x1_sg U52436 ( .A(\yHat[5][17] ), .B(n46631), .X(n39542) );
  nand_x1_sg U52437 ( .A(n39544), .B(n39545), .X(n1883) );
  nand_x1_sg U52438 ( .A(\yHat[5][18] ), .B(n46626), .X(n39544) );
  nand_x1_sg U52439 ( .A(n39546), .B(n39547), .X(n1882) );
  nand_x1_sg U52440 ( .A(\yHat[5][19] ), .B(n40520), .X(n39546) );
  nand_x1_sg U52441 ( .A(n39548), .B(n39549), .X(n1881) );
  nand_x1_sg U52442 ( .A(\yHat[6][0] ), .B(n46631), .X(n39548) );
  nand_x1_sg U52443 ( .A(n39550), .B(n39551), .X(n1880) );
  nand_x1_sg U52444 ( .A(\yHat[6][1] ), .B(n40520), .X(n39550) );
  nand_x1_sg U52445 ( .A(n39552), .B(n39553), .X(n1879) );
  nand_x1_sg U52446 ( .A(\yHat[6][2] ), .B(n46631), .X(n39552) );
  nand_x1_sg U52447 ( .A(n39554), .B(n39555), .X(n1878) );
  nand_x1_sg U52448 ( .A(\yHat[6][3] ), .B(n46632), .X(n39554) );
  nand_x1_sg U52449 ( .A(n39556), .B(n39557), .X(n1877) );
  nand_x1_sg U52450 ( .A(\yHat[6][4] ), .B(n46626), .X(n39556) );
  nand_x1_sg U52451 ( .A(n39558), .B(n39559), .X(n1876) );
  nand_x1_sg U52452 ( .A(\yHat[6][5] ), .B(n46632), .X(n39558) );
  nand_x1_sg U52453 ( .A(n39560), .B(n39561), .X(n1875) );
  nand_x1_sg U52454 ( .A(\yHat[6][6] ), .B(n46635), .X(n39560) );
  nand_x1_sg U52455 ( .A(n39562), .B(n39563), .X(n1874) );
  nand_x1_sg U52456 ( .A(\yHat[6][7] ), .B(n46634), .X(n39562) );
  nand_x1_sg U52457 ( .A(n39564), .B(n39565), .X(n1873) );
  nand_x1_sg U52458 ( .A(\yHat[6][8] ), .B(n46626), .X(n39564) );
  nand_x1_sg U52459 ( .A(n39566), .B(n39567), .X(n1872) );
  nand_x1_sg U52460 ( .A(\yHat[6][9] ), .B(n46632), .X(n39566) );
  nand_x1_sg U52461 ( .A(n39568), .B(n39569), .X(n1871) );
  nand_x1_sg U52462 ( .A(\yHat[6][10] ), .B(n46626), .X(n39568) );
  nand_x1_sg U52463 ( .A(n39570), .B(n39571), .X(n1870) );
  nand_x1_sg U52464 ( .A(\yHat[6][11] ), .B(n40520), .X(n39570) );
  nand_x1_sg U52465 ( .A(n39572), .B(n39573), .X(n1869) );
  nand_x1_sg U52466 ( .A(\yHat[6][12] ), .B(n40523), .X(n39572) );
  nand_x1_sg U52467 ( .A(n39574), .B(n39575), .X(n1868) );
  nand_x1_sg U52468 ( .A(\yHat[6][13] ), .B(n46634), .X(n39574) );
  nand_x1_sg U52469 ( .A(n39576), .B(n39577), .X(n1867) );
  nand_x1_sg U52470 ( .A(\yHat[6][14] ), .B(n46626), .X(n39576) );
  nand_x1_sg U52471 ( .A(n39578), .B(n39579), .X(n1866) );
  nand_x1_sg U52472 ( .A(\yHat[6][15] ), .B(n46632), .X(n39578) );
  nand_x1_sg U52473 ( .A(n39580), .B(n39581), .X(n1865) );
  nand_x1_sg U52474 ( .A(\yHat[6][16] ), .B(n46634), .X(n39580) );
  nand_x1_sg U52475 ( .A(n39582), .B(n39583), .X(n1864) );
  nand_x1_sg U52476 ( .A(\yHat[6][17] ), .B(n40520), .X(n39582) );
  nand_x1_sg U52477 ( .A(n39584), .B(n39585), .X(n1863) );
  nand_x1_sg U52478 ( .A(\yHat[6][18] ), .B(n46631), .X(n39584) );
  nand_x1_sg U52479 ( .A(n39586), .B(n39587), .X(n1862) );
  nand_x1_sg U52480 ( .A(\yHat[6][19] ), .B(n40521), .X(n39586) );
  nand_x1_sg U52481 ( .A(n39588), .B(n39589), .X(n1861) );
  nand_x1_sg U52482 ( .A(\yHat[7][0] ), .B(n46626), .X(n39588) );
  nand_x1_sg U52483 ( .A(n39590), .B(n39591), .X(n1860) );
  nand_x1_sg U52484 ( .A(\yHat[7][1] ), .B(n40524), .X(n39590) );
  nand_x1_sg U52485 ( .A(n39592), .B(n39593), .X(n1859) );
  nand_x1_sg U52486 ( .A(\yHat[7][2] ), .B(n40520), .X(n39592) );
  nand_x1_sg U52487 ( .A(n39594), .B(n39595), .X(n1858) );
  nand_x1_sg U52488 ( .A(\yHat[7][3] ), .B(n46631), .X(n39594) );
  nand_x1_sg U52489 ( .A(n39596), .B(n39597), .X(n1857) );
  nand_x1_sg U52490 ( .A(\yHat[7][4] ), .B(n46626), .X(n39596) );
  nand_x1_sg U52491 ( .A(n39598), .B(n39599), .X(n1856) );
  nand_x1_sg U52492 ( .A(\yHat[7][5] ), .B(n46626), .X(n39598) );
  nand_x1_sg U52493 ( .A(n39600), .B(n39601), .X(n1855) );
  nand_x1_sg U52494 ( .A(\yHat[7][6] ), .B(n40521), .X(n39600) );
  nand_x1_sg U52495 ( .A(n39602), .B(n39603), .X(n1854) );
  nand_x1_sg U52496 ( .A(\yHat[7][7] ), .B(n40520), .X(n39602) );
  nand_x1_sg U52497 ( .A(n39604), .B(n39605), .X(n1853) );
  nand_x1_sg U52498 ( .A(\yHat[7][8] ), .B(n46635), .X(n39604) );
  nand_x1_sg U52499 ( .A(n39606), .B(n39607), .X(n1852) );
  nand_x1_sg U52500 ( .A(\yHat[7][9] ), .B(n46632), .X(n39606) );
  nand_x1_sg U52501 ( .A(n39608), .B(n39609), .X(n1851) );
  nand_x1_sg U52502 ( .A(\yHat[7][10] ), .B(n46635), .X(n39608) );
  nand_x1_sg U52503 ( .A(n39610), .B(n39611), .X(n1850) );
  nand_x1_sg U52504 ( .A(\yHat[7][11] ), .B(n46626), .X(n39610) );
  nand_x1_sg U52505 ( .A(n39612), .B(n39613), .X(n1849) );
  nand_x1_sg U52506 ( .A(\yHat[7][12] ), .B(n40520), .X(n39612) );
  nand_x1_sg U52507 ( .A(n39614), .B(n39615), .X(n1848) );
  nand_x1_sg U52508 ( .A(\yHat[7][13] ), .B(n46626), .X(n39614) );
  nand_x1_sg U52509 ( .A(n39616), .B(n39617), .X(n1847) );
  nand_x1_sg U52510 ( .A(\yHat[7][14] ), .B(n46640), .X(n39616) );
  nand_x1_sg U52511 ( .A(n39618), .B(n39619), .X(n1846) );
  nand_x1_sg U52512 ( .A(\yHat[7][15] ), .B(n40524), .X(n39618) );
  nand_x1_sg U52513 ( .A(n39620), .B(n39621), .X(n1845) );
  nand_x1_sg U52514 ( .A(\yHat[7][16] ), .B(n46632), .X(n39620) );
  nand_x1_sg U52515 ( .A(n39622), .B(n39623), .X(n1844) );
  nand_x1_sg U52516 ( .A(\yHat[7][17] ), .B(n46634), .X(n39622) );
  nand_x1_sg U52517 ( .A(n39624), .B(n39625), .X(n1843) );
  nand_x1_sg U52518 ( .A(\yHat[7][18] ), .B(n46631), .X(n39624) );
  nand_x1_sg U52519 ( .A(n39626), .B(n39627), .X(n1842) );
  nand_x1_sg U52520 ( .A(\yHat[7][19] ), .B(n46634), .X(n39626) );
  nand_x1_sg U52521 ( .A(n39628), .B(n39629), .X(n1841) );
  nand_x1_sg U52522 ( .A(\yHat[8][0] ), .B(n46632), .X(n39628) );
  nand_x1_sg U52523 ( .A(n39630), .B(n39631), .X(n1840) );
  nand_x1_sg U52524 ( .A(\yHat[8][1] ), .B(n46638), .X(n39630) );
  nand_x1_sg U52525 ( .A(n39632), .B(n39633), .X(n1839) );
  nand_x1_sg U52526 ( .A(\yHat[8][2] ), .B(n46632), .X(n39632) );
  nand_x1_sg U52527 ( .A(n39634), .B(n39635), .X(n1838) );
  nand_x1_sg U52528 ( .A(\yHat[8][3] ), .B(n40521), .X(n39634) );
  nand_x1_sg U52529 ( .A(n39636), .B(n39637), .X(n1837) );
  nand_x1_sg U52530 ( .A(\yHat[8][4] ), .B(n46638), .X(n39636) );
  nand_x1_sg U52531 ( .A(n39638), .B(n39639), .X(n1836) );
  nand_x1_sg U52532 ( .A(\yHat[8][5] ), .B(n46632), .X(n39638) );
  nand_x1_sg U52533 ( .A(n39640), .B(n39641), .X(n1835) );
  nand_x1_sg U52534 ( .A(\yHat[8][6] ), .B(n46626), .X(n39640) );
  nand_x1_sg U52535 ( .A(n39642), .B(n39643), .X(n1834) );
  nand_x1_sg U52536 ( .A(\yHat[8][7] ), .B(n46626), .X(n39642) );
  nand_x1_sg U52537 ( .A(n39644), .B(n39645), .X(n1833) );
  nand_x1_sg U52538 ( .A(\yHat[8][8] ), .B(n46626), .X(n39644) );
  nand_x1_sg U52539 ( .A(n39646), .B(n39647), .X(n1832) );
  nand_x1_sg U52540 ( .A(\yHat[8][9] ), .B(n46626), .X(n39646) );
  nand_x1_sg U52541 ( .A(n39648), .B(n39649), .X(n1831) );
  nand_x1_sg U52542 ( .A(\yHat[8][10] ), .B(n46626), .X(n39648) );
  nand_x1_sg U52543 ( .A(n39650), .B(n39651), .X(n1830) );
  nand_x1_sg U52544 ( .A(\yHat[8][11] ), .B(n46626), .X(n39650) );
  nand_x1_sg U52545 ( .A(n39652), .B(n39653), .X(n1829) );
  nand_x1_sg U52546 ( .A(\yHat[8][12] ), .B(n46626), .X(n39652) );
  nand_x1_sg U52547 ( .A(n39654), .B(n39655), .X(n1828) );
  nand_x1_sg U52548 ( .A(\yHat[8][13] ), .B(n46626), .X(n39654) );
  nand_x1_sg U52549 ( .A(n39656), .B(n39657), .X(n1827) );
  nand_x1_sg U52550 ( .A(\yHat[8][14] ), .B(n46626), .X(n39656) );
  nand_x1_sg U52551 ( .A(n39658), .B(n39659), .X(n1826) );
  nand_x1_sg U52552 ( .A(\yHat[8][15] ), .B(n46626), .X(n39658) );
  nand_x1_sg U52553 ( .A(n39660), .B(n39661), .X(n1825) );
  nand_x1_sg U52554 ( .A(\yHat[8][16] ), .B(n46635), .X(n39660) );
  nand_x1_sg U52555 ( .A(n39662), .B(n39663), .X(n1824) );
  nand_x1_sg U52556 ( .A(\yHat[8][17] ), .B(n40523), .X(n39662) );
  nand_x1_sg U52557 ( .A(n39664), .B(n39665), .X(n1823) );
  nand_x1_sg U52558 ( .A(\yHat[8][18] ), .B(n46634), .X(n39664) );
  nand_x1_sg U52559 ( .A(n39666), .B(n39667), .X(n1822) );
  nand_x1_sg U52560 ( .A(\yHat[8][19] ), .B(n46626), .X(n39666) );
  nand_x1_sg U52561 ( .A(n39668), .B(n39669), .X(n1821) );
  nand_x1_sg U52562 ( .A(\yHat[9][0] ), .B(n46632), .X(n39668) );
  nand_x1_sg U52563 ( .A(n39670), .B(n39671), .X(n1820) );
  nand_x1_sg U52564 ( .A(\yHat[9][1] ), .B(n40520), .X(n39670) );
  nand_x1_sg U52565 ( .A(n39672), .B(n39673), .X(n1819) );
  nand_x1_sg U52566 ( .A(\yHat[9][2] ), .B(n40521), .X(n39672) );
  nand_x1_sg U52567 ( .A(n39674), .B(n39675), .X(n1818) );
  nand_x1_sg U52568 ( .A(\yHat[9][3] ), .B(n40520), .X(n39674) );
  nand_x1_sg U52569 ( .A(n39676), .B(n39677), .X(n1817) );
  nand_x1_sg U52570 ( .A(\yHat[9][4] ), .B(n46631), .X(n39676) );
  nand_x1_sg U52571 ( .A(n39678), .B(n39679), .X(n1816) );
  nand_x1_sg U52572 ( .A(\yHat[9][5] ), .B(n40524), .X(n39678) );
  nand_x1_sg U52573 ( .A(n39680), .B(n39681), .X(n1815) );
  nand_x1_sg U52574 ( .A(\yHat[9][6] ), .B(n46634), .X(n39680) );
  nand_x1_sg U52575 ( .A(n39682), .B(n39683), .X(n1814) );
  nand_x1_sg U52576 ( .A(\yHat[9][7] ), .B(n40523), .X(n39682) );
  nand_x1_sg U52577 ( .A(n39684), .B(n39685), .X(n1813) );
  nand_x1_sg U52578 ( .A(\yHat[9][8] ), .B(n46634), .X(n39684) );
  nand_x1_sg U52579 ( .A(n39686), .B(n39687), .X(n1812) );
  nand_x1_sg U52580 ( .A(\yHat[9][9] ), .B(n46635), .X(n39686) );
  nand_x1_sg U52581 ( .A(n39688), .B(n39689), .X(n1811) );
  nand_x1_sg U52582 ( .A(\yHat[9][10] ), .B(n46626), .X(n39688) );
  nand_x1_sg U52583 ( .A(n39690), .B(n39691), .X(n1810) );
  nand_x1_sg U52584 ( .A(\yHat[9][11] ), .B(n46632), .X(n39690) );
  nand_x1_sg U52585 ( .A(n39692), .B(n39693), .X(n1809) );
  nand_x1_sg U52586 ( .A(\yHat[9][12] ), .B(n40521), .X(n39692) );
  nand_x1_sg U52587 ( .A(n39694), .B(n39695), .X(n1808) );
  nand_x1_sg U52588 ( .A(\yHat[9][13] ), .B(n46631), .X(n39694) );
  nand_x1_sg U52589 ( .A(n39696), .B(n39697), .X(n1807) );
  nand_x1_sg U52590 ( .A(\yHat[9][14] ), .B(n46632), .X(n39696) );
  nand_x1_sg U52591 ( .A(n39698), .B(n39699), .X(n1806) );
  nand_x1_sg U52592 ( .A(\yHat[9][15] ), .B(n46626), .X(n39698) );
  nand_x1_sg U52593 ( .A(n39700), .B(n39701), .X(n1805) );
  nand_x1_sg U52594 ( .A(\yHat[9][16] ), .B(n46635), .X(n39700) );
  nand_x1_sg U52595 ( .A(n39702), .B(n39703), .X(n1804) );
  nand_x1_sg U52596 ( .A(\yHat[9][17] ), .B(n40524), .X(n39702) );
  nand_x1_sg U52597 ( .A(n39704), .B(n39705), .X(n1803) );
  nand_x1_sg U52598 ( .A(\yHat[9][18] ), .B(n46634), .X(n39704) );
  nand_x1_sg U52599 ( .A(n39706), .B(n39707), .X(n1802) );
  nand_x1_sg U52600 ( .A(\yHat[9][19] ), .B(n46635), .X(n39706) );
  nand_x1_sg U52601 ( .A(n39708), .B(n39709), .X(n1801) );
  nand_x1_sg U52602 ( .A(\yHat[10][0] ), .B(n40523), .X(n39708) );
  nand_x1_sg U52603 ( .A(n39710), .B(n39711), .X(n1800) );
  nand_x1_sg U52604 ( .A(\yHat[10][1] ), .B(n46634), .X(n39710) );
  nand_x1_sg U52605 ( .A(n39712), .B(n39713), .X(n1799) );
  nand_x1_sg U52606 ( .A(\yHat[10][2] ), .B(n46635), .X(n39712) );
  nand_x1_sg U52607 ( .A(n39714), .B(n39715), .X(n1798) );
  nand_x1_sg U52608 ( .A(\yHat[10][3] ), .B(n40520), .X(n39714) );
  nand_x1_sg U52609 ( .A(n39716), .B(n39717), .X(n1797) );
  nand_x1_sg U52610 ( .A(\yHat[10][4] ), .B(n40521), .X(n39716) );
  nand_x1_sg U52611 ( .A(n39718), .B(n39719), .X(n1796) );
  nand_x1_sg U52612 ( .A(\yHat[10][5] ), .B(n46635), .X(n39718) );
  nand_x1_sg U52613 ( .A(n39720), .B(n39721), .X(n1795) );
  nand_x1_sg U52614 ( .A(\yHat[10][6] ), .B(n40524), .X(n39720) );
  nand_x1_sg U52615 ( .A(n39722), .B(n39723), .X(n1794) );
  nand_x1_sg U52616 ( .A(\yHat[10][7] ), .B(n46634), .X(n39722) );
  nand_x1_sg U52617 ( .A(n39724), .B(n39725), .X(n1793) );
  nand_x1_sg U52618 ( .A(\yHat[10][8] ), .B(n46626), .X(n39724) );
  nand_x1_sg U52619 ( .A(n39726), .B(n39727), .X(n1792) );
  nand_x1_sg U52620 ( .A(\yHat[10][9] ), .B(n46632), .X(n39726) );
  nand_x1_sg U52621 ( .A(n39728), .B(n39729), .X(n1791) );
  nand_x1_sg U52622 ( .A(\yHat[10][10] ), .B(n46631), .X(n39728) );
  nand_x1_sg U52623 ( .A(n39730), .B(n39731), .X(n1790) );
  nand_x1_sg U52624 ( .A(\yHat[10][11] ), .B(n46631), .X(n39730) );
  nand_x1_sg U52625 ( .A(n39732), .B(n39733), .X(n1789) );
  nand_x1_sg U52626 ( .A(\yHat[10][12] ), .B(n40520), .X(n39732) );
  nand_x1_sg U52627 ( .A(n39734), .B(n39735), .X(n1788) );
  nand_x1_sg U52628 ( .A(\yHat[10][13] ), .B(n46631), .X(n39734) );
  nand_x1_sg U52629 ( .A(n39736), .B(n39737), .X(n1787) );
  nand_x1_sg U52630 ( .A(\yHat[10][14] ), .B(n46635), .X(n39736) );
  nand_x1_sg U52631 ( .A(n39738), .B(n39739), .X(n1786) );
  nand_x1_sg U52632 ( .A(\yHat[10][15] ), .B(n40523), .X(n39738) );
  nand_x1_sg U52633 ( .A(n39740), .B(n39741), .X(n1785) );
  nand_x1_sg U52634 ( .A(\yHat[10][16] ), .B(n46634), .X(n39740) );
  nand_x1_sg U52635 ( .A(n39742), .B(n39743), .X(n1784) );
  nand_x1_sg U52636 ( .A(\yHat[10][17] ), .B(n46626), .X(n39742) );
  nand_x1_sg U52637 ( .A(n39744), .B(n39745), .X(n1783) );
  nand_x1_sg U52638 ( .A(\yHat[10][18] ), .B(n46632), .X(n39744) );
  nand_x1_sg U52639 ( .A(n39746), .B(n39747), .X(n1782) );
  nand_x1_sg U52640 ( .A(\yHat[10][19] ), .B(n40520), .X(n39746) );
  nand_x1_sg U52641 ( .A(n39748), .B(n39749), .X(n1781) );
  nand_x1_sg U52642 ( .A(\yHat[11][0] ), .B(n46631), .X(n39748) );
  nand_x1_sg U52643 ( .A(n39750), .B(n39751), .X(n1780) );
  nand_x1_sg U52644 ( .A(\yHat[11][1] ), .B(n46634), .X(n39750) );
  nand_x1_sg U52645 ( .A(n39752), .B(n39753), .X(n1779) );
  nand_x1_sg U52646 ( .A(\yHat[11][2] ), .B(n46635), .X(n39752) );
  nand_x1_sg U52647 ( .A(n39754), .B(n39755), .X(n1778) );
  nand_x1_sg U52648 ( .A(\yHat[11][3] ), .B(n40523), .X(n39754) );
  nand_x1_sg U52649 ( .A(n39756), .B(n39757), .X(n1777) );
  nand_x1_sg U52650 ( .A(\yHat[11][4] ), .B(n46626), .X(n39756) );
  nand_x1_sg U52651 ( .A(n39758), .B(n39759), .X(n1776) );
  nand_x1_sg U52652 ( .A(\yHat[11][5] ), .B(n46634), .X(n39758) );
  nand_x1_sg U52653 ( .A(n39760), .B(n39761), .X(n1775) );
  nand_x1_sg U52654 ( .A(\yHat[11][6] ), .B(n46631), .X(n39760) );
  nand_x1_sg U52655 ( .A(n39762), .B(n39763), .X(n1774) );
  nand_x1_sg U52656 ( .A(\yHat[11][7] ), .B(n46632), .X(n39762) );
  nand_x1_sg U52657 ( .A(n39764), .B(n39765), .X(n1773) );
  nand_x1_sg U52658 ( .A(\yHat[11][8] ), .B(n46634), .X(n39764) );
  nand_x1_sg U52659 ( .A(n39766), .B(n39767), .X(n1772) );
  nand_x1_sg U52660 ( .A(\yHat[11][9] ), .B(n46632), .X(n39766) );
  nand_x1_sg U52661 ( .A(n39768), .B(n39769), .X(n1771) );
  nand_x1_sg U52662 ( .A(\yHat[11][10] ), .B(n46635), .X(n39768) );
  nand_x1_sg U52663 ( .A(n39770), .B(n39771), .X(n1770) );
  nand_x1_sg U52664 ( .A(\yHat[11][11] ), .B(n46634), .X(n39770) );
  nand_x1_sg U52665 ( .A(n39772), .B(n39773), .X(n1769) );
  nand_x1_sg U52666 ( .A(\yHat[11][12] ), .B(n46631), .X(n39772) );
  nand_x1_sg U52667 ( .A(n39774), .B(n39775), .X(n1768) );
  nand_x1_sg U52668 ( .A(\yHat[11][13] ), .B(n40520), .X(n39774) );
  nand_x1_sg U52669 ( .A(n39776), .B(n39777), .X(n1767) );
  nand_x1_sg U52670 ( .A(\yHat[11][14] ), .B(n46631), .X(n39776) );
  nand_x1_sg U52671 ( .A(n39778), .B(n39779), .X(n1766) );
  nand_x1_sg U52672 ( .A(\yHat[11][15] ), .B(n40523), .X(n39778) );
  nand_x1_sg U52673 ( .A(n39780), .B(n39781), .X(n1765) );
  nand_x1_sg U52674 ( .A(\yHat[11][16] ), .B(n40524), .X(n39780) );
  nand_x1_sg U52675 ( .A(n39782), .B(n39783), .X(n1764) );
  nand_x1_sg U52676 ( .A(\yHat[11][17] ), .B(n46626), .X(n39782) );
  nand_x1_sg U52677 ( .A(n39784), .B(n39785), .X(n1763) );
  nand_x1_sg U52678 ( .A(\yHat[11][18] ), .B(n40521), .X(n39784) );
  nand_x1_sg U52679 ( .A(n39786), .B(n39787), .X(n1762) );
  nand_x1_sg U52680 ( .A(\yHat[11][19] ), .B(n46631), .X(n39786) );
  nand_x1_sg U52681 ( .A(n39788), .B(n39789), .X(n1761) );
  nand_x1_sg U52682 ( .A(\yHat[12][0] ), .B(n46626), .X(n39788) );
  nand_x1_sg U52683 ( .A(n39790), .B(n39791), .X(n1760) );
  nand_x1_sg U52684 ( .A(\yHat[12][1] ), .B(n46626), .X(n39790) );
  nand_x1_sg U52685 ( .A(n39792), .B(n39793), .X(n1759) );
  nand_x1_sg U52686 ( .A(\yHat[12][2] ), .B(n46632), .X(n39792) );
  nand_x1_sg U52687 ( .A(n39794), .B(n39795), .X(n1758) );
  nand_x1_sg U52688 ( .A(\yHat[12][3] ), .B(n46626), .X(n39794) );
  nand_x1_sg U52689 ( .A(n39796), .B(n39797), .X(n1757) );
  nand_x1_sg U52690 ( .A(\yHat[12][4] ), .B(n40520), .X(n39796) );
  nand_x1_sg U52691 ( .A(n39798), .B(n39799), .X(n1756) );
  nand_x1_sg U52692 ( .A(\yHat[12][5] ), .B(n40524), .X(n39798) );
  nand_x1_sg U52693 ( .A(n39800), .B(n39801), .X(n1755) );
  nand_x1_sg U52694 ( .A(\yHat[12][6] ), .B(n46632), .X(n39800) );
  nand_x1_sg U52695 ( .A(n39802), .B(n39803), .X(n1754) );
  nand_x1_sg U52696 ( .A(\yHat[12][7] ), .B(n46632), .X(n39802) );
  nand_x1_sg U52697 ( .A(n39804), .B(n39805), .X(n1753) );
  nand_x1_sg U52698 ( .A(\yHat[12][8] ), .B(n40521), .X(n39804) );
  nand_x1_sg U52699 ( .A(n39806), .B(n39807), .X(n1752) );
  nand_x1_sg U52700 ( .A(\yHat[12][9] ), .B(n46632), .X(n39806) );
  nand_x1_sg U52701 ( .A(n39808), .B(n39809), .X(n1751) );
  nand_x1_sg U52702 ( .A(\yHat[12][10] ), .B(n46635), .X(n39808) );
  nand_x1_sg U52703 ( .A(n39810), .B(n39811), .X(n1750) );
  nand_x1_sg U52704 ( .A(\yHat[12][11] ), .B(n46631), .X(n39810) );
  nand_x1_sg U52705 ( .A(n39812), .B(n39813), .X(n1749) );
  nand_x1_sg U52706 ( .A(\yHat[12][12] ), .B(n46635), .X(n39812) );
  nand_x1_sg U52707 ( .A(n39814), .B(n39815), .X(n1748) );
  nand_x1_sg U52708 ( .A(\yHat[12][13] ), .B(n46634), .X(n39814) );
  nand_x1_sg U52709 ( .A(n39816), .B(n39817), .X(n1747) );
  nand_x1_sg U52710 ( .A(\yHat[12][14] ), .B(n46635), .X(n39816) );
  nand_x1_sg U52711 ( .A(n39818), .B(n39819), .X(n1746) );
  nand_x1_sg U52712 ( .A(\yHat[12][15] ), .B(n40523), .X(n39818) );
  nand_x1_sg U52713 ( .A(n39820), .B(n39821), .X(n1745) );
  nand_x1_sg U52714 ( .A(\yHat[12][16] ), .B(n46631), .X(n39820) );
  nand_x1_sg U52715 ( .A(n39822), .B(n39823), .X(n1744) );
  nand_x1_sg U52716 ( .A(\yHat[12][17] ), .B(n46632), .X(n39822) );
  nand_x1_sg U52717 ( .A(n39824), .B(n39825), .X(n1743) );
  nand_x1_sg U52718 ( .A(\yHat[12][18] ), .B(n46631), .X(n39824) );
  nand_x1_sg U52719 ( .A(n39826), .B(n39827), .X(n1742) );
  nand_x1_sg U52720 ( .A(\yHat[12][19] ), .B(n46626), .X(n39826) );
  nand_x1_sg U52721 ( .A(n39828), .B(n39829), .X(n1741) );
  nand_x1_sg U52722 ( .A(\yHat[13][0] ), .B(n46632), .X(n39828) );
  nand_x1_sg U52723 ( .A(n39830), .B(n39831), .X(n1740) );
  nand_x1_sg U52724 ( .A(\yHat[13][1] ), .B(n46626), .X(n39830) );
  nand_x1_sg U52725 ( .A(n39832), .B(n39833), .X(n1739) );
  nand_x1_sg U52726 ( .A(\yHat[13][2] ), .B(n40523), .X(n39832) );
  nand_x1_sg U52727 ( .A(n39834), .B(n39835), .X(n1738) );
  nand_x1_sg U52728 ( .A(\yHat[13][3] ), .B(n40523), .X(n39834) );
  nand_x1_sg U52729 ( .A(n39836), .B(n39837), .X(n1737) );
  nand_x1_sg U52730 ( .A(\yHat[13][4] ), .B(n40520), .X(n39836) );
  nand_x1_sg U52731 ( .A(n39838), .B(n39839), .X(n1736) );
  nand_x1_sg U52732 ( .A(\yHat[13][5] ), .B(n46635), .X(n39838) );
  nand_x1_sg U52733 ( .A(n39840), .B(n39841), .X(n1735) );
  nand_x1_sg U52734 ( .A(\yHat[13][6] ), .B(n46634), .X(n39840) );
  nand_x1_sg U52735 ( .A(n39842), .B(n39843), .X(n1734) );
  nand_x1_sg U52736 ( .A(\yHat[13][7] ), .B(n40521), .X(n39842) );
  nand_x1_sg U52737 ( .A(n39844), .B(n39845), .X(n1733) );
  nand_x1_sg U52738 ( .A(\yHat[13][8] ), .B(n46632), .X(n39844) );
  nand_x1_sg U52739 ( .A(n39846), .B(n39847), .X(n1732) );
  nand_x1_sg U52740 ( .A(\yHat[13][9] ), .B(n46626), .X(n39846) );
  nand_x1_sg U52741 ( .A(n39848), .B(n39849), .X(n1731) );
  nand_x1_sg U52742 ( .A(\yHat[13][10] ), .B(n40524), .X(n39848) );
  nand_x1_sg U52743 ( .A(n39850), .B(n39851), .X(n1730) );
  nand_x1_sg U52744 ( .A(\yHat[13][11] ), .B(n46635), .X(n39850) );
  nand_x1_sg U52745 ( .A(n39852), .B(n39853), .X(n1729) );
  nand_x1_sg U52746 ( .A(\yHat[13][12] ), .B(n46634), .X(n39852) );
  nand_x1_sg U52747 ( .A(n39854), .B(n39855), .X(n1728) );
  nand_x1_sg U52748 ( .A(\yHat[13][13] ), .B(n46631), .X(n39854) );
  nand_x1_sg U52749 ( .A(n39856), .B(n39857), .X(n1727) );
  nand_x1_sg U52750 ( .A(\yHat[13][14] ), .B(n46635), .X(n39856) );
  nand_x1_sg U52751 ( .A(n39858), .B(n39859), .X(n1726) );
  nand_x1_sg U52752 ( .A(\yHat[13][15] ), .B(n46634), .X(n39858) );
  nand_x1_sg U52753 ( .A(n39860), .B(n39861), .X(n1725) );
  nand_x1_sg U52754 ( .A(\yHat[13][16] ), .B(n46626), .X(n39860) );
  nand_x1_sg U52755 ( .A(n39862), .B(n39863), .X(n1724) );
  nand_x1_sg U52756 ( .A(\yHat[13][17] ), .B(n46632), .X(n39862) );
  nand_x1_sg U52757 ( .A(n39864), .B(n39865), .X(n1723) );
  nand_x1_sg U52758 ( .A(\yHat[13][18] ), .B(n46632), .X(n39864) );
  nand_x1_sg U52759 ( .A(n39866), .B(n39867), .X(n1722) );
  nand_x1_sg U52760 ( .A(\yHat[13][19] ), .B(n46626), .X(n39866) );
  nand_x1_sg U52761 ( .A(n39868), .B(n39869), .X(n1721) );
  nand_x1_sg U52762 ( .A(\yHat[14][0] ), .B(n46632), .X(n39868) );
  nand_x1_sg U52763 ( .A(n39870), .B(n39871), .X(n1720) );
  nand_x1_sg U52764 ( .A(\yHat[14][1] ), .B(n40521), .X(n39870) );
  nand_x1_sg U52765 ( .A(n39872), .B(n39873), .X(n1719) );
  nand_x1_sg U52766 ( .A(\yHat[14][2] ), .B(n46626), .X(n39872) );
  nand_x1_sg U52767 ( .A(n39874), .B(n39875), .X(n1718) );
  nand_x1_sg U52768 ( .A(\yHat[14][3] ), .B(n40524), .X(n39874) );
  nand_x1_sg U52769 ( .A(n39876), .B(n39877), .X(n1717) );
  nand_x1_sg U52770 ( .A(\yHat[14][4] ), .B(n40524), .X(n39876) );
  nand_x1_sg U52771 ( .A(n39878), .B(n39879), .X(n1716) );
  nand_x1_sg U52772 ( .A(\yHat[14][5] ), .B(n46635), .X(n39878) );
  nand_x1_sg U52773 ( .A(n39880), .B(n39881), .X(n1715) );
  nand_x1_sg U52774 ( .A(\yHat[14][6] ), .B(n46634), .X(n39880) );
  nand_x1_sg U52775 ( .A(n39882), .B(n39883), .X(n1714) );
  nand_x1_sg U52776 ( .A(\yHat[14][7] ), .B(n46635), .X(n39882) );
  nand_x1_sg U52777 ( .A(n39884), .B(n39885), .X(n1713) );
  nand_x1_sg U52778 ( .A(\yHat[14][8] ), .B(n46634), .X(n39884) );
  nand_x1_sg U52779 ( .A(n39886), .B(n39887), .X(n1712) );
  nand_x1_sg U52780 ( .A(\yHat[14][9] ), .B(n46626), .X(n39886) );
  nand_x1_sg U52781 ( .A(n39888), .B(n39889), .X(n1711) );
  nand_x1_sg U52782 ( .A(\yHat[14][10] ), .B(n40524), .X(n39888) );
  nand_x1_sg U52783 ( .A(n39890), .B(n39891), .X(n1710) );
  nand_x1_sg U52784 ( .A(\yHat[14][11] ), .B(n46631), .X(n39890) );
  nand_x1_sg U52785 ( .A(n39892), .B(n39893), .X(n1709) );
  nand_x1_sg U52786 ( .A(\yHat[14][12] ), .B(n46632), .X(n39892) );
  nand_x1_sg U52787 ( .A(n39894), .B(n39895), .X(n1708) );
  nand_x1_sg U52788 ( .A(\yHat[14][13] ), .B(n46632), .X(n39894) );
  nand_x1_sg U52789 ( .A(n39896), .B(n39897), .X(n1707) );
  nand_x1_sg U52790 ( .A(\yHat[14][14] ), .B(n46626), .X(n39896) );
  nand_x1_sg U52791 ( .A(n39898), .B(n39899), .X(n1706) );
  nand_x1_sg U52792 ( .A(\yHat[14][15] ), .B(n46632), .X(n39898) );
  nand_x1_sg U52793 ( .A(n39900), .B(n39901), .X(n1705) );
  nand_x1_sg U52794 ( .A(\yHat[14][16] ), .B(n46632), .X(n39900) );
  nand_x1_sg U52795 ( .A(n39902), .B(n39903), .X(n1704) );
  nand_x1_sg U52796 ( .A(\yHat[14][17] ), .B(n46635), .X(n39902) );
  nand_x1_sg U52797 ( .A(n39904), .B(n39905), .X(n1703) );
  nand_x1_sg U52798 ( .A(\yHat[14][18] ), .B(n46634), .X(n39904) );
  nand_x1_sg U52799 ( .A(n39906), .B(n39907), .X(n1702) );
  nand_x1_sg U52800 ( .A(\yHat[14][19] ), .B(n40523), .X(n39906) );
  nand_x1_sg U52801 ( .A(n39908), .B(n39909), .X(n1681) );
  nand_x1_sg U52802 ( .A(\y[0][0] ), .B(n46631), .X(n39908) );
  nand_x1_sg U52803 ( .A(n39910), .B(n39911), .X(n1680) );
  nand_x1_sg U52804 ( .A(\y[0][1] ), .B(n46627), .X(n39910) );
  nand_x1_sg U52805 ( .A(n39912), .B(n39913), .X(n1679) );
  nand_x1_sg U52806 ( .A(\y[0][2] ), .B(n46635), .X(n39912) );
  nand_x1_sg U52807 ( .A(n39914), .B(n39915), .X(n1678) );
  nand_x1_sg U52808 ( .A(\y[0][3] ), .B(n46635), .X(n39914) );
  nand_x1_sg U52809 ( .A(n39916), .B(n39917), .X(n1677) );
  nand_x1_sg U52810 ( .A(\y[0][4] ), .B(n40523), .X(n39916) );
  nand_x1_sg U52811 ( .A(n39918), .B(n39919), .X(n1676) );
  nand_x1_sg U52812 ( .A(\y[0][5] ), .B(n46631), .X(n39918) );
  nand_x1_sg U52813 ( .A(n39920), .B(n39921), .X(n1675) );
  nand_x1_sg U52814 ( .A(\y[0][6] ), .B(n46629), .X(n39920) );
  nand_x1_sg U52815 ( .A(n39922), .B(n39923), .X(n1674) );
  nand_x1_sg U52816 ( .A(\y[0][7] ), .B(n46629), .X(n39922) );
  nand_x1_sg U52817 ( .A(n39924), .B(n39925), .X(n1673) );
  nand_x1_sg U52818 ( .A(\y[0][8] ), .B(n46629), .X(n39924) );
  nand_x1_sg U52819 ( .A(n39926), .B(n39927), .X(n1672) );
  nand_x1_sg U52820 ( .A(\y[0][9] ), .B(n46629), .X(n39926) );
  nand_x1_sg U52821 ( .A(n39928), .B(n39929), .X(n1671) );
  nand_x1_sg U52822 ( .A(\y[0][10] ), .B(n46629), .X(n39928) );
  nand_x1_sg U52823 ( .A(n39930), .B(n39931), .X(n1670) );
  nand_x1_sg U52824 ( .A(\y[0][11] ), .B(n46629), .X(n39930) );
  nand_x1_sg U52825 ( .A(n39932), .B(n39933), .X(n1669) );
  nand_x1_sg U52826 ( .A(\y[0][12] ), .B(n46629), .X(n39932) );
  nand_x1_sg U52827 ( .A(n39934), .B(n39935), .X(n1668) );
  nand_x1_sg U52828 ( .A(\y[0][13] ), .B(n46629), .X(n39934) );
  nand_x1_sg U52829 ( .A(n39936), .B(n39937), .X(n1667) );
  nand_x1_sg U52830 ( .A(\y[0][14] ), .B(n46629), .X(n39936) );
  nand_x1_sg U52831 ( .A(n39938), .B(n39939), .X(n1666) );
  nand_x1_sg U52832 ( .A(\y[0][15] ), .B(n40521), .X(n39938) );
  nand_x1_sg U52833 ( .A(n39940), .B(n39941), .X(n1665) );
  nand_x1_sg U52834 ( .A(\y[0][16] ), .B(n40520), .X(n39940) );
  nand_x1_sg U52835 ( .A(n39942), .B(n39943), .X(n1664) );
  nand_x1_sg U52836 ( .A(\y[0][17] ), .B(n40521), .X(n39942) );
  nand_x1_sg U52837 ( .A(n39944), .B(n39945), .X(n1663) );
  nand_x1_sg U52838 ( .A(\y[0][18] ), .B(n40520), .X(n39944) );
  nand_x1_sg U52839 ( .A(n39946), .B(n39947), .X(n1662) );
  nand_x1_sg U52840 ( .A(\y[0][19] ), .B(n40521), .X(n39946) );
  nand_x1_sg U52841 ( .A(n39948), .B(n39949), .X(n1661) );
  nand_x1_sg U52842 ( .A(\y[1][0] ), .B(n40520), .X(n39948) );
  nand_x1_sg U52843 ( .A(n39950), .B(n39951), .X(n1660) );
  nand_x1_sg U52844 ( .A(\y[1][1] ), .B(n40521), .X(n39950) );
  nand_x1_sg U52845 ( .A(n39952), .B(n39953), .X(n1659) );
  nand_x1_sg U52846 ( .A(\y[1][2] ), .B(n40520), .X(n39952) );
  nand_x1_sg U52847 ( .A(n39954), .B(n39955), .X(n1658) );
  nand_x1_sg U52848 ( .A(\y[1][3] ), .B(n40521), .X(n39954) );
  nand_x1_sg U52849 ( .A(n39956), .B(n39957), .X(n1657) );
  nand_x1_sg U52850 ( .A(\y[1][4] ), .B(n46631), .X(n39956) );
  nand_x1_sg U52851 ( .A(n39958), .B(n39959), .X(n1656) );
  nand_x1_sg U52852 ( .A(\y[1][5] ), .B(n46631), .X(n39958) );
  nand_x1_sg U52853 ( .A(n39960), .B(n39961), .X(n1655) );
  nand_x1_sg U52854 ( .A(\y[1][6] ), .B(n46631), .X(n39960) );
  nand_x1_sg U52855 ( .A(n39962), .B(n39963), .X(n1654) );
  nand_x1_sg U52856 ( .A(\y[1][7] ), .B(n46631), .X(n39962) );
  nand_x1_sg U52857 ( .A(n39964), .B(n39965), .X(n1653) );
  nand_x1_sg U52858 ( .A(\y[1][8] ), .B(n46631), .X(n39964) );
  nand_x1_sg U52859 ( .A(n39966), .B(n39967), .X(n1652) );
  nand_x1_sg U52860 ( .A(\y[1][9] ), .B(n46631), .X(n39966) );
  nand_x1_sg U52861 ( .A(n39968), .B(n39969), .X(n1651) );
  nand_x1_sg U52862 ( .A(\y[1][10] ), .B(n46631), .X(n39968) );
  nand_x1_sg U52863 ( .A(n39970), .B(n39971), .X(n1650) );
  nand_x1_sg U52864 ( .A(\y[1][11] ), .B(n46631), .X(n39970) );
  nand_x1_sg U52865 ( .A(n39972), .B(n39973), .X(n1649) );
  nand_x1_sg U52866 ( .A(\y[1][12] ), .B(n46631), .X(n39972) );
  nand_x1_sg U52867 ( .A(n39974), .B(n39975), .X(n1648) );
  nand_x1_sg U52868 ( .A(\y[1][13] ), .B(n40520), .X(n39974) );
  nand_x1_sg U52869 ( .A(n39976), .B(n39977), .X(n1647) );
  nand_x1_sg U52870 ( .A(\y[1][14] ), .B(n46631), .X(n39976) );
  nand_x1_sg U52871 ( .A(n39978), .B(n39979), .X(n1646) );
  nand_x1_sg U52872 ( .A(\y[1][15] ), .B(n40521), .X(n39978) );
  nand_x1_sg U52873 ( .A(n39980), .B(n39981), .X(n1645) );
  nand_x1_sg U52874 ( .A(\y[1][16] ), .B(n46631), .X(n39980) );
  nand_x1_sg U52875 ( .A(n39982), .B(n39983), .X(n1644) );
  nand_x1_sg U52876 ( .A(\y[1][17] ), .B(n46631), .X(n39982) );
  nand_x1_sg U52877 ( .A(n39984), .B(n39985), .X(n1643) );
  nand_x1_sg U52878 ( .A(\y[1][18] ), .B(n40520), .X(n39984) );
  nand_x1_sg U52879 ( .A(n39986), .B(n39987), .X(n1642) );
  nand_x1_sg U52880 ( .A(\y[1][19] ), .B(n40521), .X(n39986) );
  nand_x1_sg U52881 ( .A(n39988), .B(n39989), .X(n1641) );
  nand_x1_sg U52882 ( .A(\y[2][0] ), .B(n46631), .X(n39988) );
  nand_x1_sg U52883 ( .A(n39990), .B(n39991), .X(n1640) );
  nand_x1_sg U52884 ( .A(\y[2][1] ), .B(n40520), .X(n39990) );
  nand_x1_sg U52885 ( .A(n39992), .B(n39993), .X(n1639) );
  nand_x1_sg U52886 ( .A(\y[2][2] ), .B(n46631), .X(n39992) );
  nand_x1_sg U52887 ( .A(n39994), .B(n39995), .X(n1638) );
  nand_x1_sg U52888 ( .A(\y[2][3] ), .B(n40520), .X(n39994) );
  nand_x1_sg U52889 ( .A(n39996), .B(n39997), .X(n1637) );
  nand_x1_sg U52890 ( .A(\y[2][4] ), .B(n46631), .X(n39996) );
  nand_x1_sg U52891 ( .A(n39998), .B(n39999), .X(n1636) );
  nand_x1_sg U52892 ( .A(\y[2][5] ), .B(n40521), .X(n39998) );
  nand_x1_sg U52893 ( .A(n40000), .B(n40001), .X(n1635) );
  nand_x1_sg U52894 ( .A(\y[2][6] ), .B(n40520), .X(n40000) );
  nand_x1_sg U52895 ( .A(n40002), .B(n40003), .X(n1634) );
  nand_x1_sg U52896 ( .A(\y[2][7] ), .B(n46631), .X(n40002) );
  nand_x1_sg U52897 ( .A(n40004), .B(n40005), .X(n1633) );
  nand_x1_sg U52898 ( .A(\y[2][8] ), .B(n46631), .X(n40004) );
  nand_x1_sg U52899 ( .A(n40006), .B(n40007), .X(n1632) );
  nand_x1_sg U52900 ( .A(\y[2][9] ), .B(n40521), .X(n40006) );
  nand_x1_sg U52901 ( .A(n40008), .B(n40009), .X(n1631) );
  nand_x1_sg U52902 ( .A(\y[2][10] ), .B(n46631), .X(n40008) );
  nand_x1_sg U52903 ( .A(n40010), .B(n40011), .X(n1630) );
  nand_x1_sg U52904 ( .A(\y[2][11] ), .B(n46632), .X(n40010) );
  nand_x1_sg U52905 ( .A(n40012), .B(n40013), .X(n1629) );
  nand_x1_sg U52906 ( .A(\y[2][12] ), .B(n40524), .X(n40012) );
  nand_x1_sg U52907 ( .A(n40014), .B(n40015), .X(n1628) );
  nand_x1_sg U52908 ( .A(\y[2][13] ), .B(n46629), .X(n40014) );
  nand_x1_sg U52909 ( .A(n40016), .B(n40017), .X(n1627) );
  nand_x1_sg U52910 ( .A(\y[2][14] ), .B(n46634), .X(n40016) );
  nand_x1_sg U52911 ( .A(n40018), .B(n40019), .X(n1626) );
  nand_x1_sg U52912 ( .A(\y[2][15] ), .B(n46634), .X(n40018) );
  nand_x1_sg U52913 ( .A(n40020), .B(n40021), .X(n1625) );
  nand_x1_sg U52914 ( .A(\y[2][16] ), .B(n40523), .X(n40020) );
  nand_x1_sg U52915 ( .A(n40022), .B(n40023), .X(n1624) );
  nand_x1_sg U52916 ( .A(\y[2][17] ), .B(n46632), .X(n40022) );
  nand_x1_sg U52917 ( .A(n40024), .B(n40025), .X(n1623) );
  nand_x1_sg U52918 ( .A(\y[2][18] ), .B(n46626), .X(n40024) );
  nand_x1_sg U52919 ( .A(n40026), .B(n40027), .X(n1622) );
  nand_x1_sg U52920 ( .A(\y[2][19] ), .B(n40520), .X(n40026) );
  nand_x1_sg U52921 ( .A(n40028), .B(n40029), .X(n1621) );
  nand_x1_sg U52922 ( .A(\y[3][0] ), .B(n40524), .X(n40028) );
  nand_x1_sg U52923 ( .A(n40030), .B(n40031), .X(n1620) );
  nand_x1_sg U52924 ( .A(\y[3][1] ), .B(n40523), .X(n40030) );
  nand_x1_sg U52925 ( .A(n40032), .B(n40033), .X(n1619) );
  nand_x1_sg U52926 ( .A(\y[3][2] ), .B(n40524), .X(n40032) );
  nand_x1_sg U52927 ( .A(n40034), .B(n40035), .X(n1618) );
  nand_x1_sg U52928 ( .A(\y[3][3] ), .B(n40523), .X(n40034) );
  nand_x1_sg U52929 ( .A(n40036), .B(n40037), .X(n1617) );
  nand_x1_sg U52930 ( .A(\y[3][4] ), .B(n40524), .X(n40036) );
  nand_x1_sg U52931 ( .A(n40038), .B(n40039), .X(n1616) );
  nand_x1_sg U52932 ( .A(\y[3][5] ), .B(n40523), .X(n40038) );
  nand_x1_sg U52933 ( .A(n40040), .B(n40041), .X(n1615) );
  nand_x1_sg U52934 ( .A(\y[3][6] ), .B(n40524), .X(n40040) );
  nand_x1_sg U52935 ( .A(n40042), .B(n40043), .X(n1614) );
  nand_x1_sg U52936 ( .A(\y[3][7] ), .B(n40523), .X(n40042) );
  nand_x1_sg U52937 ( .A(n40044), .B(n40045), .X(n1613) );
  nand_x1_sg U52938 ( .A(\y[3][8] ), .B(n40524), .X(n40044) );
  nand_x1_sg U52939 ( .A(n40046), .B(n40047), .X(n1612) );
  nand_x1_sg U52940 ( .A(\y[3][9] ), .B(n46632), .X(n40046) );
  nand_x1_sg U52941 ( .A(n40048), .B(n40049), .X(n1611) );
  nand_x1_sg U52942 ( .A(\y[3][10] ), .B(n46628), .X(n40048) );
  nand_x1_sg U52943 ( .A(n40050), .B(n40051), .X(n1610) );
  nand_x1_sg U52944 ( .A(\y[3][11] ), .B(n40524), .X(n40050) );
  nand_x1_sg U52945 ( .A(n40052), .B(n40053), .X(n1609) );
  nand_x1_sg U52946 ( .A(\y[3][12] ), .B(n46626), .X(n40052) );
  nand_x1_sg U52947 ( .A(n40054), .B(n40055), .X(n1608) );
  nand_x1_sg U52948 ( .A(\y[3][13] ), .B(n40523), .X(n40054) );
  nand_x1_sg U52949 ( .A(n40056), .B(n40057), .X(n1607) );
  nand_x1_sg U52950 ( .A(\y[3][14] ), .B(n46626), .X(n40056) );
  nand_x1_sg U52951 ( .A(n40058), .B(n40059), .X(n1606) );
  nand_x1_sg U52952 ( .A(\y[3][15] ), .B(n46638), .X(n40058) );
  nand_x1_sg U52953 ( .A(n40060), .B(n40061), .X(n1605) );
  nand_x1_sg U52954 ( .A(\y[3][16] ), .B(n46635), .X(n40060) );
  nand_x1_sg U52955 ( .A(n40062), .B(n40063), .X(n1604) );
  nand_x1_sg U52956 ( .A(\y[3][17] ), .B(n46627), .X(n40062) );
  nand_x1_sg U52957 ( .A(n40064), .B(n40065), .X(n1603) );
  nand_x1_sg U52958 ( .A(\y[3][18] ), .B(n46628), .X(n40064) );
  nand_x1_sg U52959 ( .A(n40066), .B(n40067), .X(n1602) );
  nand_x1_sg U52960 ( .A(\y[3][19] ), .B(n46627), .X(n40066) );
  nand_x1_sg U52961 ( .A(n40068), .B(n40069), .X(n1601) );
  nand_x1_sg U52962 ( .A(\y[4][0] ), .B(n46628), .X(n40068) );
  nand_x1_sg U52963 ( .A(n40070), .B(n40071), .X(n1600) );
  nand_x1_sg U52964 ( .A(\y[4][1] ), .B(n46634), .X(n40070) );
  nand_x1_sg U52965 ( .A(n40072), .B(n40073), .X(n1599) );
  nand_x1_sg U52966 ( .A(\y[4][2] ), .B(n46634), .X(n40072) );
  nand_x1_sg U52967 ( .A(n40074), .B(n40075), .X(n1598) );
  nand_x1_sg U52968 ( .A(\y[4][3] ), .B(n46629), .X(n40074) );
  nand_x1_sg U52969 ( .A(n40076), .B(n40077), .X(n1597) );
  nand_x1_sg U52970 ( .A(\y[4][4] ), .B(n40524), .X(n40076) );
  nand_x1_sg U52971 ( .A(n40078), .B(n40079), .X(n1596) );
  nand_x1_sg U52972 ( .A(\y[4][5] ), .B(n46632), .X(n40078) );
  nand_x1_sg U52973 ( .A(n40080), .B(n40081), .X(n1595) );
  nand_x1_sg U52974 ( .A(\y[4][6] ), .B(n46631), .X(n40080) );
  nand_x1_sg U52975 ( .A(n40082), .B(n40083), .X(n1594) );
  nand_x1_sg U52976 ( .A(\y[4][7] ), .B(n46635), .X(n40082) );
  nand_x1_sg U52977 ( .A(n40084), .B(n40085), .X(n1593) );
  nand_x1_sg U52978 ( .A(\y[4][8] ), .B(n40523), .X(n40084) );
  nand_x1_sg U52979 ( .A(n40086), .B(n40087), .X(n1592) );
  nand_x1_sg U52980 ( .A(\y[4][9] ), .B(n46634), .X(n40086) );
  nand_x1_sg U52981 ( .A(n40088), .B(n40089), .X(n1591) );
  nand_x1_sg U52982 ( .A(\y[4][10] ), .B(n46626), .X(n40088) );
  nand_x1_sg U52983 ( .A(n40090), .B(n40091), .X(n1590) );
  nand_x1_sg U52984 ( .A(\y[4][11] ), .B(n46632), .X(n40090) );
  nand_x1_sg U52985 ( .A(n40092), .B(n40093), .X(n1589) );
  nand_x1_sg U52986 ( .A(\y[4][12] ), .B(n40521), .X(n40092) );
  nand_x1_sg U52987 ( .A(n40094), .B(n40095), .X(n1588) );
  nand_x1_sg U52988 ( .A(\y[4][13] ), .B(n46631), .X(n40094) );
  nand_x1_sg U52989 ( .A(n40096), .B(n40097), .X(n1587) );
  nand_x1_sg U52990 ( .A(\y[4][14] ), .B(n46631), .X(n40096) );
  nand_x1_sg U52991 ( .A(n40098), .B(n40099), .X(n1586) );
  nand_x1_sg U52992 ( .A(\y[4][15] ), .B(n40521), .X(n40098) );
  nand_x1_sg U52993 ( .A(n40100), .B(n40101), .X(n1585) );
  nand_x1_sg U52994 ( .A(\y[4][16] ), .B(n40521), .X(n40100) );
  nand_x1_sg U52995 ( .A(n40102), .B(n40103), .X(n1584) );
  nand_x1_sg U52996 ( .A(\y[4][17] ), .B(n46626), .X(n40102) );
  nand_x1_sg U52997 ( .A(n40104), .B(n40105), .X(n1583) );
  nand_x1_sg U52998 ( .A(\y[4][18] ), .B(n46635), .X(n40104) );
  nand_x1_sg U52999 ( .A(n40106), .B(n40107), .X(n1582) );
  nand_x1_sg U53000 ( .A(\y[4][19] ), .B(n46638), .X(n40106) );
  nand_x1_sg U53001 ( .A(n40108), .B(n40109), .X(n1581) );
  nand_x1_sg U53002 ( .A(\y[5][0] ), .B(n40524), .X(n40108) );
  nand_x1_sg U53003 ( .A(n40110), .B(n40111), .X(n1580) );
  nand_x1_sg U53004 ( .A(\y[5][1] ), .B(n40524), .X(n40110) );
  nand_x1_sg U53005 ( .A(n40112), .B(n40113), .X(n1579) );
  nand_x1_sg U53006 ( .A(\y[5][2] ), .B(n40523), .X(n40112) );
  nand_x1_sg U53007 ( .A(n40114), .B(n40115), .X(n1578) );
  nand_x1_sg U53008 ( .A(\y[5][3] ), .B(n46634), .X(n40114) );
  nand_x1_sg U53009 ( .A(n40116), .B(n40117), .X(n1577) );
  nand_x1_sg U53010 ( .A(\y[5][4] ), .B(n46632), .X(n40116) );
  nand_x1_sg U53011 ( .A(n40118), .B(n40119), .X(n1576) );
  nand_x1_sg U53012 ( .A(\y[5][5] ), .B(n46632), .X(n40118) );
  nand_x1_sg U53013 ( .A(n40120), .B(n40121), .X(n1575) );
  nand_x1_sg U53014 ( .A(\y[5][6] ), .B(n46632), .X(n40120) );
  nand_x1_sg U53015 ( .A(n40122), .B(n40123), .X(n1574) );
  nand_x1_sg U53016 ( .A(\y[5][7] ), .B(n46632), .X(n40122) );
  nand_x1_sg U53017 ( .A(n40124), .B(n40125), .X(n1573) );
  nand_x1_sg U53018 ( .A(\y[5][8] ), .B(n46632), .X(n40124) );
  nand_x1_sg U53019 ( .A(n40126), .B(n40127), .X(n1572) );
  nand_x1_sg U53020 ( .A(\y[5][9] ), .B(n46632), .X(n40126) );
  nand_x1_sg U53021 ( .A(n40128), .B(n40129), .X(n1571) );
  nand_x1_sg U53022 ( .A(\y[5][10] ), .B(n46632), .X(n40128) );
  nand_x1_sg U53023 ( .A(n40130), .B(n40131), .X(n1570) );
  nand_x1_sg U53024 ( .A(\y[5][11] ), .B(n46632), .X(n40130) );
  nand_x1_sg U53025 ( .A(n40132), .B(n40133), .X(n1569) );
  nand_x1_sg U53026 ( .A(\y[5][12] ), .B(n46632), .X(n40132) );
  nand_x1_sg U53027 ( .A(n40134), .B(n40135), .X(n1568) );
  nand_x1_sg U53028 ( .A(\y[5][13] ), .B(n46635), .X(n40134) );
  nand_x1_sg U53029 ( .A(n40136), .B(n40137), .X(n1567) );
  nand_x1_sg U53030 ( .A(\y[5][14] ), .B(n40520), .X(n40136) );
  nand_x1_sg U53031 ( .A(n40138), .B(n40139), .X(n1566) );
  nand_x1_sg U53032 ( .A(\y[5][15] ), .B(n46638), .X(n40138) );
  nand_x1_sg U53033 ( .A(n40140), .B(n40141), .X(n1565) );
  nand_x1_sg U53034 ( .A(\y[5][16] ), .B(n40520), .X(n40140) );
  nand_x1_sg U53035 ( .A(n40142), .B(n40143), .X(n1564) );
  nand_x1_sg U53036 ( .A(\y[5][17] ), .B(n46638), .X(n40142) );
  nand_x1_sg U53037 ( .A(n40144), .B(n40145), .X(n1563) );
  nand_x1_sg U53038 ( .A(\y[5][18] ), .B(n40524), .X(n40144) );
  nand_x1_sg U53039 ( .A(n40146), .B(n40147), .X(n1562) );
  nand_x1_sg U53040 ( .A(\y[5][19] ), .B(n46638), .X(n40146) );
  nand_x1_sg U53041 ( .A(n40148), .B(n40149), .X(n1561) );
  nand_x1_sg U53042 ( .A(\y[6][0] ), .B(n40523), .X(n40148) );
  nand_x1_sg U53043 ( .A(n40150), .B(n40151), .X(n1560) );
  nand_x1_sg U53044 ( .A(\y[6][1] ), .B(n46626), .X(n40150) );
  nand_x1_sg U53045 ( .A(n40152), .B(n40153), .X(n1559) );
  nand_x1_sg U53046 ( .A(\y[6][2] ), .B(n40520), .X(n40152) );
  nand_x1_sg U53047 ( .A(n40154), .B(n40155), .X(n1558) );
  nand_x1_sg U53048 ( .A(\y[6][3] ), .B(n46635), .X(n40154) );
  nand_x1_sg U53049 ( .A(n40156), .B(n40157), .X(n1557) );
  nand_x1_sg U53050 ( .A(\y[6][4] ), .B(n46635), .X(n40156) );
  nand_x1_sg U53051 ( .A(n40158), .B(n40159), .X(n1556) );
  nand_x1_sg U53052 ( .A(\y[6][5] ), .B(n46634), .X(n40158) );
  nand_x1_sg U53053 ( .A(n40160), .B(n40161), .X(n1555) );
  nand_x1_sg U53054 ( .A(\y[6][6] ), .B(n46626), .X(n40160) );
  nand_x1_sg U53055 ( .A(n40162), .B(n40163), .X(n1554) );
  nand_x1_sg U53056 ( .A(\y[6][7] ), .B(n46631), .X(n40162) );
  nand_x1_sg U53057 ( .A(n40164), .B(n40165), .X(n1553) );
  nand_x1_sg U53058 ( .A(\y[6][8] ), .B(n40524), .X(n40164) );
  nand_x1_sg U53059 ( .A(n40166), .B(n40167), .X(n1552) );
  nand_x1_sg U53060 ( .A(\y[6][9] ), .B(n46635), .X(n40166) );
  nand_x1_sg U53061 ( .A(n40168), .B(n40169), .X(n1551) );
  nand_x1_sg U53062 ( .A(\y[6][10] ), .B(n46634), .X(n40168) );
  nand_x1_sg U53063 ( .A(n40170), .B(n40171), .X(n1550) );
  nand_x1_sg U53064 ( .A(\y[6][11] ), .B(n46632), .X(n40170) );
  nand_x1_sg U53065 ( .A(n40172), .B(n40173), .X(n1549) );
  nand_x1_sg U53066 ( .A(\y[6][12] ), .B(n46634), .X(n40172) );
  nand_x1_sg U53067 ( .A(n40174), .B(n40175), .X(n1548) );
  nand_x1_sg U53068 ( .A(\y[6][13] ), .B(n40523), .X(n40174) );
  nand_x1_sg U53069 ( .A(n40176), .B(n40177), .X(n1547) );
  nand_x1_sg U53070 ( .A(\y[6][14] ), .B(n46626), .X(n40176) );
  nand_x1_sg U53071 ( .A(n40178), .B(n40179), .X(n1546) );
  nand_x1_sg U53072 ( .A(\y[6][15] ), .B(n46632), .X(n40178) );
  nand_x1_sg U53073 ( .A(n40180), .B(n40181), .X(n1545) );
  nand_x1_sg U53074 ( .A(\y[6][16] ), .B(n46632), .X(n40180) );
  nand_x1_sg U53075 ( .A(n40182), .B(n40183), .X(n1544) );
  nand_x1_sg U53076 ( .A(\y[6][17] ), .B(n46635), .X(n40182) );
  nand_x1_sg U53077 ( .A(n40184), .B(n40185), .X(n1543) );
  nand_x1_sg U53078 ( .A(\y[6][18] ), .B(n46635), .X(n40184) );
  nand_x1_sg U53079 ( .A(n40186), .B(n40187), .X(n1542) );
  nand_x1_sg U53080 ( .A(\y[6][19] ), .B(n46626), .X(n40186) );
  nand_x1_sg U53081 ( .A(n40188), .B(n40189), .X(n1541) );
  nand_x1_sg U53082 ( .A(\y[7][0] ), .B(n46631), .X(n40188) );
  nand_x1_sg U53083 ( .A(n40190), .B(n40191), .X(n1540) );
  nand_x1_sg U53084 ( .A(\y[7][1] ), .B(n40524), .X(n40190) );
  nand_x1_sg U53085 ( .A(n40192), .B(n40193), .X(n1539) );
  nand_x1_sg U53086 ( .A(\y[7][2] ), .B(n46635), .X(n40192) );
  nand_x1_sg U53087 ( .A(n40194), .B(n40195), .X(n1538) );
  nand_x1_sg U53088 ( .A(\y[7][3] ), .B(n46634), .X(n40194) );
  nand_x1_sg U53089 ( .A(n40196), .B(n40197), .X(n1537) );
  nand_x1_sg U53090 ( .A(\y[7][4] ), .B(n46640), .X(n40196) );
  nand_x1_sg U53091 ( .A(n40198), .B(n40199), .X(n1536) );
  nand_x1_sg U53092 ( .A(\y[7][5] ), .B(n40523), .X(n40198) );
  nand_x1_sg U53093 ( .A(n40200), .B(n40201), .X(n1535) );
  nand_x1_sg U53094 ( .A(\y[7][6] ), .B(n46635), .X(n40200) );
  nand_x1_sg U53095 ( .A(n40202), .B(n40203), .X(n1534) );
  nand_x1_sg U53096 ( .A(\y[7][7] ), .B(n46634), .X(n40202) );
  nand_x1_sg U53097 ( .A(n40204), .B(n40205), .X(n1533) );
  nand_x1_sg U53098 ( .A(\y[7][8] ), .B(n46631), .X(n40204) );
  nand_x1_sg U53099 ( .A(n40206), .B(n40207), .X(n1532) );
  nand_x1_sg U53100 ( .A(\y[7][9] ), .B(n40521), .X(n40206) );
  nand_x1_sg U53101 ( .A(n40208), .B(n40209), .X(n1531) );
  nand_x1_sg U53102 ( .A(\y[7][10] ), .B(n46634), .X(n40208) );
  nand_x1_sg U53103 ( .A(n40210), .B(n40211), .X(n1530) );
  nand_x1_sg U53104 ( .A(\y[7][11] ), .B(n46631), .X(n40210) );
  nand_x1_sg U53105 ( .A(n40212), .B(n40213), .X(n1529) );
  nand_x1_sg U53106 ( .A(\y[7][12] ), .B(n46632), .X(n40212) );
  nand_x1_sg U53107 ( .A(n40214), .B(n40215), .X(n1528) );
  nand_x1_sg U53108 ( .A(\y[7][13] ), .B(n46632), .X(n40214) );
  nand_x1_sg U53109 ( .A(n40216), .B(n40217), .X(n1527) );
  nand_x1_sg U53110 ( .A(\y[7][14] ), .B(n46634), .X(n40216) );
  nand_x1_sg U53111 ( .A(n40218), .B(n40219), .X(n1526) );
  nand_x1_sg U53112 ( .A(\y[7][15] ), .B(n46632), .X(n40218) );
  nand_x1_sg U53113 ( .A(n40220), .B(n40221), .X(n1525) );
  nand_x1_sg U53114 ( .A(\y[7][16] ), .B(n46635), .X(n40220) );
  nand_x1_sg U53115 ( .A(n40222), .B(n40223), .X(n1524) );
  nand_x1_sg U53116 ( .A(\y[7][17] ), .B(n46626), .X(n40222) );
  nand_x1_sg U53117 ( .A(n40224), .B(n40225), .X(n1523) );
  nand_x1_sg U53118 ( .A(\y[7][18] ), .B(n46632), .X(n40224) );
  nand_x1_sg U53119 ( .A(n40226), .B(n40227), .X(n1522) );
  nand_x1_sg U53120 ( .A(\y[7][19] ), .B(n46634), .X(n40226) );
  nand_x1_sg U53121 ( .A(n40228), .B(n40229), .X(n1521) );
  nand_x1_sg U53122 ( .A(\y[8][0] ), .B(n40521), .X(n40228) );
  nand_x1_sg U53123 ( .A(n40230), .B(n40231), .X(n1520) );
  nand_x1_sg U53124 ( .A(\y[8][1] ), .B(n46631), .X(n40230) );
  nand_x1_sg U53125 ( .A(n40232), .B(n40233), .X(n1519) );
  nand_x1_sg U53126 ( .A(\y[8][2] ), .B(n46635), .X(n40232) );
  nand_x1_sg U53127 ( .A(n40234), .B(n40235), .X(n1518) );
  nand_x1_sg U53128 ( .A(\y[8][3] ), .B(n46626), .X(n40234) );
  nand_x1_sg U53129 ( .A(n40236), .B(n40237), .X(n1517) );
  nand_x1_sg U53130 ( .A(\y[8][4] ), .B(n46631), .X(n40236) );
  nand_x1_sg U53131 ( .A(n40238), .B(n40239), .X(n1516) );
  nand_x1_sg U53132 ( .A(\y[8][5] ), .B(n40523), .X(n40238) );
  nand_x1_sg U53133 ( .A(n40240), .B(n40241), .X(n1515) );
  nand_x1_sg U53134 ( .A(\y[8][6] ), .B(n40524), .X(n40240) );
  nand_x1_sg U53135 ( .A(n40242), .B(n40243), .X(n1514) );
  nand_x1_sg U53136 ( .A(\y[8][7] ), .B(n46635), .X(n40242) );
  nand_x1_sg U53137 ( .A(n40244), .B(n40245), .X(n1513) );
  nand_x1_sg U53138 ( .A(\y[8][8] ), .B(n46634), .X(n40244) );
  nand_x1_sg U53139 ( .A(n40246), .B(n40247), .X(n1512) );
  nand_x1_sg U53140 ( .A(\y[8][9] ), .B(n40521), .X(n40246) );
  nand_x1_sg U53141 ( .A(n40248), .B(n40249), .X(n1511) );
  nand_x1_sg U53142 ( .A(\y[8][10] ), .B(n40523), .X(n40248) );
  nand_x1_sg U53143 ( .A(n40250), .B(n40251), .X(n1510) );
  nand_x1_sg U53144 ( .A(\y[8][11] ), .B(n46635), .X(n40250) );
  nand_x1_sg U53145 ( .A(n40252), .B(n40253), .X(n1509) );
  nand_x1_sg U53146 ( .A(\y[8][12] ), .B(n46634), .X(n40252) );
  nand_x1_sg U53147 ( .A(n40254), .B(n40255), .X(n1508) );
  nand_x1_sg U53148 ( .A(\y[8][13] ), .B(n46634), .X(n40254) );
  nand_x1_sg U53149 ( .A(n40256), .B(n40257), .X(n1507) );
  nand_x1_sg U53150 ( .A(\y[8][14] ), .B(n46631), .X(n40256) );
  nand_x1_sg U53151 ( .A(n40258), .B(n40259), .X(n1506) );
  nand_x1_sg U53152 ( .A(\y[8][15] ), .B(n40523), .X(n40258) );
  nand_x1_sg U53153 ( .A(n40260), .B(n40261), .X(n1505) );
  nand_x1_sg U53154 ( .A(\y[8][16] ), .B(n46632), .X(n40260) );
  nand_x1_sg U53155 ( .A(n40262), .B(n40263), .X(n1504) );
  nand_x1_sg U53156 ( .A(\y[8][17] ), .B(n40520), .X(n40262) );
  nand_x1_sg U53157 ( .A(n40264), .B(n40265), .X(n1503) );
  nand_x1_sg U53158 ( .A(\y[8][18] ), .B(n46635), .X(n40264) );
  nand_x1_sg U53159 ( .A(n40266), .B(n40267), .X(n1502) );
  nand_x1_sg U53160 ( .A(\y[8][19] ), .B(n46626), .X(n40266) );
  nand_x1_sg U53161 ( .A(n40268), .B(n40269), .X(n1501) );
  nand_x1_sg U53162 ( .A(\y[9][0] ), .B(n46632), .X(n40268) );
  nand_x1_sg U53163 ( .A(n40270), .B(n40271), .X(n1500) );
  nand_x1_sg U53164 ( .A(\y[9][1] ), .B(n46632), .X(n40270) );
  nand_x1_sg U53165 ( .A(n40272), .B(n40273), .X(n1499) );
  nand_x1_sg U53166 ( .A(\y[9][2] ), .B(n46635), .X(n40272) );
  nand_x1_sg U53167 ( .A(n40274), .B(n40275), .X(n1498) );
  nand_x1_sg U53168 ( .A(\y[9][3] ), .B(n46634), .X(n40274) );
  nand_x1_sg U53169 ( .A(n40276), .B(n40277), .X(n1497) );
  nand_x1_sg U53170 ( .A(\y[9][4] ), .B(n40520), .X(n40276) );
  nand_x1_sg U53171 ( .A(n40278), .B(n40279), .X(n1496) );
  nand_x1_sg U53172 ( .A(\y[9][5] ), .B(n46631), .X(n40278) );
  nand_x1_sg U53173 ( .A(n40280), .B(n40281), .X(n1495) );
  nand_x1_sg U53174 ( .A(\y[9][6] ), .B(n40521), .X(n40280) );
  nand_x1_sg U53175 ( .A(n40282), .B(n40283), .X(n1494) );
  nand_x1_sg U53176 ( .A(\y[9][7] ), .B(n40523), .X(n40282) );
  nand_x1_sg U53177 ( .A(n40284), .B(n40285), .X(n1493) );
  nand_x1_sg U53178 ( .A(\y[9][8] ), .B(n46631), .X(n40284) );
  nand_x1_sg U53179 ( .A(n40286), .B(n40287), .X(n1492) );
  nand_x1_sg U53180 ( .A(\y[9][9] ), .B(n46635), .X(n40286) );
  nand_x1_sg U53181 ( .A(n40288), .B(n40289), .X(n1491) );
  nand_x1_sg U53182 ( .A(\y[9][10] ), .B(n46634), .X(n40288) );
  nand_x1_sg U53183 ( .A(n40290), .B(n40291), .X(n1490) );
  nand_x1_sg U53184 ( .A(\y[9][11] ), .B(n40524), .X(n40290) );
  nand_x1_sg U53185 ( .A(n40292), .B(n40293), .X(n1489) );
  nand_x1_sg U53186 ( .A(\y[9][12] ), .B(n46632), .X(n40292) );
  nand_x1_sg U53187 ( .A(n40294), .B(n40295), .X(n1488) );
  nand_x1_sg U53188 ( .A(\y[9][13] ), .B(n46626), .X(n40294) );
  nand_x1_sg U53189 ( .A(n40296), .B(n40297), .X(n1487) );
  nand_x1_sg U53190 ( .A(\y[9][14] ), .B(n46626), .X(n40296) );
  nand_x1_sg U53191 ( .A(n40298), .B(n40299), .X(n1486) );
  nand_x1_sg U53192 ( .A(\y[9][15] ), .B(n40521), .X(n40298) );
  nand_x1_sg U53193 ( .A(n40300), .B(n40301), .X(n1485) );
  nand_x1_sg U53194 ( .A(\y[9][16] ), .B(n46631), .X(n40300) );
  nand_x1_sg U53195 ( .A(n40302), .B(n40303), .X(n1484) );
  nand_x1_sg U53196 ( .A(\y[9][17] ), .B(n46626), .X(n40302) );
  nand_x1_sg U53197 ( .A(n40304), .B(n40305), .X(n1483) );
  nand_x1_sg U53198 ( .A(\y[9][18] ), .B(n46632), .X(n40304) );
  nand_x1_sg U53199 ( .A(n40306), .B(n40307), .X(n1482) );
  nand_x1_sg U53200 ( .A(\y[9][19] ), .B(n40524), .X(n40306) );
  nand_x1_sg U53201 ( .A(n40308), .B(n40309), .X(n1481) );
  nand_x1_sg U53202 ( .A(\y[10][0] ), .B(n46635), .X(n40308) );
  nand_x1_sg U53203 ( .A(n40310), .B(n40311), .X(n1480) );
  nand_x1_sg U53204 ( .A(\y[10][1] ), .B(n46634), .X(n40310) );
  nand_x1_sg U53205 ( .A(n40312), .B(n40313), .X(n1479) );
  nand_x1_sg U53206 ( .A(\y[10][2] ), .B(n40523), .X(n40312) );
  nand_x1_sg U53207 ( .A(n40314), .B(n40315), .X(n1478) );
  nand_x1_sg U53208 ( .A(\y[10][3] ), .B(n40520), .X(n40314) );
  nand_x1_sg U53209 ( .A(n40316), .B(n40317), .X(n1477) );
  nand_x1_sg U53210 ( .A(\y[10][4] ), .B(n46635), .X(n40316) );
  nand_x1_sg U53211 ( .A(n40318), .B(n40319), .X(n1476) );
  nand_x1_sg U53212 ( .A(\y[10][5] ), .B(n46634), .X(n40318) );
  nand_x1_sg U53213 ( .A(n40320), .B(n40321), .X(n1475) );
  nand_x1_sg U53214 ( .A(\y[10][6] ), .B(n46631), .X(n40320) );
  nand_x1_sg U53215 ( .A(n40322), .B(n40323), .X(n1474) );
  nand_x1_sg U53216 ( .A(\y[10][7] ), .B(n40521), .X(n40322) );
  nand_x1_sg U53217 ( .A(n40324), .B(n40325), .X(n1473) );
  nand_x1_sg U53218 ( .A(\y[10][8] ), .B(n46631), .X(n40324) );
  nand_x1_sg U53219 ( .A(n40326), .B(n40327), .X(n1472) );
  nand_x1_sg U53220 ( .A(\y[10][9] ), .B(n46626), .X(n40326) );
  nand_x1_sg U53221 ( .A(n40328), .B(n40329), .X(n1471) );
  nand_x1_sg U53222 ( .A(\y[10][10] ), .B(n40521), .X(n40328) );
  nand_x1_sg U53223 ( .A(n40330), .B(n40331), .X(n1470) );
  nand_x1_sg U53224 ( .A(\y[10][11] ), .B(n46631), .X(n40330) );
  nand_x1_sg U53225 ( .A(n40332), .B(n40333), .X(n1469) );
  nand_x1_sg U53226 ( .A(\y[10][12] ), .B(n46635), .X(n40332) );
  nand_x1_sg U53227 ( .A(n40334), .B(n40335), .X(n1468) );
  nand_x1_sg U53228 ( .A(\y[10][13] ), .B(n40521), .X(n40334) );
  nand_x1_sg U53229 ( .A(n40336), .B(n40337), .X(n1467) );
  nand_x1_sg U53230 ( .A(\y[10][14] ), .B(n46632), .X(n40336) );
  nand_x1_sg U53231 ( .A(n40338), .B(n40339), .X(n1466) );
  nand_x1_sg U53232 ( .A(\y[10][15] ), .B(n46631), .X(n40338) );
  nand_x1_sg U53233 ( .A(n40340), .B(n40341), .X(n1465) );
  nand_x1_sg U53234 ( .A(\y[10][16] ), .B(n40521), .X(n40340) );
  nand_x1_sg U53235 ( .A(n40342), .B(n40343), .X(n1464) );
  nand_x1_sg U53236 ( .A(\y[10][17] ), .B(n40523), .X(n40342) );
  nand_x1_sg U53237 ( .A(n40344), .B(n40345), .X(n1463) );
  nand_x1_sg U53238 ( .A(\y[10][18] ), .B(n46631), .X(n40344) );
  nand_x1_sg U53239 ( .A(n40346), .B(n40347), .X(n1462) );
  nand_x1_sg U53240 ( .A(\y[10][19] ), .B(n40520), .X(n40346) );
  nand_x1_sg U53241 ( .A(n40348), .B(n40349), .X(n1461) );
  nand_x1_sg U53242 ( .A(\y[11][0] ), .B(n46626), .X(n40348) );
  nand_x1_sg U53243 ( .A(n40350), .B(n40351), .X(n1460) );
  nand_x1_sg U53244 ( .A(\y[11][1] ), .B(n46632), .X(n40350) );
  nand_x1_sg U53245 ( .A(n40352), .B(n40353), .X(n1459) );
  nand_x1_sg U53246 ( .A(\y[11][2] ), .B(n40523), .X(n40352) );
  nand_x1_sg U53247 ( .A(n40354), .B(n40355), .X(n1458) );
  nand_x1_sg U53248 ( .A(\y[11][3] ), .B(n46635), .X(n40354) );
  nand_x1_sg U53249 ( .A(n40356), .B(n40357), .X(n1457) );
  nand_x1_sg U53250 ( .A(\y[11][4] ), .B(n46634), .X(n40356) );
  nand_x1_sg U53251 ( .A(n40358), .B(n40359), .X(n1456) );
  nand_x1_sg U53252 ( .A(\y[11][5] ), .B(n46626), .X(n40358) );
  nand_x1_sg U53253 ( .A(n40360), .B(n40361), .X(n1455) );
  nand_x1_sg U53254 ( .A(\y[11][6] ), .B(n40520), .X(n40360) );
  nand_x1_sg U53255 ( .A(n40362), .B(n40363), .X(n1454) );
  nand_x1_sg U53256 ( .A(\y[11][7] ), .B(n40520), .X(n40362) );
  nand_x1_sg U53257 ( .A(n40364), .B(n40365), .X(n1453) );
  nand_x1_sg U53258 ( .A(\y[11][8] ), .B(n46626), .X(n40364) );
  nand_x1_sg U53259 ( .A(n40366), .B(n40367), .X(n1452) );
  nand_x1_sg U53260 ( .A(\y[11][9] ), .B(n46632), .X(n40366) );
  nand_x1_sg U53261 ( .A(n40368), .B(n40369), .X(n1451) );
  nand_x1_sg U53262 ( .A(\y[11][10] ), .B(n40524), .X(n40368) );
  nand_x1_sg U53263 ( .A(n40370), .B(n40371), .X(n1450) );
  nand_x1_sg U53264 ( .A(\y[11][11] ), .B(n46635), .X(n40370) );
  nand_x1_sg U53265 ( .A(n40372), .B(n40373), .X(n1449) );
  nand_x1_sg U53266 ( .A(\y[11][12] ), .B(n46635), .X(n40372) );
  nand_x1_sg U53267 ( .A(n40374), .B(n40375), .X(n1448) );
  nand_x1_sg U53268 ( .A(\y[11][13] ), .B(n46634), .X(n40374) );
  nand_x1_sg U53269 ( .A(n40376), .B(n40377), .X(n1447) );
  nand_x1_sg U53270 ( .A(\y[11][14] ), .B(n40521), .X(n40376) );
  nand_x1_sg U53271 ( .A(n40378), .B(n40379), .X(n1446) );
  nand_x1_sg U53272 ( .A(\y[11][15] ), .B(n46631), .X(n40378) );
  nand_x1_sg U53273 ( .A(n40380), .B(n40381), .X(n1445) );
  nand_x1_sg U53274 ( .A(\y[11][16] ), .B(n46631), .X(n40380) );
  nand_x1_sg U53275 ( .A(n40382), .B(n40383), .X(n1444) );
  nand_x1_sg U53276 ( .A(\y[11][17] ), .B(n46626), .X(n40382) );
  nand_x1_sg U53277 ( .A(n40384), .B(n40385), .X(n1443) );
  nand_x1_sg U53278 ( .A(\y[11][18] ), .B(n40520), .X(n40384) );
  nand_x1_sg U53279 ( .A(n40386), .B(n40387), .X(n1442) );
  nand_x1_sg U53280 ( .A(\y[11][19] ), .B(n46631), .X(n40386) );
  nand_x1_sg U53281 ( .A(n40388), .B(n40389), .X(n1441) );
  nand_x1_sg U53282 ( .A(\y[12][0] ), .B(n40524), .X(n40388) );
  nand_x1_sg U53283 ( .A(n40390), .B(n40391), .X(n1440) );
  nand_x1_sg U53284 ( .A(\y[12][1] ), .B(n46626), .X(n40390) );
  nand_x1_sg U53285 ( .A(n40392), .B(n40393), .X(n1439) );
  nand_x1_sg U53286 ( .A(\y[12][2] ), .B(n46632), .X(n40392) );
  nand_x1_sg U53287 ( .A(n40394), .B(n40395), .X(n1438) );
  nand_x1_sg U53288 ( .A(\y[12][3] ), .B(n46631), .X(n40394) );
  nand_x1_sg U53289 ( .A(n40396), .B(n40397), .X(n1437) );
  nand_x1_sg U53290 ( .A(\y[12][4] ), .B(n46634), .X(n40396) );
  nand_x1_sg U53291 ( .A(n40398), .B(n40399), .X(n1436) );
  nand_x1_sg U53292 ( .A(\y[12][5] ), .B(n46626), .X(n40398) );
  nand_x1_sg U53293 ( .A(n40400), .B(n40401), .X(n1435) );
  nand_x1_sg U53294 ( .A(\y[12][6] ), .B(n46632), .X(n40400) );
  nand_x1_sg U53295 ( .A(n40402), .B(n40403), .X(n1434) );
  nand_x1_sg U53296 ( .A(\y[12][7] ), .B(n46634), .X(n40402) );
  nand_x1_sg U53297 ( .A(n40404), .B(n40405), .X(n1433) );
  nand_x1_sg U53298 ( .A(\y[12][8] ), .B(n40521), .X(n40404) );
  nand_x1_sg U53299 ( .A(n40406), .B(n40407), .X(n1432) );
  nand_x1_sg U53300 ( .A(\y[12][9] ), .B(n46629), .X(n40406) );
  nand_x1_sg U53301 ( .A(n40408), .B(n40409), .X(n1431) );
  nand_x1_sg U53302 ( .A(\y[12][10] ), .B(n46632), .X(n40408) );
  nand_x1_sg U53303 ( .A(n40410), .B(n40411), .X(n1430) );
  nand_x1_sg U53304 ( .A(\y[12][11] ), .B(n46634), .X(n40410) );
  nand_x1_sg U53305 ( .A(n40412), .B(n40413), .X(n1429) );
  nand_x1_sg U53306 ( .A(\y[12][12] ), .B(n46626), .X(n40412) );
  nand_x1_sg U53307 ( .A(n40414), .B(n40415), .X(n1428) );
  nand_x1_sg U53308 ( .A(\y[12][13] ), .B(n46634), .X(n40414) );
  nand_x1_sg U53309 ( .A(n40416), .B(n40417), .X(n1427) );
  nand_x1_sg U53310 ( .A(\y[12][14] ), .B(n46634), .X(n40416) );
  nand_x1_sg U53311 ( .A(n40418), .B(n40419), .X(n1426) );
  nand_x1_sg U53312 ( .A(\y[12][15] ), .B(n46634), .X(n40418) );
  nand_x1_sg U53313 ( .A(n40420), .B(n40421), .X(n1425) );
  nand_x1_sg U53314 ( .A(\y[12][16] ), .B(n46634), .X(n40420) );
  nand_x1_sg U53315 ( .A(n40422), .B(n40423), .X(n1424) );
  nand_x1_sg U53316 ( .A(\y[12][17] ), .B(n46634), .X(n40422) );
  nand_x1_sg U53317 ( .A(n40424), .B(n40425), .X(n1423) );
  nand_x1_sg U53318 ( .A(\y[12][18] ), .B(n46634), .X(n40424) );
  nand_x1_sg U53319 ( .A(n40426), .B(n40427), .X(n1422) );
  nand_x1_sg U53320 ( .A(\y[12][19] ), .B(n46634), .X(n40426) );
  nand_x1_sg U53321 ( .A(n40428), .B(n40429), .X(n1421) );
  nand_x1_sg U53322 ( .A(\y[13][0] ), .B(n46634), .X(n40428) );
  nand_x1_sg U53323 ( .A(n40430), .B(n40431), .X(n1420) );
  nand_x1_sg U53324 ( .A(\y[13][1] ), .B(n46634), .X(n40430) );
  nand_x1_sg U53325 ( .A(n40432), .B(n40433), .X(n1419) );
  nand_x1_sg U53326 ( .A(\y[13][2] ), .B(n46635), .X(n40432) );
  nand_x1_sg U53327 ( .A(n40434), .B(n40435), .X(n1418) );
  nand_x1_sg U53328 ( .A(\y[13][3] ), .B(n46634), .X(n40434) );
  nand_x1_sg U53329 ( .A(n40436), .B(n40437), .X(n1417) );
  nand_x1_sg U53330 ( .A(\y[13][4] ), .B(n40521), .X(n40436) );
  nand_x1_sg U53331 ( .A(n40438), .B(n40439), .X(n1416) );
  nand_x1_sg U53332 ( .A(\y[13][5] ), .B(n46631), .X(n40438) );
  nand_x1_sg U53333 ( .A(n40440), .B(n40441), .X(n1415) );
  nand_x1_sg U53334 ( .A(\y[13][6] ), .B(n46626), .X(n40440) );
  nand_x1_sg U53335 ( .A(n40442), .B(n40443), .X(n1414) );
  nand_x1_sg U53336 ( .A(\y[13][7] ), .B(n46638), .X(n40442) );
  nand_x1_sg U53337 ( .A(n40444), .B(n40445), .X(n1413) );
  nand_x1_sg U53338 ( .A(\y[13][8] ), .B(n46632), .X(n40444) );
  nand_x1_sg U53339 ( .A(n40446), .B(n40447), .X(n1412) );
  nand_x1_sg U53340 ( .A(\y[13][9] ), .B(n46638), .X(n40446) );
  nand_x1_sg U53341 ( .A(n40448), .B(n40449), .X(n1411) );
  nand_x1_sg U53342 ( .A(\y[13][10] ), .B(n46638), .X(n40448) );
  nand_x1_sg U53343 ( .A(n40450), .B(n40451), .X(n1410) );
  nand_x1_sg U53344 ( .A(\y[13][11] ), .B(n46632), .X(n40450) );
  nand_x1_sg U53345 ( .A(n40452), .B(n40453), .X(n1409) );
  nand_x1_sg U53346 ( .A(\y[13][12] ), .B(n40524), .X(n40452) );
  nand_x1_sg U53347 ( .A(n40454), .B(n40455), .X(n1408) );
  nand_x1_sg U53348 ( .A(\y[13][13] ), .B(n46635), .X(n40454) );
  nand_x1_sg U53349 ( .A(n40456), .B(n40457), .X(n1407) );
  nand_x1_sg U53350 ( .A(\y[13][14] ), .B(n46626), .X(n40456) );
  nand_x1_sg U53351 ( .A(n40458), .B(n40459), .X(n1406) );
  nand_x1_sg U53352 ( .A(\y[13][15] ), .B(n46632), .X(n40458) );
  nand_x1_sg U53353 ( .A(n40460), .B(n40461), .X(n1405) );
  nand_x1_sg U53354 ( .A(\y[13][16] ), .B(n40523), .X(n40460) );
  nand_x1_sg U53355 ( .A(n40462), .B(n40463), .X(n1404) );
  nand_x1_sg U53356 ( .A(\y[13][17] ), .B(n46635), .X(n40462) );
  nand_x1_sg U53357 ( .A(n40464), .B(n40465), .X(n1403) );
  nand_x1_sg U53358 ( .A(\y[13][18] ), .B(n46634), .X(n40464) );
  nand_x1_sg U53359 ( .A(n40466), .B(n40467), .X(n1402) );
  nand_x1_sg U53360 ( .A(\y[13][19] ), .B(n46626), .X(n40466) );
  nand_x1_sg U53361 ( .A(n40468), .B(n40469), .X(n1401) );
  nand_x1_sg U53362 ( .A(\y[14][0] ), .B(n46627), .X(n40468) );
  nand_x1_sg U53363 ( .A(n40470), .B(n40471), .X(n1400) );
  nand_x1_sg U53364 ( .A(\y[14][1] ), .B(n46627), .X(n40470) );
  nand_x1_sg U53365 ( .A(n40472), .B(n40473), .X(n1399) );
  nand_x1_sg U53366 ( .A(\y[14][2] ), .B(n46627), .X(n40472) );
  nand_x1_sg U53367 ( .A(n40474), .B(n40475), .X(n1398) );
  nand_x1_sg U53368 ( .A(\y[14][3] ), .B(n46627), .X(n40474) );
  nand_x1_sg U53369 ( .A(n40476), .B(n40477), .X(n1397) );
  nand_x1_sg U53370 ( .A(\y[14][4] ), .B(n46627), .X(n40476) );
  nand_x1_sg U53371 ( .A(n40478), .B(n40479), .X(n1396) );
  nand_x1_sg U53372 ( .A(\y[14][5] ), .B(n46627), .X(n40478) );
  nand_x1_sg U53373 ( .A(n40480), .B(n40481), .X(n1395) );
  nand_x1_sg U53374 ( .A(\y[14][6] ), .B(n46627), .X(n40480) );
  nand_x1_sg U53375 ( .A(n40482), .B(n40483), .X(n1394) );
  nand_x1_sg U53376 ( .A(\y[14][7] ), .B(n46627), .X(n40482) );
  nand_x1_sg U53377 ( .A(n40484), .B(n40485), .X(n1393) );
  nand_x1_sg U53378 ( .A(\y[14][8] ), .B(n46627), .X(n40484) );
  nand_x1_sg U53379 ( .A(n40486), .B(n40487), .X(n1392) );
  nand_x1_sg U53380 ( .A(\y[14][9] ), .B(n46628), .X(n40486) );
  nand_x1_sg U53381 ( .A(n40488), .B(n40489), .X(n1391) );
  nand_x1_sg U53382 ( .A(\y[14][10] ), .B(n46628), .X(n40488) );
  nand_x1_sg U53383 ( .A(n40490), .B(n40491), .X(n1390) );
  nand_x1_sg U53384 ( .A(\y[14][11] ), .B(n46628), .X(n40490) );
  nand_x1_sg U53385 ( .A(n40492), .B(n40493), .X(n1389) );
  nand_x1_sg U53386 ( .A(\y[14][12] ), .B(n46628), .X(n40492) );
  nand_x1_sg U53387 ( .A(n40494), .B(n40495), .X(n1388) );
  nand_x1_sg U53388 ( .A(\y[14][13] ), .B(n46628), .X(n40494) );
  nand_x1_sg U53389 ( .A(n40496), .B(n40497), .X(n1387) );
  nand_x1_sg U53390 ( .A(\y[14][14] ), .B(n46628), .X(n40496) );
  nand_x1_sg U53391 ( .A(n40498), .B(n40499), .X(n1386) );
  nand_x1_sg U53392 ( .A(\y[14][15] ), .B(n46628), .X(n40498) );
  nand_x1_sg U53393 ( .A(n40500), .B(n40501), .X(n1385) );
  nand_x1_sg U53394 ( .A(\y[14][16] ), .B(n46628), .X(n40500) );
  nand_x1_sg U53395 ( .A(n40502), .B(n40503), .X(n1384) );
  nand_x1_sg U53396 ( .A(\y[14][17] ), .B(n46628), .X(n40502) );
  nand_x1_sg U53397 ( .A(n40504), .B(n40505), .X(n1383) );
  nand_x1_sg U53398 ( .A(\y[14][18] ), .B(n46632), .X(n40504) );
  nand_x1_sg U53399 ( .A(n40506), .B(n40507), .X(n1382) );
  nand_x1_sg U53400 ( .A(\y[14][19] ), .B(n40523), .X(n40506) );
  nand_x1_sg U53401 ( .A(n40508), .B(n40509), .X(n1361) );
  nand_x1_sg U53402 ( .A(num[0]), .B(n46631), .X(n40508) );
  nand_x1_sg U53403 ( .A(n46647), .B(n46582), .X(n40509) );
  nand_x1_sg U53404 ( .A(n40510), .B(n40511), .X(n1360) );
  nand_x1_sg U53405 ( .A(num[1]), .B(n40520), .X(n40510) );
  nand_x1_sg U53406 ( .A(n40512), .B(n40513), .X(n1359) );
  nand_x1_sg U53407 ( .A(num[2]), .B(n46626), .X(n40512) );
  nand_x1_sg U53408 ( .A(n40514), .B(n40515), .X(n1358) );
  nand_x1_sg U53409 ( .A(num[3]), .B(n40524), .X(n40514) );
  nand_x1_sg U53410 ( .A(n46653), .B(n46584), .X(n40515) );
  nand_x1_sg U53411 ( .A(n39293), .B(n39294), .X(n40517) );
  nand_x1_sg U53412 ( .A(n39295), .B(n46576), .X(n39294) );
  nand_x1_sg U53413 ( .A(n39298), .B(n39299), .X(n40518) );
  nand_x4_sg U53414 ( .A(n29276), .B(n29277), .X(n29199) );
  nand_x4_sg U53415 ( .A(n28715), .B(n28716), .X(n28638) );
  nand_x4_sg U53416 ( .A(n28157), .B(n28158), .X(n28080) );
  nand_x4_sg U53417 ( .A(n28436), .B(n28437), .X(n28359) );
  nand_x4_sg U53418 ( .A(n27888), .B(n27889), .X(n27823) );
  nand_x4_sg U53419 ( .A(n27330), .B(n27331), .X(n27265) );
  nand_x4_sg U53420 ( .A(n26493), .B(n26494), .X(n26428) );
  nand_x2_sg U53421 ( .A(n42843), .B(n29287), .X(n29286) );
  nand_x2_sg U53422 ( .A(n42845), .B(n28726), .X(n28725) );
  nand_x2_sg U53423 ( .A(n42847), .B(n28168), .X(n28167) );
  nand_x2_sg U53424 ( .A(n46031), .B(n51549), .X(n25929) );
  inv_x2_sg U53425 ( .A(n43748), .X(n43749) );
  inv_x2_sg U53426 ( .A(n43750), .X(n43751) );
  inv_x2_sg U53427 ( .A(n43752), .X(n43753) );
  inv_x4_sg U53428 ( .A(n12509), .X(n51949) );
  nor_x4_sg U53429 ( .A(n12218), .B(n12030), .X(n12509) );
  inv_x4_sg U53430 ( .A(n11743), .X(n51647) );
  nor_x4_sg U53431 ( .A(n46533), .B(n11394), .X(n11743) );
  nand_x4_sg U53432 ( .A(n27038), .B(n27039), .X(n26961) );
  nand_x2_sg U53433 ( .A(n43749), .B(n27881), .X(n27880) );
  nand_x2_sg U53434 ( .A(n43751), .B(n27323), .X(n27322) );
  nand_x2_sg U53435 ( .A(n43753), .B(n26486), .X(n26485) );
  nand_x2_sg U53436 ( .A(n45989), .B(n54909), .X(n29283) );
  nand_x2_sg U53437 ( .A(n45991), .B(n54341), .X(n28722) );
  nand_x2_sg U53438 ( .A(n45993), .B(n53776), .X(n28164) );
  nand_x4_sg U53439 ( .A(n25658), .B(n25659), .X(n25594) );
  nand_x4_sg U53440 ( .A(n25934), .B(n25935), .X(n25869) );
  nor_x4_sg U53441 ( .A(n11638), .B(n51560), .X(n11689) );
  inv_x4_sg U53442 ( .A(n43754), .X(n43755) );
  inv_x2_sg U53443 ( .A(n43756), .X(n43757) );
  inv_x2_sg U53444 ( .A(n43758), .X(n43759) );
  inv_x2_sg U53445 ( .A(n43760), .X(n43761) );
  inv_x2_sg U53446 ( .A(n43762), .X(n43763) );
  inv_x2_sg U53447 ( .A(n43764), .X(n43765) );
  inv_x4_sg U53448 ( .A(n43766), .X(n43767) );
  inv_x4_sg U53449 ( .A(n43768), .X(n43769) );
  nor_x2_sg U53450 ( .A(n46232), .B(n51377), .X(n25467) );
  inv_x4_sg U53451 ( .A(n17203), .X(n53595) );
  nor_x4_sg U53452 ( .A(n46377), .B(n16854), .X(n17203) );
  inv_x4_sg U53453 ( .A(n15637), .X(n53037) );
  nor_x4_sg U53454 ( .A(n46421), .B(n15288), .X(n15637) );
  inv_x4_sg U53455 ( .A(n14084), .X(n52480) );
  nor_x4_sg U53456 ( .A(n13735), .B(n46469), .X(n14084) );
  inv_x4_sg U53457 ( .A(n13304), .X(n52203) );
  nor_x4_sg U53458 ( .A(n46489), .B(n12955), .X(n13304) );
  inv_x4_sg U53459 ( .A(n16983), .X(n53614) );
  nor_x4_sg U53460 ( .A(n16898), .B(n46389), .X(n16983) );
  inv_x4_sg U53461 ( .A(n15417), .X(n53056) );
  nor_x4_sg U53462 ( .A(n15332), .B(n46433), .X(n15417) );
  inv_x4_sg U53463 ( .A(n13084), .X(n52222) );
  nor_x4_sg U53464 ( .A(n12999), .B(n46501), .X(n13084) );
  inv_x4_sg U53465 ( .A(n21065), .X(n55013) );
  nor_x4_sg U53466 ( .A(n54947), .B(n20717), .X(n21065) );
  inv_x4_sg U53467 ( .A(n19521), .X(n54445) );
  nor_x4_sg U53468 ( .A(n54379), .B(n19173), .X(n19521) );
  inv_x4_sg U53469 ( .A(n17976), .X(n53880) );
  nor_x4_sg U53470 ( .A(n53814), .B(n17628), .X(n17976) );
  inv_x4_sg U53471 ( .A(n16198), .X(n53335) );
  nor_x4_sg U53472 ( .A(n16113), .B(n46411), .X(n16198) );
  inv_x4_sg U53473 ( .A(n11523), .X(n51666) );
  nor_x4_sg U53474 ( .A(n11438), .B(n46545), .X(n11523) );
  inv_x4_sg U53475 ( .A(n21614), .X(n55313) );
  nor_x4_sg U53476 ( .A(n21532), .B(n46254), .X(n21614) );
  inv_x4_sg U53477 ( .A(n20069), .X(n54745) );
  nor_x4_sg U53478 ( .A(n19987), .B(n46299), .X(n20069) );
  inv_x4_sg U53479 ( .A(n13864), .X(n52499) );
  nor_x4_sg U53480 ( .A(n13779), .B(n46479), .X(n13864) );
  inv_x4_sg U53481 ( .A(n20845), .X(n55031) );
  nor_x4_sg U53482 ( .A(n20762), .B(n46274), .X(n20845) );
  inv_x4_sg U53483 ( .A(n19301), .X(n54463) );
  nor_x4_sg U53484 ( .A(n19218), .B(n46319), .X(n19301) );
  inv_x4_sg U53485 ( .A(n17756), .X(n53898) );
  nor_x4_sg U53486 ( .A(n17673), .B(n46366), .X(n17756) );
  nand_x2_sg U53487 ( .A(n44717), .B(n46200), .X(n29620) );
  nand_x4_sg U53488 ( .A(n27876), .B(n27877), .X(n27799) );
  nand_x4_sg U53489 ( .A(n27318), .B(n27319), .X(n27241) );
  nand_x4_sg U53490 ( .A(n26481), .B(n26482), .X(n26404) );
  nand_x2_sg U53491 ( .A(n43759), .B(n28441), .X(n28440) );
  nand_x4_sg U53492 ( .A(n51302), .B(n25643), .X(n25564) );
  nand_x2_sg U53493 ( .A(n45985), .B(n54041), .X(n28454) );
  nand_x4_sg U53494 ( .A(n28727), .B(n28728), .X(n28662) );
  nand_x4_sg U53495 ( .A(n28169), .B(n28170), .X(n28104) );
  nand_x4_sg U53496 ( .A(n29288), .B(n29289), .X(n29223) );
  nand_x2_sg U53497 ( .A(n43761), .B(n27887), .X(n27886) );
  nand_x2_sg U53498 ( .A(n43763), .B(n27329), .X(n27328) );
  nand_x2_sg U53499 ( .A(n43765), .B(n26492), .X(n26491) );
  nand_x4_sg U53500 ( .A(n29008), .B(n29009), .X(n28946) );
  nand_x2_sg U53501 ( .A(n45293), .B(n26210), .X(n26209) );
  nand_x4_sg U53502 ( .A(n29569), .B(n29570), .X(n29507) );
  nand_x2_sg U53503 ( .A(n45301), .B(n27605), .X(n27604) );
  nand_x4_sg U53504 ( .A(n25652), .B(n25653), .X(n25582) );
  nand_x2_sg U53505 ( .A(n43757), .B(n25927), .X(n25926) );
  nor_x4_sg U53506 ( .A(n17099), .B(n53509), .X(n17148) );
  nor_x4_sg U53507 ( .A(n15533), .B(n52951), .X(n15582) );
  nor_x4_sg U53508 ( .A(n13200), .B(n52117), .X(n13249) );
  nor_x4_sg U53509 ( .A(n14547), .B(n46456), .X(n14545) );
  nor_x4_sg U53510 ( .A(n17162), .B(n46389), .X(n17160) );
  nor_x4_sg U53511 ( .A(n15596), .B(n46433), .X(n15594) );
  nor_x4_sg U53512 ( .A(n14043), .B(n46479), .X(n14041) );
  nor_x4_sg U53513 ( .A(n13263), .B(n46501), .X(n13261) );
  nor_x4_sg U53514 ( .A(n54921), .B(n46274), .X(n20566) );
  nor_x4_sg U53515 ( .A(n54353), .B(n46319), .X(n19022) );
  nor_x4_sg U53516 ( .A(n53788), .B(n46366), .X(n17477) );
  nor_x4_sg U53517 ( .A(n46477), .B(n46485), .X(n13507) );
  inv_x4_sg U53518 ( .A(n43770), .X(n43771) );
  nor_x4_sg U53519 ( .A(n46514), .B(n46523), .X(n12099) );
  nor_x4_sg U53520 ( .A(n46533), .B(n46545), .X(n11319) );
  nor_x4_sg U53521 ( .A(n51560), .B(n46533), .X(n11475) );
  nor_x4_sg U53522 ( .A(n54097), .B(n46337), .X(n18476) );
  inv_x4_sg U53523 ( .A(n44817), .X(n52681) );
  inv_x4_sg U53524 ( .A(n43772), .X(n43773) );
  inv_x2_sg U53525 ( .A(n43774), .X(n43775) );
  inv_x2_sg U53526 ( .A(n43776), .X(n43777) );
  inv_x2_sg U53527 ( .A(n43778), .X(n43779) );
  inv_x2_sg U53528 ( .A(n43780), .X(n43781) );
  inv_x2_sg U53529 ( .A(n55373), .X(n43782) );
  inv_x4_sg U53530 ( .A(n21707), .X(n55373) );
  inv_x2_sg U53531 ( .A(n52832), .X(n43783) );
  inv_x4_sg U53532 ( .A(n14728), .X(n52832) );
  nor_x8_sg U53533 ( .A(n29383), .B(n55344), .X(n29390) );
  nor_x8_sg U53534 ( .A(n29101), .B(n55059), .X(n29108) );
  nor_x8_sg U53535 ( .A(n28542), .B(n54491), .X(n28549) );
  inv_x4_sg U53536 ( .A(n43785), .X(n43786) );
  inv_x4_sg U53537 ( .A(n43787), .X(n43788) );
  inv_x4_sg U53538 ( .A(n43789), .X(n43790) );
  inv_x4_sg U53539 ( .A(n43791), .X(n43792) );
  inv_x4_sg U53540 ( .A(n43793), .X(n43794) );
  inv_x4_sg U53541 ( .A(n43795), .X(n43796) );
  nor_x2_sg U53542 ( .A(n46216), .B(n53641), .X(n27714) );
  nor_x2_sg U53543 ( .A(n46220), .B(n53083), .X(n27154) );
  nor_x2_sg U53544 ( .A(n46226), .B(n52249), .X(n26318) );
  inv_x4_sg U53545 ( .A(n16404), .X(n53337) );
  nor_x4_sg U53546 ( .A(n15925), .B(n16113), .X(n16404) );
  inv_x4_sg U53547 ( .A(n10946), .X(n51391) );
  nor_x4_sg U53548 ( .A(n10660), .B(n10518), .X(n10946) );
  inv_x4_sg U53549 ( .A(n12523), .X(n51928) );
  nor_x4_sg U53550 ( .A(n12174), .B(n46514), .X(n12523) );
  inv_x4_sg U53551 ( .A(n16417), .X(n53316) );
  nor_x4_sg U53552 ( .A(n46402), .B(n16069), .X(n16417) );
  inv_x4_sg U53553 ( .A(n12303), .X(n51947) );
  nor_x4_sg U53554 ( .A(n12218), .B(n46523), .X(n12303) );
  inv_x4_sg U53555 ( .A(n14634), .X(n52795) );
  nor_x4_sg U53556 ( .A(n14627), .B(n46452), .X(n14634) );
  inv_x4_sg U53557 ( .A(n19520), .X(n54518) );
  nor_x4_sg U53558 ( .A(n19401), .B(n46317), .X(n19520) );
  nor_x4_sg U53559 ( .A(n21774), .B(n46255), .X(n21613) );
  inv_x4_sg U53560 ( .A(n13863), .X(n52516) );
  nor_x4_sg U53561 ( .A(n13856), .B(n46480), .X(n13863) );
  inv_x4_sg U53562 ( .A(n20844), .X(n55049) );
  nor_x4_sg U53563 ( .A(n20837), .B(n46275), .X(n20844) );
  nor_x2_sg U53564 ( .A(n46195), .B(n46582), .X(n29619) );
  nand_x2_sg U53565 ( .A(n45283), .B(n27046), .X(n27045) );
  nand_x4_sg U53566 ( .A(n25922), .B(n25923), .X(n25845) );
  nand_x2_sg U53567 ( .A(n43775), .B(n29281), .X(n29280) );
  nand_x2_sg U53568 ( .A(n43777), .B(n28720), .X(n28719) );
  nand_x2_sg U53569 ( .A(n43779), .B(n28162), .X(n28161) );
  nand_x4_sg U53570 ( .A(n27891), .B(n27892), .X(n27829) );
  nand_x4_sg U53571 ( .A(n27333), .B(n27334), .X(n27271) );
  nand_x4_sg U53572 ( .A(n26496), .B(n26497), .X(n26434) );
  nand_x4_sg U53573 ( .A(n26774), .B(n26775), .X(n26712) );
  nand_x4_sg U53574 ( .A(n26217), .B(n26218), .X(n26155) );
  nand_x4_sg U53575 ( .A(n27612), .B(n27613), .X(n27550) );
  nand_x4_sg U53576 ( .A(n28730), .B(n28731), .X(n28668) );
  nand_x4_sg U53577 ( .A(n28172), .B(n28173), .X(n28110) );
  nand_x4_sg U53578 ( .A(n29291), .B(n29292), .X(n29229) );
  nand_x4_sg U53579 ( .A(n27053), .B(n27054), .X(n26991) );
  nand_x2_sg U53580 ( .A(n45995), .B(n53498), .X(n27883) );
  nand_x2_sg U53581 ( .A(n45997), .B(n52940), .X(n27325) );
  nand_x2_sg U53582 ( .A(n45999), .B(n52106), .X(n26488) );
  nand_x4_sg U53583 ( .A(n25937), .B(n25938), .X(n25875) );
  inv_x4_sg U53584 ( .A(n43797), .X(n43798) );
  nor_x4_sg U53585 ( .A(n16894), .B(n46389), .X(n16892) );
  nor_x4_sg U53586 ( .A(n16109), .B(n46411), .X(n16107) );
  nor_x4_sg U53587 ( .A(n15328), .B(n46433), .X(n15326) );
  nor_x4_sg U53588 ( .A(n12995), .B(n46501), .X(n12993) );
  nor_x4_sg U53589 ( .A(n11434), .B(n46545), .X(n11432) );
  nor_x4_sg U53590 ( .A(n21025), .B(n46274), .X(n21023) );
  nor_x4_sg U53591 ( .A(n19481), .B(n46319), .X(n19479) );
  nor_x4_sg U53592 ( .A(n17936), .B(n46366), .X(n17934) );
  nor_x4_sg U53593 ( .A(n14815), .B(n46456), .X(n14813) );
  nor_x4_sg U53594 ( .A(n46272), .B(n46281), .X(n20495) );
  nor_x4_sg U53595 ( .A(n46317), .B(n46326), .X(n18951) );
  nor_x4_sg U53596 ( .A(n46364), .B(n46373), .X(n17406) );
  nor_x4_sg U53597 ( .A(n13775), .B(n46469), .X(n14132) );
  nor_x4_sg U53598 ( .A(n20613), .B(n20685), .X(n20909) );
  nor_x4_sg U53599 ( .A(n19069), .B(n19141), .X(n19365) );
  nor_x4_sg U53600 ( .A(n17524), .B(n17596), .X(n17820) );
  nor_x4_sg U53601 ( .A(n15517), .B(n46434), .X(n15532) );
  nor_x4_sg U53602 ( .A(n13184), .B(n46502), .X(n13199) );
  inv_x4_sg U53603 ( .A(n43799), .X(n43800) );
  nor_x4_sg U53604 ( .A(n46377), .B(n46389), .X(n16779) );
  nor_x4_sg U53605 ( .A(n46421), .B(n46433), .X(n15213) );
  nor_x4_sg U53606 ( .A(n46489), .B(n46501), .X(n12880) );
  nor_x4_sg U53607 ( .A(n46568), .B(n46573), .X(n10395) );
  nor_x4_sg U53608 ( .A(n46381), .B(n46383), .X(n16816) );
  nor_x4_sg U53609 ( .A(n46425), .B(n46427), .X(n15250) );
  nor_x4_sg U53610 ( .A(n46493), .B(n46495), .X(n12917) );
  nor_x4_sg U53611 ( .A(n53509), .B(n46377), .X(n16935) );
  nor_x4_sg U53612 ( .A(n52951), .B(n46421), .X(n15369) );
  nor_x4_sg U53613 ( .A(n52117), .B(n46489), .X(n13036) );
  nor_x4_sg U53614 ( .A(n54947), .B(n54921), .X(n20796) );
  nor_x4_sg U53615 ( .A(n54379), .B(n54353), .X(n19252) );
  nor_x4_sg U53616 ( .A(n53814), .B(n53788), .X(n17707) );
  nor_x2_sg U53617 ( .A(n26973), .B(n51068), .X(n27043) );
  inv_x4_sg U53618 ( .A(n46149), .X(n51068) );
  inv_x4_sg U53619 ( .A(n43801), .X(n43802) );
  inv_x2_sg U53620 ( .A(n54805), .X(n43803) );
  inv_x4_sg U53621 ( .A(n20162), .X(n54805) );
  nor_x8_sg U53622 ( .A(n26851), .B(n52763), .X(n26858) );
  nor_x8_sg U53623 ( .A(n25456), .B(n51377), .X(n25464) );
  nor_x4_sg U53624 ( .A(n46469), .B(n46479), .X(n13660) );
  nor_x4_sg U53625 ( .A(n46409), .B(n46411), .X(n15868) );
  nor_x4_sg U53626 ( .A(n46521), .B(n46523), .X(n11973) );
  inv_x2_sg U53627 ( .A(reg_num[3]), .X(n44716) );
  inv_x2_sg U53628 ( .A(n8785), .X(n44284) );
  inv_x4_sg U53629 ( .A(n43804), .X(n43805) );
  nor_x2_sg U53630 ( .A(n52833), .B(n52760), .X(n14850) );
  nor_x2_sg U53631 ( .A(n50972), .B(n25576), .X(n25647) );
  nor_x2_sg U53632 ( .A(n26694), .B(n51049), .X(n26763) );
  nor_x2_sg U53633 ( .A(n51238), .B(n29489), .X(n29558) );
  nor_x2_sg U53634 ( .A(n51200), .B(n28928), .X(n28997) );
  nor_x2_sg U53635 ( .A(n51106), .B(n27532), .X(n27601) );
  nor_x2_sg U53636 ( .A(n51010), .B(n26137), .X(n26206) );
  inv_x4_sg U53637 ( .A(n43806), .X(n43807) );
  inv_x4_sg U53638 ( .A(n43808), .X(n43809) );
  nor_x4_sg U53639 ( .A(n39300), .B(n46672), .X(n11830) );
  inv_x4_sg U53640 ( .A(n43810), .X(n43811) );
  inv_x4_sg U53641 ( .A(n43814), .X(n43815) );
  inv_x4_sg U53642 ( .A(n43816), .X(n43817) );
  inv_x4_sg U53643 ( .A(n43818), .X(n43819) );
  inv_x4_sg U53644 ( .A(n43820), .X(n43821) );
  inv_x4_sg U53645 ( .A(n43822), .X(n43823) );
  inv_x4_sg U53646 ( .A(n43824), .X(n43825) );
  inv_x4_sg U53647 ( .A(n43826), .X(n43827) );
  inv_x4_sg U53648 ( .A(n43828), .X(n43829) );
  inv_x4_sg U53649 ( .A(n43830), .X(n43831) );
  inv_x4_sg U53650 ( .A(n43832), .X(n43833) );
  inv_x4_sg U53651 ( .A(n43834), .X(n43835) );
  nand_x2_sg U53652 ( .A(n29148), .B(n44169), .X(n29146) );
  nor_x2_sg U53653 ( .A(n46224), .B(n52525), .X(n26597) );
  nor_x2_sg U53654 ( .A(n46232), .B(n51418), .X(n25481) );
  nor_x2_sg U53655 ( .A(n14793), .B(n52887), .X(n14795) );
  inv_x4_sg U53656 ( .A(n21822), .X(n55315) );
  nor_x4_sg U53657 ( .A(n21532), .B(n46246), .X(n21822) );
  inv_x4_sg U53658 ( .A(n20277), .X(n54747) );
  nor_x4_sg U53659 ( .A(n19987), .B(n46291), .X(n20277) );
  inv_x4_sg U53660 ( .A(n18731), .X(n54180) );
  nor_x4_sg U53661 ( .A(n18442), .B(n46335), .X(n18731) );
  inv_x4_sg U53662 ( .A(n17189), .X(n53616) );
  nor_x4_sg U53663 ( .A(n46381), .B(n16898), .X(n17189) );
  inv_x4_sg U53664 ( .A(n15623), .X(n53058) );
  nor_x4_sg U53665 ( .A(n46425), .B(n15332), .X(n15623) );
  inv_x4_sg U53666 ( .A(n13290), .X(n52224) );
  nor_x4_sg U53667 ( .A(n46493), .B(n12999), .X(n13290) );
  inv_x4_sg U53668 ( .A(n43836), .X(n43837) );
  inv_x4_sg U53669 ( .A(n43838), .X(n43839) );
  inv_x4_sg U53670 ( .A(n43840), .X(n43841) );
  inv_x4_sg U53671 ( .A(n43842), .X(n43843) );
  inv_x4_sg U53672 ( .A(n14083), .X(n52563) );
  nor_x4_sg U53673 ( .A(n13964), .B(n46477), .X(n14083) );
  inv_x4_sg U53674 ( .A(n21064), .X(n55086) );
  nor_x4_sg U53675 ( .A(n20945), .B(n46272), .X(n21064) );
  inv_x4_sg U53676 ( .A(n17975), .X(n53953) );
  nor_x4_sg U53677 ( .A(n17856), .B(n46364), .X(n17975) );
  inv_x4_sg U53678 ( .A(n14855), .X(n52760) );
  nor_x4_sg U53679 ( .A(n14507), .B(n46445), .X(n14855) );
  nor_x4_sg U53680 ( .A(n16190), .B(n46407), .X(n16197) );
  nor_x4_sg U53681 ( .A(n11515), .B(n46546), .X(n11522) );
  nor_x4_sg U53682 ( .A(n20229), .B(n46300), .X(n20068) );
  inv_x4_sg U53683 ( .A(n19300), .X(n54481) );
  nor_x4_sg U53684 ( .A(n19293), .B(n46320), .X(n19300) );
  inv_x4_sg U53685 ( .A(n17755), .X(n53916) );
  nor_x4_sg U53686 ( .A(n17748), .B(n46367), .X(n17755) );
  inv_x4_sg U53687 ( .A(n10831), .X(n51413) );
  nor_x4_sg U53688 ( .A(n46568), .B(n46555), .X(n10831) );
  inv_x4_sg U53689 ( .A(n10293), .X(n51262) );
  nand_x4_sg U53690 ( .A(n51261), .B(n51257), .X(n10293) );
  nand_x4_sg U53691 ( .A(n55248), .B(n45459), .X(n21323) );
  nand_x4_sg U53692 ( .A(n54680), .B(n45463), .X(n19778) );
  nand_x4_sg U53693 ( .A(n53269), .B(n45471), .X(n15898) );
  nand_x4_sg U53694 ( .A(n51882), .B(n45481), .X(n12003) );
  nand_x4_sg U53695 ( .A(n11325), .B(n11324), .X(n11322) );
  nand_x4_sg U53696 ( .A(n44909), .B(n55426), .X(n29525) );
  nand_x4_sg U53697 ( .A(n44911), .B(n55406), .X(n29531) );
  nand_x4_sg U53698 ( .A(n44923), .B(n55141), .X(n29247) );
  nand_x4_sg U53699 ( .A(n44925), .B(n55121), .X(n29253) );
  nand_x4_sg U53700 ( .A(n44937), .B(n54858), .X(n28964) );
  nand_x4_sg U53701 ( .A(n44939), .B(n54838), .X(n28970) );
  nand_x4_sg U53702 ( .A(n44951), .B(n54573), .X(n28686) );
  nand_x4_sg U53703 ( .A(n44953), .B(n54553), .X(n28692) );
  nand_x4_sg U53704 ( .A(n44965), .B(n54290), .X(n28407) );
  nand_x4_sg U53705 ( .A(n44967), .B(n54271), .X(n28413) );
  nand_x4_sg U53706 ( .A(n44983), .B(n54008), .X(n28128) );
  nand_x4_sg U53707 ( .A(n44985), .B(n53988), .X(n28134) );
  nand_x4_sg U53708 ( .A(n44997), .B(n53727), .X(n27847) );
  nand_x4_sg U53709 ( .A(n44999), .B(n53708), .X(n27853) );
  nand_x4_sg U53710 ( .A(n45027), .B(n53169), .X(n27289) );
  nand_x4_sg U53711 ( .A(n45029), .B(n53150), .X(n27295) );
  nand_x4_sg U53712 ( .A(n45041), .B(n52888), .X(n27009) );
  nand_x4_sg U53713 ( .A(n45043), .B(n52868), .X(n27015) );
  nand_x4_sg U53714 ( .A(n45055), .B(n52610), .X(n26730) );
  nand_x4_sg U53715 ( .A(n45057), .B(n52591), .X(n26736) );
  nand_x4_sg U53716 ( .A(n45069), .B(n52335), .X(n26452) );
  nand_x4_sg U53717 ( .A(n45071), .B(n52316), .X(n26458) );
  nand_x4_sg U53718 ( .A(n45083), .B(n52058), .X(n26173) );
  nand_x4_sg U53719 ( .A(n45085), .B(n52040), .X(n26179) );
  nand_x4_sg U53720 ( .A(n45099), .B(n51778), .X(n25893) );
  nand_x4_sg U53721 ( .A(n45101), .B(n51759), .X(n25899) );
  nand_x4_sg U53722 ( .A(n45011), .B(n53447), .X(n27568) );
  nand_x4_sg U53723 ( .A(n45013), .B(n53428), .X(n27574) );
  nand_x4_sg U53724 ( .A(n16000), .B(n15999), .X(n15997) );
  nand_x4_sg U53725 ( .A(n45145), .B(n51479), .X(n25618) );
  nand_x4_sg U53726 ( .A(n45201), .B(n54122), .X(n28354) );
  nand_x4_sg U53727 ( .A(n45203), .B(n55254), .X(n29472) );
  nand_x4_sg U53728 ( .A(n45205), .B(n54686), .X(n28911) );
  nand_x4_sg U53729 ( .A(n45207), .B(n51332), .X(n25559) );
  nor_x2_sg U53730 ( .A(n55460), .B(n55462), .X(n29616) );
  nand_x2_sg U53731 ( .A(n55469), .B(n26358), .X(n27195) );
  nand_x4_sg U53732 ( .A(n52415), .B(n26759), .X(n26682) );
  nand_x4_sg U53733 ( .A(n26768), .B(n26769), .X(n26700) );
  nand_x4_sg U53734 ( .A(n29563), .B(n29564), .X(n29495) );
  nand_x4_sg U53735 ( .A(n29002), .B(n29003), .X(n28934) );
  nand_x4_sg U53736 ( .A(n27047), .B(n27048), .X(n26979) );
  nand_x4_sg U53737 ( .A(n28442), .B(n28443), .X(n28371) );
  nand_x4_sg U53738 ( .A(n55224), .B(n29554), .X(n29477) );
  nand_x4_sg U53739 ( .A(n54656), .B(n28993), .X(n28916) );
  nand_x4_sg U53740 ( .A(n53249), .B(n27597), .X(n27520) );
  nand_x4_sg U53741 ( .A(n51863), .B(n26202), .X(n26125) );
  nand_x4_sg U53742 ( .A(n26211), .B(n26212), .X(n26143) );
  nand_x4_sg U53743 ( .A(n27606), .B(n27607), .X(n27538) );
  nand_x2_sg U53744 ( .A(n45327), .B(n25651), .X(n25650) );
  nand_x2_sg U53745 ( .A(n43781), .B(n25933), .X(n25932) );
  nor_x4_sg U53746 ( .A(n46248), .B(n21653), .X(n21782) );
  inv_x4_sg U53747 ( .A(n43844), .X(n43845) );
  nor_x4_sg U53748 ( .A(n20884), .B(n54921), .X(n21011) );
  nor_x4_sg U53749 ( .A(n46293), .B(n20108), .X(n20237) );
  inv_x4_sg U53750 ( .A(n43846), .X(n43847) );
  nor_x4_sg U53751 ( .A(n19340), .B(n54353), .X(n19467) );
  nor_x4_sg U53752 ( .A(n17795), .B(n53788), .X(n17922) );
  nor_x4_sg U53753 ( .A(n14674), .B(n46449), .X(n14801) );
  nor_x4_sg U53754 ( .A(n13980), .B(n46473), .X(n14029) );
  nor_x4_sg U53755 ( .A(n46344), .B(n46353), .X(n18177) );
  nor_x4_sg U53756 ( .A(n14411), .B(n46447), .X(n14699) );
  nor_x4_sg U53757 ( .A(n17083), .B(n46390), .X(n17098) );
  inv_x4_sg U53758 ( .A(n44789), .X(n51291) );
  inv_x4_sg U53759 ( .A(n44791), .X(n53238) );
  inv_x4_sg U53760 ( .A(n44795), .X(n51852) );
  nor_x4_sg U53761 ( .A(n20685), .B(n46268), .X(n20683) );
  nor_x4_sg U53762 ( .A(n19141), .B(n46313), .X(n19139) );
  nor_x4_sg U53763 ( .A(n17596), .B(n46360), .X(n17594) );
  nor_x4_sg U53764 ( .A(n15925), .B(n53227), .X(n16031) );
  nor_x4_sg U53765 ( .A(n12030), .B(n51839), .X(n12136) );
  nor_x4_sg U53766 ( .A(n46469), .B(n46473), .X(n13816) );
  nor_x4_sg U53767 ( .A(n46404), .B(n46402), .X(n16150) );
  inv_x4_sg U53768 ( .A(n44839), .X(n52404) );
  inv_x4_sg U53769 ( .A(n44859), .X(n55213) );
  inv_x4_sg U53770 ( .A(n44861), .X(n54645) );
  inv_x2_sg U53771 ( .A(n54247), .X(n43848) );
  inv_x4_sg U53772 ( .A(n18616), .X(n54247) );
  nor_x8_sg U53773 ( .A(n28822), .B(n54776), .X(n28829) );
  nor_x8_sg U53774 ( .A(n27984), .B(n53926), .X(n27991) );
  nor_x8_sg U53775 ( .A(n25442), .B(n51334), .X(n25449) );
  nor_x4_sg U53776 ( .A(n46537), .B(n46546), .X(n11239) );
  inv_x4_sg U53777 ( .A(n43849), .X(n43850) );
  inv_x2_sg U53778 ( .A(\reg_y[14][19] ), .X(n45602) );
  inv_x2_sg U53779 ( .A(\reg_y[11][19] ), .X(n45608) );
  inv_x2_sg U53780 ( .A(\reg_y[7][19] ), .X(n45616) );
  inv_x2_sg U53781 ( .A(\reg_y[2][19] ), .X(n45626) );
  inv_x2_sg U53782 ( .A(\reg_y[1][19] ), .X(n45628) );
  inv_x2_sg U53783 ( .A(\reg_y[0][19] ), .X(n45630) );
  inv_x2_sg U53784 ( .A(\reg_y[8][6] ), .X(n45220) );
  inv_x2_sg U53785 ( .A(\reg_y[6][6] ), .X(n45222) );
  inv_x2_sg U53786 ( .A(\reg_y[3][6] ), .X(n45224) );
  inv_x2_sg U53787 ( .A(\reg_yHat[8][7] ), .X(n44314) );
  inv_x2_sg U53788 ( .A(\reg_yHat[6][7] ), .X(n44316) );
  inv_x2_sg U53789 ( .A(\reg_yHat[3][7] ), .X(n44318) );
  inv_x2_sg U53790 ( .A(\reg_yHat[13][5] ), .X(n44802) );
  inv_x2_sg U53791 ( .A(\reg_yHat[11][5] ), .X(n44804) );
  inv_x2_sg U53792 ( .A(\reg_yHat[9][5] ), .X(n44806) );
  inv_x2_sg U53793 ( .A(\reg_y[5][6] ), .X(n44816) );
  inv_x2_sg U53794 ( .A(\reg_y[11][4] ), .X(n46056) );
  inv_x2_sg U53795 ( .A(\reg_y[9][4] ), .X(n46058) );
  inv_x2_sg U53796 ( .A(\reg_y[13][4] ), .X(n46060) );
  inv_x4_sg U53797 ( .A(n43851), .X(n43852) );
  inv_x4_sg U53798 ( .A(n43853), .X(n43854) );
  nor_x4_sg U53799 ( .A(n29626), .B(n26078), .X(n9399) );
  nand_x4_sg U53800 ( .A(n29627), .B(n46582), .X(n29626) );
  nor_x4_sg U53801 ( .A(n29632), .B(n15726), .X(n9403) );
  nand_x4_sg U53802 ( .A(n46583), .B(n55457), .X(n29632) );
  inv_x4_sg U53803 ( .A(n43855), .X(n43856) );
  nor_x2_sg U53804 ( .A(n55512), .B(n46200), .X(n20380) );
  inv_x4_sg U53805 ( .A(n21925), .X(n55790) );
  inv_x4_sg U53806 ( .A(n43857), .X(n43858) );
  inv_x4_sg U53807 ( .A(n43859), .X(n43860) );
  inv_x4_sg U53808 ( .A(n43861), .X(n43862) );
  inv_x4_sg U53809 ( .A(n43863), .X(n43864) );
  inv_x4_sg U53810 ( .A(n43871), .X(n43872) );
  inv_x2_sg U53811 ( .A(n43873), .X(n43874) );
  inv_x4_sg U53812 ( .A(n43875), .X(n43876) );
  inv_x2_sg U53813 ( .A(n43877), .X(n43878) );
  nand_x4_sg U53814 ( .A(n26164), .B(n51811), .X(n11952) );
  nand_x4_sg U53815 ( .A(n27559), .B(n53199), .X(n15847) );
  inv_x4_sg U53816 ( .A(n43879), .X(n43880) );
  inv_x2_sg U53817 ( .A(n43881), .X(n43882) );
  nand_x4_sg U53818 ( .A(n29238), .B(n54890), .X(n20521) );
  nand_x4_sg U53819 ( .A(n28677), .B(n54322), .X(n18977) );
  nand_x4_sg U53820 ( .A(n28119), .B(n53757), .X(n17432) );
  inv_x4_sg U53821 ( .A(n43883), .X(n43884) );
  inv_x2_sg U53822 ( .A(n43885), .X(n43886) );
  inv_x4_sg U53823 ( .A(n43887), .X(n43888) );
  inv_x2_sg U53824 ( .A(n43889), .X(n43890) );
  inv_x4_sg U53825 ( .A(n43891), .X(n43892) );
  inv_x2_sg U53826 ( .A(n43893), .X(n43894) );
  inv_x4_sg U53827 ( .A(n43895), .X(n43896) );
  inv_x2_sg U53828 ( .A(n43897), .X(n43898) );
  nand_x4_sg U53829 ( .A(n27838), .B(n53479), .X(n16624) );
  nand_x4_sg U53830 ( .A(n27280), .B(n52921), .X(n15058) );
  nand_x4_sg U53831 ( .A(n26443), .B(n52087), .X(n12725) );
  nand_x4_sg U53832 ( .A(n25884), .B(n51529), .X(n11164) );
  nand_x4_sg U53833 ( .A(n25851), .B(n46202), .X(n46201) );
  inv_x4_sg U53834 ( .A(state[1]), .X(n55796) );
  inv_x4_sg U53835 ( .A(n43899), .X(n43900) );
  inv_x4_sg U53836 ( .A(n43901), .X(n43902) );
  inv_x4_sg U53837 ( .A(n43903), .X(n43904) );
  inv_x4_sg U53838 ( .A(n43905), .X(n43906) );
  inv_x4_sg U53839 ( .A(n43907), .X(n43908) );
  inv_x4_sg U53840 ( .A(n43909), .X(n43910) );
  inv_x4_sg U53841 ( .A(n43911), .X(n43912) );
  inv_x4_sg U53842 ( .A(n43913), .X(n43914) );
  inv_x4_sg U53843 ( .A(n43915), .X(n43916) );
  inv_x4_sg U53844 ( .A(n43917), .X(n43918) );
  inv_x4_sg U53845 ( .A(n43919), .X(n43920) );
  inv_x4_sg U53846 ( .A(n43921), .X(n43922) );
  inv_x4_sg U53847 ( .A(n43923), .X(n43924) );
  inv_x4_sg U53848 ( .A(n43925), .X(n43926) );
  inv_x4_sg U53849 ( .A(n43927), .X(n43928) );
  inv_x4_sg U53850 ( .A(n43929), .X(n43930) );
  inv_x4_sg U53851 ( .A(n43931), .X(n43932) );
  inv_x4_sg U53852 ( .A(n43933), .X(n43934) );
  nor_x4_sg U53853 ( .A(n16854), .B(n46387), .X(n16943) );
  nor_x4_sg U53854 ( .A(n15288), .B(n46431), .X(n15377) );
  nor_x4_sg U53855 ( .A(n12955), .B(n46499), .X(n13044) );
  nor_x4_sg U53856 ( .A(n11314), .B(n11313), .X(n11308) );
  nor_x4_sg U53857 ( .A(n51587), .B(n11315), .X(n11313) );
  nor_x4_sg U53858 ( .A(n51560), .B(n51606), .X(n11315) );
  inv_x4_sg U53859 ( .A(n10608), .X(n51359) );
  nand_x8_sg U53860 ( .A(n27697), .B(n16975), .X(n27704) );
  nor_x8_sg U53861 ( .A(n27690), .B(n53598), .X(n27697) );
  nand_x8_sg U53862 ( .A(n27137), .B(n15409), .X(n27144) );
  nor_x8_sg U53863 ( .A(n27130), .B(n53040), .X(n27137) );
  nand_x8_sg U53864 ( .A(n26301), .B(n13076), .X(n26308) );
  nor_x8_sg U53865 ( .A(n26294), .B(n52206), .X(n26301) );
  nor_x2_sg U53866 ( .A(n15880), .B(n15881), .X(n15879) );
  nor_x4_sg U53867 ( .A(n15887), .B(n43257), .X(n15880) );
  nand_x4_sg U53868 ( .A(n53240), .B(n46417), .X(n15881) );
  nand_x4_sg U53869 ( .A(n52406), .B(n46484), .X(n13547) );
  nor_x2_sg U53870 ( .A(n11985), .B(n11986), .X(n11984) );
  nor_x4_sg U53871 ( .A(n11992), .B(n43263), .X(n11985) );
  nand_x4_sg U53872 ( .A(n51854), .B(n46529), .X(n11986) );
  nor_x2_sg U53873 ( .A(n14691), .B(n14692), .X(n14690) );
  nor_x2_sg U53874 ( .A(n10838), .B(n51406), .X(n10837) );
  inv_x4_sg U53875 ( .A(n21051), .X(n55033) );
  nor_x4_sg U53876 ( .A(n20685), .B(n20762), .X(n21051) );
  inv_x4_sg U53877 ( .A(n19507), .X(n54465) );
  nor_x4_sg U53878 ( .A(n19141), .B(n19218), .X(n19507) );
  inv_x4_sg U53879 ( .A(n17962), .X(n53900) );
  nor_x4_sg U53880 ( .A(n17596), .B(n17673), .X(n17962) );
  inv_x4_sg U53881 ( .A(n14841), .X(n52780) );
  nor_x4_sg U53882 ( .A(n14552), .B(n46447), .X(n14841) );
  inv_x4_sg U53883 ( .A(n14070), .X(n52501) );
  nor_x4_sg U53884 ( .A(n13779), .B(n46471), .X(n14070) );
  inv_x4_sg U53885 ( .A(n11729), .X(n51668) );
  nor_x4_sg U53886 ( .A(n46537), .B(n11438), .X(n11729) );
  inv_x1_sg U53887 ( .A(n17287), .X(n53732) );
  inv_x1_sg U53888 ( .A(n15721), .X(n53174) );
  inv_x1_sg U53889 ( .A(n14168), .X(n52615) );
  inv_x1_sg U53890 ( .A(n13388), .X(n52340) );
  inv_x1_sg U53891 ( .A(n12606), .X(n52063) );
  inv_x1_sg U53892 ( .A(n16504), .X(n53451) );
  inv_x4_sg U53893 ( .A(n43935), .X(n43936) );
  inv_x4_sg U53894 ( .A(n43937), .X(n43938) );
  inv_x4_sg U53895 ( .A(n17202), .X(n53680) );
  nor_x4_sg U53896 ( .A(n17083), .B(n46387), .X(n17202) );
  inv_x4_sg U53897 ( .A(n15636), .X(n53122) );
  nor_x4_sg U53898 ( .A(n15517), .B(n46431), .X(n15636) );
  inv_x4_sg U53899 ( .A(n13303), .X(n52288) );
  nor_x4_sg U53900 ( .A(n13184), .B(n46499), .X(n13303) );
  inv_x4_sg U53901 ( .A(n16416), .X(n53403) );
  nor_x4_sg U53902 ( .A(n16299), .B(n46409), .X(n16416) );
  inv_x1_sg U53903 ( .A(n12565), .X(n52014) );
  inv_x4_sg U53904 ( .A(n12302), .X(n51964) );
  nor_x4_sg U53905 ( .A(n12295), .B(n46519), .X(n12302) );
  inv_x4_sg U53906 ( .A(n14854), .X(n52833) );
  nor_x4_sg U53907 ( .A(n14735), .B(n46454), .X(n14854) );
  inv_x4_sg U53908 ( .A(n20539), .X(n54937) );
  nand_x4_sg U53909 ( .A(n44363), .B(n20531), .X(n20539) );
  inv_x4_sg U53910 ( .A(n18995), .X(n54369) );
  nand_x4_sg U53911 ( .A(n44365), .B(n18987), .X(n18995) );
  inv_x4_sg U53912 ( .A(n17450), .X(n53804) );
  nand_x4_sg U53913 ( .A(n44367), .B(n17442), .X(n17450) );
  nand_x1_sg U53914 ( .A(n54930), .B(n20846), .X(n43939) );
  nand_x1_sg U53915 ( .A(n54930), .B(n20846), .X(n20841) );
  inv_x4_sg U53916 ( .A(n20546), .X(n54930) );
  nand_x1_sg U53917 ( .A(n54362), .B(n19302), .X(n43940) );
  nand_x1_sg U53918 ( .A(n54362), .B(n19302), .X(n19297) );
  inv_x4_sg U53919 ( .A(n19002), .X(n54362) );
  nand_x1_sg U53920 ( .A(n53797), .B(n17757), .X(n43941) );
  nand_x1_sg U53921 ( .A(n53797), .B(n17757), .X(n17752) );
  inv_x4_sg U53922 ( .A(n17457), .X(n53797) );
  inv_x4_sg U53923 ( .A(n18523), .X(n54199) );
  nor_x4_sg U53924 ( .A(n18574), .B(n46341), .X(n18523) );
  nor_x1_sg U53925 ( .A(n28459), .B(n21152), .X(n29149) );
  inv_x8_sg U53926 ( .A(n11048), .X(n51476) );
  nor_x4_sg U53927 ( .A(n10923), .B(n46570), .X(n11048) );
  nand_x4_sg U53928 ( .A(n52716), .B(n45475), .X(n14343) );
  nand_x4_sg U53929 ( .A(n51326), .B(n45485), .X(n10451) );
  inv_x1_sg U53930 ( .A(n16946), .X(n53643) );
  inv_x1_sg U53931 ( .A(n15380), .X(n53085) );
  inv_x1_sg U53932 ( .A(n13047), .X(n52251) );
  nand_x4_sg U53933 ( .A(n16652), .B(n16653), .X(n16643) );
  nand_x4_sg U53934 ( .A(n15086), .B(n15087), .X(n15077) );
  nand_x4_sg U53935 ( .A(n12753), .B(n12754), .X(n12744) );
  nand_x4_sg U53936 ( .A(n11192), .B(n11193), .X(n11183) );
  nand_x2_sg U53937 ( .A(n45273), .B(n26767), .X(n26766) );
  nand_x2_sg U53938 ( .A(n45277), .B(n29562), .X(n29561) );
  nand_x2_sg U53939 ( .A(n45279), .B(n29001), .X(n29000) );
  inv_x4_sg U53940 ( .A(n21756), .X(n55411) );
  inv_x4_sg U53941 ( .A(n20986), .X(n55126) );
  inv_x4_sg U53942 ( .A(n20211), .X(n54843) );
  inv_x4_sg U53943 ( .A(n19442), .X(n54558) );
  inv_x4_sg U53944 ( .A(n43942), .X(n43943) );
  inv_x4_sg U53945 ( .A(n18666), .X(n54276) );
  inv_x4_sg U53946 ( .A(n17897), .X(n53993) );
  inv_x4_sg U53947 ( .A(n14776), .X(n52873) );
  nor_x4_sg U53948 ( .A(n46516), .B(n12344), .X(n12468) );
  inv_x4_sg U53949 ( .A(n11664), .X(n51764) );
  nor_x4_sg U53950 ( .A(n16239), .B(n46404), .X(n16363) );
  nor_x4_sg U53951 ( .A(n46563), .B(n10782), .X(n10908) );
  nand_x4_sg U53952 ( .A(n46241), .B(n21686), .X(n21683) );
  nand_x4_sg U53953 ( .A(n46286), .B(n20141), .X(n20138) );
  inv_x4_sg U53954 ( .A(n16904), .X(n53623) );
  inv_x4_sg U53955 ( .A(n15338), .X(n53065) );
  inv_x4_sg U53956 ( .A(n13785), .X(n52508) );
  inv_x4_sg U53957 ( .A(n13005), .X(n52231) );
  inv_x4_sg U53958 ( .A(n12224), .X(n51956) );
  nor_x4_sg U53959 ( .A(n46387), .B(n46396), .X(n16621) );
  nor_x4_sg U53960 ( .A(n46431), .B(n46440), .X(n15055) );
  nor_x4_sg U53961 ( .A(n46499), .B(n46508), .X(n12722) );
  nor_x4_sg U53962 ( .A(n18705), .B(n46346), .X(n18703) );
  nor_x4_sg U53963 ( .A(n46270), .B(n46281), .X(n20504) );
  nor_x4_sg U53964 ( .A(n46315), .B(n46326), .X(n18960) );
  nor_x4_sg U53965 ( .A(n46362), .B(n46373), .X(n17415) );
  nor_x4_sg U53966 ( .A(n46242), .B(n46246), .X(n21678) );
  nor_x4_sg U53967 ( .A(n46287), .B(n46291), .X(n20133) );
  nor_x4_sg U53968 ( .A(n46559), .B(n10518), .X(n10807) );
  inv_x4_sg U53969 ( .A(n43944), .X(n43945) );
  nor_x4_sg U53970 ( .A(n44687), .B(n55138), .X(n20448) );
  inv_x4_sg U53971 ( .A(n43946), .X(n43947) );
  nor_x4_sg U53972 ( .A(n44689), .B(n54570), .X(n18904) );
  inv_x4_sg U53973 ( .A(n43948), .X(n43949) );
  nor_x4_sg U53974 ( .A(n44691), .B(n54005), .X(n17359) );
  inv_x4_sg U53975 ( .A(n43950), .X(n43951) );
  nor_x4_sg U53976 ( .A(n44693), .B(n52885), .X(n14240) );
  nor_x2_sg U53977 ( .A(n55277), .B(n21670), .X(n21669) );
  inv_x4_sg U53978 ( .A(n21674), .X(n55277) );
  nor_x2_sg U53979 ( .A(n54709), .B(n20125), .X(n20124) );
  inv_x4_sg U53980 ( .A(n20129), .X(n54709) );
  inv_x4_sg U53981 ( .A(n43952), .X(n43953) );
  nor_x2_sg U53982 ( .A(n40798), .B(out_L1[7]), .X(n32108) );
  nor_x2_sg U53983 ( .A(n40797), .B(out_L2[7]), .X(n24442) );
  inv_x4_sg U53984 ( .A(n43954), .X(n43955) );
  inv_x4_sg U53985 ( .A(n43956), .X(n43957) );
  inv_x4_sg U53986 ( .A(n43958), .X(n43959) );
  inv_x4_sg U53987 ( .A(n43960), .X(n43961) );
  inv_x4_sg U53988 ( .A(n43962), .X(n43963) );
  inv_x4_sg U53989 ( .A(n43964), .X(n43965) );
  inv_x4_sg U53990 ( .A(n43966), .X(n43967) );
  inv_x4_sg U53991 ( .A(n43968), .X(n43969) );
  inv_x4_sg U53992 ( .A(n43970), .X(n43971) );
  inv_x4_sg U53993 ( .A(n43972), .X(n43973) );
  inv_x4_sg U53994 ( .A(n46131), .X(n50973) );
  inv_x4_sg U53995 ( .A(n46119), .X(n51050) );
  inv_x4_sg U53996 ( .A(n46121), .X(n51239) );
  inv_x4_sg U53997 ( .A(n46123), .X(n51201) );
  inv_x4_sg U53998 ( .A(n46125), .X(n51107) );
  inv_x4_sg U53999 ( .A(n44837), .X(n54047) );
  inv_x4_sg U54000 ( .A(n46127), .X(n51011) );
  nor_x4_sg U54001 ( .A(n46471), .B(n52391), .X(n13697) );
  nand_x4_sg U54002 ( .A(n52525), .B(n46484), .X(n13904) );
  inv_x2_sg U54003 ( .A(n18069), .X(n43974) );
  nand_x8_sg U54004 ( .A(n46345), .B(n46352), .X(n18069) );
  inv_x2_sg U54005 ( .A(n14178), .X(n43975) );
  nand_x8_sg U54006 ( .A(n52648), .B(n46462), .X(n14178) );
  inv_x2_sg U54007 ( .A(n55085), .X(n43976) );
  inv_x4_sg U54008 ( .A(n20938), .X(n55085) );
  inv_x2_sg U54009 ( .A(n54517), .X(n43977) );
  inv_x4_sg U54010 ( .A(n19394), .X(n54517) );
  inv_x2_sg U54011 ( .A(n53952), .X(n43978) );
  inv_x4_sg U54012 ( .A(n17849), .X(n53952) );
  inv_x2_sg U54013 ( .A(n52556), .X(n43979) );
  inv_x4_sg U54014 ( .A(n13957), .X(n52556) );
  inv_x2_sg U54015 ( .A(n51732), .X(n43980) );
  inv_x4_sg U54016 ( .A(n11616), .X(n51732) );
  nor_x8_sg U54017 ( .A(n28264), .B(n54209), .X(n28271) );
  nor_x4_sg U54018 ( .A(n46381), .B(n46390), .X(n16699) );
  nor_x4_sg U54019 ( .A(n46425), .B(n46434), .X(n15133) );
  nor_x4_sg U54020 ( .A(n46493), .B(n46502), .X(n12800) );
  nor_x4_sg U54021 ( .A(n46543), .B(n46552), .X(n11161) );
  inv_x4_sg U54022 ( .A(n43981), .X(n43982) );
  inv_x4_sg U54023 ( .A(n43983), .X(n43984) );
  inv_x4_sg U54024 ( .A(n43985), .X(n43986) );
  inv_x4_sg U54025 ( .A(n43987), .X(n43988) );
  inv_x4_sg U54026 ( .A(n43989), .X(n43990) );
  inv_x4_sg U54027 ( .A(n43991), .X(n43992) );
  inv_x4_sg U54028 ( .A(n43993), .X(n43994) );
  inv_x4_sg U54029 ( .A(n43995), .X(n43996) );
  inv_x2_sg U54030 ( .A(\reg_y[13][19] ), .X(n45604) );
  inv_x2_sg U54031 ( .A(\reg_y[12][19] ), .X(n45606) );
  inv_x2_sg U54032 ( .A(\reg_y[10][19] ), .X(n45610) );
  inv_x2_sg U54033 ( .A(\reg_y[9][19] ), .X(n45612) );
  inv_x2_sg U54034 ( .A(\reg_y[8][19] ), .X(n45614) );
  inv_x2_sg U54035 ( .A(\reg_y[6][19] ), .X(n45618) );
  inv_x2_sg U54036 ( .A(\reg_y[5][19] ), .X(n45620) );
  inv_x2_sg U54037 ( .A(\reg_y[4][19] ), .X(n45622) );
  inv_x2_sg U54038 ( .A(\reg_y[3][19] ), .X(n45624) );
  inv_x2_sg U54039 ( .A(\reg_yHat[14][19] ), .X(n44758) );
  inv_x2_sg U54040 ( .A(\reg_yHat[11][19] ), .X(n44764) );
  inv_x2_sg U54041 ( .A(\reg_yHat[7][19] ), .X(n44772) );
  inv_x2_sg U54042 ( .A(\reg_yHat[2][19] ), .X(n44782) );
  inv_x2_sg U54043 ( .A(\reg_yHat[1][19] ), .X(n44784) );
  inv_x2_sg U54044 ( .A(\reg_yHat[0][19] ), .X(n44786) );
  inv_x2_sg U54045 ( .A(\reg_y[0][6] ), .X(n44788) );
  inv_x2_sg U54046 ( .A(\reg_y[7][6] ), .X(n44790) );
  inv_x2_sg U54047 ( .A(\reg_yHat[8][6] ), .X(n44308) );
  inv_x2_sg U54048 ( .A(\reg_yHat[6][6] ), .X(n44310) );
  inv_x2_sg U54049 ( .A(\reg_yHat[3][6] ), .X(n44312) );
  inv_x2_sg U54050 ( .A(\reg_y[1][6] ), .X(n46034) );
  inv_x2_sg U54051 ( .A(\reg_y[2][6] ), .X(n44794) );
  inv_x2_sg U54052 ( .A(\reg_y[13][7] ), .X(n45976) );
  inv_x2_sg U54053 ( .A(\reg_y[11][7] ), .X(n45978) );
  inv_x2_sg U54054 ( .A(\reg_y[9][7] ), .X(n45980) );
  inv_x2_sg U54055 ( .A(\reg_y[10][7] ), .X(n45210) );
  inv_x2_sg U54056 ( .A(\reg_y[8][7] ), .X(n45212) );
  inv_x2_sg U54057 ( .A(\reg_y[6][7] ), .X(n45214) );
  inv_x2_sg U54058 ( .A(\reg_y[3][7] ), .X(n45216) );
  inv_x2_sg U54059 ( .A(\reg_y[10][5] ), .X(n45218) );
  nand_x2_sg U54060 ( .A(n13728), .B(n13663), .X(n13727) );
  nand_x4_sg U54061 ( .A(n13666), .B(n13665), .X(n13663) );
  inv_x2_sg U54062 ( .A(\reg_y[13][6] ), .X(n46036) );
  inv_x2_sg U54063 ( .A(\reg_y[11][6] ), .X(n46038) );
  inv_x2_sg U54064 ( .A(\reg_y[9][6] ), .X(n46040) );
  inv_x2_sg U54065 ( .A(\reg_y[10][1] ), .X(n44814) );
  inv_x2_sg U54066 ( .A(\reg_yHat[1][5] ), .X(n44818) );
  inv_x2_sg U54067 ( .A(\reg_yHat[8][5] ), .X(n44820) );
  inv_x2_sg U54068 ( .A(\reg_yHat[6][5] ), .X(n44822) );
  inv_x2_sg U54069 ( .A(\reg_yHat[3][5] ), .X(n44824) );
  inv_x2_sg U54070 ( .A(\reg_y[13][1] ), .X(n44826) );
  inv_x2_sg U54071 ( .A(\reg_y[11][1] ), .X(n44828) );
  inv_x2_sg U54072 ( .A(\reg_y[9][1] ), .X(n44830) );
  inv_x2_sg U54073 ( .A(\reg_y[10][6] ), .X(n46042) );
  inv_x2_sg U54074 ( .A(\reg_y[10][3] ), .X(n45208) );
  inv_x2_sg U54075 ( .A(\reg_y[1][1] ), .X(n44834) );
  inv_x2_sg U54076 ( .A(\reg_y[8][4] ), .X(n46044) );
  inv_x2_sg U54077 ( .A(\reg_y[6][4] ), .X(n46046) );
  inv_x2_sg U54078 ( .A(\reg_y[3][4] ), .X(n46048) );
  inv_x2_sg U54079 ( .A(\reg_y[4][6] ), .X(n44838) );
  inv_x2_sg U54080 ( .A(\reg_y[8][1] ), .X(n44840) );
  inv_x2_sg U54081 ( .A(\reg_y[6][1] ), .X(n44842) );
  inv_x2_sg U54082 ( .A(\reg_y[3][1] ), .X(n44844) );
  inv_x2_sg U54083 ( .A(\reg_y[7][1] ), .X(n44846) );
  inv_x2_sg U54084 ( .A(\reg_y[4][1] ), .X(n44854) );
  inv_x2_sg U54085 ( .A(\reg_y[2][1] ), .X(n44856) );
  inv_x2_sg U54086 ( .A(\reg_y[8][3] ), .X(n46050) );
  inv_x2_sg U54087 ( .A(\reg_y[6][3] ), .X(n46052) );
  inv_x2_sg U54088 ( .A(\reg_y[3][3] ), .X(n46054) );
  inv_x2_sg U54089 ( .A(\reg_y[14][6] ), .X(n44858) );
  inv_x2_sg U54090 ( .A(\reg_y[12][6] ), .X(n44860) );
  inv_x2_sg U54091 ( .A(\reg_y[12][1] ), .X(n44862) );
  inv_x2_sg U54092 ( .A(\reg_y[0][1] ), .X(n44864) );
  inv_x2_sg U54093 ( .A(\reg_y[5][1] ), .X(n44866) );
  inv_x2_sg U54094 ( .A(\reg_y[14][17] ), .X(n45646) );
  inv_x2_sg U54095 ( .A(\reg_y[14][16] ), .X(n45648) );
  inv_x2_sg U54096 ( .A(\reg_y[14][15] ), .X(n45650) );
  inv_x2_sg U54097 ( .A(\reg_y[14][12] ), .X(n45652) );
  inv_x2_sg U54098 ( .A(\reg_y[14][11] ), .X(n45654) );
  inv_x2_sg U54099 ( .A(\reg_y[14][10] ), .X(n45656) );
  inv_x2_sg U54100 ( .A(\reg_y[14][8] ), .X(n45658) );
  inv_x2_sg U54101 ( .A(\reg_y[13][17] ), .X(n45660) );
  inv_x2_sg U54102 ( .A(\reg_y[13][16] ), .X(n45662) );
  inv_x2_sg U54103 ( .A(\reg_y[13][15] ), .X(n45664) );
  inv_x2_sg U54104 ( .A(\reg_y[13][13] ), .X(n45666) );
  inv_x2_sg U54105 ( .A(\reg_y[13][11] ), .X(n45668) );
  inv_x2_sg U54106 ( .A(\reg_y[13][10] ), .X(n45670) );
  inv_x2_sg U54107 ( .A(\reg_y[13][8] ), .X(n45672) );
  inv_x2_sg U54108 ( .A(\reg_y[12][17] ), .X(n45674) );
  inv_x2_sg U54109 ( .A(\reg_y[12][16] ), .X(n45676) );
  inv_x2_sg U54110 ( .A(\reg_y[12][15] ), .X(n45678) );
  inv_x2_sg U54111 ( .A(\reg_y[12][12] ), .X(n45680) );
  inv_x2_sg U54112 ( .A(\reg_y[12][11] ), .X(n45682) );
  inv_x2_sg U54113 ( .A(\reg_y[12][10] ), .X(n45684) );
  inv_x2_sg U54114 ( .A(\reg_y[12][8] ), .X(n45686) );
  inv_x2_sg U54115 ( .A(\reg_y[11][17] ), .X(n45688) );
  inv_x2_sg U54116 ( .A(\reg_y[11][16] ), .X(n45690) );
  inv_x2_sg U54117 ( .A(\reg_y[11][15] ), .X(n45692) );
  inv_x2_sg U54118 ( .A(\reg_y[11][13] ), .X(n45694) );
  inv_x2_sg U54119 ( .A(\reg_y[11][11] ), .X(n45696) );
  inv_x2_sg U54120 ( .A(\reg_y[11][10] ), .X(n45698) );
  inv_x2_sg U54121 ( .A(\reg_y[11][8] ), .X(n45700) );
  inv_x2_sg U54122 ( .A(\reg_y[10][17] ), .X(n45702) );
  inv_x2_sg U54123 ( .A(\reg_y[10][16] ), .X(n45704) );
  inv_x2_sg U54124 ( .A(\reg_y[10][15] ), .X(n45706) );
  inv_x2_sg U54125 ( .A(\reg_y[10][14] ), .X(n45708) );
  inv_x2_sg U54126 ( .A(\reg_y[10][13] ), .X(n45710) );
  inv_x2_sg U54127 ( .A(\reg_y[10][12] ), .X(n45712) );
  inv_x2_sg U54128 ( .A(\reg_y[10][11] ), .X(n45714) );
  inv_x2_sg U54129 ( .A(\reg_y[10][10] ), .X(n45716) );
  inv_x2_sg U54130 ( .A(\reg_y[10][8] ), .X(n45718) );
  inv_x2_sg U54131 ( .A(\reg_y[9][17] ), .X(n45720) );
  inv_x2_sg U54132 ( .A(\reg_y[9][16] ), .X(n45722) );
  inv_x2_sg U54133 ( .A(\reg_y[9][15] ), .X(n45724) );
  inv_x2_sg U54134 ( .A(\reg_y[9][13] ), .X(n45726) );
  inv_x2_sg U54135 ( .A(\reg_y[9][11] ), .X(n45728) );
  inv_x2_sg U54136 ( .A(\reg_y[9][10] ), .X(n45730) );
  inv_x2_sg U54137 ( .A(\reg_y[9][8] ), .X(n45732) );
  inv_x2_sg U54138 ( .A(\reg_y[8][17] ), .X(n45734) );
  inv_x2_sg U54139 ( .A(\reg_y[8][16] ), .X(n45736) );
  inv_x2_sg U54140 ( .A(\reg_y[8][15] ), .X(n45738) );
  inv_x2_sg U54141 ( .A(\reg_y[8][14] ), .X(n45740) );
  inv_x2_sg U54142 ( .A(\reg_y[8][12] ), .X(n45742) );
  inv_x2_sg U54143 ( .A(\reg_y[8][10] ), .X(n45744) );
  inv_x2_sg U54144 ( .A(\reg_y[8][8] ), .X(n45746) );
  inv_x2_sg U54145 ( .A(\reg_y[7][17] ), .X(n45748) );
  inv_x2_sg U54146 ( .A(\reg_y[7][16] ), .X(n45750) );
  inv_x2_sg U54147 ( .A(\reg_y[7][15] ), .X(n45752) );
  inv_x2_sg U54148 ( .A(\reg_y[7][14] ), .X(n45754) );
  inv_x2_sg U54149 ( .A(\reg_y[7][12] ), .X(n45756) );
  inv_x2_sg U54150 ( .A(\reg_y[7][11] ), .X(n45758) );
  inv_x2_sg U54151 ( .A(\reg_y[7][10] ), .X(n45760) );
  inv_x2_sg U54152 ( .A(\reg_y[7][8] ), .X(n45762) );
  inv_x2_sg U54153 ( .A(\reg_y[6][17] ), .X(n45764) );
  inv_x2_sg U54154 ( .A(\reg_y[6][16] ), .X(n45766) );
  inv_x2_sg U54155 ( .A(\reg_y[6][15] ), .X(n45768) );
  inv_x2_sg U54156 ( .A(\reg_y[6][14] ), .X(n45770) );
  inv_x2_sg U54157 ( .A(\reg_y[6][12] ), .X(n45772) );
  inv_x2_sg U54158 ( .A(\reg_y[6][10] ), .X(n45774) );
  inv_x2_sg U54159 ( .A(\reg_y[6][8] ), .X(n45776) );
  inv_x2_sg U54160 ( .A(\reg_y[5][17] ), .X(n45778) );
  inv_x2_sg U54161 ( .A(\reg_y[5][16] ), .X(n45780) );
  inv_x2_sg U54162 ( .A(\reg_y[5][15] ), .X(n45782) );
  inv_x2_sg U54163 ( .A(\reg_y[5][13] ), .X(n45784) );
  inv_x2_sg U54164 ( .A(\reg_y[5][11] ), .X(n45786) );
  inv_x2_sg U54165 ( .A(\reg_y[5][10] ), .X(n45788) );
  inv_x2_sg U54166 ( .A(\reg_y[5][8] ), .X(n45790) );
  inv_x2_sg U54167 ( .A(\reg_y[4][17] ), .X(n45792) );
  inv_x2_sg U54168 ( .A(\reg_y[4][16] ), .X(n45794) );
  inv_x2_sg U54169 ( .A(\reg_y[4][15] ), .X(n45796) );
  inv_x2_sg U54170 ( .A(\reg_y[4][14] ), .X(n45798) );
  inv_x2_sg U54171 ( .A(\reg_y[4][12] ), .X(n45800) );
  inv_x2_sg U54172 ( .A(\reg_y[4][10] ), .X(n45802) );
  inv_x2_sg U54173 ( .A(\reg_y[4][8] ), .X(n45804) );
  inv_x2_sg U54174 ( .A(\reg_y[3][17] ), .X(n45806) );
  inv_x2_sg U54175 ( .A(\reg_y[3][16] ), .X(n45808) );
  inv_x2_sg U54176 ( .A(\reg_y[3][15] ), .X(n45810) );
  inv_x2_sg U54177 ( .A(\reg_y[3][14] ), .X(n45812) );
  inv_x2_sg U54178 ( .A(\reg_y[3][12] ), .X(n45814) );
  inv_x2_sg U54179 ( .A(\reg_y[3][10] ), .X(n45816) );
  inv_x2_sg U54180 ( .A(\reg_y[3][8] ), .X(n45818) );
  inv_x2_sg U54181 ( .A(\reg_y[2][17] ), .X(n45820) );
  inv_x2_sg U54182 ( .A(\reg_y[2][16] ), .X(n45822) );
  inv_x2_sg U54183 ( .A(\reg_y[2][15] ), .X(n45824) );
  inv_x2_sg U54184 ( .A(\reg_y[2][14] ), .X(n45826) );
  inv_x2_sg U54185 ( .A(\reg_y[2][12] ), .X(n45828) );
  inv_x2_sg U54186 ( .A(\reg_y[2][11] ), .X(n45830) );
  inv_x2_sg U54187 ( .A(\reg_y[2][10] ), .X(n45832) );
  inv_x2_sg U54188 ( .A(\reg_y[2][8] ), .X(n45834) );
  inv_x2_sg U54189 ( .A(\reg_y[1][17] ), .X(n45836) );
  inv_x2_sg U54190 ( .A(\reg_y[1][16] ), .X(n45838) );
  inv_x2_sg U54191 ( .A(\reg_y[1][15] ), .X(n45840) );
  inv_x2_sg U54192 ( .A(\reg_y[1][14] ), .X(n45842) );
  inv_x2_sg U54193 ( .A(\reg_y[1][12] ), .X(n45844) );
  inv_x2_sg U54194 ( .A(\reg_y[1][11] ), .X(n45846) );
  inv_x2_sg U54195 ( .A(\reg_y[1][10] ), .X(n45848) );
  inv_x2_sg U54196 ( .A(\reg_y[1][8] ), .X(n45850) );
  inv_x2_sg U54197 ( .A(\reg_y[0][15] ), .X(n45852) );
  inv_x2_sg U54198 ( .A(\reg_y[0][14] ), .X(n45854) );
  inv_x2_sg U54199 ( .A(\reg_y[0][12] ), .X(n45856) );
  inv_x2_sg U54200 ( .A(\reg_y[0][11] ), .X(n45858) );
  inv_x2_sg U54201 ( .A(\reg_y[0][10] ), .X(n45860) );
  inv_x2_sg U54202 ( .A(\reg_y[0][8] ), .X(n45862) );
  inv_x2_sg U54203 ( .A(\reg_y[0][17] ), .X(n45864) );
  inv_x2_sg U54204 ( .A(\reg_y[5][14] ), .X(n45866) );
  inv_x2_sg U54205 ( .A(\reg_y[13][14] ), .X(n45868) );
  inv_x2_sg U54206 ( .A(\reg_y[11][14] ), .X(n45870) );
  inv_x2_sg U54207 ( .A(\reg_y[9][14] ), .X(n45872) );
  inv_x2_sg U54208 ( .A(\reg_y[4][11] ), .X(n45874) );
  inv_x2_sg U54209 ( .A(\reg_y[8][11] ), .X(n45876) );
  inv_x2_sg U54210 ( .A(\reg_y[6][11] ), .X(n45878) );
  inv_x2_sg U54211 ( .A(\reg_y[3][11] ), .X(n45880) );
  inv_x2_sg U54212 ( .A(\reg_y[0][16] ), .X(n45882) );
  inv_x2_sg U54213 ( .A(\reg_y[1][13] ), .X(n45884) );
  inv_x2_sg U54214 ( .A(\reg_y[14][13] ), .X(n45886) );
  inv_x2_sg U54215 ( .A(\reg_y[12][13] ), .X(n45888) );
  inv_x2_sg U54216 ( .A(\reg_y[2][13] ), .X(n45890) );
  inv_x2_sg U54217 ( .A(\reg_y[14][14] ), .X(n45892) );
  inv_x2_sg U54218 ( .A(\reg_y[12][14] ), .X(n45894) );
  inv_x2_sg U54219 ( .A(\reg_y[1][9] ), .X(n45896) );
  inv_x2_sg U54220 ( .A(\reg_y[14][1] ), .X(n44874) );
  inv_x2_sg U54221 ( .A(\reg_y[7][13] ), .X(n45898) );
  inv_x2_sg U54222 ( .A(\reg_y[4][13] ), .X(n45900) );
  inv_x2_sg U54223 ( .A(\reg_y[8][9] ), .X(n45902) );
  inv_x2_sg U54224 ( .A(\reg_y[6][9] ), .X(n45904) );
  inv_x2_sg U54225 ( .A(\reg_y[3][9] ), .X(n45906) );
  inv_x2_sg U54226 ( .A(\reg_y[4][9] ), .X(n45908) );
  inv_x2_sg U54227 ( .A(\reg_y[1][3] ), .X(n46062) );
  inv_x2_sg U54228 ( .A(\reg_y[2][9] ), .X(n45910) );
  inv_x2_sg U54229 ( .A(\reg_y[8][13] ), .X(n45912) );
  inv_x2_sg U54230 ( .A(\reg_y[6][13] ), .X(n45914) );
  inv_x2_sg U54231 ( .A(\reg_y[3][13] ), .X(n45916) );
  inv_x2_sg U54232 ( .A(\reg_y[11][3] ), .X(n46064) );
  inv_x2_sg U54233 ( .A(\reg_y[9][3] ), .X(n46066) );
  inv_x2_sg U54234 ( .A(\reg_y[13][3] ), .X(n46068) );
  inv_x2_sg U54235 ( .A(\reg_y[7][9] ), .X(n45918) );
  inv_x2_sg U54236 ( .A(\reg_y[4][3] ), .X(n46070) );
  inv_x2_sg U54237 ( .A(\reg_y[0][13] ), .X(n45920) );
  inv_x2_sg U54238 ( .A(\reg_y[5][12] ), .X(n45922) );
  inv_x2_sg U54239 ( .A(\reg_y[13][12] ), .X(n45924) );
  inv_x2_sg U54240 ( .A(\reg_y[11][12] ), .X(n45926) );
  inv_x2_sg U54241 ( .A(\reg_y[9][12] ), .X(n45928) );
  inv_x2_sg U54242 ( .A(\reg_y[13][9] ), .X(n45930) );
  inv_x2_sg U54243 ( .A(\reg_y[11][9] ), .X(n45932) );
  inv_x2_sg U54244 ( .A(\reg_y[9][9] ), .X(n45934) );
  inv_x2_sg U54245 ( .A(\reg_y[5][9] ), .X(n45936) );
  inv_x2_sg U54246 ( .A(\reg_y[2][3] ), .X(n46072) );
  inv_x2_sg U54247 ( .A(\reg_y[10][9] ), .X(n45938) );
  inv_x2_sg U54248 ( .A(\reg_y[7][3] ), .X(n46074) );
  inv_x2_sg U54249 ( .A(\reg_y[1][4] ), .X(n46076) );
  inv_x2_sg U54250 ( .A(\reg_y[14][9] ), .X(n45940) );
  inv_x2_sg U54251 ( .A(\reg_y[12][9] ), .X(n45942) );
  inv_x2_sg U54252 ( .A(\reg_y[0][9] ), .X(n45944) );
  inv_x2_sg U54253 ( .A(\reg_y[12][3] ), .X(n46078) );
  inv_x2_sg U54254 ( .A(\reg_y[14][3] ), .X(n46080) );
  inv_x2_sg U54255 ( .A(\reg_y[5][3] ), .X(n46082) );
  inv_x2_sg U54256 ( .A(\reg_y[0][3] ), .X(n46084) );
  inv_x2_sg U54257 ( .A(\reg_y[4][0] ), .X(n45946) );
  inv_x2_sg U54258 ( .A(\reg_y[1][7] ), .X(n46028) );
  nor_x1_sg U54259 ( .A(n25227), .B(n25228), .X(n25225) );
  nor_x1_sg U54260 ( .A(n10119), .B(n10120), .X(n10117) );
  nor_x1_sg U54261 ( .A(n18685), .B(n46335), .X(n18684) );
  nor_x2_sg U54262 ( .A(n18683), .B(n54289), .X(n18685) );
  nor_x1_sg U54263 ( .A(n40888), .B(n12030), .X(n12460) );
  nor_x1_sg U54264 ( .A(n11683), .B(n46537), .X(n11682) );
  nor_x2_sg U54265 ( .A(n11681), .B(n51777), .X(n11683) );
  nor_x1_sg U54266 ( .A(n40886), .B(n15925), .X(n16355) );
  inv_x4_sg U54267 ( .A(n43997), .X(n43998) );
  nand_x4_sg U54268 ( .A(n43998), .B(n18083), .X(n18081) );
  nor_x2_sg U54269 ( .A(n18187), .B(n18188), .X(n18186) );
  nor_x2_sg U54270 ( .A(n45284), .B(n46143), .X(n27546) );
  nor_x2_sg U54271 ( .A(n45308), .B(n46169), .X(n26987) );
  nand_x4_sg U54272 ( .A(n21648), .B(n21649), .X(n21581) );
  nand_x4_sg U54273 ( .A(n20103), .B(n20104), .X(n20036) );
  nand_x4_sg U54274 ( .A(n12339), .B(n12340), .X(n12270) );
  inv_x4_sg U54275 ( .A(n16507), .X(n55792) );
  inv_x4_sg U54276 ( .A(n43999), .X(n44000) );
  inv_x4_sg U54277 ( .A(n44001), .X(n44002) );
  inv_x4_sg U54278 ( .A(n44003), .X(n44004) );
  nand_x4_sg U54279 ( .A(n28398), .B(n54041), .X(n18184) );
  inv_x4_sg U54280 ( .A(n44005), .X(n44006) );
  inv_x2_sg U54281 ( .A(n44007), .X(n44008) );
  inv_x4_sg U54282 ( .A(n44009), .X(n44010) );
  inv_x2_sg U54283 ( .A(n44011), .X(n44012) );
  inv_x4_sg U54284 ( .A(n44013), .X(n44014) );
  inv_x2_sg U54285 ( .A(n44015), .X(n44016) );
  inv_x4_sg U54286 ( .A(n44017), .X(n44018) );
  inv_x2_sg U54287 ( .A(n44019), .X(n44020) );
  inv_x2_sg U54288 ( .A(n44023), .X(n44024) );
  inv_x2_sg U54289 ( .A(n44027), .X(n44028) );
  inv_x4_sg U54290 ( .A(n44029), .X(n44030) );
  inv_x2_sg U54291 ( .A(n44031), .X(n44032) );
  nand_x4_sg U54292 ( .A(n27000), .B(n52640), .X(n14295) );
  nand_x4_sg U54293 ( .A(n28955), .B(n54606), .X(n19730) );
  nand_x4_sg U54294 ( .A(n29516), .B(n55174), .X(n21275) );
  nand_x4_sg U54295 ( .A(n25603), .B(n51253), .X(n10403) );
  inv_x4_sg U54296 ( .A(n44033), .X(n44034) );
  inv_x4_sg U54297 ( .A(n44035), .X(n44036) );
  inv_x4_sg U54298 ( .A(n44037), .X(n44038) );
  inv_x4_sg U54299 ( .A(n44039), .X(n44040) );
  inv_x4_sg U54300 ( .A(n44041), .X(n44042) );
  inv_x4_sg U54301 ( .A(n44043), .X(n44044) );
  inv_x4_sg U54302 ( .A(n44045), .X(n44046) );
  inv_x4_sg U54303 ( .A(n44047), .X(n44048) );
  inv_x4_sg U54304 ( .A(n44049), .X(n44050) );
  inv_x4_sg U54305 ( .A(n44051), .X(n44052) );
  inv_x4_sg U54306 ( .A(n44053), .X(n44054) );
  inv_x4_sg U54307 ( .A(n44055), .X(n44056) );
  inv_x4_sg U54308 ( .A(n44057), .X(n44058) );
  inv_x4_sg U54309 ( .A(n44059), .X(n44060) );
  inv_x4_sg U54310 ( .A(n44061), .X(n44062) );
  inv_x4_sg U54311 ( .A(n44063), .X(n44064) );
  nor_x4_sg U54312 ( .A(n16190), .B(n46406), .X(n16477) );
  inv_x4_sg U54313 ( .A(n44065), .X(n44066) );
  inv_x4_sg U54314 ( .A(n44067), .X(n44068) );
  inv_x4_sg U54315 ( .A(n44069), .X(n44070) );
  inv_x4_sg U54316 ( .A(n44071), .X(n44072) );
  inv_x4_sg U54317 ( .A(n21315), .X(n55199) );
  nor_x4_sg U54318 ( .A(n46250), .B(n46254), .X(n21315) );
  inv_x4_sg U54319 ( .A(n19770), .X(n54631) );
  nor_x4_sg U54320 ( .A(n46295), .B(n46299), .X(n19770) );
  inv_x4_sg U54321 ( .A(n21885), .X(n55316) );
  nor_x4_sg U54322 ( .A(n21532), .B(n46250), .X(n21885) );
  inv_x4_sg U54323 ( .A(n20340), .X(n54748) );
  nor_x4_sg U54324 ( .A(n19987), .B(n46295), .X(n20340) );
  inv_x4_sg U54325 ( .A(n18796), .X(n54181) );
  nor_x4_sg U54326 ( .A(n18442), .B(n46340), .X(n18796) );
  nand_x8_sg U54327 ( .A(n46333), .B(n46345), .X(n18329) );
  inv_x4_sg U54328 ( .A(n44073), .X(n44074) );
  nor_x4_sg U54329 ( .A(n15989), .B(n15988), .X(n15983) );
  nor_x4_sg U54330 ( .A(n53262), .B(n15990), .X(n15988) );
  nor_x4_sg U54331 ( .A(n46404), .B(n53274), .X(n15990) );
  nor_x4_sg U54332 ( .A(n12094), .B(n12093), .X(n12088) );
  nor_x4_sg U54333 ( .A(n51875), .B(n12095), .X(n12093) );
  nor_x4_sg U54334 ( .A(n46516), .B(n51887), .X(n12095) );
  inv_x4_sg U54335 ( .A(n44075), .X(n44076) );
  nor_x4_sg U54336 ( .A(n16845), .B(n53592), .X(n16838) );
  inv_x4_sg U54337 ( .A(n16846), .X(n53592) );
  nand_x2_sg U54338 ( .A(n16847), .B(n16782), .X(n16846) );
  nand_x4_sg U54339 ( .A(n16785), .B(n16784), .X(n16782) );
  inv_x4_sg U54340 ( .A(n16061), .X(n53312) );
  nand_x2_sg U54341 ( .A(n16062), .B(n15997), .X(n16061) );
  nor_x4_sg U54342 ( .A(n15279), .B(n53034), .X(n15272) );
  inv_x4_sg U54343 ( .A(n15280), .X(n53034) );
  nand_x2_sg U54344 ( .A(n15281), .B(n15216), .X(n15280) );
  nand_x4_sg U54345 ( .A(n15219), .B(n15218), .X(n15216) );
  nor_x4_sg U54346 ( .A(n12946), .B(n52200), .X(n12939) );
  inv_x4_sg U54347 ( .A(n12947), .X(n52200) );
  nand_x2_sg U54348 ( .A(n12948), .B(n12883), .X(n12947) );
  nand_x4_sg U54349 ( .A(n12886), .B(n12885), .X(n12883) );
  nor_x4_sg U54350 ( .A(n12165), .B(n51924), .X(n12158) );
  inv_x4_sg U54351 ( .A(n12166), .X(n51924) );
  nand_x2_sg U54352 ( .A(n12167), .B(n12102), .X(n12166) );
  nand_x4_sg U54353 ( .A(n12105), .B(n12104), .X(n12102) );
  inv_x4_sg U54354 ( .A(n11386), .X(n51644) );
  nand_x2_sg U54355 ( .A(n11387), .B(n11322), .X(n11386) );
  inv_x4_sg U54356 ( .A(n21480), .X(n55281) );
  inv_x4_sg U54357 ( .A(n19935), .X(n54713) );
  inv_x4_sg U54358 ( .A(n18390), .X(n54148) );
  inv_x4_sg U54359 ( .A(n20610), .X(n54974) );
  inv_x4_sg U54360 ( .A(n19066), .X(n54406) );
  inv_x4_sg U54361 ( .A(n17521), .X(n53841) );
  inv_x4_sg U54362 ( .A(n13627), .X(n52443) );
  nor_x4_sg U54363 ( .A(n55512), .B(n26078), .X(n12609) );
  nand_x8_sg U54364 ( .A(n29376), .B(n21774), .X(n29383) );
  nor_x8_sg U54365 ( .A(n29368), .B(n55299), .X(n29376) );
  nand_x8_sg U54366 ( .A(n29094), .B(n20837), .X(n29101) );
  nor_x8_sg U54367 ( .A(n29087), .B(n55016), .X(n29094) );
  nand_x8_sg U54368 ( .A(n28815), .B(n20229), .X(n28822) );
  nor_x8_sg U54369 ( .A(n28807), .B(n54731), .X(n28815) );
  nand_x8_sg U54370 ( .A(n28535), .B(n19293), .X(n28542) );
  nor_x8_sg U54371 ( .A(n28528), .B(n54448), .X(n28535) );
  nand_x8_sg U54372 ( .A(n27977), .B(n17748), .X(n27984) );
  nor_x8_sg U54373 ( .A(n27970), .B(n53883), .X(n27977) );
  nor_x8_sg U54374 ( .A(n26865), .B(n52806), .X(n26872) );
  nand_x8_sg U54375 ( .A(n26858), .B(n14627), .X(n26865) );
  nand_x8_sg U54376 ( .A(n26580), .B(n13856), .X(n26587) );
  nor_x8_sg U54377 ( .A(n26573), .B(n52483), .X(n26580) );
  nand_x8_sg U54378 ( .A(n25464), .B(n46555), .X(n25471) );
  inv_x4_sg U54379 ( .A(n14791), .X(n52887) );
  nor_x4_sg U54380 ( .A(n14815), .B(n46452), .X(n14791) );
  nor_x4_sg U54381 ( .A(n18330), .B(n54097), .X(n18291) );
  nand_x4_sg U54382 ( .A(n46348), .B(n18198), .X(n18330) );
  nor_x4_sg U54383 ( .A(n55794), .B(n39300), .X(n39297) );
  inv_x4_sg U54384 ( .A(n39301), .X(n55794) );
  nor_x2_sg U54385 ( .A(n55795), .B(n39296), .X(n39301) );
  inv_x4_sg U54386 ( .A(n39303), .X(n55795) );
  nor_x4_sg U54387 ( .A(n46242), .B(n46248), .X(n21663) );
  nor_x4_sg U54388 ( .A(n46287), .B(n46293), .X(n20118) );
  nand_x2_sg U54389 ( .A(n21787), .B(n55442), .X(n29543) );
  nor_x2_sg U54390 ( .A(n21787), .B(n55442), .X(n21784) );
  inv_x4_sg U54391 ( .A(n21786), .X(n55442) );
  nand_x2_sg U54392 ( .A(n21016), .B(n55158), .X(n29265) );
  nor_x2_sg U54393 ( .A(n21016), .B(n55158), .X(n21013) );
  inv_x4_sg U54394 ( .A(n21015), .X(n55158) );
  nand_x2_sg U54395 ( .A(n20242), .B(n54874), .X(n28982) );
  nor_x2_sg U54396 ( .A(n20242), .B(n54874), .X(n20239) );
  inv_x4_sg U54397 ( .A(n20241), .X(n54874) );
  nand_x2_sg U54398 ( .A(n19472), .B(n54590), .X(n28704) );
  nor_x2_sg U54399 ( .A(n19472), .B(n54590), .X(n19469) );
  inv_x4_sg U54400 ( .A(n19471), .X(n54590) );
  nand_x2_sg U54401 ( .A(n18696), .B(n54306), .X(n28425) );
  nor_x2_sg U54402 ( .A(n18696), .B(n54306), .X(n18693) );
  inv_x4_sg U54403 ( .A(n18695), .X(n54306) );
  nand_x2_sg U54404 ( .A(n17927), .B(n54025), .X(n28146) );
  nor_x2_sg U54405 ( .A(n17927), .B(n54025), .X(n17924) );
  inv_x4_sg U54406 ( .A(n17926), .X(n54025) );
  nand_x2_sg U54407 ( .A(n17153), .B(n53741), .X(n27865) );
  nor_x2_sg U54408 ( .A(n17153), .B(n53741), .X(n17150) );
  inv_x4_sg U54409 ( .A(n17152), .X(n53741) );
  nand_x2_sg U54410 ( .A(n16368), .B(n53463), .X(n27586) );
  nor_x2_sg U54411 ( .A(n16368), .B(n53463), .X(n16365) );
  inv_x4_sg U54412 ( .A(n16367), .X(n53463) );
  nand_x2_sg U54413 ( .A(n15587), .B(n53183), .X(n27307) );
  nor_x2_sg U54414 ( .A(n15587), .B(n53183), .X(n15584) );
  inv_x4_sg U54415 ( .A(n15586), .X(n53183) );
  nand_x2_sg U54416 ( .A(n14806), .B(n52905), .X(n27027) );
  nor_x2_sg U54417 ( .A(n14806), .B(n52905), .X(n14803) );
  inv_x4_sg U54418 ( .A(n14805), .X(n52905) );
  nand_x2_sg U54419 ( .A(n14034), .B(n52624), .X(n26748) );
  nor_x2_sg U54420 ( .A(n14034), .B(n52624), .X(n14031) );
  inv_x4_sg U54421 ( .A(n14033), .X(n52624) );
  nand_x2_sg U54422 ( .A(n13254), .B(n52349), .X(n26470) );
  nor_x2_sg U54423 ( .A(n13254), .B(n52349), .X(n13251) );
  inv_x4_sg U54424 ( .A(n13253), .X(n52349) );
  nand_x2_sg U54425 ( .A(n12473), .B(n52071), .X(n26191) );
  nor_x2_sg U54426 ( .A(n12473), .B(n52071), .X(n12470) );
  inv_x4_sg U54427 ( .A(n12472), .X(n52071) );
  nand_x2_sg U54428 ( .A(n11694), .B(n51795), .X(n25911) );
  nor_x2_sg U54429 ( .A(n11694), .B(n51795), .X(n11691) );
  inv_x4_sg U54430 ( .A(n11693), .X(n51795) );
  nor_x4_sg U54431 ( .A(n14411), .B(n46449), .X(n14684) );
  nor_x4_sg U54432 ( .A(n46559), .B(n46570), .X(n10552) );
  nor_x4_sg U54433 ( .A(n46200), .B(n46582), .X(n29018) );
  nand_x2_sg U54434 ( .A(n26075), .B(n45421), .X(n26073) );
  nor_x2_sg U54435 ( .A(n51938), .B(n12197), .X(n12196) );
  inv_x4_sg U54436 ( .A(n12251), .X(n51938) );
  inv_x1_sg U54437 ( .A(n10835), .X(n51466) );
  inv_x4_sg U54438 ( .A(n44077), .X(n44078) );
  inv_x4_sg U54439 ( .A(n44079), .X(n44080) );
  inv_x4_sg U54440 ( .A(n44081), .X(n44082) );
  inv_x4_sg U54441 ( .A(n10435), .X(n51295) );
  nand_x4_sg U54442 ( .A(n44369), .B(n10427), .X(n10435) );
  inv_x1_sg U54443 ( .A(n14689), .X(n52840) );
  inv_x4_sg U54444 ( .A(n12522), .X(n52011) );
  nor_x4_sg U54445 ( .A(n12404), .B(n46521), .X(n12522) );
  inv_x4_sg U54446 ( .A(n14635), .X(n52778) );
  nor_x4_sg U54447 ( .A(n14552), .B(n46456), .X(n14635) );
  inv_x4_sg U54448 ( .A(n18524), .X(n54178) );
  nor_x4_sg U54449 ( .A(n18442), .B(n46346), .X(n18524) );
  nand_x4_sg U54450 ( .A(n53215), .B(n15845), .X(n15851) );
  nand_x4_sg U54451 ( .A(n52379), .B(n13512), .X(n13517) );
  nand_x4_sg U54452 ( .A(n51827), .B(n11950), .X(n11956) );
  inv_x1_sg U54453 ( .A(n20899), .X(n55093) );
  inv_x1_sg U54454 ( .A(n19355), .X(n54525) );
  inv_x1_sg U54455 ( .A(n17810), .X(n53960) );
  inv_x1_sg U54456 ( .A(n21706), .X(n55394) );
  inv_x1_sg U54457 ( .A(n20161), .X(n54826) );
  inv_x1_sg U54458 ( .A(n18615), .X(n54259) );
  inv_x1_sg U54459 ( .A(n12396), .X(n52028) );
  inv_x1_sg U54460 ( .A(n16291), .X(n53415) );
  nand_x4_sg U54461 ( .A(n54117), .B(n18247), .X(n18232) );
  inv_x4_sg U54462 ( .A(n17181), .X(n53688) );
  nand_x4_sg U54463 ( .A(n53687), .B(n17222), .X(n17181) );
  inv_x4_sg U54464 ( .A(n15615), .X(n53130) );
  nand_x4_sg U54465 ( .A(n53129), .B(n15656), .X(n15615) );
  inv_x4_sg U54466 ( .A(n13282), .X(n52296) );
  nand_x4_sg U54467 ( .A(n52295), .B(n13323), .X(n13282) );
  inv_x4_sg U54468 ( .A(n12501), .X(n52020) );
  nand_x4_sg U54469 ( .A(n52019), .B(n12542), .X(n12501) );
  inv_x4_sg U54470 ( .A(n21207), .X(n55329) );
  nand_x4_sg U54471 ( .A(n21198), .B(n21252), .X(n21207) );
  inv_x4_sg U54472 ( .A(n20434), .X(n55047) );
  nand_x4_sg U54473 ( .A(n20425), .B(n20480), .X(n20434) );
  inv_x4_sg U54474 ( .A(n19662), .X(n54761) );
  nand_x4_sg U54475 ( .A(n19653), .B(n19707), .X(n19662) );
  inv_x4_sg U54476 ( .A(n18890), .X(n54479) );
  nand_x4_sg U54477 ( .A(n18881), .B(n18936), .X(n18890) );
  inv_x4_sg U54478 ( .A(n18117), .X(n54194) );
  nand_x4_sg U54479 ( .A(n18108), .B(n18162), .X(n18117) );
  inv_x4_sg U54480 ( .A(n17345), .X(n53914) );
  nand_x4_sg U54481 ( .A(n17336), .B(n17391), .X(n17345) );
  inv_x4_sg U54482 ( .A(n16562), .X(n53630) );
  nand_x4_sg U54483 ( .A(n16553), .B(n16607), .X(n16562) );
  inv_x4_sg U54484 ( .A(n15780), .X(n53351) );
  nand_x4_sg U54485 ( .A(n15771), .B(n15825), .X(n15780) );
  inv_x4_sg U54486 ( .A(n14996), .X(n53072) );
  nand_x4_sg U54487 ( .A(n14987), .B(n15041), .X(n14996) );
  inv_x4_sg U54488 ( .A(n14226), .X(n52794) );
  nand_x4_sg U54489 ( .A(n14217), .B(n14272), .X(n14226) );
  inv_x4_sg U54490 ( .A(n13447), .X(n52515) );
  nand_x4_sg U54491 ( .A(n13438), .B(n13492), .X(n13447) );
  inv_x4_sg U54492 ( .A(n12663), .X(n52238) );
  nand_x4_sg U54493 ( .A(n12654), .B(n12708), .X(n12663) );
  inv_x4_sg U54494 ( .A(n11885), .X(n51963) );
  nand_x4_sg U54495 ( .A(n11876), .B(n11930), .X(n11885) );
  inv_x4_sg U54496 ( .A(n11102), .X(n51682) );
  nand_x4_sg U54497 ( .A(n11093), .B(n11147), .X(n11102) );
  inv_x4_sg U54498 ( .A(n10334), .X(n51405) );
  nand_x4_sg U54499 ( .A(n10325), .B(n10380), .X(n10334) );
  nand_x4_sg U54500 ( .A(n53518), .B(n16984), .X(n16979) );
  inv_x4_sg U54501 ( .A(n16676), .X(n53518) );
  nand_x4_sg U54502 ( .A(n52960), .B(n15418), .X(n15413) );
  inv_x4_sg U54503 ( .A(n15110), .X(n52960) );
  nand_x4_sg U54504 ( .A(n52126), .B(n13085), .X(n13080) );
  inv_x4_sg U54505 ( .A(n12777), .X(n52126) );
  nand_x4_sg U54506 ( .A(n51569), .B(n11524), .X(n11519) );
  inv_x4_sg U54507 ( .A(n11216), .X(n51569) );
  inv_x4_sg U54508 ( .A(n16421), .X(n53441) );
  inv_x4_sg U54509 ( .A(n10963), .X(n51492) );
  nor_x4_sg U54510 ( .A(n18654), .B(n46337), .X(n18691) );
  inv_x4_sg U54511 ( .A(n44407), .X(n53692) );
  inv_x4_sg U54512 ( .A(n44409), .X(n53134) );
  inv_x4_sg U54513 ( .A(n44411), .X(n52575) );
  inv_x4_sg U54514 ( .A(n44413), .X(n52300) );
  nor_x2_sg U54515 ( .A(n40771), .B(n50824), .X(n23069) );
  inv_x4_sg U54516 ( .A(n22819), .X(n50824) );
  inv_x4_sg U54517 ( .A(n21878), .X(n55305) );
  inv_x4_sg U54518 ( .A(n20333), .X(n54737) );
  nor_x4_sg U54519 ( .A(n21527), .B(n46254), .X(n21525) );
  nor_x4_sg U54520 ( .A(n20757), .B(n46274), .X(n20755) );
  nor_x4_sg U54521 ( .A(n19982), .B(n46299), .X(n19980) );
  nor_x4_sg U54522 ( .A(n19213), .B(n46319), .X(n19211) );
  inv_x4_sg U54523 ( .A(n18787), .X(n54171) );
  nor_x4_sg U54524 ( .A(n17668), .B(n46366), .X(n17666) );
  nor_x4_sg U54525 ( .A(n13775), .B(n46479), .X(n13773) );
  inv_x4_sg U54526 ( .A(n11000), .X(n51383) );
  nand_x4_sg U54527 ( .A(n51435), .B(n46569), .X(n11020) );
  inv_x4_sg U54528 ( .A(n16119), .X(n53344) );
  inv_x4_sg U54529 ( .A(n11444), .X(n51675) );
  inv_x4_sg U54530 ( .A(n16972), .X(n53621) );
  nor_x4_sg U54531 ( .A(n16975), .B(n46396), .X(n16972) );
  inv_x4_sg U54532 ( .A(n15406), .X(n53063) );
  nor_x4_sg U54533 ( .A(n15409), .B(n46440), .X(n15406) );
  inv_x4_sg U54534 ( .A(n13853), .X(n52506) );
  nor_x4_sg U54535 ( .A(n13856), .B(n46485), .X(n13853) );
  inv_x4_sg U54536 ( .A(n13073), .X(n52229) );
  nor_x4_sg U54537 ( .A(n13076), .B(n46508), .X(n13073) );
  inv_x4_sg U54538 ( .A(n12292), .X(n51954) );
  nor_x4_sg U54539 ( .A(n12295), .B(n46528), .X(n12292) );
  nor_x2_sg U54540 ( .A(n51460), .B(n11002), .X(n11010) );
  inv_x4_sg U54541 ( .A(n44503), .X(n51460) );
  nor_x2_sg U54542 ( .A(n53605), .B(n16877), .X(n16876) );
  inv_x4_sg U54543 ( .A(n16931), .X(n53605) );
  nor_x2_sg U54544 ( .A(n53047), .B(n15311), .X(n15310) );
  inv_x4_sg U54545 ( .A(n15365), .X(n53047) );
  nor_x2_sg U54546 ( .A(n52490), .B(n13758), .X(n13757) );
  inv_x4_sg U54547 ( .A(n13812), .X(n52490) );
  nor_x2_sg U54548 ( .A(n52213), .B(n12978), .X(n12977) );
  inv_x4_sg U54549 ( .A(n13032), .X(n52213) );
  nor_x2_sg U54550 ( .A(n55300), .B(n21510), .X(n21509) );
  inv_x4_sg U54551 ( .A(n21562), .X(n55300) );
  nor_x2_sg U54552 ( .A(n54732), .B(n19965), .X(n19964) );
  inv_x4_sg U54553 ( .A(n20017), .X(n54732) );
  nor_x2_sg U54554 ( .A(n52764), .B(n14530), .X(n14529) );
  inv_x4_sg U54555 ( .A(n14582), .X(n52764) );
  nor_x4_sg U54556 ( .A(n21796), .B(n46254), .X(n21794) );
  nor_x4_sg U54557 ( .A(n20251), .B(n46299), .X(n20249) );
  nor_x4_sg U54558 ( .A(n12482), .B(n46523), .X(n12480) );
  nor_x4_sg U54559 ( .A(n46449), .B(n46456), .X(n14354) );
  nor_x4_sg U54560 ( .A(n46297), .B(n46306), .X(n19722) );
  nor_x4_sg U54561 ( .A(n46409), .B(n46416), .X(n15840) );
  nor_x4_sg U54562 ( .A(n46377), .B(n16894), .X(n17251) );
  nor_x4_sg U54563 ( .A(n46421), .B(n15328), .X(n15685) );
  nor_x4_sg U54564 ( .A(n46489), .B(n12995), .X(n13352) );
  inv_x4_sg U54565 ( .A(n21797), .X(n55387) );
  inv_x4_sg U54566 ( .A(n21026), .X(n55102) );
  inv_x4_sg U54567 ( .A(n20252), .X(n54819) );
  inv_x4_sg U54568 ( .A(n19482), .X(n54534) );
  inv_x4_sg U54569 ( .A(n18706), .X(n54251) );
  inv_x4_sg U54570 ( .A(n17937), .X(n53969) );
  inv_x4_sg U54571 ( .A(n14816), .X(n52849) );
  inv_x4_sg U54572 ( .A(n11704), .X(n51739) );
  inv_x4_sg U54573 ( .A(n21845), .X(n55417) );
  inv_x4_sg U54574 ( .A(n20300), .X(n54849) );
  inv_x4_sg U54575 ( .A(n18754), .X(n54282) );
  nor_x4_sg U54576 ( .A(n16378), .B(n46411), .X(n16376) );
  nor_x2_sg U54577 ( .A(n12339), .B(n12342), .X(n12341) );
  nor_x4_sg U54578 ( .A(n12344), .B(n46528), .X(n12342) );
  inv_x4_sg U54579 ( .A(n44083), .X(n44084) );
  inv_x4_sg U54580 ( .A(n44085), .X(n44086) );
  inv_x4_sg U54581 ( .A(n44087), .X(n44088) );
  inv_x4_sg U54582 ( .A(n44089), .X(n44090) );
  inv_x4_sg U54583 ( .A(n44091), .X(n44092) );
  inv_x4_sg U54584 ( .A(n44093), .X(n44094) );
  inv_x4_sg U54585 ( .A(n44095), .X(n44096) );
  inv_x4_sg U54586 ( .A(n11752), .X(n51770) );
  nor_x2_sg U54587 ( .A(n54074), .B(n54062), .X(n18185) );
  inv_x4_sg U54588 ( .A(n18188), .X(n54062) );
  nor_x2_sg U54589 ( .A(n52674), .B(n52665), .X(n14296) );
  inv_x4_sg U54590 ( .A(n14299), .X(n52665) );
  nor_x2_sg U54591 ( .A(n20879), .B(n20882), .X(n20881) );
  nor_x4_sg U54592 ( .A(n20884), .B(n46281), .X(n20882) );
  nor_x2_sg U54593 ( .A(n19335), .B(n19338), .X(n19337) );
  nor_x4_sg U54594 ( .A(n19340), .B(n46326), .X(n19338) );
  nor_x2_sg U54595 ( .A(n17790), .B(n17793), .X(n17792) );
  nor_x4_sg U54596 ( .A(n17795), .B(n46373), .X(n17793) );
  nor_x2_sg U54597 ( .A(n16234), .B(n16237), .X(n16236) );
  nor_x4_sg U54598 ( .A(n16239), .B(n46416), .X(n16237) );
  nor_x2_sg U54599 ( .A(n10777), .B(n10780), .X(n10779) );
  nor_x4_sg U54600 ( .A(n10782), .B(n46573), .X(n10780) );
  nor_x2_sg U54601 ( .A(n21648), .B(n21651), .X(n21650) );
  nor_x4_sg U54602 ( .A(n21653), .B(n46261), .X(n21651) );
  nor_x2_sg U54603 ( .A(n20103), .B(n20106), .X(n20105) );
  nor_x4_sg U54604 ( .A(n20108), .B(n46306), .X(n20106) );
  nor_x2_sg U54605 ( .A(n53569), .B(n53560), .X(n16808) );
  inv_x4_sg U54606 ( .A(n16810), .X(n53560) );
  nor_x2_sg U54607 ( .A(n53011), .B(n53002), .X(n15242) );
  inv_x4_sg U54608 ( .A(n15244), .X(n53002) );
  nor_x2_sg U54609 ( .A(n52452), .B(n52442), .X(n13689) );
  inv_x4_sg U54610 ( .A(n13691), .X(n52442) );
  nor_x2_sg U54611 ( .A(n52177), .B(n52168), .X(n12909) );
  inv_x4_sg U54612 ( .A(n12911), .X(n52168) );
  inv_x4_sg U54613 ( .A(n15960), .X(n53274) );
  inv_x4_sg U54614 ( .A(n12065), .X(n51887) );
  nor_x2_sg U54615 ( .A(n55004), .B(n54968), .X(n20650) );
  inv_x4_sg U54616 ( .A(n20653), .X(n54968) );
  nor_x2_sg U54617 ( .A(n54436), .B(n54400), .X(n19106) );
  inv_x4_sg U54618 ( .A(n19109), .X(n54400) );
  nor_x2_sg U54619 ( .A(n53871), .B(n53835), .X(n17561) );
  inv_x4_sg U54620 ( .A(n17564), .X(n53835) );
  nor_x2_sg U54621 ( .A(n52751), .B(n52708), .X(n14441) );
  inv_x4_sg U54622 ( .A(n14444), .X(n52708) );
  nor_x2_sg U54623 ( .A(n51160), .B(n45271), .X(n28384) );
  inv_x4_sg U54624 ( .A(n46117), .X(n51160) );
  nor_x4_sg U54625 ( .A(n46252), .B(n46261), .X(n21267) );
  nor_x4_sg U54626 ( .A(n46454), .B(n46463), .X(n14287) );
  inv_x4_sg U54627 ( .A(n16357), .X(n53424) );
  nor_x4_sg U54628 ( .A(n46331), .B(n46353), .X(n18300) );
  inv_x4_sg U54629 ( .A(n17120), .X(n53733) );
  inv_x4_sg U54630 ( .A(n15554), .X(n53175) );
  inv_x4_sg U54631 ( .A(n14001), .X(n52616) );
  inv_x4_sg U54632 ( .A(n13221), .X(n52341) );
  inv_x4_sg U54633 ( .A(n12440), .X(n52064) );
  inv_x4_sg U54634 ( .A(n16335), .X(n53452) );
  nor_x4_sg U54635 ( .A(n46246), .B(n55202), .X(n21454) );
  nor_x4_sg U54636 ( .A(n46291), .B(n54634), .X(n19909) );
  nor_x4_sg U54637 ( .A(n46335), .B(n54070), .X(n18364) );
  nor_x4_sg U54638 ( .A(n46447), .B(n52670), .X(n14474) );
  nor_x4_sg U54639 ( .A(n46537), .B(n46539), .X(n11356) );
  nor_x4_sg U54640 ( .A(n10518), .B(n51280), .X(n10582) );
  nor_x4_sg U54641 ( .A(n46516), .B(n46514), .X(n12255) );
  nand_x4_sg U54642 ( .A(n53641), .B(n46395), .X(n17023) );
  nand_x4_sg U54643 ( .A(n53083), .B(n46439), .X(n15457) );
  nand_x4_sg U54644 ( .A(n52249), .B(n46507), .X(n13124) );
  nand_x4_sg U54645 ( .A(n51693), .B(n46551), .X(n11563) );
  inv_x8_sg U54646 ( .A(n11638), .X(n51693) );
  inv_x1_sg U54647 ( .A(n11018), .X(n51415) );
  nand_x4_sg U54648 ( .A(n10880), .B(n11040), .X(n10961) );
  nand_x4_sg U54649 ( .A(n10879), .B(n44379), .X(n10880) );
  inv_x4_sg U54650 ( .A(n20716), .X(n55002) );
  nor_x4_sg U54651 ( .A(n20717), .B(n46281), .X(n20716) );
  inv_x4_sg U54652 ( .A(n19172), .X(n54434) );
  nor_x4_sg U54653 ( .A(n19173), .B(n46326), .X(n19172) );
  inv_x4_sg U54654 ( .A(n17627), .X(n53869) );
  nor_x4_sg U54655 ( .A(n17628), .B(n46373), .X(n17627) );
  inv_x4_sg U54656 ( .A(n14506), .X(n52749) );
  nor_x4_sg U54657 ( .A(n14507), .B(n46463), .X(n14506) );
  inv_x4_sg U54658 ( .A(n44097), .X(n44098) );
  inv_x4_sg U54659 ( .A(n44099), .X(n44100) );
  nand_x4_sg U54660 ( .A(n18525), .B(n54078), .X(n18520) );
  inv_x4_sg U54661 ( .A(n18223), .X(n54078) );
  nor_x4_sg U54662 ( .A(n46379), .B(n46389), .X(n16785) );
  nor_x4_sg U54663 ( .A(n46423), .B(n46433), .X(n15219) );
  nor_x4_sg U54664 ( .A(n46491), .B(n46501), .X(n12886) );
  nor_x4_sg U54665 ( .A(n46535), .B(n46545), .X(n11325) );
  nor_x4_sg U54666 ( .A(n46467), .B(n46479), .X(n13666) );
  nor_x2_sg U54667 ( .A(n10286), .B(n51257), .X(n10285) );
  inv_x4_sg U54668 ( .A(n10283), .X(n51257) );
  nor_x2_sg U54669 ( .A(n51104), .B(n45285), .X(n27545) );
  inv_x4_sg U54670 ( .A(n46143), .X(n51104) );
  inv_x4_sg U54671 ( .A(n44101), .X(n44102) );
  nand_x4_sg U54672 ( .A(n44102), .B(n11659), .X(n11660) );
  nor_x2_sg U54673 ( .A(n51066), .B(n45309), .X(n26986) );
  inv_x4_sg U54674 ( .A(n46169), .X(n51066) );
  inv_x4_sg U54675 ( .A(n44103), .X(n44104) );
  inv_x4_sg U54676 ( .A(n44105), .X(n44106) );
  nor_x4_sg U54677 ( .A(n46400), .B(n46411), .X(n16000) );
  inv_x4_sg U54678 ( .A(n21345), .X(n55236) );
  inv_x4_sg U54679 ( .A(n19800), .X(n54668) );
  inv_x4_sg U54680 ( .A(n13590), .X(n52426) );
  inv_x4_sg U54681 ( .A(n12025), .X(n51874) );
  inv_x2_sg U54682 ( .A(\reg_yHat[13][19] ), .X(n44760) );
  inv_x2_sg U54683 ( .A(\reg_yHat[12][19] ), .X(n44762) );
  inv_x2_sg U54684 ( .A(\reg_yHat[10][19] ), .X(n44766) );
  inv_x2_sg U54685 ( .A(\reg_yHat[9][19] ), .X(n44768) );
  inv_x2_sg U54686 ( .A(\reg_yHat[8][19] ), .X(n44770) );
  inv_x2_sg U54687 ( .A(\reg_yHat[6][19] ), .X(n44774) );
  inv_x2_sg U54688 ( .A(\reg_yHat[5][19] ), .X(n44776) );
  inv_x2_sg U54689 ( .A(\reg_yHat[4][19] ), .X(n44778) );
  inv_x2_sg U54690 ( .A(\reg_yHat[3][19] ), .X(n44780) );
  inv_x2_sg U54691 ( .A(\reg_yHat[1][6] ), .X(n44792) );
  inv_x2_sg U54692 ( .A(\reg_yHat[0][6] ), .X(n45634) );
  inv_x2_sg U54693 ( .A(\reg_yHat[7][6] ), .X(n45636) );
  inv_x2_sg U54694 ( .A(\reg_yHat[2][6] ), .X(n45638) );
  inv_x2_sg U54695 ( .A(\reg_yHat[13][7] ), .X(n44796) );
  inv_x2_sg U54696 ( .A(\reg_yHat[11][7] ), .X(n44798) );
  inv_x2_sg U54697 ( .A(\reg_yHat[9][7] ), .X(n44800) );
  inv_x2_sg U54698 ( .A(\reg_yHat[10][7] ), .X(n45982) );
  inv_x2_sg U54699 ( .A(\reg_y[4][7] ), .X(n45226) );
  inv_x2_sg U54700 ( .A(\reg_yHat[13][6] ), .X(n44808) );
  inv_x2_sg U54701 ( .A(\reg_yHat[11][6] ), .X(n44810) );
  inv_x2_sg U54702 ( .A(\reg_yHat[9][6] ), .X(n44812) );
  inv_x2_sg U54703 ( .A(\reg_yHat[10][1] ), .X(n45984) );
  inv_x2_sg U54704 ( .A(\reg_y[14][7] ), .X(n45228) );
  inv_x2_sg U54705 ( .A(\reg_y[12][7] ), .X(n45230) );
  inv_x2_sg U54706 ( .A(\reg_y[7][7] ), .X(n45232) );
  inv_x2_sg U54707 ( .A(\reg_y[10][0] ), .X(n45552) );
  inv_x2_sg U54708 ( .A(\reg_y[2][7] ), .X(n45234) );
  inv_x2_sg U54709 ( .A(\reg_yHat[10][5] ), .X(n45986) );
  inv_x2_sg U54710 ( .A(\reg_y[0][7] ), .X(n45236) );
  inv_x2_sg U54711 ( .A(\reg_yHat[10][6] ), .X(n44832) );
  inv_x2_sg U54712 ( .A(\reg_y[10][2] ), .X(n44836) );
  inv_x2_sg U54713 ( .A(\reg_y[2][0] ), .X(n45554) );
  inv_x2_sg U54714 ( .A(\reg_yHat[4][6] ), .X(n45640) );
  inv_x2_sg U54715 ( .A(\reg_y[7][0] ), .X(n45556) );
  inv_x2_sg U54716 ( .A(\reg_y[13][5] ), .X(n45988) );
  inv_x2_sg U54717 ( .A(\reg_y[11][5] ), .X(n45990) );
  inv_x2_sg U54718 ( .A(\reg_y[9][5] ), .X(n45992) );
  inv_x2_sg U54719 ( .A(\reg_y[13][0] ), .X(n45558) );
  inv_x2_sg U54720 ( .A(\reg_y[11][0] ), .X(n45560) );
  inv_x2_sg U54721 ( .A(\reg_y[9][0] ), .X(n45562) );
  inv_x2_sg U54722 ( .A(\reg_yHat[8][4] ), .X(n44848) );
  inv_x2_sg U54723 ( .A(\reg_yHat[6][4] ), .X(n44850) );
  inv_x2_sg U54724 ( .A(\reg_yHat[3][4] ), .X(n44852) );
  inv_x2_sg U54725 ( .A(\reg_yHat[14][6] ), .X(n45642) );
  inv_x2_sg U54726 ( .A(\reg_yHat[12][6] ), .X(n45644) );
  nor_x2_sg U54727 ( .A(n21436), .B(n44423), .X(n21473) );
  nor_x2_sg U54728 ( .A(n19891), .B(n44425), .X(n19928) );
  nor_x2_sg U54729 ( .A(n10564), .B(n44427), .X(n10601) );
  inv_x2_sg U54730 ( .A(\reg_yHat[14][17] ), .X(n44908) );
  inv_x2_sg U54731 ( .A(\reg_yHat[14][16] ), .X(n44910) );
  inv_x2_sg U54732 ( .A(\reg_yHat[14][15] ), .X(n44912) );
  inv_x2_sg U54733 ( .A(\reg_yHat[14][12] ), .X(n44914) );
  inv_x2_sg U54734 ( .A(\reg_yHat[14][11] ), .X(n44916) );
  inv_x2_sg U54735 ( .A(\reg_yHat[14][10] ), .X(n44918) );
  inv_x2_sg U54736 ( .A(\reg_yHat[14][8] ), .X(n44920) );
  inv_x2_sg U54737 ( .A(\reg_yHat[13][17] ), .X(n44922) );
  inv_x2_sg U54738 ( .A(\reg_yHat[13][16] ), .X(n44924) );
  inv_x2_sg U54739 ( .A(\reg_yHat[13][15] ), .X(n44926) );
  inv_x2_sg U54740 ( .A(\reg_yHat[13][13] ), .X(n44928) );
  inv_x2_sg U54741 ( .A(\reg_yHat[13][11] ), .X(n44930) );
  inv_x2_sg U54742 ( .A(\reg_yHat[13][10] ), .X(n44932) );
  inv_x2_sg U54743 ( .A(\reg_yHat[13][8] ), .X(n44934) );
  inv_x2_sg U54744 ( .A(\reg_yHat[12][17] ), .X(n44936) );
  inv_x2_sg U54745 ( .A(\reg_yHat[12][16] ), .X(n44938) );
  inv_x2_sg U54746 ( .A(\reg_yHat[12][15] ), .X(n44940) );
  inv_x2_sg U54747 ( .A(\reg_yHat[12][12] ), .X(n44942) );
  inv_x2_sg U54748 ( .A(\reg_yHat[12][11] ), .X(n44944) );
  inv_x2_sg U54749 ( .A(\reg_yHat[12][10] ), .X(n44946) );
  inv_x2_sg U54750 ( .A(\reg_yHat[12][8] ), .X(n44948) );
  inv_x2_sg U54751 ( .A(\reg_yHat[11][17] ), .X(n44950) );
  inv_x2_sg U54752 ( .A(\reg_yHat[11][16] ), .X(n44952) );
  inv_x2_sg U54753 ( .A(\reg_yHat[11][15] ), .X(n44954) );
  inv_x2_sg U54754 ( .A(\reg_yHat[11][13] ), .X(n44956) );
  inv_x2_sg U54755 ( .A(\reg_yHat[11][11] ), .X(n44958) );
  inv_x2_sg U54756 ( .A(\reg_yHat[11][10] ), .X(n44960) );
  inv_x2_sg U54757 ( .A(\reg_yHat[11][8] ), .X(n44962) );
  inv_x2_sg U54758 ( .A(\reg_yHat[10][17] ), .X(n44964) );
  inv_x2_sg U54759 ( .A(\reg_yHat[10][16] ), .X(n44966) );
  inv_x2_sg U54760 ( .A(\reg_yHat[10][15] ), .X(n44968) );
  inv_x2_sg U54761 ( .A(\reg_yHat[10][14] ), .X(n44970) );
  inv_x2_sg U54762 ( .A(\reg_yHat[10][13] ), .X(n44972) );
  inv_x2_sg U54763 ( .A(\reg_yHat[10][12] ), .X(n44974) );
  inv_x2_sg U54764 ( .A(\reg_yHat[10][11] ), .X(n44976) );
  inv_x2_sg U54765 ( .A(\reg_yHat[10][10] ), .X(n44978) );
  inv_x2_sg U54766 ( .A(\reg_yHat[10][8] ), .X(n44980) );
  inv_x2_sg U54767 ( .A(\reg_yHat[9][17] ), .X(n44982) );
  inv_x2_sg U54768 ( .A(\reg_yHat[9][16] ), .X(n44984) );
  inv_x2_sg U54769 ( .A(\reg_yHat[9][15] ), .X(n44986) );
  inv_x2_sg U54770 ( .A(\reg_yHat[9][13] ), .X(n44988) );
  inv_x2_sg U54771 ( .A(\reg_yHat[9][11] ), .X(n44990) );
  inv_x2_sg U54772 ( .A(\reg_yHat[9][10] ), .X(n44992) );
  inv_x2_sg U54773 ( .A(\reg_yHat[9][8] ), .X(n44994) );
  inv_x2_sg U54774 ( .A(\reg_yHat[8][17] ), .X(n44996) );
  inv_x2_sg U54775 ( .A(\reg_yHat[8][16] ), .X(n44998) );
  inv_x2_sg U54776 ( .A(\reg_yHat[8][15] ), .X(n45000) );
  inv_x2_sg U54777 ( .A(\reg_yHat[8][14] ), .X(n45002) );
  inv_x2_sg U54778 ( .A(\reg_yHat[8][12] ), .X(n45004) );
  inv_x2_sg U54779 ( .A(\reg_yHat[8][10] ), .X(n45006) );
  inv_x2_sg U54780 ( .A(\reg_yHat[8][8] ), .X(n45008) );
  inv_x2_sg U54781 ( .A(\reg_yHat[7][17] ), .X(n45010) );
  inv_x2_sg U54782 ( .A(\reg_yHat[7][16] ), .X(n45012) );
  inv_x2_sg U54783 ( .A(\reg_yHat[7][15] ), .X(n45014) );
  inv_x2_sg U54784 ( .A(\reg_yHat[7][14] ), .X(n45016) );
  inv_x2_sg U54785 ( .A(\reg_yHat[7][12] ), .X(n45018) );
  inv_x2_sg U54786 ( .A(\reg_yHat[7][11] ), .X(n45020) );
  inv_x2_sg U54787 ( .A(\reg_yHat[7][10] ), .X(n45022) );
  inv_x2_sg U54788 ( .A(\reg_yHat[7][8] ), .X(n45024) );
  inv_x2_sg U54789 ( .A(\reg_yHat[6][17] ), .X(n45026) );
  inv_x2_sg U54790 ( .A(\reg_yHat[6][16] ), .X(n45028) );
  inv_x2_sg U54791 ( .A(\reg_yHat[6][15] ), .X(n45030) );
  inv_x2_sg U54792 ( .A(\reg_yHat[6][14] ), .X(n45032) );
  inv_x2_sg U54793 ( .A(\reg_yHat[6][12] ), .X(n45034) );
  inv_x2_sg U54794 ( .A(\reg_yHat[6][10] ), .X(n45036) );
  inv_x2_sg U54795 ( .A(\reg_yHat[6][8] ), .X(n45038) );
  inv_x2_sg U54796 ( .A(\reg_yHat[5][17] ), .X(n45040) );
  inv_x2_sg U54797 ( .A(\reg_yHat[5][16] ), .X(n45042) );
  inv_x2_sg U54798 ( .A(\reg_yHat[5][15] ), .X(n45044) );
  inv_x2_sg U54799 ( .A(\reg_yHat[5][13] ), .X(n45046) );
  inv_x2_sg U54800 ( .A(\reg_yHat[5][11] ), .X(n45048) );
  inv_x2_sg U54801 ( .A(\reg_yHat[5][10] ), .X(n45050) );
  inv_x2_sg U54802 ( .A(\reg_yHat[5][8] ), .X(n45052) );
  inv_x2_sg U54803 ( .A(\reg_yHat[4][17] ), .X(n45054) );
  inv_x2_sg U54804 ( .A(\reg_yHat[4][16] ), .X(n45056) );
  inv_x2_sg U54805 ( .A(\reg_yHat[4][15] ), .X(n45058) );
  inv_x2_sg U54806 ( .A(\reg_yHat[4][14] ), .X(n45060) );
  inv_x2_sg U54807 ( .A(\reg_yHat[4][12] ), .X(n45062) );
  inv_x2_sg U54808 ( .A(\reg_yHat[4][10] ), .X(n45064) );
  inv_x2_sg U54809 ( .A(\reg_yHat[4][8] ), .X(n45066) );
  inv_x2_sg U54810 ( .A(\reg_yHat[3][17] ), .X(n45068) );
  inv_x2_sg U54811 ( .A(\reg_yHat[3][16] ), .X(n45070) );
  inv_x2_sg U54812 ( .A(\reg_yHat[3][15] ), .X(n45072) );
  inv_x2_sg U54813 ( .A(\reg_yHat[3][14] ), .X(n45074) );
  inv_x2_sg U54814 ( .A(\reg_yHat[3][12] ), .X(n45076) );
  inv_x2_sg U54815 ( .A(\reg_yHat[3][10] ), .X(n45078) );
  inv_x2_sg U54816 ( .A(\reg_yHat[3][8] ), .X(n45080) );
  inv_x2_sg U54817 ( .A(\reg_yHat[2][17] ), .X(n45082) );
  inv_x2_sg U54818 ( .A(\reg_yHat[2][16] ), .X(n45084) );
  inv_x2_sg U54819 ( .A(\reg_yHat[2][15] ), .X(n45086) );
  inv_x2_sg U54820 ( .A(\reg_yHat[2][14] ), .X(n45088) );
  inv_x2_sg U54821 ( .A(\reg_yHat[2][12] ), .X(n45090) );
  inv_x2_sg U54822 ( .A(\reg_yHat[2][11] ), .X(n45092) );
  inv_x2_sg U54823 ( .A(\reg_yHat[2][10] ), .X(n45094) );
  inv_x2_sg U54824 ( .A(\reg_yHat[2][8] ), .X(n45096) );
  inv_x2_sg U54825 ( .A(\reg_yHat[1][17] ), .X(n45098) );
  inv_x2_sg U54826 ( .A(\reg_yHat[1][16] ), .X(n45100) );
  inv_x2_sg U54827 ( .A(\reg_yHat[1][15] ), .X(n45102) );
  inv_x2_sg U54828 ( .A(\reg_yHat[1][14] ), .X(n45104) );
  inv_x2_sg U54829 ( .A(\reg_yHat[1][12] ), .X(n45106) );
  inv_x2_sg U54830 ( .A(\reg_yHat[1][11] ), .X(n45108) );
  inv_x2_sg U54831 ( .A(\reg_yHat[1][10] ), .X(n45110) );
  inv_x2_sg U54832 ( .A(\reg_yHat[1][8] ), .X(n45112) );
  inv_x2_sg U54833 ( .A(\reg_yHat[0][15] ), .X(n45114) );
  inv_x2_sg U54834 ( .A(\reg_yHat[0][14] ), .X(n45116) );
  inv_x2_sg U54835 ( .A(\reg_yHat[0][12] ), .X(n45118) );
  inv_x2_sg U54836 ( .A(\reg_yHat[0][11] ), .X(n45120) );
  inv_x2_sg U54837 ( .A(\reg_yHat[0][10] ), .X(n45122) );
  inv_x2_sg U54838 ( .A(\reg_yHat[0][8] ), .X(n45124) );
  inv_x2_sg U54839 ( .A(\reg_yHat[0][17] ), .X(n45126) );
  inv_x2_sg U54840 ( .A(\reg_yHat[5][14] ), .X(n45128) );
  inv_x2_sg U54841 ( .A(\reg_yHat[13][14] ), .X(n45130) );
  inv_x2_sg U54842 ( .A(\reg_yHat[11][14] ), .X(n45132) );
  inv_x2_sg U54843 ( .A(\reg_yHat[9][14] ), .X(n45134) );
  inv_x2_sg U54844 ( .A(\reg_yHat[4][11] ), .X(n45136) );
  inv_x2_sg U54845 ( .A(\reg_yHat[8][11] ), .X(n45138) );
  inv_x2_sg U54846 ( .A(\reg_yHat[6][11] ), .X(n45140) );
  inv_x2_sg U54847 ( .A(\reg_yHat[3][11] ), .X(n45142) );
  inv_x2_sg U54848 ( .A(\reg_yHat[0][16] ), .X(n45144) );
  inv_x2_sg U54849 ( .A(\reg_yHat[1][13] ), .X(n45146) );
  inv_x2_sg U54850 ( .A(\reg_yHat[14][13] ), .X(n45148) );
  inv_x2_sg U54851 ( .A(\reg_yHat[12][13] ), .X(n45150) );
  inv_x2_sg U54852 ( .A(\reg_y[8][0] ), .X(n45564) );
  inv_x2_sg U54853 ( .A(\reg_y[6][0] ), .X(n45566) );
  inv_x2_sg U54854 ( .A(\reg_y[3][0] ), .X(n45568) );
  inv_x2_sg U54855 ( .A(\reg_y[1][0] ), .X(n45570) );
  inv_x2_sg U54856 ( .A(\reg_yHat[2][13] ), .X(n45152) );
  inv_x2_sg U54857 ( .A(\reg_yHat[8][3] ), .X(n44868) );
  inv_x2_sg U54858 ( .A(\reg_yHat[6][3] ), .X(n44870) );
  inv_x2_sg U54859 ( .A(\reg_yHat[3][3] ), .X(n44872) );
  inv_x2_sg U54860 ( .A(\reg_y[5][0] ), .X(n45572) );
  inv_x2_sg U54861 ( .A(\reg_y[12][0] ), .X(n45574) );
  inv_x2_sg U54862 ( .A(\reg_yHat[14][14] ), .X(n45154) );
  inv_x2_sg U54863 ( .A(\reg_yHat[12][14] ), .X(n45156) );
  inv_x2_sg U54864 ( .A(\reg_y[8][5] ), .X(n45994) );
  inv_x2_sg U54865 ( .A(\reg_y[6][5] ), .X(n45996) );
  inv_x2_sg U54866 ( .A(\reg_y[3][5] ), .X(n45998) );
  inv_x2_sg U54867 ( .A(\reg_yHat[1][9] ), .X(n45158) );
  inv_x2_sg U54868 ( .A(\reg_yHat[7][13] ), .X(n45160) );
  inv_x2_sg U54869 ( .A(\reg_yHat[4][13] ), .X(n45162) );
  inv_x2_sg U54870 ( .A(\reg_yHat[8][9] ), .X(n45164) );
  inv_x2_sg U54871 ( .A(\reg_yHat[6][9] ), .X(n45166) );
  inv_x2_sg U54872 ( .A(\reg_yHat[3][9] ), .X(n45168) );
  inv_x2_sg U54873 ( .A(\reg_yHat[4][9] ), .X(n45170) );
  inv_x2_sg U54874 ( .A(\reg_yHat[2][9] ), .X(n45172) );
  inv_x2_sg U54875 ( .A(\reg_y[14][0] ), .X(n45576) );
  inv_x2_sg U54876 ( .A(\reg_yHat[8][13] ), .X(n45174) );
  inv_x2_sg U54877 ( .A(\reg_yHat[6][13] ), .X(n45176) );
  inv_x2_sg U54878 ( .A(\reg_yHat[3][13] ), .X(n45178) );
  inv_x2_sg U54879 ( .A(\reg_y[0][0] ), .X(n45578) );
  inv_x2_sg U54880 ( .A(\reg_yHat[7][9] ), .X(n45180) );
  inv_x2_sg U54881 ( .A(\reg_yHat[13][1] ), .X(n46000) );
  inv_x2_sg U54882 ( .A(\reg_yHat[11][1] ), .X(n46002) );
  inv_x2_sg U54883 ( .A(\reg_yHat[9][1] ), .X(n46004) );
  inv_x2_sg U54884 ( .A(\reg_yHat[4][3] ), .X(n44876) );
  inv_x2_sg U54885 ( .A(\reg_yHat[8][1] ), .X(n46006) );
  inv_x2_sg U54886 ( .A(\reg_yHat[6][1] ), .X(n46008) );
  inv_x2_sg U54887 ( .A(\reg_yHat[3][1] ), .X(n46010) );
  inv_x2_sg U54888 ( .A(\reg_yHat[0][13] ), .X(n45182) );
  inv_x2_sg U54889 ( .A(\reg_yHat[5][12] ), .X(n45184) );
  inv_x2_sg U54890 ( .A(\reg_yHat[13][12] ), .X(n45186) );
  inv_x2_sg U54891 ( .A(\reg_yHat[11][12] ), .X(n45188) );
  inv_x2_sg U54892 ( .A(\reg_yHat[9][12] ), .X(n45190) );
  inv_x2_sg U54893 ( .A(\reg_yHat[11][4] ), .X(n44878) );
  inv_x2_sg U54894 ( .A(\reg_yHat[9][4] ), .X(n44880) );
  inv_x2_sg U54895 ( .A(\reg_yHat[13][4] ), .X(n44882) );
  inv_x2_sg U54896 ( .A(\reg_yHat[13][9] ), .X(n45192) );
  inv_x2_sg U54897 ( .A(\reg_yHat[11][9] ), .X(n45194) );
  inv_x2_sg U54898 ( .A(\reg_yHat[9][9] ), .X(n45196) );
  inv_x2_sg U54899 ( .A(\reg_yHat[5][9] ), .X(n45198) );
  inv_x2_sg U54900 ( .A(\reg_yHat[2][3] ), .X(n44884) );
  inv_x2_sg U54901 ( .A(\reg_yHat[10][9] ), .X(n45200) );
  inv_x2_sg U54902 ( .A(\reg_yHat[7][1] ), .X(n46012) );
  inv_x2_sg U54903 ( .A(\reg_yHat[7][3] ), .X(n44886) );
  inv_x2_sg U54904 ( .A(\reg_yHat[4][1] ), .X(n46014) );
  inv_x2_sg U54905 ( .A(\reg_yHat[11][3] ), .X(n44888) );
  inv_x2_sg U54906 ( .A(\reg_yHat[9][3] ), .X(n44890) );
  inv_x2_sg U54907 ( .A(\reg_yHat[13][3] ), .X(n44892) );
  inv_x2_sg U54908 ( .A(\reg_yHat[14][9] ), .X(n45202) );
  inv_x2_sg U54909 ( .A(\reg_yHat[12][9] ), .X(n45204) );
  inv_x2_sg U54910 ( .A(\reg_yHat[2][1] ), .X(n46016) );
  inv_x2_sg U54911 ( .A(\reg_yHat[1][1] ), .X(n46018) );
  inv_x2_sg U54912 ( .A(\reg_yHat[0][9] ), .X(n45206) );
  inv_x2_sg U54913 ( .A(\reg_yHat[12][3] ), .X(n44894) );
  inv_x2_sg U54914 ( .A(\reg_yHat[1][3] ), .X(n44896) );
  inv_x2_sg U54915 ( .A(\reg_yHat[12][1] ), .X(n46020) );
  inv_x2_sg U54916 ( .A(\reg_yHat[14][3] ), .X(n44898) );
  inv_x2_sg U54917 ( .A(\reg_yHat[5][1] ), .X(n46022) );
  inv_x2_sg U54918 ( .A(\reg_yHat[14][1] ), .X(n46024) );
  inv_x2_sg U54919 ( .A(\reg_yHat[0][1] ), .X(n46026) );
  inv_x2_sg U54920 ( .A(\reg_yHat[5][3] ), .X(n44900) );
  inv_x2_sg U54921 ( .A(\reg_yHat[0][3] ), .X(n44902) );
  inv_x2_sg U54922 ( .A(\reg_yHat[1][4] ), .X(n44904) );
  inv_x2_sg U54923 ( .A(\reg_yHat[1][7] ), .X(n44906) );
  inv_x2_sg U54924 ( .A(\reg_y[1][5] ), .X(n46030) );
  inv_x4_sg U54925 ( .A(n44107), .X(n44108) );
  nor_x2_sg U54926 ( .A(n18099), .B(n54120), .X(n18097) );
  inv_x4_sg U54927 ( .A(n18100), .X(n54120) );
  inv_x4_sg U54928 ( .A(n44109), .X(n44110) );
  nor_x2_sg U54929 ( .A(n16569), .B(n53671), .X(n16567) );
  inv_x4_sg U54930 ( .A(n16570), .X(n53671) );
  inv_x4_sg U54931 ( .A(n44111), .X(n44112) );
  nor_x2_sg U54932 ( .A(n16565), .B(n53651), .X(n16563) );
  inv_x4_sg U54933 ( .A(n16566), .X(n53651) );
  inv_x4_sg U54934 ( .A(n44113), .X(n44114) );
  nor_x2_sg U54935 ( .A(n15787), .B(n53392), .X(n15785) );
  inv_x4_sg U54936 ( .A(n15788), .X(n53392) );
  inv_x4_sg U54937 ( .A(n44115), .X(n44116) );
  nor_x2_sg U54938 ( .A(n15783), .B(n53373), .X(n15781) );
  inv_x4_sg U54939 ( .A(n15784), .X(n53373) );
  inv_x4_sg U54940 ( .A(n44117), .X(n44118) );
  nor_x2_sg U54941 ( .A(n15003), .B(n53113), .X(n15001) );
  inv_x4_sg U54942 ( .A(n15004), .X(n53113) );
  inv_x4_sg U54943 ( .A(n44119), .X(n44120) );
  nor_x2_sg U54944 ( .A(n14999), .B(n53093), .X(n14997) );
  inv_x4_sg U54945 ( .A(n15000), .X(n53093) );
  inv_x4_sg U54946 ( .A(n44121), .X(n44122) );
  nor_x2_sg U54947 ( .A(n13454), .B(n52554), .X(n13452) );
  inv_x4_sg U54948 ( .A(n13455), .X(n52554) );
  inv_x4_sg U54949 ( .A(n44123), .X(n44124) );
  nor_x2_sg U54950 ( .A(n13450), .B(n52535), .X(n13448) );
  inv_x4_sg U54951 ( .A(n13451), .X(n52535) );
  inv_x4_sg U54952 ( .A(n44125), .X(n44126) );
  nor_x2_sg U54953 ( .A(n12670), .B(n52279), .X(n12668) );
  inv_x4_sg U54954 ( .A(n12671), .X(n52279) );
  inv_x4_sg U54955 ( .A(n44127), .X(n44128) );
  nor_x2_sg U54956 ( .A(n12666), .B(n52259), .X(n12664) );
  inv_x4_sg U54957 ( .A(n12667), .X(n52259) );
  inv_x4_sg U54958 ( .A(n44129), .X(n44130) );
  nor_x2_sg U54959 ( .A(n11892), .B(n52003), .X(n11890) );
  inv_x4_sg U54960 ( .A(n11893), .X(n52003) );
  inv_x4_sg U54961 ( .A(n44131), .X(n44132) );
  nor_x2_sg U54962 ( .A(n11888), .B(n51984), .X(n11886) );
  inv_x4_sg U54963 ( .A(n11889), .X(n51984) );
  inv_x4_sg U54964 ( .A(n44133), .X(n44134) );
  nor_x2_sg U54965 ( .A(n11109), .B(n51725), .X(n11107) );
  inv_x4_sg U54966 ( .A(n11110), .X(n51725) );
  inv_x4_sg U54967 ( .A(n44135), .X(n44136) );
  nor_x2_sg U54968 ( .A(n11105), .B(n51703), .X(n11103) );
  inv_x4_sg U54969 ( .A(n11106), .X(n51703) );
  nor_x1_sg U54970 ( .A(n25178), .B(n25179), .X(n25176) );
  nor_x1_sg U54971 ( .A(n24503), .B(n24504), .X(n24500) );
  nor_x1_sg U54972 ( .A(n10070), .B(n10071), .X(n10068) );
  nor_x1_sg U54973 ( .A(n9389), .B(n9390), .X(n9386) );
  inv_x4_sg U54974 ( .A(n44137), .X(n44138) );
  nor_x2_sg U54975 ( .A(n21273), .B(n21272), .X(n21270) );
  inv_x4_sg U54976 ( .A(n44139), .X(n44140) );
  nor_x2_sg U54977 ( .A(n10401), .B(n10400), .X(n10398) );
  nor_x1_sg U54978 ( .A(n21776), .B(n46246), .X(n21775) );
  nor_x2_sg U54979 ( .A(n21773), .B(n55425), .X(n21776) );
  nor_x1_sg U54980 ( .A(n21005), .B(n20685), .X(n21004) );
  nor_x2_sg U54981 ( .A(n21003), .B(n55140), .X(n21005) );
  nor_x1_sg U54982 ( .A(n20231), .B(n46291), .X(n20230) );
  nor_x2_sg U54983 ( .A(n20228), .B(n54857), .X(n20231) );
  nor_x1_sg U54984 ( .A(n19461), .B(n19141), .X(n19460) );
  nor_x2_sg U54985 ( .A(n19459), .B(n54572), .X(n19461) );
  nor_x1_sg U54986 ( .A(n17916), .B(n17596), .X(n17915) );
  nor_x2_sg U54987 ( .A(n17914), .B(n54007), .X(n17916) );
  nor_x1_sg U54988 ( .A(n40878), .B(n46381), .X(n17140) );
  nor_x1_sg U54989 ( .A(n40876), .B(n46425), .X(n15574) );
  nor_x1_sg U54990 ( .A(n14795), .B(n46447), .X(n14794) );
  nor_x1_sg U54991 ( .A(n40874), .B(n46471), .X(n14021) );
  nor_x1_sg U54992 ( .A(n40872), .B(n46493), .X(n13241) );
  inv_x1_sg U54993 ( .A(n16665), .X(n53541) );
  nor_x2_sg U54994 ( .A(n16682), .B(n16681), .X(n16679) );
  nand_x4_sg U54995 ( .A(n16689), .B(n16690), .X(n16681) );
  inv_x1_sg U54996 ( .A(n15099), .X(n52983) );
  nor_x2_sg U54997 ( .A(n15116), .B(n15115), .X(n15113) );
  nand_x4_sg U54998 ( .A(n15123), .B(n15124), .X(n15115) );
  inv_x1_sg U54999 ( .A(n12766), .X(n52149) );
  nor_x2_sg U55000 ( .A(n12783), .B(n12782), .X(n12780) );
  nand_x4_sg U55001 ( .A(n12790), .B(n12791), .X(n12782) );
  inv_x1_sg U55002 ( .A(n11205), .X(n51591) );
  nor_x2_sg U55003 ( .A(n11222), .B(n11221), .X(n11219) );
  nand_x4_sg U55004 ( .A(n11229), .B(n11230), .X(n11221) );
  inv_x4_sg U55005 ( .A(n44141), .X(n44142) );
  nor_x2_sg U55006 ( .A(n53657), .B(n16992), .X(n16989) );
  inv_x4_sg U55007 ( .A(n44143), .X(n44144) );
  nor_x2_sg U55008 ( .A(n53099), .B(n15426), .X(n15423) );
  inv_x4_sg U55009 ( .A(n44145), .X(n44146) );
  nor_x2_sg U55010 ( .A(n52541), .B(n13873), .X(n13870) );
  inv_x4_sg U55011 ( .A(n44147), .X(n44148) );
  nor_x2_sg U55012 ( .A(n52265), .B(n13093), .X(n13090) );
  inv_x4_sg U55013 ( .A(n44149), .X(n44150) );
  nor_x2_sg U55014 ( .A(n51709), .B(n11532), .X(n11529) );
  inv_x4_sg U55015 ( .A(n44151), .X(n44152) );
  nor_x2_sg U55016 ( .A(n51900), .B(n51891), .X(n12128) );
  inv_x4_sg U55017 ( .A(n12130), .X(n51891) );
  nor_x2_sg U55018 ( .A(n51105), .B(n45301), .X(n27539) );
  inv_x4_sg U55019 ( .A(n46161), .X(n51105) );
  nor_x2_sg U55020 ( .A(n45300), .B(n46161), .X(n27540) );
  nor_x2_sg U55021 ( .A(n51009), .B(n45293), .X(n26144) );
  inv_x4_sg U55022 ( .A(n46153), .X(n51009) );
  nor_x2_sg U55023 ( .A(n45292), .B(n46153), .X(n26145) );
  nor_x2_sg U55024 ( .A(n51048), .B(n45273), .X(n26701) );
  inv_x4_sg U55025 ( .A(n46129), .X(n51048) );
  nor_x2_sg U55026 ( .A(n45272), .B(n46129), .X(n26702) );
  nor_x2_sg U55027 ( .A(n51237), .B(n45277), .X(n29496) );
  inv_x4_sg U55028 ( .A(n46135), .X(n51237) );
  nor_x2_sg U55029 ( .A(n45276), .B(n46135), .X(n29497) );
  nor_x2_sg U55030 ( .A(n51199), .B(n45279), .X(n28935) );
  inv_x4_sg U55031 ( .A(n46137), .X(n51199) );
  nor_x2_sg U55032 ( .A(n45278), .B(n46137), .X(n28936) );
  nor_x2_sg U55033 ( .A(n51067), .B(n45283), .X(n26980) );
  inv_x4_sg U55034 ( .A(n46141), .X(n51067) );
  nor_x2_sg U55035 ( .A(n45282), .B(n46141), .X(n26981) );
  nor_x2_sg U55036 ( .A(n50970), .B(n45275), .X(n25589) );
  inv_x4_sg U55037 ( .A(n46133), .X(n50970) );
  nor_x2_sg U55038 ( .A(n45274), .B(n46133), .X(n25590) );
  nor_x2_sg U55039 ( .A(n51008), .B(n45281), .X(n26150) );
  inv_x4_sg U55040 ( .A(n46139), .X(n51008) );
  nor_x2_sg U55041 ( .A(n45280), .B(n46139), .X(n26151) );
  nor_x2_sg U55042 ( .A(n51236), .B(n45287), .X(n29502) );
  inv_x4_sg U55043 ( .A(n46145), .X(n51236) );
  nor_x2_sg U55044 ( .A(n45286), .B(n46145), .X(n29503) );
  nor_x2_sg U55045 ( .A(n51198), .B(n45289), .X(n28941) );
  inv_x4_sg U55046 ( .A(n46147), .X(n51198) );
  nor_x2_sg U55047 ( .A(n45288), .B(n46147), .X(n28942) );
  nor_x2_sg U55048 ( .A(n51047), .B(n45291), .X(n26707) );
  inv_x4_sg U55049 ( .A(n46151), .X(n51047) );
  nor_x2_sg U55050 ( .A(n45290), .B(n46151), .X(n26708) );
  nor_x2_sg U55051 ( .A(n50971), .B(n45327), .X(n25583) );
  inv_x4_sg U55052 ( .A(n46187), .X(n50971) );
  nor_x2_sg U55053 ( .A(n45326), .B(n46187), .X(n25584) );
  nand_x4_sg U55054 ( .A(n9406), .B(n46200), .X(n29607) );
  inv_x4_sg U55055 ( .A(n18826), .X(n54142) );
  nor_x2_sg U55056 ( .A(n44457), .B(n20551), .X(n20548) );
  nor_x2_sg U55057 ( .A(n44459), .B(n19007), .X(n19004) );
  nor_x2_sg U55058 ( .A(n44461), .B(n17462), .X(n17459) );
  nand_x4_sg U55059 ( .A(n44034), .B(n20982), .X(n20980) );
  nand_x4_sg U55060 ( .A(n44036), .B(n19438), .X(n19436) );
  nand_x4_sg U55061 ( .A(n44038), .B(n17893), .X(n17891) );
  inv_x4_sg U55062 ( .A(n44157), .X(n44158) );
  inv_x4_sg U55063 ( .A(n44159), .X(n44160) );
  inv_x4_sg U55064 ( .A(n44161), .X(n44162) );
  inv_x4_sg U55065 ( .A(n44163), .X(n44164) );
  inv_x4_sg U55066 ( .A(n44165), .X(n44166) );
  inv_x4_sg U55067 ( .A(n44167), .X(n44168) );
  inv_x4_sg U55068 ( .A(n55783), .X(n44169) );
  inv_x4_sg U55069 ( .A(n44170), .X(n44171) );
  inv_x4_sg U55070 ( .A(n44172), .X(n44173) );
  nor_x2_sg U55071 ( .A(n55512), .B(n46584), .X(n15724) );
  inv_x4_sg U55072 ( .A(n44174), .X(n44175) );
  inv_x4_sg U55073 ( .A(n13391), .X(n55787) );
  nor_x2_sg U55074 ( .A(n21299), .B(n21300), .X(n21298) );
  nor_x4_sg U55075 ( .A(n55191), .B(n21296), .X(n21300) );
  inv_x4_sg U55076 ( .A(n21297), .X(n55191) );
  nor_x2_sg U55077 ( .A(n19754), .B(n19755), .X(n19753) );
  nor_x4_sg U55078 ( .A(n54623), .B(n19751), .X(n19755) );
  inv_x4_sg U55079 ( .A(n19752), .X(n54623) );
  inv_x4_sg U55080 ( .A(n44176), .X(n44177) );
  inv_x4_sg U55081 ( .A(n44178), .X(n44179) );
  inv_x4_sg U55082 ( .A(n44180), .X(n44181) );
  inv_x4_sg U55083 ( .A(n44182), .X(n44183) );
  inv_x4_sg U55084 ( .A(n44184), .X(n44185) );
  inv_x4_sg U55085 ( .A(n44186), .X(n44187) );
  inv_x4_sg U55086 ( .A(n44188), .X(n44189) );
  inv_x4_sg U55087 ( .A(n44190), .X(n44191) );
  inv_x4_sg U55088 ( .A(n44192), .X(n44193) );
  nand_x4_sg U55089 ( .A(n41344), .B(n41174), .X(n13413) );
  inv_x4_sg U55090 ( .A(n44194), .X(n44195) );
  inv_x4_sg U55091 ( .A(n44196), .X(n44197) );
  inv_x4_sg U55092 ( .A(n44198), .X(n44199) );
  inv_x4_sg U55093 ( .A(n14327), .X(n52685) );
  inv_x4_sg U55094 ( .A(n44200), .X(n44201) );
  inv_x4_sg U55095 ( .A(n44202), .X(n44203) );
  inv_x4_sg U55096 ( .A(n44204), .X(n44205) );
  inv_x4_sg U55097 ( .A(n44206), .X(n44207) );
  inv_x4_sg U55098 ( .A(n44208), .X(n44209) );
  inv_x4_sg U55099 ( .A(n44210), .X(n44211) );
  inv_x4_sg U55100 ( .A(n44212), .X(n44213) );
  inv_x4_sg U55101 ( .A(n44214), .X(n44215) );
  inv_x4_sg U55102 ( .A(n18637), .X(n54240) );
  inv_x4_sg U55103 ( .A(n46195), .X(n55459) );
  inv_x4_sg U55104 ( .A(n44216), .X(n44217) );
  inv_x4_sg U55105 ( .A(n44218), .X(n44219) );
  inv_x4_sg U55106 ( .A(n44220), .X(n44221) );
  inv_x4_sg U55107 ( .A(n44222), .X(n44223) );
  inv_x4_sg U55108 ( .A(n44224), .X(n44225) );
  inv_x4_sg U55109 ( .A(n44226), .X(n44227) );
  inv_x4_sg U55110 ( .A(n44228), .X(n44229) );
  inv_x4_sg U55111 ( .A(n44230), .X(n44231) );
  inv_x4_sg U55112 ( .A(n44232), .X(n44233) );
  inv_x4_sg U55113 ( .A(n44234), .X(n44235) );
  inv_x4_sg U55114 ( .A(n44236), .X(n44237) );
  inv_x4_sg U55115 ( .A(n44238), .X(n44239) );
  inv_x4_sg U55116 ( .A(n44240), .X(n44241) );
  inv_x4_sg U55117 ( .A(n44242), .X(n44243) );
  inv_x4_sg U55118 ( .A(n44244), .X(n44245) );
  inv_x4_sg U55119 ( .A(n44246), .X(n44247) );
  nor_x4_sg U55120 ( .A(n13735), .B(n46477), .X(n13824) );
  nor_x4_sg U55121 ( .A(n11394), .B(n46543), .X(n11483) );
  nor_x4_sg U55122 ( .A(n16897), .B(n16898), .X(n16883) );
  nand_x4_sg U55123 ( .A(n46395), .B(n16842), .X(n16897) );
  nor_x4_sg U55124 ( .A(n15331), .B(n15332), .X(n15317) );
  nand_x4_sg U55125 ( .A(n46439), .B(n15276), .X(n15331) );
  nor_x4_sg U55126 ( .A(n12998), .B(n12999), .X(n12984) );
  nand_x4_sg U55127 ( .A(n46507), .B(n12943), .X(n12998) );
  nor_x4_sg U55128 ( .A(n11437), .B(n11438), .X(n11423) );
  nand_x4_sg U55129 ( .A(n46551), .B(n11382), .X(n11437) );
  nor_x4_sg U55130 ( .A(n20717), .B(n46272), .X(n20804) );
  nor_x4_sg U55131 ( .A(n19173), .B(n46317), .X(n19260) );
  nor_x4_sg U55132 ( .A(n17628), .B(n46364), .X(n17715) );
  nor_x4_sg U55133 ( .A(n14507), .B(n46454), .X(n14594) );
  inv_x4_sg U55134 ( .A(n44248), .X(n44249) );
  nor_x2_sg U55135 ( .A(n50984), .B(n45241), .X(n25664) );
  inv_x4_sg U55136 ( .A(n46087), .X(n50984) );
  nor_x2_sg U55137 ( .A(n45240), .B(n46087), .X(n25665) );
  nor_x4_sg U55138 ( .A(n13726), .B(n52477), .X(n13719) );
  inv_x4_sg U55139 ( .A(n13727), .X(n52477) );
  inv_x4_sg U55140 ( .A(n44250), .X(n44251) );
  nor_x2_sg U55141 ( .A(n51215), .B(n45295), .X(n29236) );
  inv_x4_sg U55142 ( .A(n46155), .X(n51215) );
  nor_x2_sg U55143 ( .A(n45294), .B(n46155), .X(n29237) );
  inv_x4_sg U55144 ( .A(n44252), .X(n44253) );
  nor_x2_sg U55145 ( .A(n51177), .B(n45297), .X(n28675) );
  inv_x4_sg U55146 ( .A(n46157), .X(n51177) );
  nor_x2_sg U55147 ( .A(n45296), .B(n46157), .X(n28676) );
  inv_x4_sg U55148 ( .A(n44254), .X(n44255) );
  nor_x2_sg U55149 ( .A(n51140), .B(n45299), .X(n28117) );
  inv_x4_sg U55150 ( .A(n46159), .X(n51140) );
  nor_x2_sg U55151 ( .A(n45298), .B(n46159), .X(n28118) );
  inv_x4_sg U55152 ( .A(n44256), .X(n44257) );
  nor_x2_sg U55153 ( .A(n50968), .B(n45303), .X(n25601) );
  inv_x4_sg U55154 ( .A(n46163), .X(n50968) );
  nor_x2_sg U55155 ( .A(n45302), .B(n46163), .X(n25602) );
  inv_x4_sg U55156 ( .A(n44258), .X(n44259) );
  nor_x2_sg U55157 ( .A(n50987), .B(n45305), .X(n25882) );
  inv_x4_sg U55158 ( .A(n46165), .X(n50987) );
  nor_x2_sg U55159 ( .A(n45304), .B(n46165), .X(n25883) );
  inv_x4_sg U55160 ( .A(n44260), .X(n44261) );
  nor_x2_sg U55161 ( .A(n51102), .B(n45307), .X(n27557) );
  inv_x4_sg U55162 ( .A(n46167), .X(n51102) );
  nor_x2_sg U55163 ( .A(n45306), .B(n46167), .X(n27558) );
  inv_x4_sg U55164 ( .A(n44262), .X(n44263) );
  nor_x2_sg U55165 ( .A(n51196), .B(n45311), .X(n28953) );
  inv_x4_sg U55166 ( .A(n46171), .X(n51196) );
  nor_x2_sg U55167 ( .A(n45310), .B(n46171), .X(n28954) );
  inv_x4_sg U55168 ( .A(n44264), .X(n44265) );
  nor_x2_sg U55169 ( .A(n51064), .B(n45313), .X(n26998) );
  inv_x4_sg U55170 ( .A(n46173), .X(n51064) );
  nor_x2_sg U55171 ( .A(n45312), .B(n46173), .X(n26999) );
  inv_x4_sg U55172 ( .A(n44266), .X(n44267) );
  nor_x2_sg U55173 ( .A(n51234), .B(n45315), .X(n29514) );
  inv_x4_sg U55174 ( .A(n46175), .X(n51234) );
  nor_x2_sg U55175 ( .A(n45314), .B(n46175), .X(n29515) );
  inv_x4_sg U55176 ( .A(n44268), .X(n44269) );
  nor_x2_sg U55177 ( .A(n51045), .B(n45317), .X(n26719) );
  inv_x4_sg U55178 ( .A(n46177), .X(n51045) );
  nor_x2_sg U55179 ( .A(n45316), .B(n46177), .X(n26720) );
  inv_x4_sg U55180 ( .A(n44270), .X(n44271) );
  nor_x2_sg U55181 ( .A(n51121), .B(n45319), .X(n27836) );
  inv_x4_sg U55182 ( .A(n46179), .X(n51121) );
  nor_x2_sg U55183 ( .A(n45318), .B(n46179), .X(n27837) );
  inv_x4_sg U55184 ( .A(n44272), .X(n44273) );
  nor_x2_sg U55185 ( .A(n51083), .B(n45321), .X(n27278) );
  inv_x4_sg U55186 ( .A(n46181), .X(n51083) );
  nor_x2_sg U55187 ( .A(n45320), .B(n46181), .X(n27279) );
  inv_x4_sg U55188 ( .A(n44274), .X(n44275) );
  nor_x2_sg U55189 ( .A(n51025), .B(n45323), .X(n26441) );
  inv_x4_sg U55190 ( .A(n46183), .X(n51025) );
  nor_x2_sg U55191 ( .A(n45322), .B(n46183), .X(n26442) );
  inv_x4_sg U55192 ( .A(n44276), .X(n44277) );
  nor_x2_sg U55193 ( .A(n51006), .B(n45325), .X(n26162) );
  inv_x4_sg U55194 ( .A(n46185), .X(n51006) );
  nor_x2_sg U55195 ( .A(n45324), .B(n46185), .X(n26163) );
  nor_x2_sg U55196 ( .A(n54053), .B(n46193), .X(n28391) );
  inv_x4_sg U55197 ( .A(n45209), .X(n54053) );
  inv_x4_sg U55198 ( .A(n15739), .X(n53209) );
  inv_x4_sg U55199 ( .A(n11844), .X(n51821) );
  inv_x4_sg U55200 ( .A(n13406), .X(n52373) );
  inv_x4_sg U55201 ( .A(n19621), .X(n54616) );
  inv_x4_sg U55202 ( .A(n18076), .X(n54051) );
  nand_x4_sg U55203 ( .A(n54050), .B(n54045), .X(n18076) );
  inv_x4_sg U55204 ( .A(n44278), .X(n44279) );
  inv_x4_sg U55205 ( .A(n44280), .X(n44281) );
  inv_x4_sg U55206 ( .A(n44282), .X(n44283) );
  inv_x4_sg U55207 ( .A(n21166), .X(n55184) );
  inv_x4_sg U55208 ( .A(n14185), .X(n52650) );
  nand_x4_sg U55209 ( .A(n52649), .B(n52644), .X(n14185) );
  inv_x4_sg U55210 ( .A(n16746), .X(n53561) );
  inv_x4_sg U55211 ( .A(n15961), .X(n53279) );
  inv_x4_sg U55212 ( .A(n15180), .X(n53003) );
  inv_x4_sg U55213 ( .A(n12847), .X(n52169) );
  inv_x4_sg U55214 ( .A(n12066), .X(n51892) );
  inv_x4_sg U55215 ( .A(n11286), .X(n51611) );
  inv_x4_sg U55216 ( .A(n44284), .X(n44285) );
  nor_x2_sg U55217 ( .A(n51043), .B(n45947), .X(n26721) );
  inv_x4_sg U55218 ( .A(n45581), .X(n51043) );
  inv_x8_sg U55219 ( .A(n45948), .X(n45949) );
  inv_x8_sg U55220 ( .A(n45950), .X(n45951) );
  inv_x8_sg U55221 ( .A(n45952), .X(n45953) );
  inv_x8_sg U55222 ( .A(n45954), .X(n45955) );
  inv_x8_sg U55223 ( .A(n45956), .X(n45957) );
  inv_x8_sg U55224 ( .A(n45958), .X(n45959) );
  inv_x8_sg U55225 ( .A(n45960), .X(n45961) );
  inv_x8_sg U55226 ( .A(n45962), .X(n45963) );
  inv_x8_sg U55227 ( .A(n45964), .X(n45965) );
  inv_x8_sg U55228 ( .A(n45966), .X(n45967) );
  inv_x8_sg U55229 ( .A(n45968), .X(n45969) );
  inv_x8_sg U55230 ( .A(n45970), .X(n45971) );
  inv_x8_sg U55231 ( .A(n45972), .X(n45973) );
  inv_x8_sg U55232 ( .A(n45974), .X(n45975) );
  inv_x4_sg U55233 ( .A(n31737), .X(n49284) );
  inv_x4_sg U55234 ( .A(n30590), .X(n49290) );
  inv_x4_sg U55235 ( .A(n22924), .X(n50149) );
  inv_x4_sg U55236 ( .A(n24071), .X(n50143) );
  inv_x4_sg U55237 ( .A(n29721), .X(n49294) );
  inv_x4_sg U55238 ( .A(n22056), .X(n50153) );
  nand_x8_sg U55239 ( .A(n28257), .B(n18574), .X(n28264) );
  nor_x8_sg U55240 ( .A(n28249), .B(n54165), .X(n28257) );
  nand_x8_sg U55241 ( .A(n29390), .B(n21714), .X(n29397) );
  nand_x8_sg U55242 ( .A(n29108), .B(n20945), .X(n29115) );
  nand_x8_sg U55243 ( .A(n28829), .B(n20169), .X(n28836) );
  nand_x8_sg U55244 ( .A(n28549), .B(n19401), .X(n28556) );
  nand_x8_sg U55245 ( .A(n27991), .B(n17856), .X(n27998) );
  nand_x8_sg U55246 ( .A(n26872), .B(n14735), .X(n26879) );
  inv_x4_sg U55247 ( .A(n44286), .X(n44287) );
  nor_x4_sg U55248 ( .A(n44287), .B(n50729), .X(n23537) );
  inv_x4_sg U55249 ( .A(n23724), .X(n50729) );
  inv_x4_sg U55250 ( .A(n44288), .X(n44289) );
  nor_x4_sg U55251 ( .A(n44289), .B(n50794), .X(n23106) );
  inv_x4_sg U55252 ( .A(n23329), .X(n50794) );
  inv_x4_sg U55253 ( .A(n44290), .X(n44291) );
  nor_x4_sg U55254 ( .A(n44291), .B(n49870), .X(n31203) );
  inv_x4_sg U55255 ( .A(n31390), .X(n49870) );
  inv_x4_sg U55256 ( .A(n44292), .X(n44293) );
  nor_x4_sg U55257 ( .A(n44293), .B(n49935), .X(n30772) );
  inv_x4_sg U55258 ( .A(n30995), .X(n49935) );
  inv_x4_sg U55259 ( .A(n44294), .X(n44295) );
  inv_x4_sg U55260 ( .A(n44296), .X(n44297) );
  nor_x4_sg U55261 ( .A(n44297), .B(n44295), .X(n32107) );
  inv_x4_sg U55262 ( .A(n44298), .X(n44299) );
  inv_x4_sg U55263 ( .A(n44300), .X(n44301) );
  nor_x4_sg U55264 ( .A(n44301), .B(n44299), .X(n24441) );
  inv_x4_sg U55265 ( .A(n18681), .X(n54289) );
  nor_x4_sg U55266 ( .A(n18705), .B(n46341), .X(n18681) );
  inv_x4_sg U55267 ( .A(n11679), .X(n51777) );
  nor_x4_sg U55268 ( .A(n11703), .B(n46546), .X(n11679) );
  inv_x4_sg U55269 ( .A(n21419), .X(n55237) );
  nand_x2_sg U55270 ( .A(n21420), .B(n21290), .X(n21419) );
  inv_x4_sg U55271 ( .A(n19874), .X(n54669) );
  nand_x2_sg U55272 ( .A(n19875), .B(n19745), .X(n19874) );
  nor_x4_sg U55273 ( .A(n14440), .B(n46445), .X(n14400) );
  nand_x4_sg U55274 ( .A(n46458), .B(n14310), .X(n14440) );
  inv_x4_sg U55275 ( .A(n20648), .X(n54948) );
  nand_x2_sg U55276 ( .A(n20649), .B(n20520), .X(n20648) );
  inv_x4_sg U55277 ( .A(n19104), .X(n54380) );
  nand_x2_sg U55278 ( .A(n19105), .B(n18976), .X(n19104) );
  inv_x4_sg U55279 ( .A(n17559), .X(n53815) );
  nand_x2_sg U55280 ( .A(n17560), .B(n17431), .X(n17559) );
  nor_x4_sg U55281 ( .A(n21025), .B(n46281), .X(n21106) );
  nor_x4_sg U55282 ( .A(n19481), .B(n46326), .X(n19562) );
  nor_x4_sg U55283 ( .A(n17936), .B(n46373), .X(n18017) );
  nor_x4_sg U55284 ( .A(n14815), .B(n46463), .X(n14896) );
  nor_x4_sg U55285 ( .A(n46250), .B(n46242), .X(n21536) );
  nor_x4_sg U55286 ( .A(n46295), .B(n46287), .X(n19991) );
  nor_x4_sg U55287 ( .A(n46559), .B(n46565), .X(n10664) );
  nor_x4_sg U55288 ( .A(n46331), .B(n46337), .X(n18571) );
  nor_x4_sg U55289 ( .A(n46559), .B(n46563), .X(n10792) );
  nor_x4_sg U55290 ( .A(n21418), .B(n21417), .X(n21441) );
  nor_x4_sg U55291 ( .A(n20646), .B(n20647), .X(n20670) );
  nor_x4_sg U55292 ( .A(n19873), .B(n19872), .X(n19896) );
  nor_x4_sg U55293 ( .A(n19102), .B(n19103), .X(n19126) );
  nor_x4_sg U55294 ( .A(n18329), .B(n18327), .X(n18351) );
  nor_x4_sg U55295 ( .A(n17557), .B(n17558), .X(n17581) );
  nor_x4_sg U55296 ( .A(n14438), .B(n14439), .X(n14461) );
  nor_x4_sg U55297 ( .A(n46467), .B(n46475), .X(n13783) );
  nor_x4_sg U55298 ( .A(n15925), .B(n16069), .X(n16457) );
  nor_x4_sg U55299 ( .A(n46377), .B(n46387), .X(n16851) );
  nor_x4_sg U55300 ( .A(n46421), .B(n46431), .X(n15285) );
  nor_x4_sg U55301 ( .A(n46489), .B(n46499), .X(n12952) );
  nor_x4_sg U55302 ( .A(n46533), .B(n46543), .X(n11391) );
  nor_x4_sg U55303 ( .A(n12174), .B(n12030), .X(n12554) );
  nor_x4_sg U55304 ( .A(n46521), .B(n46514), .X(n12171) );
  nor_x2_sg U55305 ( .A(n21423), .B(n21424), .X(n21421) );
  nor_x4_sg U55306 ( .A(n46242), .B(n46254), .X(n21424) );
  nor_x2_sg U55307 ( .A(n19878), .B(n19879), .X(n19876) );
  nor_x4_sg U55308 ( .A(n46287), .B(n46299), .X(n19879) );
  nor_x4_sg U55309 ( .A(n54097), .B(n46344), .X(n18395) );
  nor_x4_sg U55310 ( .A(n46561), .B(n46568), .X(n10613) );
  nor_x4_sg U55311 ( .A(n13980), .B(n46477), .X(n14111) );
  inv_x4_sg U55312 ( .A(n44302), .X(n44303) );
  nor_x4_sg U55313 ( .A(n49872), .B(n44303), .X(n30731) );
  inv_x4_sg U55314 ( .A(n30957), .X(n49872) );
  inv_x4_sg U55315 ( .A(n44304), .X(n44305) );
  nor_x4_sg U55316 ( .A(n50731), .B(n44305), .X(n23065) );
  inv_x4_sg U55317 ( .A(n23291), .X(n50731) );
  nor_x4_sg U55318 ( .A(n46297), .B(n46300), .X(n19729) );
  nand_x4_sg U55319 ( .A(n21274), .B(n42627), .X(n21273) );
  nor_x4_sg U55320 ( .A(n46252), .B(n46255), .X(n21274) );
  nand_x4_sg U55321 ( .A(n51261), .B(n10402), .X(n10389) );
  nand_x4_sg U55322 ( .A(n10402), .B(n10389), .X(n10401) );
  nor_x4_sg U55323 ( .A(n46568), .B(n46566), .X(n10402) );
  inv_x2_sg U55324 ( .A(n17072), .X(n53638) );
  nor_x4_sg U55325 ( .A(n16975), .B(n46387), .X(n17072) );
  inv_x2_sg U55326 ( .A(n15506), .X(n53080) );
  nor_x4_sg U55327 ( .A(n15409), .B(n46431), .X(n15506) );
  inv_x2_sg U55328 ( .A(n13173), .X(n52246) );
  nor_x4_sg U55329 ( .A(n13076), .B(n46499), .X(n13173) );
  inv_x2_sg U55330 ( .A(n12393), .X(n51971) );
  nor_x4_sg U55331 ( .A(n12295), .B(n46521), .X(n12393) );
  nor_x4_sg U55332 ( .A(n29575), .B(n29576), .X(n21787) );
  nor_x4_sg U55333 ( .A(n51250), .B(n45243), .X(n29575) );
  inv_x4_sg U55334 ( .A(n46089), .X(n51250) );
  nor_x4_sg U55335 ( .A(n55443), .B(n46089), .X(n29576) );
  inv_x4_sg U55336 ( .A(n45243), .X(n55443) );
  nor_x4_sg U55337 ( .A(n29297), .B(n29298), .X(n21016) );
  nor_x4_sg U55338 ( .A(n51231), .B(n45251), .X(n29297) );
  inv_x4_sg U55339 ( .A(n46097), .X(n51231) );
  nor_x4_sg U55340 ( .A(n55159), .B(n46097), .X(n29298) );
  inv_x4_sg U55341 ( .A(n45251), .X(n55159) );
  nor_x4_sg U55342 ( .A(n29014), .B(n29015), .X(n20242) );
  nor_x4_sg U55343 ( .A(n51212), .B(n45245), .X(n29014) );
  inv_x4_sg U55344 ( .A(n46091), .X(n51212) );
  nor_x4_sg U55345 ( .A(n54875), .B(n46091), .X(n29015) );
  inv_x4_sg U55346 ( .A(n45245), .X(n54875) );
  nor_x4_sg U55347 ( .A(n28736), .B(n28737), .X(n19472) );
  nor_x4_sg U55348 ( .A(n51193), .B(n45253), .X(n28736) );
  inv_x4_sg U55349 ( .A(n46099), .X(n51193) );
  nor_x4_sg U55350 ( .A(n54591), .B(n46099), .X(n28737) );
  inv_x4_sg U55351 ( .A(n45253), .X(n54591) );
  nor_x4_sg U55352 ( .A(n28457), .B(n28458), .X(n18696) );
  nor_x4_sg U55353 ( .A(n51174), .B(n45247), .X(n28457) );
  inv_x4_sg U55354 ( .A(n46093), .X(n51174) );
  nor_x4_sg U55355 ( .A(n54307), .B(n46093), .X(n28458) );
  inv_x4_sg U55356 ( .A(n45247), .X(n54307) );
  nor_x4_sg U55357 ( .A(n28178), .B(n28179), .X(n17927) );
  nor_x4_sg U55358 ( .A(n51156), .B(n45255), .X(n28178) );
  inv_x4_sg U55359 ( .A(n46101), .X(n51156) );
  nor_x4_sg U55360 ( .A(n54026), .B(n46101), .X(n28179) );
  inv_x4_sg U55361 ( .A(n45255), .X(n54026) );
  nor_x4_sg U55362 ( .A(n27897), .B(n27898), .X(n17153) );
  nor_x4_sg U55363 ( .A(n51137), .B(n45265), .X(n27897) );
  inv_x4_sg U55364 ( .A(n46111), .X(n51137) );
  nor_x4_sg U55365 ( .A(n53742), .B(n46111), .X(n27898) );
  inv_x4_sg U55366 ( .A(n45265), .X(n53742) );
  nor_x4_sg U55367 ( .A(n27339), .B(n27340), .X(n15587) );
  nor_x4_sg U55368 ( .A(n51099), .B(n45267), .X(n27339) );
  inv_x4_sg U55369 ( .A(n46113), .X(n51099) );
  nor_x4_sg U55370 ( .A(n53184), .B(n46113), .X(n27340) );
  inv_x4_sg U55371 ( .A(n45267), .X(n53184) );
  nor_x4_sg U55372 ( .A(n27059), .B(n27060), .X(n14806) );
  nor_x4_sg U55373 ( .A(n51080), .B(n45249), .X(n27059) );
  inv_x4_sg U55374 ( .A(n46095), .X(n51080) );
  nor_x4_sg U55375 ( .A(n52906), .B(n46095), .X(n27060) );
  inv_x4_sg U55376 ( .A(n45249), .X(n52906) );
  nor_x4_sg U55377 ( .A(n26780), .B(n26781), .X(n14034) );
  nor_x4_sg U55378 ( .A(n51061), .B(n45261), .X(n26780) );
  inv_x4_sg U55379 ( .A(n46107), .X(n51061) );
  nor_x4_sg U55380 ( .A(n52625), .B(n46107), .X(n26781) );
  inv_x4_sg U55381 ( .A(n45261), .X(n52625) );
  nor_x4_sg U55382 ( .A(n26502), .B(n26503), .X(n13254) );
  nor_x4_sg U55383 ( .A(n51041), .B(n45269), .X(n26502) );
  inv_x4_sg U55384 ( .A(n46115), .X(n51041) );
  nor_x4_sg U55385 ( .A(n52350), .B(n46115), .X(n26503) );
  inv_x4_sg U55386 ( .A(n45269), .X(n52350) );
  nor_x4_sg U55387 ( .A(n26223), .B(n26224), .X(n12473) );
  nor_x4_sg U55388 ( .A(n51022), .B(n45263), .X(n26223) );
  inv_x4_sg U55389 ( .A(n46109), .X(n51022) );
  nor_x4_sg U55390 ( .A(n52072), .B(n46109), .X(n26224) );
  inv_x4_sg U55391 ( .A(n45263), .X(n52072) );
  nor_x4_sg U55392 ( .A(n25943), .B(n25944), .X(n11694) );
  nor_x4_sg U55393 ( .A(n51003), .B(n45259), .X(n25943) );
  inv_x4_sg U55394 ( .A(n46105), .X(n51003) );
  nor_x4_sg U55395 ( .A(n51796), .B(n46105), .X(n25944) );
  inv_x4_sg U55396 ( .A(n45259), .X(n51796) );
  nor_x4_sg U55397 ( .A(n27618), .B(n27619), .X(n16368) );
  nor_x4_sg U55398 ( .A(n51118), .B(n45257), .X(n27618) );
  inv_x4_sg U55399 ( .A(n46103), .X(n51118) );
  nor_x4_sg U55400 ( .A(n53464), .B(n46103), .X(n27619) );
  inv_x4_sg U55401 ( .A(n45257), .X(n53464) );
  nor_x4_sg U55402 ( .A(n39302), .B(n55797), .X(n39296) );
  nand_x4_sg U55403 ( .A(n55796), .B(done), .X(n39302) );
  inv_x4_sg U55404 ( .A(state[0]), .X(n55797) );
  inv_x4_sg U55405 ( .A(n44306), .X(n44307) );
  nor_x4_sg U55406 ( .A(n10543), .B(n44307), .X(n10508) );
  nor_x4_sg U55407 ( .A(n10546), .B(n51321), .X(n10543) );
  nor_x4_sg U55408 ( .A(n25471), .B(n51418), .X(n25478) );
  inv_x8_sg U55409 ( .A(n10782), .X(n51418) );
  inv_x4_sg U55410 ( .A(n44308), .X(n44309) );
  inv_x4_sg U55411 ( .A(n44309), .X(n51125) );
  inv_x4_sg U55412 ( .A(n44310), .X(n44311) );
  inv_x4_sg U55413 ( .A(n44311), .X(n51087) );
  inv_x4_sg U55414 ( .A(n44312), .X(n44313) );
  inv_x4_sg U55415 ( .A(n44313), .X(n51029) );
  inv_x4_sg U55416 ( .A(n44314), .X(n44315) );
  inv_x4_sg U55417 ( .A(n44315), .X(n51126) );
  inv_x4_sg U55418 ( .A(n44316), .X(n44317) );
  inv_x4_sg U55419 ( .A(n44317), .X(n51088) );
  inv_x4_sg U55420 ( .A(n44318), .X(n44319) );
  inv_x4_sg U55421 ( .A(n44319), .X(n51030) );
  nor_x4_sg U55422 ( .A(n13662), .B(n46469), .X(n13625) );
  nand_x4_sg U55423 ( .A(n46481), .B(n13530), .X(n13662) );
  inv_x4_sg U55424 ( .A(n26966), .X(n44320) );
  inv_x2_sg U55425 ( .A(n44322), .X(n44323) );
  nor_x2_sg U55426 ( .A(n52668), .B(n46149), .X(n27041) );
  nor_x2_sg U55427 ( .A(n46200), .B(n55457), .X(n29603) );
  nor_x2_sg U55428 ( .A(n55457), .B(n55458), .X(n30163) );
  nor_x2_sg U55429 ( .A(n46584), .B(n55457), .X(n29595) );
  inv_x8_sg U55430 ( .A(n46582), .X(n55457) );
  inv_x8_sg U55431 ( .A(n29617), .X(n55462) );
  nand_x8_sg U55432 ( .A(n29151), .B(n29620), .X(n29617) );
  nor_x2_sg U55433 ( .A(n54144), .B(n18579), .X(n18578) );
  nand_x4_sg U55434 ( .A(n54124), .B(n54070), .X(n18579) );
  nor_x2_sg U55435 ( .A(n51355), .B(n10799), .X(n10798) );
  inv_x4_sg U55436 ( .A(n10803), .X(n51355) );
  nor_x2_sg U55437 ( .A(n46232), .B(n46569), .X(n25402) );
  nand_x4_sg U55438 ( .A(n55215), .B(n46260), .X(n21306) );
  nand_x4_sg U55439 ( .A(n54647), .B(n46305), .X(n19761) );
  nand_x4_sg U55440 ( .A(n52683), .B(n46462), .X(n14326) );
  nor_x2_sg U55441 ( .A(n10433), .B(n10434), .X(n10432) );
  nor_x4_sg U55442 ( .A(n43261), .B(n43259), .X(n10433) );
  nand_x4_sg U55443 ( .A(n51293), .B(n46574), .X(n10434) );
  inv_x1_sg U55444 ( .A(n31257), .X(n49310) );
  nand_x2_sg U55445 ( .A(n49329), .B(n31257), .X(n31256) );
  inv_x1_sg U55446 ( .A(n23591), .X(n50169) );
  nand_x2_sg U55447 ( .A(n50188), .B(n23591), .X(n23590) );
  inv_x4_sg U55448 ( .A(n11742), .X(n51733) );
  nor_x4_sg U55449 ( .A(n11623), .B(n46543), .X(n11742) );
  inv_x4_sg U55450 ( .A(n16982), .X(n53631) );
  nor_x4_sg U55451 ( .A(n16975), .B(n46390), .X(n16982) );
  inv_x4_sg U55452 ( .A(n15416), .X(n53073) );
  nor_x4_sg U55453 ( .A(n15409), .B(n46434), .X(n15416) );
  inv_x4_sg U55454 ( .A(n13083), .X(n52239) );
  nor_x4_sg U55455 ( .A(n13076), .B(n46502), .X(n13083) );
  inv_x4_sg U55456 ( .A(n44324), .X(n44325) );
  inv_x4_sg U55457 ( .A(n44326), .X(n44327) );
  nand_x4_sg U55458 ( .A(n55210), .B(n21615), .X(n21610) );
  nor_x4_sg U55459 ( .A(n21532), .B(n46244), .X(n21615) );
  nand_x4_sg U55460 ( .A(n54642), .B(n20070), .X(n20065) );
  nor_x4_sg U55461 ( .A(n19987), .B(n46289), .X(n20070) );
  nand_x4_sg U55462 ( .A(n51288), .B(n10744), .X(n10739) );
  nor_x4_sg U55463 ( .A(n46561), .B(n10660), .X(n10744) );
  inv_x1_sg U55464 ( .A(n16254), .X(n53397) );
  inv_x1_sg U55465 ( .A(n11615), .X(n51746) );
  nor_x1_sg U55466 ( .A(n46611), .B(n12609), .X(n26076) );
  inv_x4_sg U55467 ( .A(n44328), .X(n44329) );
  inv_x4_sg U55468 ( .A(n14062), .X(n52571) );
  nand_x4_sg U55469 ( .A(n52570), .B(n14103), .X(n14062) );
  nand_x1_sg U55470 ( .A(n32018), .B(n32021), .X(n32046) );
  nand_x1_sg U55471 ( .A(n24352), .B(n24355), .X(n24380) );
  nand_x2_sg U55472 ( .A(n16726), .B(n16725), .X(n16722) );
  nand_x2_sg U55473 ( .A(n15160), .B(n15159), .X(n15156) );
  nand_x2_sg U55474 ( .A(n12827), .B(n12826), .X(n12823) );
  nand_x4_sg U55475 ( .A(n52838), .B(n14746), .X(n14705) );
  nand_x4_sg U55476 ( .A(n55091), .B(n20956), .X(n20915) );
  nand_x4_sg U55477 ( .A(n54523), .B(n19412), .X(n19371) );
  nand_x4_sg U55478 ( .A(n53958), .B(n17867), .X(n17826) );
  nor_x8_sg U55479 ( .A(n39300), .B(n46582), .X(n26079) );
  nor_x2_sg U55480 ( .A(n49742), .B(n49733), .X(n31806) );
  inv_x4_sg U55481 ( .A(n31698), .X(n49742) );
  nor_x2_sg U55482 ( .A(n49833), .B(n49791), .X(n31509) );
  inv_x4_sg U55483 ( .A(n31374), .X(n49833) );
  nor_x2_sg U55484 ( .A(n49879), .B(n49836), .X(n31338) );
  inv_x4_sg U55485 ( .A(n31184), .X(n49879) );
  nor_x2_sg U55486 ( .A(n49925), .B(n49882), .X(n31148) );
  inv_x4_sg U55487 ( .A(n30979), .X(n49925) );
  nor_x2_sg U55488 ( .A(n49969), .B(n49928), .X(n30943) );
  inv_x4_sg U55489 ( .A(n30753), .X(n49969) );
  nor_x2_sg U55490 ( .A(n50013), .B(n49972), .X(n30717) );
  inv_x4_sg U55491 ( .A(n30498), .X(n50013) );
  nor_x2_sg U55492 ( .A(n50057), .B(n50016), .X(n30462) );
  inv_x4_sg U55493 ( .A(n30227), .X(n50057) );
  inv_x4_sg U55494 ( .A(n44330), .X(n44331) );
  inv_x4_sg U55495 ( .A(n44332), .X(n44333) );
  nor_x2_sg U55496 ( .A(n50601), .B(n50592), .X(n24140) );
  inv_x4_sg U55497 ( .A(n24032), .X(n50601) );
  nor_x2_sg U55498 ( .A(n50692), .B(n50650), .X(n23843) );
  inv_x4_sg U55499 ( .A(n23708), .X(n50692) );
  nor_x2_sg U55500 ( .A(n50784), .B(n50741), .X(n23482) );
  inv_x4_sg U55501 ( .A(n23313), .X(n50784) );
  nor_x2_sg U55502 ( .A(n50872), .B(n50831), .X(n23051) );
  inv_x4_sg U55503 ( .A(n22832), .X(n50872) );
  nor_x2_sg U55504 ( .A(n50916), .B(n50875), .X(n22796) );
  inv_x4_sg U55505 ( .A(n22561), .X(n50916) );
  nor_x2_sg U55506 ( .A(n53434), .B(n16338), .X(n16337) );
  inv_x4_sg U55507 ( .A(n16339), .X(n53434) );
  nor_x2_sg U55508 ( .A(n51485), .B(n10883), .X(n10882) );
  inv_x4_sg U55509 ( .A(n10884), .X(n51485) );
  nor_x2_sg U55510 ( .A(n40772), .B(n49921), .X(n30961) );
  inv_x4_sg U55511 ( .A(n30740), .X(n49921) );
  nor_x2_sg U55512 ( .A(n50738), .B(n50695), .X(n23672) );
  inv_x4_sg U55513 ( .A(n23518), .X(n50738) );
  nor_x2_sg U55514 ( .A(n50828), .B(n50787), .X(n23277) );
  inv_x4_sg U55515 ( .A(n23087), .X(n50828) );
  inv_x4_sg U55516 ( .A(n10570), .X(n51347) );
  nand_x4_sg U55517 ( .A(n46558), .B(n10815), .X(n10813) );
  inv_x4_sg U55518 ( .A(n20766), .X(n55040) );
  inv_x4_sg U55519 ( .A(n19222), .X(n54472) );
  inv_x4_sg U55520 ( .A(n17677), .X(n53907) );
  inv_x4_sg U55521 ( .A(n14556), .X(n52787) );
  nor_x2_sg U55522 ( .A(n49788), .B(n49745), .X(n31662) );
  inv_x4_sg U55523 ( .A(n31545), .X(n49788) );
  nor_x2_sg U55524 ( .A(n50647), .B(n50604), .X(n23996) );
  inv_x4_sg U55525 ( .A(n23879), .X(n50647) );
  nor_x2_sg U55526 ( .A(n51657), .B(n11417), .X(n11416) );
  inv_x4_sg U55527 ( .A(n11471), .X(n51657) );
  nor_x2_sg U55528 ( .A(n53326), .B(n16092), .X(n16091) );
  inv_x4_sg U55529 ( .A(n16146), .X(n53326) );
  nor_x2_sg U55530 ( .A(n55017), .B(n20740), .X(n20739) );
  inv_x4_sg U55531 ( .A(n20792), .X(n55017) );
  nor_x2_sg U55532 ( .A(n54449), .B(n19196), .X(n19195) );
  inv_x4_sg U55533 ( .A(n19248), .X(n54449) );
  nor_x2_sg U55534 ( .A(n54166), .B(n18420), .X(n18419) );
  inv_x4_sg U55535 ( .A(n18472), .X(n54166) );
  nor_x2_sg U55536 ( .A(n53884), .B(n17651), .X(n17650) );
  inv_x4_sg U55537 ( .A(n17703), .X(n53884) );
  nor_x2_sg U55538 ( .A(n51378), .B(n10638), .X(n10637) );
  inv_x4_sg U55539 ( .A(n10690), .X(n51378) );
  nor_x4_sg U55540 ( .A(n11703), .B(n46545), .X(n11701) );
  nor_x4_sg U55541 ( .A(n46337), .B(n46346), .X(n18244) );
  nor_x4_sg U55542 ( .A(n46563), .B(n46570), .X(n10462) );
  nor_x4_sg U55543 ( .A(n12214), .B(n46514), .X(n12570) );
  nor_x4_sg U55544 ( .A(n46521), .B(n46528), .X(n11945) );
  nor_x4_sg U55545 ( .A(n10919), .B(n46570), .X(n10917) );
  nor_x4_sg U55546 ( .A(n46331), .B(n46335), .X(n18587) );
  inv_x4_sg U55547 ( .A(n21823), .X(n55429) );
  inv_x4_sg U55548 ( .A(n21052), .X(n55144) );
  inv_x4_sg U55549 ( .A(n20278), .X(n54861) );
  inv_x4_sg U55550 ( .A(n19508), .X(n54576) );
  inv_x4_sg U55551 ( .A(n18732), .X(n54293) );
  inv_x4_sg U55552 ( .A(n17963), .X(n54011) );
  inv_x4_sg U55553 ( .A(n17190), .X(n53730) );
  inv_x4_sg U55554 ( .A(n15624), .X(n53172) );
  inv_x4_sg U55555 ( .A(n14842), .X(n52891) );
  inv_x4_sg U55556 ( .A(n14071), .X(n52613) );
  inv_x4_sg U55557 ( .A(n13291), .X(n52338) );
  inv_x4_sg U55558 ( .A(n12510), .X(n52061) );
  inv_x4_sg U55559 ( .A(n11730), .X(n51781) );
  nor_x2_sg U55560 ( .A(n53521), .B(n16667), .X(n16666) );
  inv_x4_sg U55561 ( .A(n16671), .X(n53521) );
  nor_x2_sg U55562 ( .A(n52963), .B(n15101), .X(n15100) );
  inv_x4_sg U55563 ( .A(n15105), .X(n52963) );
  nor_x2_sg U55564 ( .A(n52129), .B(n12768), .X(n12767) );
  inv_x4_sg U55565 ( .A(n12772), .X(n52129) );
  nor_x2_sg U55566 ( .A(n51572), .B(n11207), .X(n11206) );
  inv_x4_sg U55567 ( .A(n11211), .X(n51572) );
  nor_x4_sg U55568 ( .A(n13964), .B(n46480), .X(n13979) );
  inv_x4_sg U55569 ( .A(n21074), .X(n55132) );
  inv_x4_sg U55570 ( .A(n19530), .X(n54564) );
  inv_x4_sg U55571 ( .A(n17985), .X(n53999) );
  inv_x4_sg U55572 ( .A(n14864), .X(n52879) );
  inv_x4_sg U55573 ( .A(n18187), .X(n54074) );
  nor_x2_sg U55574 ( .A(n14669), .B(n14672), .X(n14671) );
  nor_x4_sg U55575 ( .A(n14674), .B(n46463), .X(n14672) );
  inv_x4_sg U55576 ( .A(n32077), .X(n49320) );
  inv_x4_sg U55577 ( .A(n24411), .X(n50179) );
  inv_x4_sg U55578 ( .A(n44334), .X(n44335) );
  inv_x4_sg U55579 ( .A(n44336), .X(n44337) );
  inv_x4_sg U55580 ( .A(n44338), .X(n44339) );
  inv_x4_sg U55581 ( .A(n44340), .X(n44341) );
  inv_x4_sg U55582 ( .A(n11285), .X(n51606) );
  inv_x4_sg U55583 ( .A(n12022), .X(n51905) );
  nor_x4_sg U55584 ( .A(n46248), .B(n46244), .X(n21566) );
  nor_x4_sg U55585 ( .A(n46293), .B(n46289), .X(n20021) );
  nor_x4_sg U55586 ( .A(n46445), .B(n46449), .X(n14586) );
  nand_x4_sg U55587 ( .A(n44342), .B(n21253), .X(n21198) );
  nand_x4_sg U55588 ( .A(n44343), .B(n20481), .X(n20425) );
  nand_x4_sg U55589 ( .A(n44344), .B(n19708), .X(n19653) );
  nand_x4_sg U55590 ( .A(n44345), .B(n18937), .X(n18881) );
  nand_x4_sg U55591 ( .A(n44346), .B(n18163), .X(n18108) );
  nand_x4_sg U55592 ( .A(n44347), .B(n17392), .X(n17336) );
  nand_x4_sg U55593 ( .A(n44348), .B(n16608), .X(n16553) );
  nand_x4_sg U55594 ( .A(n44349), .B(n15826), .X(n15771) );
  nand_x4_sg U55595 ( .A(n44350), .B(n15042), .X(n14987) );
  nand_x4_sg U55596 ( .A(n44351), .B(n14273), .X(n14217) );
  nand_x4_sg U55597 ( .A(n44352), .B(n13493), .X(n13438) );
  nand_x4_sg U55598 ( .A(n44353), .B(n12709), .X(n12654) );
  nand_x4_sg U55599 ( .A(n44354), .B(n11931), .X(n11876) );
  nand_x4_sg U55600 ( .A(n44355), .B(n11148), .X(n11093) );
  nand_x4_sg U55601 ( .A(n44356), .B(n10381), .X(n10325) );
  nand_x4_sg U55602 ( .A(n52433), .B(n45477), .X(n13564) );
  inv_x2_sg U55603 ( .A(n53673), .X(n44357) );
  inv_x4_sg U55604 ( .A(n17076), .X(n53673) );
  inv_x2_sg U55605 ( .A(n53402), .X(n44358) );
  inv_x4_sg U55606 ( .A(n16292), .X(n53402) );
  inv_x2_sg U55607 ( .A(n53115), .X(n44359) );
  inv_x4_sg U55608 ( .A(n15510), .X(n53115) );
  inv_x2_sg U55609 ( .A(n52281), .X(n44360) );
  inv_x4_sg U55610 ( .A(n13177), .X(n52281) );
  inv_x2_sg U55611 ( .A(n52010), .X(n44361) );
  inv_x4_sg U55612 ( .A(n12397), .X(n52010) );
  inv_x4_sg U55613 ( .A(n44362), .X(n44363) );
  nand_x4_sg U55614 ( .A(n46269), .B(n46276), .X(n20528) );
  inv_x4_sg U55615 ( .A(n44364), .X(n44365) );
  nand_x4_sg U55616 ( .A(n46314), .B(n46321), .X(n18984) );
  inv_x4_sg U55617 ( .A(n44366), .X(n44367) );
  nand_x4_sg U55618 ( .A(n46361), .B(n46368), .X(n17439) );
  nand_x4_sg U55619 ( .A(n14320), .B(n14319), .X(n14327) );
  nor_x2_sg U55620 ( .A(n14319), .B(n14320), .X(n14318) );
  nor_x4_sg U55621 ( .A(n52658), .B(n14316), .X(n14320) );
  inv_x4_sg U55622 ( .A(n16266), .X(n53375) );
  nor_x4_sg U55623 ( .A(n16239), .B(n46407), .X(n16266) );
  inv_x4_sg U55624 ( .A(n44368), .X(n44369) );
  nand_x4_sg U55625 ( .A(n46564), .B(n46572), .X(n10424) );
  inv_x4_sg U55626 ( .A(n44370), .X(n44371) );
  inv_x4_sg U55627 ( .A(n44372), .X(n44373) );
  nor_x2_sg U55628 ( .A(n40794), .B(n8477), .X(n32097) );
  nor_x2_sg U55629 ( .A(n40793), .B(n8777), .X(n24431) );
  nor_x2_sg U55630 ( .A(n15732), .B(n53203), .X(n15731) );
  nand_x4_sg U55631 ( .A(n53208), .B(n53203), .X(n15739) );
  inv_x4_sg U55632 ( .A(n15729), .X(n53203) );
  nor_x2_sg U55633 ( .A(n11837), .B(n51815), .X(n11836) );
  nand_x4_sg U55634 ( .A(n51820), .B(n51815), .X(n11844) );
  inv_x4_sg U55635 ( .A(n11834), .X(n51815) );
  nor_x2_sg U55636 ( .A(n13399), .B(n52368), .X(n13398) );
  nand_x4_sg U55637 ( .A(n52372), .B(n52368), .X(n13406) );
  inv_x4_sg U55638 ( .A(n13396), .X(n52368) );
  nor_x2_sg U55639 ( .A(n19614), .B(n54610), .X(n19613) );
  nand_x4_sg U55640 ( .A(n54615), .B(n54610), .X(n19621) );
  inv_x4_sg U55641 ( .A(n19611), .X(n54610) );
  nor_x2_sg U55642 ( .A(n18069), .B(n54045), .X(n18068) );
  inv_x4_sg U55643 ( .A(n18066), .X(n54045) );
  nor_x2_sg U55644 ( .A(n21159), .B(n55178), .X(n21158) );
  nand_x4_sg U55645 ( .A(n55183), .B(n55178), .X(n21166) );
  inv_x4_sg U55646 ( .A(n21156), .X(n55178) );
  nor_x2_sg U55647 ( .A(n14178), .B(n52644), .X(n14177) );
  inv_x4_sg U55648 ( .A(n14175), .X(n52644) );
  inv_x4_sg U55649 ( .A(n44374), .X(n44375) );
  nand_x4_sg U55650 ( .A(n44375), .B(n21752), .X(n21750) );
  inv_x4_sg U55651 ( .A(n44376), .X(n44377) );
  nand_x4_sg U55652 ( .A(n44377), .B(n20207), .X(n20205) );
  inv_x4_sg U55653 ( .A(n44378), .X(n44379) );
  inv_x4_sg U55654 ( .A(n25415), .X(n51270) );
  nand_x4_sg U55655 ( .A(n10858), .B(n51321), .X(n10815) );
  inv_x4_sg U55656 ( .A(n10545), .X(n51321) );
  inv_x4_sg U55657 ( .A(n44380), .X(n44381) );
  inv_x4_sg U55658 ( .A(n44382), .X(n44383) );
  inv_x4_sg U55659 ( .A(n44384), .X(n44385) );
  nor_x4_sg U55660 ( .A(n46512), .B(n46523), .X(n12105) );
  inv_x4_sg U55661 ( .A(n15920), .X(n53261) );
  inv_x4_sg U55662 ( .A(n14365), .X(n52703) );
  inv_x4_sg U55663 ( .A(n10473), .X(n51314) );
  inv_x2_sg U55664 ( .A(\reg_yHat[5][7] ), .X(n45632) );
  inv_x2_sg U55665 ( .A(\reg_y[5][7] ), .X(n46032) );
  inv_x2_sg U55666 ( .A(\reg_yHat[4][0] ), .X(n45580) );
  inv_x4_sg U55667 ( .A(n44386), .X(n44387) );
  nor_x2_sg U55668 ( .A(n21214), .B(n55369), .X(n21212) );
  inv_x4_sg U55669 ( .A(n21215), .X(n55369) );
  inv_x4_sg U55670 ( .A(n44388), .X(n44389) );
  nor_x2_sg U55671 ( .A(n20441), .B(n55084), .X(n20439) );
  inv_x4_sg U55672 ( .A(n20442), .X(n55084) );
  inv_x4_sg U55673 ( .A(n44390), .X(n44391) );
  nor_x2_sg U55674 ( .A(n19669), .B(n54801), .X(n19667) );
  inv_x4_sg U55675 ( .A(n19670), .X(n54801) );
  inv_x4_sg U55676 ( .A(n44392), .X(n44393) );
  nor_x2_sg U55677 ( .A(n18897), .B(n54516), .X(n18895) );
  inv_x4_sg U55678 ( .A(n18898), .X(n54516) );
  inv_x4_sg U55679 ( .A(n44394), .X(n44395) );
  nor_x2_sg U55680 ( .A(n18124), .B(n54236), .X(n18122) );
  inv_x4_sg U55681 ( .A(n18125), .X(n54236) );
  inv_x4_sg U55682 ( .A(n44396), .X(n44397) );
  nor_x2_sg U55683 ( .A(n17352), .B(n53951), .X(n17350) );
  inv_x4_sg U55684 ( .A(n17353), .X(n53951) );
  inv_x4_sg U55685 ( .A(n44398), .X(n44399) );
  nor_x2_sg U55686 ( .A(n14233), .B(n52831), .X(n14231) );
  inv_x4_sg U55687 ( .A(n14234), .X(n52831) );
  inv_x4_sg U55688 ( .A(n44400), .X(n44401) );
  nor_x2_sg U55689 ( .A(n10341), .B(n51442), .X(n10339) );
  inv_x4_sg U55690 ( .A(n10342), .X(n51442) );
  inv_x4_sg U55691 ( .A(n44402), .X(n44403) );
  nor_x2_sg U55692 ( .A(n18182), .B(n18181), .X(n18179) );
  inv_x4_sg U55693 ( .A(n44404), .X(n44405) );
  nor_x2_sg U55694 ( .A(n14293), .B(n14292), .X(n14290) );
  inv_x4_sg U55695 ( .A(n44406), .X(n44407) );
  nor_x2_sg U55696 ( .A(n17092), .B(n53691), .X(n17091) );
  inv_x4_sg U55697 ( .A(n17093), .X(n53691) );
  inv_x4_sg U55698 ( .A(n44408), .X(n44409) );
  nor_x2_sg U55699 ( .A(n15526), .B(n53133), .X(n15525) );
  inv_x4_sg U55700 ( .A(n15527), .X(n53133) );
  inv_x4_sg U55701 ( .A(n44410), .X(n44411) );
  nor_x2_sg U55702 ( .A(n13973), .B(n52574), .X(n13972) );
  inv_x4_sg U55703 ( .A(n13974), .X(n52574) );
  inv_x4_sg U55704 ( .A(n44412), .X(n44413) );
  nor_x2_sg U55705 ( .A(n13193), .B(n52299), .X(n13192) );
  inv_x4_sg U55706 ( .A(n13194), .X(n52299) );
  nor_x1_sg U55707 ( .A(n29634), .B(n29635), .X(n29629) );
  inv_x2_sg U55708 ( .A(n44414), .X(n44415) );
  inv_x1_sg U55709 ( .A(n21668), .X(n55378) );
  nand_x4_sg U55710 ( .A(n55376), .B(n21725), .X(n21684) );
  inv_x2_sg U55711 ( .A(n44416), .X(n44417) );
  inv_x1_sg U55712 ( .A(n20123), .X(n54810) );
  nand_x4_sg U55713 ( .A(n54808), .B(n20180), .X(n20139) );
  inv_x1_sg U55714 ( .A(n18425), .X(n54189) );
  nor_x2_sg U55715 ( .A(n18445), .B(n18446), .X(n18443) );
  nor_x4_sg U55716 ( .A(n18515), .B(n54186), .X(n18445) );
  inv_x4_sg U55717 ( .A(n44418), .X(n44419) );
  nor_x2_sg U55718 ( .A(n53293), .B(n53278), .X(n16023) );
  inv_x4_sg U55719 ( .A(n16025), .X(n53278) );
  inv_x4_sg U55720 ( .A(n44420), .X(n44421) );
  nor_x2_sg U55721 ( .A(n51626), .B(n51610), .X(n11348) );
  inv_x4_sg U55722 ( .A(n11350), .X(n51610) );
  inv_x4_sg U55723 ( .A(n44422), .X(n44423) );
  nand_x1_sg U55724 ( .A(n44423), .B(n21436), .X(n21434) );
  inv_x4_sg U55725 ( .A(n44424), .X(n44425) );
  nand_x1_sg U55726 ( .A(n44425), .B(n19891), .X(n19889) );
  inv_x4_sg U55727 ( .A(n44426), .X(n44427) );
  nand_x1_sg U55728 ( .A(n44427), .B(n10564), .X(n10562) );
  nand_x4_sg U55729 ( .A(n44177), .B(n21633), .X(n21631) );
  nand_x4_sg U55730 ( .A(n44179), .B(n20088), .X(n20086) );
  nand_x4_sg U55731 ( .A(n44181), .B(n18543), .X(n18541) );
  nand_x4_sg U55732 ( .A(n44183), .B(n17004), .X(n17002) );
  nand_x4_sg U55733 ( .A(n44185), .B(n15438), .X(n15436) );
  nand_x4_sg U55734 ( .A(n44187), .B(n13885), .X(n13883) );
  nand_x4_sg U55735 ( .A(n44189), .B(n13105), .X(n13103) );
  nand_x4_sg U55736 ( .A(n44191), .B(n12324), .X(n12322) );
  nand_x4_sg U55737 ( .A(n44193), .B(n11544), .X(n11542) );
  inv_x4_sg U55738 ( .A(n12369), .X(n51893) );
  nor_x4_sg U55739 ( .A(n46512), .B(n12030), .X(n12369) );
  nand_x4_sg U55740 ( .A(n44213), .B(n18662), .X(n18660) );
  nand_x4_sg U55741 ( .A(n44215), .B(n14772), .X(n14770) );
  nand_x8_sg U55742 ( .A(n46576), .B(n27195), .X(n26783) );
  nor_x4_sg U55743 ( .A(n29607), .B(n29151), .X(n10266) );
  inv_x4_sg U55744 ( .A(n44428), .X(n44429) );
  nor_x2_sg U55745 ( .A(n55512), .B(n46195), .X(n18835) );
  inv_x8_sg U55746 ( .A(n26079), .X(n55512) );
  inv_x4_sg U55747 ( .A(n14171), .X(n55788) );
  nor_x2_sg U55748 ( .A(n14349), .B(n14350), .X(n14348) );
  nor_x4_sg U55749 ( .A(n42336), .B(n14334), .X(n14350) );
  nor_x2_sg U55750 ( .A(n10454), .B(n10455), .X(n10453) );
  nor_x4_sg U55751 ( .A(n41870), .B(n10442), .X(n10455) );
  inv_x4_sg U55752 ( .A(n44430), .X(n44431) );
  inv_x4_sg U55753 ( .A(n44432), .X(n44433) );
  inv_x4_sg U55754 ( .A(n44434), .X(n44435) );
  inv_x4_sg U55755 ( .A(n44436), .X(n44437) );
  inv_x4_sg U55756 ( .A(n44438), .X(n44439) );
  inv_x4_sg U55757 ( .A(n44440), .X(n44441) );
  inv_x4_sg U55758 ( .A(n44442), .X(n44443) );
  inv_x4_sg U55759 ( .A(n44444), .X(n44445) );
  inv_x4_sg U55760 ( .A(n44446), .X(n44447) );
  inv_x4_sg U55761 ( .A(n44448), .X(n44449) );
  inv_x4_sg U55762 ( .A(n44450), .X(n44451) );
  inv_x4_sg U55763 ( .A(n44452), .X(n44453) );
  inv_x4_sg U55764 ( .A(n44454), .X(n44455) );
  inv_x4_sg U55765 ( .A(n44456), .X(n44457) );
  inv_x4_sg U55766 ( .A(n44458), .X(n44459) );
  inv_x4_sg U55767 ( .A(n44460), .X(n44461) );
  nand_x8_sg U55768 ( .A(n53505), .B(n53509), .X(n27657) );
  inv_x4_sg U55769 ( .A(n27656), .X(n53505) );
  nand_x8_sg U55770 ( .A(n52947), .B(n52951), .X(n27097) );
  inv_x4_sg U55771 ( .A(n27096), .X(n52947) );
  nand_x8_sg U55772 ( .A(n52113), .B(n52117), .X(n26261) );
  inv_x4_sg U55773 ( .A(n26260), .X(n52113) );
  nand_x8_sg U55774 ( .A(n51556), .B(n51560), .X(n25702) );
  inv_x4_sg U55775 ( .A(n25701), .X(n51556) );
  inv_x4_sg U55776 ( .A(n44462), .X(n44463) );
  inv_x4_sg U55777 ( .A(n44464), .X(n44465) );
  nand_x8_sg U55778 ( .A(n54917), .B(n54921), .X(n29054) );
  inv_x4_sg U55779 ( .A(n29053), .X(n54917) );
  nand_x8_sg U55780 ( .A(n54349), .B(n54353), .X(n28495) );
  inv_x4_sg U55781 ( .A(n28494), .X(n54349) );
  nand_x8_sg U55782 ( .A(n53784), .B(n53788), .X(n27937) );
  inv_x4_sg U55783 ( .A(n27936), .X(n53784) );
  inv_x4_sg U55784 ( .A(n44466), .X(n44467) );
  inv_x4_sg U55785 ( .A(n44468), .X(n44469) );
  inv_x4_sg U55786 ( .A(n44470), .X(n44471) );
  inv_x4_sg U55787 ( .A(n44472), .X(n44473) );
  inv_x4_sg U55788 ( .A(n44474), .X(n44475) );
  inv_x4_sg U55789 ( .A(n44476), .X(n44477) );
  inv_x4_sg U55790 ( .A(n11637), .X(n51726) );
  inv_x4_sg U55791 ( .A(n44478), .X(n44479) );
  inv_x4_sg U55792 ( .A(n44480), .X(n44481) );
  inv_x4_sg U55793 ( .A(n44482), .X(n44483) );
  inv_x4_sg U55794 ( .A(n44484), .X(n44485) );
  inv_x4_sg U55795 ( .A(n44486), .X(n44487) );
  inv_x4_sg U55796 ( .A(n44488), .X(n44489) );
  inv_x4_sg U55797 ( .A(n44490), .X(n44491) );
  inv_x4_sg U55798 ( .A(n44492), .X(n44493) );
  inv_x4_sg U55799 ( .A(n44494), .X(n44495) );
  inv_x4_sg U55800 ( .A(n44496), .X(n44497) );
  inv_x4_sg U55801 ( .A(n44498), .X(n44499) );
  inv_x4_sg U55802 ( .A(n44500), .X(n44501) );
  inv_x4_sg U55803 ( .A(n44502), .X(n44503) );
  inv_x4_sg U55804 ( .A(n44504), .X(n44505) );
  inv_x4_sg U55805 ( .A(n44506), .X(n44507) );
  inv_x4_sg U55806 ( .A(n44508), .X(n44509) );
  inv_x4_sg U55807 ( .A(n44510), .X(n44511) );
  inv_x4_sg U55808 ( .A(n44512), .X(n44513) );
  inv_x4_sg U55809 ( .A(n44514), .X(n44515) );
  inv_x4_sg U55810 ( .A(n44516), .X(n44517) );
  inv_x4_sg U55811 ( .A(n44518), .X(n44519) );
  inv_x4_sg U55812 ( .A(n44520), .X(n44521) );
  inv_x4_sg U55813 ( .A(n44522), .X(n44523) );
  inv_x4_sg U55814 ( .A(n44524), .X(n44525) );
  inv_x4_sg U55815 ( .A(n44526), .X(n44527) );
  inv_x4_sg U55816 ( .A(n44528), .X(n44529) );
  inv_x4_sg U55817 ( .A(n44530), .X(n44531) );
  inv_x4_sg U55818 ( .A(n44532), .X(n44533) );
  inv_x4_sg U55819 ( .A(n44534), .X(n44535) );
  inv_x4_sg U55820 ( .A(n44536), .X(n44537) );
  inv_x4_sg U55821 ( .A(n44538), .X(n44539) );
  inv_x4_sg U55822 ( .A(n44540), .X(n44541) );
  inv_x4_sg U55823 ( .A(n44542), .X(n44543) );
  inv_x4_sg U55824 ( .A(n44544), .X(n44545) );
  inv_x4_sg U55825 ( .A(n44546), .X(n44547) );
  inv_x4_sg U55826 ( .A(n44548), .X(n44549) );
  inv_x4_sg U55827 ( .A(n44550), .X(n44551) );
  inv_x4_sg U55828 ( .A(n44552), .X(n44553) );
  inv_x4_sg U55829 ( .A(n44554), .X(n44555) );
  inv_x4_sg U55830 ( .A(n44556), .X(n44557) );
  inv_x4_sg U55831 ( .A(n44558), .X(n44559) );
  inv_x4_sg U55832 ( .A(n44560), .X(n44561) );
  inv_x4_sg U55833 ( .A(n44562), .X(n44563) );
  inv_x4_sg U55834 ( .A(n44564), .X(n44565) );
  inv_x4_sg U55835 ( .A(n44566), .X(n44567) );
  inv_x4_sg U55836 ( .A(n44568), .X(n44569) );
  inv_x4_sg U55837 ( .A(n44570), .X(n44571) );
  inv_x4_sg U55838 ( .A(n44572), .X(n44573) );
  inv_x4_sg U55839 ( .A(n44576), .X(n44577) );
  inv_x4_sg U55840 ( .A(n44578), .X(n44579) );
  inv_x4_sg U55841 ( .A(n44580), .X(n44581) );
  inv_x4_sg U55842 ( .A(n44582), .X(n44583) );
  inv_x4_sg U55843 ( .A(n44584), .X(n44585) );
  inv_x4_sg U55844 ( .A(n44586), .X(n44587) );
  inv_x4_sg U55845 ( .A(n44588), .X(n44589) );
  inv_x4_sg U55846 ( .A(n44590), .X(n44591) );
  inv_x4_sg U55847 ( .A(n44592), .X(n44593) );
  inv_x4_sg U55848 ( .A(n44594), .X(n44595) );
  inv_x4_sg U55849 ( .A(n44596), .X(n44597) );
  inv_x4_sg U55850 ( .A(n44598), .X(n44599) );
  inv_x4_sg U55851 ( .A(n44600), .X(n44601) );
  inv_x4_sg U55852 ( .A(n44602), .X(n44603) );
  inv_x4_sg U55853 ( .A(n44604), .X(n44605) );
  inv_x4_sg U55854 ( .A(n44606), .X(n44607) );
  inv_x4_sg U55855 ( .A(n44608), .X(n44609) );
  inv_x4_sg U55856 ( .A(n44610), .X(n44611) );
  inv_x4_sg U55857 ( .A(n44612), .X(n44613) );
  inv_x4_sg U55858 ( .A(n44614), .X(n44615) );
  inv_x4_sg U55859 ( .A(n44616), .X(n44617) );
  inv_x4_sg U55860 ( .A(n44618), .X(n44619) );
  inv_x4_sg U55861 ( .A(n44620), .X(n44621) );
  inv_x4_sg U55862 ( .A(n44622), .X(n44623) );
  inv_x4_sg U55863 ( .A(n44624), .X(n44625) );
  inv_x4_sg U55864 ( .A(n44626), .X(n44627) );
  inv_x4_sg U55865 ( .A(n44628), .X(n44629) );
  inv_x4_sg U55866 ( .A(n44630), .X(n44631) );
  inv_x4_sg U55867 ( .A(n44632), .X(n44633) );
  inv_x4_sg U55868 ( .A(n44634), .X(n44635) );
  inv_x4_sg U55869 ( .A(n44636), .X(n44637) );
  inv_x4_sg U55870 ( .A(n44638), .X(n44639) );
  inv_x4_sg U55871 ( .A(n44640), .X(n44641) );
  inv_x4_sg U55872 ( .A(n44642), .X(n44643) );
  inv_x4_sg U55873 ( .A(n44644), .X(n44645) );
  inv_x4_sg U55874 ( .A(n44646), .X(n44647) );
  inv_x4_sg U55875 ( .A(n44648), .X(n44649) );
  inv_x4_sg U55876 ( .A(n44650), .X(n44651) );
  inv_x4_sg U55877 ( .A(n44652), .X(n44653) );
  inv_x2_sg U55878 ( .A(n53658), .X(n44658) );
  inv_x4_sg U55879 ( .A(n16991), .X(n53657) );
  inv_x4_sg U55880 ( .A(n17039), .X(n53658) );
  inv_x2_sg U55881 ( .A(n53100), .X(n44659) );
  inv_x4_sg U55882 ( .A(n15425), .X(n53099) );
  inv_x4_sg U55883 ( .A(n15473), .X(n53100) );
  inv_x2_sg U55884 ( .A(n52542), .X(n44660) );
  inv_x4_sg U55885 ( .A(n13872), .X(n52541) );
  inv_x4_sg U55886 ( .A(n13920), .X(n52542) );
  inv_x2_sg U55887 ( .A(n52266), .X(n44661) );
  inv_x4_sg U55888 ( .A(n13092), .X(n52265) );
  inv_x4_sg U55889 ( .A(n13140), .X(n52266) );
  inv_x2_sg U55890 ( .A(n51710), .X(n44662) );
  inv_x4_sg U55891 ( .A(n11531), .X(n51709) );
  inv_x4_sg U55892 ( .A(n11579), .X(n51710) );
  inv_x2_sg U55893 ( .A(n54258), .X(n44663) );
  inv_x4_sg U55894 ( .A(n18812), .X(n54258) );
  inv_x2_sg U55895 ( .A(n51465), .X(n44664) );
  inv_x4_sg U55896 ( .A(n11025), .X(n51465) );
  inv_x2_sg U55897 ( .A(n55393), .X(n44667) );
  inv_x4_sg U55898 ( .A(n21902), .X(n55393) );
  inv_x2_sg U55899 ( .A(n54825), .X(n44668) );
  inv_x4_sg U55900 ( .A(n20357), .X(n54825) );
  nor_x4_sg U55901 ( .A(n12177), .B(n12176), .X(n12195) );
  inv_x4_sg U55902 ( .A(n44669), .X(n44670) );
  inv_x4_sg U55903 ( .A(n44671), .X(n44672) );
  inv_x4_sg U55904 ( .A(n44673), .X(n44674) );
  inv_x4_sg U55905 ( .A(n44675), .X(n44676) );
  nor_x4_sg U55906 ( .A(n16112), .B(n16113), .X(n16098) );
  nand_x4_sg U55907 ( .A(n46417), .B(n16057), .X(n16112) );
  nor_x4_sg U55908 ( .A(n13778), .B(n13779), .X(n13764) );
  nand_x4_sg U55909 ( .A(n46484), .B(n13723), .X(n13778) );
  nor_x4_sg U55910 ( .A(n12217), .B(n12218), .X(n12203) );
  nand_x4_sg U55911 ( .A(n46529), .B(n12162), .X(n12217) );
  nor_x4_sg U55912 ( .A(n16857), .B(n16856), .X(n16875) );
  nor_x4_sg U55913 ( .A(n15291), .B(n15290), .X(n15309) );
  nor_x4_sg U55914 ( .A(n12958), .B(n12957), .X(n12976) );
  nor_x4_sg U55915 ( .A(n13738), .B(n13737), .X(n13756) );
  nor_x4_sg U55916 ( .A(n46409), .B(n16069), .X(n16158) );
  inv_x2_sg U55917 ( .A(n52027), .X(n44677) );
  inv_x4_sg U55918 ( .A(n12584), .X(n52027) );
  nor_x4_sg U55919 ( .A(n10842), .B(n10843), .X(n10836) );
  nand_x4_sg U55920 ( .A(n46574), .B(n10754), .X(n10842) );
  nor_x4_sg U55921 ( .A(n16820), .B(n45539), .X(n16837) );
  nor_x4_sg U55922 ( .A(n16035), .B(n45541), .X(n16052) );
  nor_x4_sg U55923 ( .A(n15254), .B(n45543), .X(n15271) );
  nor_x4_sg U55924 ( .A(n13701), .B(n45545), .X(n13718) );
  nor_x4_sg U55925 ( .A(n12921), .B(n45547), .X(n12938) );
  nor_x4_sg U55926 ( .A(n12140), .B(n45549), .X(n12157) );
  nor_x4_sg U55927 ( .A(n11360), .B(n45551), .X(n11377) );
  inv_x4_sg U55928 ( .A(n16157), .X(n53295) );
  inv_x4_sg U55929 ( .A(n12262), .X(n51908) );
  inv_x4_sg U55930 ( .A(n16942), .X(n53566) );
  inv_x4_sg U55931 ( .A(n15376), .X(n53008) );
  inv_x4_sg U55932 ( .A(n13823), .X(n52449) );
  inv_x4_sg U55933 ( .A(n13043), .X(n52174) );
  inv_x4_sg U55934 ( .A(n44678), .X(n44679) );
  inv_x4_sg U55935 ( .A(n44680), .X(n44681) );
  inv_x4_sg U55936 ( .A(n44682), .X(n44683) );
  inv_x4_sg U55937 ( .A(n44684), .X(n44685) );
  inv_x4_sg U55938 ( .A(n44686), .X(n44687) );
  inv_x4_sg U55939 ( .A(n44688), .X(n44689) );
  inv_x4_sg U55940 ( .A(n44690), .X(n44691) );
  inv_x4_sg U55941 ( .A(n44692), .X(n44693) );
  inv_x4_sg U55942 ( .A(n12064), .X(n51875) );
  inv_x4_sg U55943 ( .A(n44694), .X(n44695) );
  inv_x4_sg U55944 ( .A(n44696), .X(n44697) );
  nor_x2_sg U55945 ( .A(n16787), .B(n16788), .X(n16786) );
  nand_x4_sg U55946 ( .A(n16818), .B(n53600), .X(n16787) );
  inv_x4_sg U55947 ( .A(n44698), .X(n44699) );
  nor_x2_sg U55948 ( .A(n16002), .B(n16003), .X(n16001) );
  nand_x4_sg U55949 ( .A(n16033), .B(n53321), .X(n16002) );
  inv_x4_sg U55950 ( .A(n44700), .X(n44701) );
  nor_x2_sg U55951 ( .A(n15221), .B(n15222), .X(n15220) );
  nand_x4_sg U55952 ( .A(n15252), .B(n53042), .X(n15221) );
  inv_x4_sg U55953 ( .A(n44702), .X(n44703) );
  nor_x2_sg U55954 ( .A(n13668), .B(n13669), .X(n13667) );
  nand_x4_sg U55955 ( .A(n13699), .B(n52485), .X(n13668) );
  inv_x4_sg U55956 ( .A(n44704), .X(n44705) );
  nor_x2_sg U55957 ( .A(n12888), .B(n12889), .X(n12887) );
  nand_x4_sg U55958 ( .A(n12919), .B(n52208), .X(n12888) );
  inv_x4_sg U55959 ( .A(n44706), .X(n44707) );
  nor_x2_sg U55960 ( .A(n12107), .B(n12108), .X(n12106) );
  nand_x4_sg U55961 ( .A(n12138), .B(n51933), .X(n12107) );
  inv_x4_sg U55962 ( .A(n44708), .X(n44709) );
  nor_x2_sg U55963 ( .A(n11327), .B(n11328), .X(n11326) );
  nand_x4_sg U55964 ( .A(n11358), .B(n51652), .X(n11327) );
  inv_x4_sg U55965 ( .A(n20710), .X(n55009) );
  inv_x4_sg U55966 ( .A(n19166), .X(n54441) );
  inv_x4_sg U55967 ( .A(n17621), .X(n53876) );
  inv_x4_sg U55968 ( .A(n14500), .X(n52756) );
  inv_x4_sg U55969 ( .A(n44710), .X(n44711) );
  nor_x4_sg U55970 ( .A(n21376), .B(n55253), .X(n21372) );
  nand_x4_sg U55971 ( .A(n55253), .B(n21376), .X(n21370) );
  nor_x4_sg U55972 ( .A(n55263), .B(n44711), .X(n21376) );
  inv_x4_sg U55973 ( .A(n21395), .X(n55263) );
  nand_x4_sg U55974 ( .A(n55256), .B(n46260), .X(n21394) );
  inv_x4_sg U55975 ( .A(n44712), .X(n44713) );
  nor_x4_sg U55976 ( .A(n19831), .B(n54685), .X(n19827) );
  nand_x4_sg U55977 ( .A(n54685), .B(n19831), .X(n19825) );
  nor_x4_sg U55978 ( .A(n54695), .B(n44713), .X(n19831) );
  inv_x4_sg U55979 ( .A(n19850), .X(n54695) );
  nand_x4_sg U55980 ( .A(n54688), .B(n46305), .X(n19849) );
  inv_x4_sg U55981 ( .A(n44714), .X(n44715) );
  nor_x4_sg U55982 ( .A(n14395), .B(n52721), .X(n14391) );
  nand_x4_sg U55983 ( .A(n52721), .B(n14395), .X(n14389) );
  nor_x4_sg U55984 ( .A(n52731), .B(n44715), .X(n14395) );
  inv_x4_sg U55985 ( .A(n14415), .X(n52731) );
  nand_x4_sg U55986 ( .A(n46443), .B(n14295), .X(n14414) );
  nor_x4_sg U55987 ( .A(n10504), .B(n51331), .X(n10500) );
  nand_x4_sg U55988 ( .A(n51331), .B(n10504), .X(n10498) );
  nor_x4_sg U55989 ( .A(n51341), .B(n10520), .X(n10504) );
  inv_x4_sg U55990 ( .A(n10523), .X(n51341) );
  nor_x4_sg U55991 ( .A(n10521), .B(n10522), .X(n10520) );
  inv_x4_sg U55992 ( .A(n29334), .X(n55200) );
  inv_x4_sg U55993 ( .A(n28773), .X(n54632) );
  inv_x4_sg U55994 ( .A(n28215), .X(n54066) );
  inv_x4_sg U55995 ( .A(n27376), .X(n53225) );
  inv_x4_sg U55996 ( .A(n26539), .X(n52389) );
  inv_x4_sg U55997 ( .A(n25979), .X(n51837) );
  inv_x4_sg U55998 ( .A(n25422), .X(n51278) );
  nand_x4_sg U55999 ( .A(n51270), .B(n46565), .X(n25422) );
  inv_x4_sg U56000 ( .A(n26817), .X(n52667) );
  inv_x4_sg U56001 ( .A(n44716), .X(n44717) );
  inv_x4_sg U56002 ( .A(n31978), .X(n49282) );
  inv_x4_sg U56003 ( .A(n24312), .X(n50141) );
  inv_x4_sg U56004 ( .A(n18216), .X(n54086) );
  inv_x4_sg U56005 ( .A(n15882), .X(n53242) );
  inv_x4_sg U56006 ( .A(n13548), .X(n52408) );
  inv_x4_sg U56007 ( .A(n11987), .X(n51856) );
  nand_x8_sg U56008 ( .A(n28271), .B(n18623), .X(n28278) );
  inv_x4_sg U56009 ( .A(n12587), .X(n51890) );
  inv_x4_sg U56010 ( .A(n15853), .X(n53215) );
  nand_x8_sg U56011 ( .A(n53214), .B(n46413), .X(n15853) );
  inv_x4_sg U56012 ( .A(n13519), .X(n52379) );
  nand_x8_sg U56013 ( .A(n52378), .B(n46481), .X(n13519) );
  inv_x4_sg U56014 ( .A(n11958), .X(n51827) );
  nand_x8_sg U56015 ( .A(n51826), .B(n46525), .X(n11958) );
  nor_x4_sg U56016 ( .A(n10759), .B(n51494), .X(n10716) );
  inv_x4_sg U56017 ( .A(n10760), .X(n51494) );
  nor_x4_sg U56018 ( .A(n45455), .B(n10762), .X(n10759) );
  nor_x4_sg U56019 ( .A(n21541), .B(n55366), .X(n21248) );
  inv_x4_sg U56020 ( .A(n21542), .X(n55366) );
  nor_x4_sg U56021 ( .A(n45389), .B(n21544), .X(n21541) );
  nor_x4_sg U56022 ( .A(n20771), .B(n55081), .X(n20476) );
  inv_x4_sg U56023 ( .A(n20772), .X(n55081) );
  nor_x4_sg U56024 ( .A(n45391), .B(n20774), .X(n20771) );
  nor_x4_sg U56025 ( .A(n19996), .B(n54798), .X(n19703) );
  inv_x4_sg U56026 ( .A(n19997), .X(n54798) );
  nor_x4_sg U56027 ( .A(n45393), .B(n19999), .X(n19996) );
  nor_x4_sg U56028 ( .A(n19227), .B(n54513), .X(n18932) );
  inv_x4_sg U56029 ( .A(n19228), .X(n54513) );
  nor_x4_sg U56030 ( .A(n45395), .B(n19230), .X(n19227) );
  nor_x4_sg U56031 ( .A(n18451), .B(n54233), .X(n18158) );
  inv_x4_sg U56032 ( .A(n18452), .X(n54233) );
  nor_x4_sg U56033 ( .A(n45397), .B(n18454), .X(n18451) );
  nor_x4_sg U56034 ( .A(n17682), .B(n53948), .X(n17387) );
  inv_x4_sg U56035 ( .A(n17683), .X(n53948) );
  nor_x4_sg U56036 ( .A(n45399), .B(n17685), .X(n17682) );
  nor_x4_sg U56037 ( .A(n14561), .B(n52828), .X(n14268) );
  inv_x4_sg U56038 ( .A(n14562), .X(n52828) );
  nor_x4_sg U56039 ( .A(n45401), .B(n14564), .X(n14561) );
  nor_x4_sg U56040 ( .A(n10669), .B(n51439), .X(n10376) );
  inv_x4_sg U56041 ( .A(n10670), .X(n51439) );
  nor_x4_sg U56042 ( .A(n45403), .B(n10672), .X(n10669) );
  inv_x4_sg U56043 ( .A(n18583), .X(n54144) );
  nor_x4_sg U56044 ( .A(n54143), .B(n46340), .X(n18583) );
  nor_x4_sg U56045 ( .A(n25371), .B(n8202), .X(n25338) );
  nor_x4_sg U56046 ( .A(n10264), .B(n8502), .X(n10230) );
  inv_x4_sg U56047 ( .A(n21001), .X(n55140) );
  nor_x4_sg U56048 ( .A(n21025), .B(n46275), .X(n21001) );
  inv_x4_sg U56049 ( .A(n19457), .X(n54572) );
  nor_x4_sg U56050 ( .A(n19481), .B(n46320), .X(n19457) );
  inv_x4_sg U56051 ( .A(n17912), .X(n54007) );
  nor_x4_sg U56052 ( .A(n17936), .B(n46367), .X(n17912) );
  inv_x4_sg U56053 ( .A(n21771), .X(n55425) );
  nor_x4_sg U56054 ( .A(n21796), .B(n46255), .X(n21771) );
  inv_x4_sg U56055 ( .A(n20226), .X(n54857) );
  nor_x4_sg U56056 ( .A(n20251), .B(n46300), .X(n20226) );
  inv_x4_sg U56057 ( .A(n29241), .X(n54890) );
  nor_x4_sg U56058 ( .A(n54889), .B(n45953), .X(n29241) );
  inv_x4_sg U56059 ( .A(n28680), .X(n54322) );
  nor_x4_sg U56060 ( .A(n54321), .B(n45955), .X(n28680) );
  inv_x4_sg U56061 ( .A(n28122), .X(n53757) );
  nor_x4_sg U56062 ( .A(n53756), .B(n45957), .X(n28122) );
  inv_x4_sg U56063 ( .A(n27562), .X(n53199) );
  nor_x4_sg U56064 ( .A(n53198), .B(n45959), .X(n27562) );
  inv_x4_sg U56065 ( .A(n26167), .X(n51811) );
  nor_x4_sg U56066 ( .A(n51810), .B(n45951), .X(n26167) );
  inv_x4_sg U56067 ( .A(n28401), .X(n54041) );
  nor_x4_sg U56068 ( .A(n54040), .B(n45949), .X(n28401) );
  inv_x4_sg U56069 ( .A(n27841), .X(n53479) );
  nor_x4_sg U56070 ( .A(n53478), .B(n45961), .X(n27841) );
  inv_x4_sg U56071 ( .A(n27283), .X(n52921) );
  nor_x4_sg U56072 ( .A(n52920), .B(n45963), .X(n27283) );
  inv_x4_sg U56073 ( .A(n26446), .X(n52087) );
  nor_x4_sg U56074 ( .A(n52086), .B(n45965), .X(n26446) );
  inv_x4_sg U56075 ( .A(n25887), .X(n51529) );
  nor_x4_sg U56076 ( .A(n51528), .B(n45967), .X(n25887) );
  inv_x4_sg U56077 ( .A(n28958), .X(n54606) );
  nor_x4_sg U56078 ( .A(n54605), .B(n45969), .X(n28958) );
  inv_x4_sg U56079 ( .A(n27003), .X(n52640) );
  nor_x4_sg U56080 ( .A(n52639), .B(n45971), .X(n27003) );
  inv_x4_sg U56081 ( .A(n25606), .X(n51253) );
  nor_x4_sg U56082 ( .A(n51252), .B(n45975), .X(n25606) );
  inv_x4_sg U56083 ( .A(n29519), .X(n55174) );
  nor_x4_sg U56084 ( .A(n55173), .B(n45973), .X(n29519) );
  inv_x4_sg U56085 ( .A(n17266), .X(n53559) );
  nand_x8_sg U56086 ( .A(n53548), .B(n16725), .X(n17266) );
  inv_x4_sg U56087 ( .A(n15700), .X(n53001) );
  nand_x8_sg U56088 ( .A(n52990), .B(n15159), .X(n15700) );
  inv_x4_sg U56089 ( .A(n14147), .X(n52441) );
  nand_x8_sg U56090 ( .A(n52430), .B(n46468), .X(n14147) );
  inv_x4_sg U56091 ( .A(n13367), .X(n52167) );
  nand_x8_sg U56092 ( .A(n52156), .B(n12826), .X(n13367) );
  inv_x4_sg U56093 ( .A(n10547), .X(n51315) );
  nand_x2_sg U56094 ( .A(n10548), .B(n10418), .X(n10547) );
  inv_x4_sg U56095 ( .A(n21521), .X(n55288) );
  inv_x4_sg U56096 ( .A(n20751), .X(n54996) );
  inv_x4_sg U56097 ( .A(n19976), .X(n54720) );
  inv_x4_sg U56098 ( .A(n19207), .X(n54428) );
  inv_x4_sg U56099 ( .A(n18431), .X(n54155) );
  inv_x4_sg U56100 ( .A(n17662), .X(n53863) );
  inv_x4_sg U56101 ( .A(n16888), .X(n53585) );
  inv_x4_sg U56102 ( .A(n16103), .X(n53305) );
  inv_x4_sg U56103 ( .A(n15322), .X(n53027) );
  inv_x4_sg U56104 ( .A(n14541), .X(n52743) );
  inv_x4_sg U56105 ( .A(n13769), .X(n52470) );
  inv_x4_sg U56106 ( .A(n12989), .X(n52193) );
  inv_x4_sg U56107 ( .A(n12208), .X(n51918) );
  inv_x4_sg U56108 ( .A(n11428), .X(n51637) );
  inv_x4_sg U56109 ( .A(n10649), .X(n51366) );
  inv_x4_sg U56110 ( .A(n11345), .X(n51620) );
  nor_x4_sg U56111 ( .A(n17162), .B(n46396), .X(n17235) );
  nor_x4_sg U56112 ( .A(n15596), .B(n46440), .X(n15669) );
  nor_x4_sg U56113 ( .A(n13263), .B(n46508), .X(n13336) );
  inv_x4_sg U56114 ( .A(n16805), .X(n53571) );
  inv_x4_sg U56115 ( .A(n16020), .X(n53287) );
  inv_x4_sg U56116 ( .A(n15239), .X(n53013) );
  inv_x4_sg U56117 ( .A(n13686), .X(n52454) );
  inv_x4_sg U56118 ( .A(n12906), .X(n52179) );
  inv_x4_sg U56119 ( .A(n12125), .X(n51902) );
  inv_x4_sg U56120 ( .A(n44718), .X(n44719) );
  nor_x4_sg U56121 ( .A(n18481), .B(n44719), .X(n18468) );
  nor_x4_sg U56122 ( .A(n18484), .B(n42603), .X(n18481) );
  nor_x4_sg U56123 ( .A(n16378), .B(n46416), .X(n16458) );
  nor_x4_sg U56124 ( .A(n55276), .B(n46246), .X(n21876) );
  nor_x4_sg U56125 ( .A(n54708), .B(n46291), .X(n20331) );
  nor_x4_sg U56126 ( .A(n54143), .B(n46335), .X(n18785) );
  inv_x8_sg U56127 ( .A(n46329), .X(n54143) );
  nor_x4_sg U56128 ( .A(n46535), .B(n51560), .X(n11573) );
  nor_x4_sg U56129 ( .A(n20613), .B(n54921), .X(n20894) );
  nor_x4_sg U56130 ( .A(n19069), .B(n54353), .X(n19350) );
  nor_x4_sg U56131 ( .A(n17524), .B(n53788), .X(n17805) );
  nor_x4_sg U56132 ( .A(n53702), .B(n16913), .X(n16569) );
  inv_x4_sg U56133 ( .A(n16602), .X(n53702) );
  nor_x4_sg U56134 ( .A(n16914), .B(n16915), .X(n16913) );
  nor_x4_sg U56135 ( .A(n53669), .B(n16862), .X(n16565) );
  inv_x4_sg U56136 ( .A(n16604), .X(n53669) );
  nor_x4_sg U56137 ( .A(n16863), .B(n16864), .X(n16862) );
  nor_x4_sg U56138 ( .A(n53421), .B(n16128), .X(n15787) );
  inv_x4_sg U56139 ( .A(n15820), .X(n53421) );
  nor_x4_sg U56140 ( .A(n16129), .B(n16130), .X(n16128) );
  nor_x4_sg U56141 ( .A(n53390), .B(n16077), .X(n15783) );
  inv_x4_sg U56142 ( .A(n15822), .X(n53390) );
  nor_x4_sg U56143 ( .A(n16078), .B(n16079), .X(n16077) );
  nor_x4_sg U56144 ( .A(n53144), .B(n15347), .X(n15003) );
  inv_x4_sg U56145 ( .A(n15036), .X(n53144) );
  nor_x4_sg U56146 ( .A(n15348), .B(n15349), .X(n15347) );
  nor_x4_sg U56147 ( .A(n53111), .B(n15296), .X(n14999) );
  inv_x4_sg U56148 ( .A(n15038), .X(n53111) );
  nor_x4_sg U56149 ( .A(n15297), .B(n15298), .X(n15296) );
  nor_x4_sg U56150 ( .A(n52585), .B(n13794), .X(n13454) );
  inv_x4_sg U56151 ( .A(n13487), .X(n52585) );
  nor_x4_sg U56152 ( .A(n13795), .B(n13796), .X(n13794) );
  nor_x4_sg U56153 ( .A(n52552), .B(n13743), .X(n13450) );
  inv_x4_sg U56154 ( .A(n13489), .X(n52552) );
  nor_x4_sg U56155 ( .A(n13744), .B(n13745), .X(n13743) );
  nor_x4_sg U56156 ( .A(n52310), .B(n13014), .X(n12670) );
  inv_x4_sg U56157 ( .A(n12703), .X(n52310) );
  nor_x4_sg U56158 ( .A(n13015), .B(n13016), .X(n13014) );
  nor_x4_sg U56159 ( .A(n52277), .B(n12963), .X(n12666) );
  inv_x4_sg U56160 ( .A(n12705), .X(n52277) );
  nor_x4_sg U56161 ( .A(n12964), .B(n12965), .X(n12963) );
  nor_x4_sg U56162 ( .A(n52035), .B(n12233), .X(n11892) );
  inv_x4_sg U56163 ( .A(n11925), .X(n52035) );
  nor_x4_sg U56164 ( .A(n12234), .B(n12235), .X(n12233) );
  nor_x4_sg U56165 ( .A(n52001), .B(n12182), .X(n11888) );
  inv_x4_sg U56166 ( .A(n11927), .X(n52001) );
  nor_x4_sg U56167 ( .A(n12183), .B(n12184), .X(n12182) );
  nor_x4_sg U56168 ( .A(n51752), .B(n11453), .X(n11109) );
  inv_x4_sg U56169 ( .A(n11142), .X(n51752) );
  nor_x4_sg U56170 ( .A(n11454), .B(n11455), .X(n11453) );
  nor_x4_sg U56171 ( .A(n51723), .B(n11402), .X(n11105) );
  inv_x4_sg U56172 ( .A(n11144), .X(n51723) );
  nor_x4_sg U56173 ( .A(n11403), .B(n11404), .X(n11402) );
  nor_x4_sg U56174 ( .A(n20685), .B(n20717), .X(n21105) );
  nor_x4_sg U56175 ( .A(n19141), .B(n19173), .X(n19561) );
  nor_x4_sg U56176 ( .A(n17596), .B(n17628), .X(n18016) );
  nor_x4_sg U56177 ( .A(n14507), .B(n46447), .X(n14895) );
  nor_x4_sg U56178 ( .A(n46406), .B(n46400), .X(n16117) );
  nor_x4_sg U56179 ( .A(n46535), .B(n46541), .X(n11442) );
  nor_x4_sg U56180 ( .A(n46537), .B(n11394), .X(n11782) );
  nor_x4_sg U56181 ( .A(n12482), .B(n46528), .X(n12555) );
  inv_x4_sg U56182 ( .A(n44720), .X(n44721) );
  nor_x4_sg U56183 ( .A(n18250), .B(n44721), .X(n18099) );
  nor_x4_sg U56184 ( .A(n18253), .B(n54134), .X(n18250) );
  nor_x4_sg U56185 ( .A(n46469), .B(n46477), .X(n13732) );
  nor_x4_sg U56186 ( .A(n14043), .B(n46485), .X(n14116) );
  nor_x4_sg U56187 ( .A(n51354), .B(n10518), .X(n10998) );
  nor_x4_sg U56188 ( .A(n46409), .B(n46402), .X(n16066) );
  nor_x4_sg U56189 ( .A(n15925), .B(n46411), .X(n15964) );
  nor_x4_sg U56190 ( .A(n46537), .B(n46545), .X(n11289) );
  nor_x4_sg U56191 ( .A(n17099), .B(n46387), .X(n17230) );
  nor_x4_sg U56192 ( .A(n15533), .B(n46431), .X(n15664) );
  nor_x4_sg U56193 ( .A(n13200), .B(n46499), .X(n13331) );
  nor_x4_sg U56194 ( .A(n46261), .B(n46242), .X(n21383) );
  nor_x4_sg U56195 ( .A(n46306), .B(n46287), .X(n19838) );
  nor_x4_sg U56196 ( .A(n46463), .B(n14411), .X(n14403) );
  nor_x4_sg U56197 ( .A(n46573), .B(n46559), .X(n10511) );
  nor_x4_sg U56198 ( .A(n46521), .B(n12344), .X(n12550) );
  inv_x4_sg U56199 ( .A(n26725), .X(n52364) );
  nor_x4_sg U56200 ( .A(n46456), .B(n14735), .X(n14886) );
  nor_x4_sg U56201 ( .A(n46274), .B(n20945), .X(n21096) );
  nor_x4_sg U56202 ( .A(n46319), .B(n19401), .X(n19552) );
  nor_x4_sg U56203 ( .A(n46366), .B(n17856), .X(n18007) );
  nor_x4_sg U56204 ( .A(n46254), .B(n21714), .X(n21867) );
  nor_x4_sg U56205 ( .A(n46299), .B(n20169), .X(n20322) );
  inv_x4_sg U56206 ( .A(n44722), .X(n44723) );
  nor_x4_sg U56207 ( .A(n49689), .B(n44723), .X(n31523) );
  inv_x4_sg U56208 ( .A(n31676), .X(n49689) );
  inv_x4_sg U56209 ( .A(n44724), .X(n44725) );
  nor_x4_sg U56210 ( .A(n50548), .B(n44725), .X(n23857) );
  inv_x4_sg U56211 ( .A(n24010), .X(n50548) );
  nand_x4_sg U56212 ( .A(n54050), .B(n18183), .X(n18171) );
  nand_x4_sg U56213 ( .A(n18183), .B(n18171), .X(n18182) );
  nor_x4_sg U56214 ( .A(n46344), .B(n46341), .X(n18183) );
  nand_x4_sg U56215 ( .A(n52649), .B(n14294), .X(n14281) );
  nand_x4_sg U56216 ( .A(n14294), .B(n14281), .X(n14293) );
  nor_x4_sg U56217 ( .A(n46454), .B(n46452), .X(n14294) );
  inv_x2_sg U56218 ( .A(n14724), .X(n52803) );
  nor_x4_sg U56219 ( .A(n14627), .B(n46454), .X(n14724) );
  inv_x2_sg U56220 ( .A(n13953), .X(n52522) );
  nor_x4_sg U56221 ( .A(n13856), .B(n46477), .X(n13953) );
  inv_x2_sg U56222 ( .A(n11612), .X(n51690) );
  nor_x4_sg U56223 ( .A(n11515), .B(n46543), .X(n11612) );
  inv_x4_sg U56224 ( .A(n44726), .X(n44727) );
  nor_x4_sg U56225 ( .A(n44727), .B(n55279), .X(n21423) );
  inv_x4_sg U56226 ( .A(n21484), .X(n55279) );
  nand_x2_sg U56227 ( .A(n21485), .B(n21486), .X(n21484) );
  nand_x4_sg U56228 ( .A(n46240), .B(n46260), .X(n21486) );
  inv_x4_sg U56229 ( .A(n44728), .X(n44729) );
  nor_x4_sg U56230 ( .A(n44729), .B(n54711), .X(n19878) );
  inv_x4_sg U56231 ( .A(n19939), .X(n54711) );
  nand_x2_sg U56232 ( .A(n19940), .B(n19941), .X(n19939) );
  nand_x4_sg U56233 ( .A(n46285), .B(n46305), .X(n19941) );
  inv_x4_sg U56234 ( .A(n9600), .X(n50748) );
  inv_x4_sg U56235 ( .A(n9503), .X(n50838) );
  inv_x4_sg U56236 ( .A(n24708), .X(n49889) );
  inv_x4_sg U56237 ( .A(n24611), .X(n49979) );
  nor_x4_sg U56238 ( .A(n20762), .B(n54947), .X(n20846) );
  nor_x4_sg U56239 ( .A(n19218), .B(n54379), .X(n19302) );
  nor_x4_sg U56240 ( .A(n18442), .B(n54097), .X(n18525) );
  nor_x4_sg U56241 ( .A(n17673), .B(n53814), .X(n17757) );
  nor_x4_sg U56242 ( .A(n16898), .B(n46377), .X(n16984) );
  nor_x4_sg U56243 ( .A(n15332), .B(n46421), .X(n15418) );
  nand_x4_sg U56244 ( .A(n14636), .B(n52678), .X(n14631) );
  nor_x4_sg U56245 ( .A(n14552), .B(n46445), .X(n14636) );
  nor_x4_sg U56246 ( .A(n12999), .B(n46489), .X(n13085) );
  nor_x4_sg U56247 ( .A(n11438), .B(n46533), .X(n11524) );
  nor_x2_sg U56248 ( .A(n55242), .B(n21477), .X(n21474) );
  inv_x2_sg U56249 ( .A(n21477), .X(n55306) );
  nor_x4_sg U56250 ( .A(n21532), .B(n46261), .X(n21477) );
  nor_x2_sg U56251 ( .A(n54674), .B(n19932), .X(n19929) );
  inv_x2_sg U56252 ( .A(n19932), .X(n54738) );
  nor_x4_sg U56253 ( .A(n19987), .B(n46306), .X(n19932) );
  nor_x2_sg U56254 ( .A(n51320), .B(n10605), .X(n10602) );
  inv_x2_sg U56255 ( .A(n10605), .X(n51384) );
  nor_x4_sg U56256 ( .A(n10660), .B(n46573), .X(n10605) );
  nor_x4_sg U56257 ( .A(n11638), .B(n46546), .X(n11589) );
  nor_x4_sg U56258 ( .A(n46379), .B(n46381), .X(n17050) );
  nor_x4_sg U56259 ( .A(n46423), .B(n46425), .X(n15484) );
  nor_x4_sg U56260 ( .A(n46467), .B(n46471), .X(n13931) );
  nor_x4_sg U56261 ( .A(n46491), .B(n46493), .X(n13151) );
  inv_x4_sg U56262 ( .A(n10286), .X(n51261) );
  nand_x4_sg U56263 ( .A(n53340), .B(n53207), .X(n16295) );
  inv_x4_sg U56264 ( .A(n16190), .X(n53340) );
  nor_x4_sg U56265 ( .A(n46252), .B(n46254), .X(n21297) );
  nor_x4_sg U56266 ( .A(n46297), .B(n46299), .X(n19752) );
  inv_x4_sg U56267 ( .A(n44730), .X(n44731) );
  nor_x4_sg U56268 ( .A(n50821), .B(n44731), .X(n22538) );
  inv_x4_sg U56269 ( .A(n22810), .X(n50821) );
  inv_x4_sg U56270 ( .A(n44732), .X(n44733) );
  nor_x4_sg U56271 ( .A(n49962), .B(n44733), .X(n30204) );
  inv_x4_sg U56272 ( .A(n30476), .X(n49962) );
  nor_x4_sg U56273 ( .A(n20837), .B(n46272), .X(n20934) );
  nor_x4_sg U56274 ( .A(n19293), .B(n46317), .X(n19390) );
  nor_x4_sg U56275 ( .A(n17748), .B(n46364), .X(n17845) );
  inv_x4_sg U56276 ( .A(n44734), .X(n44735) );
  nor_x2_sg U56277 ( .A(n40773), .B(n22583), .X(n22846) );
  nor_x4_sg U56278 ( .A(n44735), .B(n50882), .X(n22583) );
  inv_x4_sg U56279 ( .A(n22848), .X(n50882) );
  inv_x4_sg U56280 ( .A(n44736), .X(n44737) );
  nor_x2_sg U56281 ( .A(n40774), .B(n30249), .X(n30512) );
  nor_x4_sg U56282 ( .A(n44737), .B(n50023), .X(n30249) );
  inv_x4_sg U56283 ( .A(n30514), .X(n50023) );
  inv_x4_sg U56284 ( .A(n44738), .X(n44739) );
  nor_x4_sg U56285 ( .A(n53533), .B(n44739), .X(n16682) );
  inv_x4_sg U56286 ( .A(n16695), .X(n53533) );
  nand_x4_sg U56287 ( .A(n16696), .B(n53532), .X(n16693) );
  inv_x4_sg U56288 ( .A(n44740), .X(n44741) );
  nor_x4_sg U56289 ( .A(n52975), .B(n44741), .X(n15116) );
  inv_x4_sg U56290 ( .A(n15129), .X(n52975) );
  nand_x4_sg U56291 ( .A(n15130), .B(n52974), .X(n15127) );
  inv_x4_sg U56292 ( .A(n44742), .X(n44743) );
  nor_x4_sg U56293 ( .A(n52141), .B(n44743), .X(n12783) );
  inv_x4_sg U56294 ( .A(n12796), .X(n52141) );
  nand_x4_sg U56295 ( .A(n12797), .B(n52140), .X(n12794) );
  inv_x4_sg U56296 ( .A(n44744), .X(n44745) );
  nor_x4_sg U56297 ( .A(n51583), .B(n44745), .X(n11222) );
  inv_x4_sg U56298 ( .A(n11235), .X(n51583) );
  nand_x4_sg U56299 ( .A(n11236), .B(n51582), .X(n11233) );
  inv_x4_sg U56300 ( .A(n23607), .X(n50260) );
  inv_x4_sg U56301 ( .A(n31273), .X(n49401) );
  inv_x4_sg U56302 ( .A(n31327), .X(n49822) );
  inv_x4_sg U56303 ( .A(n23661), .X(n50681) );
  inv_x4_sg U56304 ( .A(n44746), .X(n44747) );
  nor_x2_sg U56305 ( .A(n29586), .B(n9373), .X(n29585) );
  nor_x4_sg U56306 ( .A(n50094), .B(n44747), .X(n29586) );
  inv_x4_sg U56307 ( .A(n30196), .X(n50094) );
  nand_x2_sg U56308 ( .A(n30195), .B(n29628), .X(n30196) );
  inv_x4_sg U56309 ( .A(n44748), .X(n44749) );
  nor_x2_sg U56310 ( .A(n21936), .B(n9373), .X(n21935) );
  nor_x4_sg U56311 ( .A(n50953), .B(n44749), .X(n21936) );
  inv_x4_sg U56312 ( .A(n22530), .X(n50953) );
  nand_x2_sg U56313 ( .A(n22529), .B(n21965), .X(n22530) );
  inv_x4_sg U56314 ( .A(n44750), .X(n44751) );
  nor_x4_sg U56315 ( .A(n14436), .B(n44751), .X(n14399) );
  nor_x4_sg U56316 ( .A(n14439), .B(n52711), .X(n14436) );
  inv_x4_sg U56317 ( .A(n44752), .X(n44753) );
  nor_x4_sg U56318 ( .A(n20644), .B(n44753), .X(n20609) );
  nor_x4_sg U56319 ( .A(n20647), .B(n54971), .X(n20644) );
  inv_x4_sg U56320 ( .A(n44754), .X(n44755) );
  nor_x4_sg U56321 ( .A(n19100), .B(n44755), .X(n19065) );
  nor_x4_sg U56322 ( .A(n19103), .B(n54403), .X(n19100) );
  inv_x4_sg U56323 ( .A(n44756), .X(n44757) );
  nor_x4_sg U56324 ( .A(n17555), .B(n44757), .X(n17520) );
  nor_x4_sg U56325 ( .A(n17558), .B(n53838), .X(n17555) );
  nor_x2_sg U56326 ( .A(n46337), .B(n18290), .X(n18325) );
  nor_x4_sg U56327 ( .A(n54112), .B(n18326), .X(n18290) );
  inv_x4_sg U56328 ( .A(n18328), .X(n54112) );
  nand_x2_sg U56329 ( .A(n54105), .B(n18327), .X(n18328) );
  nor_x4_sg U56330 ( .A(n18327), .B(n54105), .X(n18326) );
  nor_x4_sg U56331 ( .A(n21415), .B(n41516), .X(n21380) );
  nor_x4_sg U56332 ( .A(n21418), .B(n55243), .X(n21415) );
  nor_x4_sg U56333 ( .A(n19870), .B(n41520), .X(n19835) );
  nor_x4_sg U56334 ( .A(n19873), .B(n54675), .X(n19870) );
  nor_x4_sg U56335 ( .A(n25367), .B(n8282), .X(n30343) );
  nor_x4_sg U56336 ( .A(n10260), .B(n8582), .X(n22677) );
  nor_x4_sg U56337 ( .A(n10241), .B(n8702), .X(n23931) );
  nor_x4_sg U56338 ( .A(n25349), .B(n8402), .X(n31597) );
  nor_x4_sg U56339 ( .A(n25385), .B(n8242), .X(n29916) );
  nor_x4_sg U56340 ( .A(n10279), .B(n8542), .X(n22251) );
  nor_x4_sg U56341 ( .A(n25348), .B(n8442), .X(n31875) );
  nor_x4_sg U56342 ( .A(n10245), .B(n8742), .X(n24209) );
  nor_x4_sg U56343 ( .A(n25360), .B(n8322), .X(n30842) );
  nor_x4_sg U56344 ( .A(n10252), .B(n8622), .X(n23176) );
  nor_x4_sg U56345 ( .A(n25352), .B(n8382), .X(n31435) );
  nor_x4_sg U56346 ( .A(n10244), .B(n8682), .X(n23769) );
  nor_x4_sg U56347 ( .A(n25364), .B(n8262), .X(n30072) );
  nor_x4_sg U56348 ( .A(n10257), .B(n8562), .X(n22407) );
  nor_x4_sg U56349 ( .A(n25353), .B(n8342), .X(n31056) );
  nor_x4_sg U56350 ( .A(n10240), .B(n8642), .X(n23390) );
  nor_x4_sg U56351 ( .A(n25386), .B(n8222), .X(n29725) );
  nor_x4_sg U56352 ( .A(n10280), .B(n8522), .X(n22060) );
  nor_x4_sg U56353 ( .A(n25363), .B(n8302), .X(n30594) );
  nor_x4_sg U56354 ( .A(n10255), .B(n8602), .X(n22928) );
  nor_x4_sg U56355 ( .A(n39300), .B(n46200), .X(n21152) );
  inv_x4_sg U56356 ( .A(n44758), .X(n44759) );
  inv_x4_sg U56357 ( .A(n44760), .X(n44761) );
  inv_x4_sg U56358 ( .A(n44762), .X(n44763) );
  inv_x4_sg U56359 ( .A(n44764), .X(n44765) );
  inv_x4_sg U56360 ( .A(n44766), .X(n44767) );
  inv_x4_sg U56361 ( .A(n44768), .X(n44769) );
  inv_x4_sg U56362 ( .A(n44770), .X(n44771) );
  inv_x4_sg U56363 ( .A(n44772), .X(n44773) );
  inv_x4_sg U56364 ( .A(n44774), .X(n44775) );
  inv_x4_sg U56365 ( .A(n44776), .X(n44777) );
  inv_x4_sg U56366 ( .A(n44778), .X(n44779) );
  inv_x4_sg U56367 ( .A(n44780), .X(n44781) );
  inv_x4_sg U56368 ( .A(n44782), .X(n44783) );
  inv_x4_sg U56369 ( .A(n44784), .X(n44785) );
  inv_x4_sg U56370 ( .A(n44786), .X(n44787) );
  nor_x4_sg U56371 ( .A(n18654), .B(n46346), .X(n18636) );
  nand_x8_sg U56372 ( .A(n29080), .B(n20717), .X(n29087) );
  nor_x8_sg U56373 ( .A(n29073), .B(n46264), .X(n29080) );
  nand_x8_sg U56374 ( .A(n28521), .B(n19173), .X(n28528) );
  nor_x8_sg U56375 ( .A(n28514), .B(n46309), .X(n28521) );
  nand_x8_sg U56376 ( .A(n27963), .B(n17628), .X(n27970) );
  nor_x8_sg U56377 ( .A(n27956), .B(n46356), .X(n27963) );
  nand_x8_sg U56378 ( .A(n27403), .B(n16069), .X(n27410) );
  nor_x8_sg U56379 ( .A(n27396), .B(n53282), .X(n27403) );
  nand_x8_sg U56380 ( .A(n26844), .B(n14507), .X(n26851) );
  nor_x8_sg U56381 ( .A(n26837), .B(n46443), .X(n26844) );
  nor_x4_sg U56382 ( .A(n27704), .B(n53641), .X(n27711) );
  inv_x8_sg U56383 ( .A(n17099), .X(n53641) );
  nor_x4_sg U56384 ( .A(n27144), .B(n53083), .X(n27151) );
  inv_x8_sg U56385 ( .A(n15533), .X(n53083) );
  nor_x4_sg U56386 ( .A(n26587), .B(n52525), .X(n26594) );
  inv_x8_sg U56387 ( .A(n13980), .X(n52525) );
  nor_x4_sg U56388 ( .A(n26308), .B(n52249), .X(n26315) );
  inv_x8_sg U56389 ( .A(n13200), .X(n52249) );
  nand_x8_sg U56390 ( .A(n25449), .B(n25459), .X(n25456) );
  inv_x4_sg U56391 ( .A(n26078), .X(n55468) );
  inv_x4_sg U56392 ( .A(n17282), .X(n53726) );
  nor_x4_sg U56393 ( .A(n17162), .B(n46390), .X(n17282) );
  inv_x4_sg U56394 ( .A(n15716), .X(n53168) );
  nor_x4_sg U56395 ( .A(n15596), .B(n46434), .X(n15716) );
  inv_x4_sg U56396 ( .A(n14163), .X(n52609) );
  nor_x4_sg U56397 ( .A(n14043), .B(n46480), .X(n14163) );
  inv_x4_sg U56398 ( .A(n13383), .X(n52334) );
  nor_x4_sg U56399 ( .A(n13263), .B(n46502), .X(n13383) );
  inv_x4_sg U56400 ( .A(n44788), .X(n44789) );
  inv_x4_sg U56401 ( .A(n44790), .X(n44791) );
  inv_x4_sg U56402 ( .A(n44792), .X(n44793) );
  inv_x4_sg U56403 ( .A(n44793), .X(n50991) );
  inv_x4_sg U56404 ( .A(n44794), .X(n44795) );
  inv_x4_sg U56405 ( .A(n44796), .X(n44797) );
  inv_x4_sg U56406 ( .A(n44797), .X(n51220) );
  inv_x4_sg U56407 ( .A(n44798), .X(n44799) );
  inv_x4_sg U56408 ( .A(n44799), .X(n51182) );
  inv_x4_sg U56409 ( .A(n44800), .X(n44801) );
  inv_x4_sg U56410 ( .A(n44801), .X(n51145) );
  inv_x4_sg U56411 ( .A(n44802), .X(n44803) );
  inv_x4_sg U56412 ( .A(n44803), .X(n51218) );
  inv_x4_sg U56413 ( .A(n44804), .X(n44805) );
  inv_x4_sg U56414 ( .A(n44805), .X(n51180) );
  inv_x4_sg U56415 ( .A(n44806), .X(n44807) );
  inv_x4_sg U56416 ( .A(n44807), .X(n51143) );
  inv_x4_sg U56417 ( .A(n44808), .X(n44809) );
  inv_x4_sg U56418 ( .A(n44809), .X(n51219) );
  inv_x4_sg U56419 ( .A(n44810), .X(n44811) );
  inv_x4_sg U56420 ( .A(n44811), .X(n51181) );
  inv_x4_sg U56421 ( .A(n44812), .X(n44813) );
  inv_x4_sg U56422 ( .A(n44813), .X(n51144) );
  inv_x4_sg U56423 ( .A(n44814), .X(n44815) );
  inv_x4_sg U56424 ( .A(n44816), .X(n44817) );
  inv_x4_sg U56425 ( .A(n44818), .X(n44819) );
  inv_x4_sg U56426 ( .A(n44819), .X(n50990) );
  inv_x4_sg U56427 ( .A(n44820), .X(n44821) );
  inv_x4_sg U56428 ( .A(n44821), .X(n51124) );
  inv_x4_sg U56429 ( .A(n44822), .X(n44823) );
  inv_x4_sg U56430 ( .A(n44823), .X(n51086) );
  inv_x4_sg U56431 ( .A(n44824), .X(n44825) );
  inv_x4_sg U56432 ( .A(n44825), .X(n51028) );
  inv_x4_sg U56433 ( .A(n44826), .X(n44827) );
  inv_x4_sg U56434 ( .A(n44828), .X(n44829) );
  inv_x4_sg U56435 ( .A(n44830), .X(n44831) );
  inv_x4_sg U56436 ( .A(n44832), .X(n44833) );
  inv_x4_sg U56437 ( .A(n44833), .X(n51162) );
  inv_x4_sg U56438 ( .A(n44834), .X(n44835) );
  inv_x4_sg U56439 ( .A(n44836), .X(n44837) );
  inv_x4_sg U56440 ( .A(n44838), .X(n44839) );
  inv_x4_sg U56441 ( .A(n44840), .X(n44841) );
  inv_x4_sg U56442 ( .A(n44842), .X(n44843) );
  inv_x4_sg U56443 ( .A(n44844), .X(n44845) );
  inv_x4_sg U56444 ( .A(n44846), .X(n44847) );
  inv_x4_sg U56445 ( .A(n44848), .X(n44849) );
  inv_x4_sg U56446 ( .A(n44849), .X(n51123) );
  inv_x4_sg U56447 ( .A(n44850), .X(n44851) );
  inv_x4_sg U56448 ( .A(n44851), .X(n51085) );
  inv_x4_sg U56449 ( .A(n44852), .X(n44853) );
  inv_x4_sg U56450 ( .A(n44853), .X(n51027) );
  inv_x4_sg U56451 ( .A(n44854), .X(n44855) );
  inv_x4_sg U56452 ( .A(n44856), .X(n44857) );
  inv_x4_sg U56453 ( .A(n44858), .X(n44859) );
  inv_x4_sg U56454 ( .A(n44860), .X(n44861) );
  inv_x4_sg U56455 ( .A(n44862), .X(n44863) );
  inv_x4_sg U56456 ( .A(n44864), .X(n44865) );
  inv_x4_sg U56457 ( .A(n44866), .X(n44867) );
  inv_x4_sg U56458 ( .A(n44868), .X(n44869) );
  inv_x4_sg U56459 ( .A(n44869), .X(n51122) );
  inv_x4_sg U56460 ( .A(n44870), .X(n44871) );
  inv_x4_sg U56461 ( .A(n44871), .X(n51084) );
  inv_x4_sg U56462 ( .A(n44872), .X(n44873) );
  inv_x4_sg U56463 ( .A(n44873), .X(n51026) );
  inv_x4_sg U56464 ( .A(n44874), .X(n44875) );
  inv_x4_sg U56465 ( .A(n44876), .X(n44877) );
  inv_x4_sg U56466 ( .A(n44877), .X(n51046) );
  inv_x4_sg U56467 ( .A(n44878), .X(n44879) );
  inv_x4_sg U56468 ( .A(n44879), .X(n51179) );
  inv_x4_sg U56469 ( .A(n44880), .X(n44881) );
  inv_x4_sg U56470 ( .A(n44881), .X(n51142) );
  inv_x4_sg U56471 ( .A(n44882), .X(n44883) );
  inv_x4_sg U56472 ( .A(n44883), .X(n51217) );
  inv_x4_sg U56473 ( .A(n44884), .X(n44885) );
  inv_x4_sg U56474 ( .A(n44885), .X(n51007) );
  inv_x4_sg U56475 ( .A(n44886), .X(n44887) );
  inv_x4_sg U56476 ( .A(n44887), .X(n51103) );
  inv_x4_sg U56477 ( .A(n44888), .X(n44889) );
  inv_x4_sg U56478 ( .A(n44889), .X(n51178) );
  inv_x4_sg U56479 ( .A(n44890), .X(n44891) );
  inv_x4_sg U56480 ( .A(n44891), .X(n51141) );
  inv_x4_sg U56481 ( .A(n44892), .X(n44893) );
  inv_x4_sg U56482 ( .A(n44893), .X(n51216) );
  inv_x4_sg U56483 ( .A(n44894), .X(n44895) );
  inv_x4_sg U56484 ( .A(n44895), .X(n51197) );
  inv_x4_sg U56485 ( .A(n44896), .X(n44897) );
  inv_x4_sg U56486 ( .A(n44897), .X(n50988) );
  inv_x4_sg U56487 ( .A(n44898), .X(n44899) );
  inv_x4_sg U56488 ( .A(n44899), .X(n51235) );
  inv_x4_sg U56489 ( .A(n44900), .X(n44901) );
  inv_x4_sg U56490 ( .A(n44901), .X(n51065) );
  inv_x4_sg U56491 ( .A(n44902), .X(n44903) );
  inv_x4_sg U56492 ( .A(n44903), .X(n50969) );
  inv_x4_sg U56493 ( .A(n44904), .X(n44905) );
  inv_x4_sg U56494 ( .A(n44905), .X(n50989) );
  inv_x4_sg U56495 ( .A(n44906), .X(n44907) );
  inv_x4_sg U56496 ( .A(n44907), .X(n50992) );
  inv_x4_sg U56497 ( .A(n44908), .X(n44909) );
  inv_x1_sg U56498 ( .A(n44909), .X(n51249) );
  inv_x4_sg U56499 ( .A(n44910), .X(n44911) );
  inv_x1_sg U56500 ( .A(n44911), .X(n51248) );
  inv_x4_sg U56501 ( .A(n44912), .X(n44913) );
  inv_x1_sg U56502 ( .A(n44913), .X(n51247) );
  inv_x4_sg U56503 ( .A(n44914), .X(n44915) );
  inv_x1_sg U56504 ( .A(n44915), .X(n51244) );
  inv_x4_sg U56505 ( .A(n44916), .X(n44917) );
  inv_x1_sg U56506 ( .A(n44917), .X(n51243) );
  inv_x4_sg U56507 ( .A(n44918), .X(n44919) );
  inv_x1_sg U56508 ( .A(n44919), .X(n51242) );
  inv_x4_sg U56509 ( .A(n44920), .X(n44921) );
  inv_x1_sg U56510 ( .A(n44921), .X(n51240) );
  inv_x4_sg U56511 ( .A(n44922), .X(n44923) );
  inv_x1_sg U56512 ( .A(n44923), .X(n51230) );
  inv_x4_sg U56513 ( .A(n44924), .X(n44925) );
  inv_x1_sg U56514 ( .A(n44925), .X(n51229) );
  inv_x4_sg U56515 ( .A(n44926), .X(n44927) );
  inv_x1_sg U56516 ( .A(n44927), .X(n51228) );
  inv_x4_sg U56517 ( .A(n44928), .X(n44929) );
  inv_x1_sg U56518 ( .A(n44929), .X(n51226) );
  inv_x4_sg U56519 ( .A(n44930), .X(n44931) );
  inv_x1_sg U56520 ( .A(n44931), .X(n51224) );
  inv_x4_sg U56521 ( .A(n44932), .X(n44933) );
  inv_x1_sg U56522 ( .A(n44933), .X(n51223) );
  inv_x4_sg U56523 ( .A(n44934), .X(n44935) );
  inv_x1_sg U56524 ( .A(n44935), .X(n51221) );
  inv_x4_sg U56525 ( .A(n44936), .X(n44937) );
  inv_x1_sg U56526 ( .A(n44937), .X(n51211) );
  inv_x4_sg U56527 ( .A(n44938), .X(n44939) );
  inv_x1_sg U56528 ( .A(n44939), .X(n51210) );
  inv_x4_sg U56529 ( .A(n44940), .X(n44941) );
  inv_x1_sg U56530 ( .A(n44941), .X(n51209) );
  inv_x4_sg U56531 ( .A(n44942), .X(n44943) );
  inv_x1_sg U56532 ( .A(n44943), .X(n51206) );
  inv_x4_sg U56533 ( .A(n44944), .X(n44945) );
  inv_x1_sg U56534 ( .A(n44945), .X(n51205) );
  inv_x4_sg U56535 ( .A(n44946), .X(n44947) );
  inv_x1_sg U56536 ( .A(n44947), .X(n51204) );
  inv_x4_sg U56537 ( .A(n44948), .X(n44949) );
  inv_x1_sg U56538 ( .A(n44949), .X(n51202) );
  inv_x4_sg U56539 ( .A(n44950), .X(n44951) );
  inv_x1_sg U56540 ( .A(n44951), .X(n51192) );
  inv_x4_sg U56541 ( .A(n44952), .X(n44953) );
  inv_x1_sg U56542 ( .A(n44953), .X(n51191) );
  inv_x4_sg U56543 ( .A(n44954), .X(n44955) );
  inv_x1_sg U56544 ( .A(n44955), .X(n51190) );
  inv_x4_sg U56545 ( .A(n44956), .X(n44957) );
  inv_x1_sg U56546 ( .A(n44957), .X(n51188) );
  inv_x4_sg U56547 ( .A(n44958), .X(n44959) );
  inv_x1_sg U56548 ( .A(n44959), .X(n51186) );
  inv_x4_sg U56549 ( .A(n44960), .X(n44961) );
  inv_x1_sg U56550 ( .A(n44961), .X(n51185) );
  inv_x4_sg U56551 ( .A(n44962), .X(n44963) );
  inv_x1_sg U56552 ( .A(n44963), .X(n51183) );
  inv_x4_sg U56553 ( .A(n44964), .X(n44965) );
  inv_x1_sg U56554 ( .A(n44965), .X(n51173) );
  inv_x4_sg U56555 ( .A(n44966), .X(n44967) );
  inv_x1_sg U56556 ( .A(n44967), .X(n51172) );
  inv_x4_sg U56557 ( .A(n44968), .X(n44969) );
  inv_x1_sg U56558 ( .A(n44969), .X(n51171) );
  inv_x4_sg U56559 ( .A(n44970), .X(n44971) );
  inv_x1_sg U56560 ( .A(n44971), .X(n51170) );
  inv_x4_sg U56561 ( .A(n44972), .X(n44973) );
  inv_x1_sg U56562 ( .A(n44973), .X(n51169) );
  inv_x4_sg U56563 ( .A(n44974), .X(n44975) );
  inv_x1_sg U56564 ( .A(n44975), .X(n51168) );
  inv_x4_sg U56565 ( .A(n44976), .X(n44977) );
  inv_x1_sg U56566 ( .A(n44977), .X(n51167) );
  inv_x4_sg U56567 ( .A(n44978), .X(n44979) );
  inv_x1_sg U56568 ( .A(n44979), .X(n51166) );
  inv_x4_sg U56569 ( .A(n44980), .X(n44981) );
  inv_x1_sg U56570 ( .A(n44981), .X(n51164) );
  inv_x4_sg U56571 ( .A(n44982), .X(n44983) );
  inv_x1_sg U56572 ( .A(n44983), .X(n51155) );
  inv_x4_sg U56573 ( .A(n44984), .X(n44985) );
  inv_x1_sg U56574 ( .A(n44985), .X(n51154) );
  inv_x4_sg U56575 ( .A(n44986), .X(n44987) );
  inv_x1_sg U56576 ( .A(n44987), .X(n51153) );
  inv_x4_sg U56577 ( .A(n44988), .X(n44989) );
  inv_x1_sg U56578 ( .A(n44989), .X(n51151) );
  inv_x4_sg U56579 ( .A(n44990), .X(n44991) );
  inv_x1_sg U56580 ( .A(n44991), .X(n51149) );
  inv_x4_sg U56581 ( .A(n44992), .X(n44993) );
  inv_x1_sg U56582 ( .A(n44993), .X(n51148) );
  inv_x4_sg U56583 ( .A(n44994), .X(n44995) );
  inv_x1_sg U56584 ( .A(n44995), .X(n51146) );
  inv_x4_sg U56585 ( .A(n44996), .X(n44997) );
  inv_x1_sg U56586 ( .A(n44997), .X(n51136) );
  inv_x4_sg U56587 ( .A(n44998), .X(n44999) );
  inv_x1_sg U56588 ( .A(n44999), .X(n51135) );
  inv_x4_sg U56589 ( .A(n45000), .X(n45001) );
  inv_x1_sg U56590 ( .A(n45001), .X(n51134) );
  inv_x4_sg U56591 ( .A(n45002), .X(n45003) );
  inv_x1_sg U56592 ( .A(n45003), .X(n51133) );
  inv_x4_sg U56593 ( .A(n45004), .X(n45005) );
  inv_x1_sg U56594 ( .A(n45005), .X(n51131) );
  inv_x4_sg U56595 ( .A(n45006), .X(n45007) );
  inv_x1_sg U56596 ( .A(n45007), .X(n51129) );
  inv_x4_sg U56597 ( .A(n45008), .X(n45009) );
  inv_x1_sg U56598 ( .A(n45009), .X(n51127) );
  inv_x4_sg U56599 ( .A(n45010), .X(n45011) );
  inv_x1_sg U56600 ( .A(n45011), .X(n51117) );
  inv_x4_sg U56601 ( .A(n45012), .X(n45013) );
  inv_x1_sg U56602 ( .A(n45013), .X(n51116) );
  inv_x4_sg U56603 ( .A(n45014), .X(n45015) );
  inv_x1_sg U56604 ( .A(n45015), .X(n51115) );
  inv_x4_sg U56605 ( .A(n45016), .X(n45017) );
  inv_x1_sg U56606 ( .A(n45017), .X(n51114) );
  inv_x4_sg U56607 ( .A(n45018), .X(n45019) );
  inv_x1_sg U56608 ( .A(n45019), .X(n51112) );
  inv_x4_sg U56609 ( .A(n45020), .X(n45021) );
  inv_x1_sg U56610 ( .A(n45021), .X(n51111) );
  inv_x4_sg U56611 ( .A(n45022), .X(n45023) );
  inv_x1_sg U56612 ( .A(n45023), .X(n51110) );
  inv_x4_sg U56613 ( .A(n45024), .X(n45025) );
  inv_x1_sg U56614 ( .A(n45025), .X(n51108) );
  inv_x4_sg U56615 ( .A(n45026), .X(n45027) );
  inv_x1_sg U56616 ( .A(n45027), .X(n51098) );
  inv_x4_sg U56617 ( .A(n45028), .X(n45029) );
  inv_x1_sg U56618 ( .A(n45029), .X(n51097) );
  inv_x4_sg U56619 ( .A(n45030), .X(n45031) );
  inv_x1_sg U56620 ( .A(n45031), .X(n51096) );
  inv_x4_sg U56621 ( .A(n45032), .X(n45033) );
  inv_x1_sg U56622 ( .A(n45033), .X(n51095) );
  inv_x4_sg U56623 ( .A(n45034), .X(n45035) );
  inv_x1_sg U56624 ( .A(n45035), .X(n51093) );
  inv_x4_sg U56625 ( .A(n45036), .X(n45037) );
  inv_x1_sg U56626 ( .A(n45037), .X(n51091) );
  inv_x4_sg U56627 ( .A(n45038), .X(n45039) );
  inv_x1_sg U56628 ( .A(n45039), .X(n51089) );
  inv_x4_sg U56629 ( .A(n45040), .X(n45041) );
  inv_x1_sg U56630 ( .A(n45041), .X(n51079) );
  inv_x4_sg U56631 ( .A(n45042), .X(n45043) );
  inv_x1_sg U56632 ( .A(n45043), .X(n51078) );
  inv_x4_sg U56633 ( .A(n45044), .X(n45045) );
  inv_x1_sg U56634 ( .A(n45045), .X(n51077) );
  inv_x4_sg U56635 ( .A(n45046), .X(n45047) );
  inv_x1_sg U56636 ( .A(n45047), .X(n51075) );
  inv_x4_sg U56637 ( .A(n45048), .X(n45049) );
  inv_x1_sg U56638 ( .A(n45049), .X(n51073) );
  inv_x4_sg U56639 ( .A(n45050), .X(n45051) );
  inv_x1_sg U56640 ( .A(n45051), .X(n51072) );
  inv_x4_sg U56641 ( .A(n45052), .X(n45053) );
  inv_x1_sg U56642 ( .A(n45053), .X(n51070) );
  inv_x4_sg U56643 ( .A(n45054), .X(n45055) );
  inv_x1_sg U56644 ( .A(n45055), .X(n51060) );
  inv_x4_sg U56645 ( .A(n45056), .X(n45057) );
  inv_x1_sg U56646 ( .A(n45057), .X(n51059) );
  inv_x4_sg U56647 ( .A(n45058), .X(n45059) );
  inv_x1_sg U56648 ( .A(n45059), .X(n51058) );
  inv_x4_sg U56649 ( .A(n45060), .X(n45061) );
  inv_x1_sg U56650 ( .A(n45061), .X(n51057) );
  inv_x4_sg U56651 ( .A(n45062), .X(n45063) );
  inv_x1_sg U56652 ( .A(n45063), .X(n51055) );
  inv_x4_sg U56653 ( .A(n45064), .X(n45065) );
  inv_x1_sg U56654 ( .A(n45065), .X(n51053) );
  inv_x4_sg U56655 ( .A(n45066), .X(n45067) );
  inv_x1_sg U56656 ( .A(n45067), .X(n51051) );
  inv_x4_sg U56657 ( .A(n45068), .X(n45069) );
  inv_x1_sg U56658 ( .A(n45069), .X(n51040) );
  inv_x4_sg U56659 ( .A(n45070), .X(n45071) );
  inv_x1_sg U56660 ( .A(n45071), .X(n51039) );
  inv_x4_sg U56661 ( .A(n45072), .X(n45073) );
  inv_x1_sg U56662 ( .A(n45073), .X(n51038) );
  inv_x4_sg U56663 ( .A(n45074), .X(n45075) );
  inv_x1_sg U56664 ( .A(n45075), .X(n51037) );
  inv_x4_sg U56665 ( .A(n45076), .X(n45077) );
  inv_x1_sg U56666 ( .A(n45077), .X(n51035) );
  inv_x4_sg U56667 ( .A(n45078), .X(n45079) );
  inv_x1_sg U56668 ( .A(n45079), .X(n51033) );
  inv_x4_sg U56669 ( .A(n45080), .X(n45081) );
  inv_x1_sg U56670 ( .A(n45081), .X(n51031) );
  inv_x4_sg U56671 ( .A(n45082), .X(n45083) );
  inv_x1_sg U56672 ( .A(n45083), .X(n51021) );
  inv_x4_sg U56673 ( .A(n45084), .X(n45085) );
  inv_x1_sg U56674 ( .A(n45085), .X(n51020) );
  inv_x4_sg U56675 ( .A(n45086), .X(n45087) );
  inv_x1_sg U56676 ( .A(n45087), .X(n51019) );
  inv_x4_sg U56677 ( .A(n45088), .X(n45089) );
  inv_x1_sg U56678 ( .A(n45089), .X(n51018) );
  inv_x4_sg U56679 ( .A(n45090), .X(n45091) );
  inv_x1_sg U56680 ( .A(n45091), .X(n51016) );
  inv_x4_sg U56681 ( .A(n45092), .X(n45093) );
  inv_x1_sg U56682 ( .A(n45093), .X(n51015) );
  inv_x4_sg U56683 ( .A(n45094), .X(n45095) );
  inv_x1_sg U56684 ( .A(n45095), .X(n51014) );
  inv_x4_sg U56685 ( .A(n45096), .X(n45097) );
  inv_x1_sg U56686 ( .A(n45097), .X(n51012) );
  inv_x4_sg U56687 ( .A(n45098), .X(n45099) );
  inv_x1_sg U56688 ( .A(n45099), .X(n51002) );
  inv_x4_sg U56689 ( .A(n45100), .X(n45101) );
  inv_x1_sg U56690 ( .A(n45101), .X(n51001) );
  inv_x4_sg U56691 ( .A(n45102), .X(n45103) );
  inv_x1_sg U56692 ( .A(n45103), .X(n51000) );
  inv_x4_sg U56693 ( .A(n45104), .X(n45105) );
  inv_x1_sg U56694 ( .A(n45105), .X(n50999) );
  inv_x4_sg U56695 ( .A(n45106), .X(n45107) );
  inv_x1_sg U56696 ( .A(n45107), .X(n50997) );
  inv_x4_sg U56697 ( .A(n45108), .X(n45109) );
  inv_x1_sg U56698 ( .A(n45109), .X(n50996) );
  inv_x4_sg U56699 ( .A(n45110), .X(n45111) );
  inv_x1_sg U56700 ( .A(n45111), .X(n50995) );
  inv_x4_sg U56701 ( .A(n45112), .X(n45113) );
  inv_x1_sg U56702 ( .A(n45113), .X(n50993) );
  inv_x4_sg U56703 ( .A(n45114), .X(n45115) );
  inv_x1_sg U56704 ( .A(n45115), .X(n50981) );
  inv_x4_sg U56705 ( .A(n45116), .X(n45117) );
  inv_x1_sg U56706 ( .A(n45117), .X(n50980) );
  inv_x4_sg U56707 ( .A(n45118), .X(n45119) );
  inv_x1_sg U56708 ( .A(n45119), .X(n50978) );
  inv_x4_sg U56709 ( .A(n45120), .X(n45121) );
  inv_x1_sg U56710 ( .A(n45121), .X(n50977) );
  inv_x4_sg U56711 ( .A(n45122), .X(n45123) );
  inv_x1_sg U56712 ( .A(n45123), .X(n50976) );
  inv_x4_sg U56713 ( .A(n45124), .X(n45125) );
  inv_x1_sg U56714 ( .A(n45125), .X(n50974) );
  inv_x4_sg U56715 ( .A(n45126), .X(n45127) );
  inv_x1_sg U56716 ( .A(n45127), .X(n50983) );
  inv_x4_sg U56717 ( .A(n45128), .X(n45129) );
  inv_x1_sg U56718 ( .A(n45129), .X(n51076) );
  inv_x4_sg U56719 ( .A(n45130), .X(n45131) );
  inv_x1_sg U56720 ( .A(n45131), .X(n51227) );
  inv_x4_sg U56721 ( .A(n45132), .X(n45133) );
  inv_x1_sg U56722 ( .A(n45133), .X(n51189) );
  inv_x4_sg U56723 ( .A(n45134), .X(n45135) );
  inv_x1_sg U56724 ( .A(n45135), .X(n51152) );
  inv_x4_sg U56725 ( .A(n45136), .X(n45137) );
  inv_x1_sg U56726 ( .A(n45137), .X(n51054) );
  inv_x4_sg U56727 ( .A(n45138), .X(n45139) );
  inv_x1_sg U56728 ( .A(n45139), .X(n51130) );
  inv_x4_sg U56729 ( .A(n45140), .X(n45141) );
  inv_x1_sg U56730 ( .A(n45141), .X(n51092) );
  inv_x4_sg U56731 ( .A(n45142), .X(n45143) );
  inv_x1_sg U56732 ( .A(n45143), .X(n51034) );
  inv_x4_sg U56733 ( .A(n45144), .X(n45145) );
  inv_x1_sg U56734 ( .A(n45145), .X(n50982) );
  inv_x4_sg U56735 ( .A(n45146), .X(n45147) );
  inv_x1_sg U56736 ( .A(n45147), .X(n50998) );
  inv_x4_sg U56737 ( .A(n45148), .X(n45149) );
  inv_x1_sg U56738 ( .A(n45149), .X(n51245) );
  inv_x4_sg U56739 ( .A(n45150), .X(n45151) );
  inv_x1_sg U56740 ( .A(n45151), .X(n51207) );
  inv_x4_sg U56741 ( .A(n45152), .X(n45153) );
  inv_x1_sg U56742 ( .A(n45153), .X(n51017) );
  inv_x4_sg U56743 ( .A(n45154), .X(n45155) );
  inv_x1_sg U56744 ( .A(n45155), .X(n51246) );
  inv_x4_sg U56745 ( .A(n45156), .X(n45157) );
  inv_x1_sg U56746 ( .A(n45157), .X(n51208) );
  inv_x4_sg U56747 ( .A(n45158), .X(n45159) );
  inv_x1_sg U56748 ( .A(n45159), .X(n50994) );
  inv_x4_sg U56749 ( .A(n45160), .X(n45161) );
  inv_x1_sg U56750 ( .A(n45161), .X(n51113) );
  inv_x4_sg U56751 ( .A(n45162), .X(n45163) );
  inv_x1_sg U56752 ( .A(n45163), .X(n51056) );
  inv_x4_sg U56753 ( .A(n45164), .X(n45165) );
  inv_x1_sg U56754 ( .A(n45165), .X(n51128) );
  inv_x4_sg U56755 ( .A(n45166), .X(n45167) );
  inv_x1_sg U56756 ( .A(n45167), .X(n51090) );
  inv_x4_sg U56757 ( .A(n45168), .X(n45169) );
  inv_x1_sg U56758 ( .A(n45169), .X(n51032) );
  inv_x4_sg U56759 ( .A(n45170), .X(n45171) );
  inv_x1_sg U56760 ( .A(n45171), .X(n51052) );
  inv_x4_sg U56761 ( .A(n45172), .X(n45173) );
  inv_x1_sg U56762 ( .A(n45173), .X(n51013) );
  inv_x4_sg U56763 ( .A(n45174), .X(n45175) );
  inv_x1_sg U56764 ( .A(n45175), .X(n51132) );
  inv_x4_sg U56765 ( .A(n45176), .X(n45177) );
  inv_x1_sg U56766 ( .A(n45177), .X(n51094) );
  inv_x4_sg U56767 ( .A(n45178), .X(n45179) );
  inv_x1_sg U56768 ( .A(n45179), .X(n51036) );
  inv_x4_sg U56769 ( .A(n45180), .X(n45181) );
  inv_x1_sg U56770 ( .A(n45181), .X(n51109) );
  inv_x4_sg U56771 ( .A(n45182), .X(n45183) );
  inv_x1_sg U56772 ( .A(n45183), .X(n50979) );
  inv_x4_sg U56773 ( .A(n45184), .X(n45185) );
  inv_x1_sg U56774 ( .A(n45185), .X(n51074) );
  inv_x4_sg U56775 ( .A(n45186), .X(n45187) );
  inv_x1_sg U56776 ( .A(n45187), .X(n51225) );
  inv_x4_sg U56777 ( .A(n45188), .X(n45189) );
  inv_x1_sg U56778 ( .A(n45189), .X(n51187) );
  inv_x4_sg U56779 ( .A(n45190), .X(n45191) );
  inv_x1_sg U56780 ( .A(n45191), .X(n51150) );
  inv_x4_sg U56781 ( .A(n45192), .X(n45193) );
  inv_x1_sg U56782 ( .A(n45193), .X(n51222) );
  inv_x4_sg U56783 ( .A(n45194), .X(n45195) );
  inv_x1_sg U56784 ( .A(n45195), .X(n51184) );
  inv_x4_sg U56785 ( .A(n45196), .X(n45197) );
  inv_x1_sg U56786 ( .A(n45197), .X(n51147) );
  inv_x4_sg U56787 ( .A(n45198), .X(n45199) );
  inv_x1_sg U56788 ( .A(n45199), .X(n51071) );
  inv_x4_sg U56789 ( .A(n45200), .X(n45201) );
  inv_x1_sg U56790 ( .A(n45201), .X(n51165) );
  inv_x4_sg U56791 ( .A(n45202), .X(n45203) );
  inv_x1_sg U56792 ( .A(n45203), .X(n51241) );
  inv_x4_sg U56793 ( .A(n45204), .X(n45205) );
  inv_x1_sg U56794 ( .A(n45205), .X(n51203) );
  inv_x4_sg U56795 ( .A(n45206), .X(n45207) );
  inv_x1_sg U56796 ( .A(n45207), .X(n50975) );
  inv_x4_sg U56797 ( .A(n45208), .X(n45209) );
  nor_x4_sg U56798 ( .A(n46568), .B(n10782), .X(n10985) );
  nor_x4_sg U56799 ( .A(n16239), .B(n46409), .X(n16444) );
  nand_x4_sg U56800 ( .A(n51899), .B(n12257), .X(n12177) );
  nor_x8_sg U56801 ( .A(n12174), .B(n46523), .X(n12257) );
  nand_x4_sg U56802 ( .A(n53568), .B(n16937), .X(n16857) );
  nor_x8_sg U56803 ( .A(n16854), .B(n46389), .X(n16937) );
  nand_x4_sg U56804 ( .A(n53010), .B(n15371), .X(n15291) );
  nor_x8_sg U56805 ( .A(n15288), .B(n46433), .X(n15371) );
  nand_x4_sg U56806 ( .A(n52176), .B(n13038), .X(n12958) );
  nor_x8_sg U56807 ( .A(n12955), .B(n46501), .X(n13038) );
  nand_x4_sg U56808 ( .A(n52451), .B(n13818), .X(n13738) );
  nor_x8_sg U56809 ( .A(n13735), .B(n46479), .X(n13818) );
  nor_x8_sg U56810 ( .A(n46473), .B(n46477), .X(n13530) );
  nand_x4_sg U56811 ( .A(n16781), .B(n16651), .X(n16744) );
  nor_x8_sg U56812 ( .A(n53509), .B(n46387), .X(n16651) );
  nand_x4_sg U56813 ( .A(n15215), .B(n15085), .X(n15178) );
  nor_x8_sg U56814 ( .A(n52951), .B(n46431), .X(n15085) );
  nand_x4_sg U56815 ( .A(n12882), .B(n12752), .X(n12845) );
  nor_x8_sg U56816 ( .A(n52117), .B(n46499), .X(n12752) );
  nand_x4_sg U56817 ( .A(n12101), .B(n11969), .X(n12064) );
  nor_x8_sg U56818 ( .A(n46521), .B(n46516), .X(n11969) );
  inv_x4_sg U56819 ( .A(n45210), .X(n45211) );
  inv_x1_sg U56820 ( .A(n45211), .X(n54095) );
  inv_x4_sg U56821 ( .A(n45212), .X(n45213) );
  inv_x1_sg U56822 ( .A(n45213), .X(n53536) );
  inv_x4_sg U56823 ( .A(n45214), .X(n45215) );
  inv_x1_sg U56824 ( .A(n45215), .X(n52978) );
  inv_x4_sg U56825 ( .A(n45216), .X(n45217) );
  inv_x1_sg U56826 ( .A(n45217), .X(n52144) );
  inv_x4_sg U56827 ( .A(n45218), .X(n45219) );
  inv_x1_sg U56828 ( .A(n45219), .X(n54068) );
  inv_x4_sg U56829 ( .A(n45220), .X(n45221) );
  inv_x4_sg U56830 ( .A(n45222), .X(n45223) );
  inv_x4_sg U56831 ( .A(n45224), .X(n45225) );
  inv_x4_sg U56832 ( .A(n45226), .X(n45227) );
  inv_x4_sg U56833 ( .A(n45228), .X(n45229) );
  inv_x4_sg U56834 ( .A(n45230), .X(n45231) );
  inv_x4_sg U56835 ( .A(n45232), .X(n45233) );
  inv_x4_sg U56836 ( .A(n45234), .X(n45235) );
  inv_x4_sg U56837 ( .A(n45236), .X(n45237) );
  inv_x4_sg U56838 ( .A(n41139), .X(n45238) );
  inv_x8_sg U56839 ( .A(n45238), .X(state[1]) );
  inv_x4_sg U56840 ( .A(n41051), .X(n45240) );
  inv_x4_sg U56841 ( .A(n41131), .X(n45242) );
  inv_x8_sg U56842 ( .A(n45242), .X(n45243) );
  inv_x4_sg U56843 ( .A(n41119), .X(n45244) );
  inv_x8_sg U56844 ( .A(n45244), .X(n45245) );
  inv_x4_sg U56845 ( .A(n41107), .X(n45246) );
  inv_x8_sg U56846 ( .A(n45246), .X(n45247) );
  inv_x4_sg U56847 ( .A(n41083), .X(n45248) );
  inv_x8_sg U56848 ( .A(n45248), .X(n45249) );
  inv_x4_sg U56849 ( .A(n41123), .X(n45250) );
  inv_x8_sg U56850 ( .A(n45250), .X(n45251) );
  inv_x4_sg U56851 ( .A(n41111), .X(n45252) );
  inv_x8_sg U56852 ( .A(n45252), .X(n45253) );
  inv_x4_sg U56853 ( .A(n41103), .X(n45254) );
  inv_x8_sg U56854 ( .A(n45254), .X(n45255) );
  inv_x4_sg U56855 ( .A(n41095), .X(n45256) );
  inv_x8_sg U56856 ( .A(n45256), .X(n45257) );
  inv_x4_sg U56857 ( .A(n41055), .X(n45258) );
  inv_x8_sg U56858 ( .A(n45258), .X(n45259) );
  inv_x4_sg U56859 ( .A(n41075), .X(n45260) );
  inv_x8_sg U56860 ( .A(n45260), .X(n45261) );
  inv_x4_sg U56861 ( .A(n41063), .X(n45262) );
  inv_x8_sg U56862 ( .A(n45262), .X(n45263) );
  inv_x4_sg U56863 ( .A(n41099), .X(n45264) );
  inv_x8_sg U56864 ( .A(n45264), .X(n45265) );
  inv_x4_sg U56865 ( .A(n41087), .X(n45266) );
  inv_x8_sg U56866 ( .A(n45266), .X(n45267) );
  inv_x4_sg U56867 ( .A(n41067), .X(n45268) );
  inv_x8_sg U56868 ( .A(n45268), .X(n45269) );
  inv_x4_sg U56869 ( .A(n41105), .X(n45270) );
  inv_x4_sg U56870 ( .A(n41073), .X(n45272) );
  inv_x4_sg U56871 ( .A(n41047), .X(n45274) );
  inv_x4_sg U56872 ( .A(n41129), .X(n45276) );
  inv_x4_sg U56873 ( .A(n41117), .X(n45278) );
  inv_x4_sg U56874 ( .A(n41059), .X(n45280) );
  inv_x4_sg U56875 ( .A(n41081), .X(n45282) );
  inv_x4_sg U56876 ( .A(n41091), .X(n45284) );
  inv_x4_sg U56877 ( .A(n41127), .X(n45286) );
  inv_x4_sg U56878 ( .A(n41115), .X(n45288) );
  inv_x4_sg U56879 ( .A(n41071), .X(n45290) );
  inv_x4_sg U56880 ( .A(n41061), .X(n45292) );
  inv_x4_sg U56881 ( .A(n41121), .X(n45294) );
  inv_x4_sg U56882 ( .A(n41109), .X(n45296) );
  inv_x4_sg U56883 ( .A(n41101), .X(n45298) );
  inv_x4_sg U56884 ( .A(n41093), .X(n45300) );
  inv_x4_sg U56885 ( .A(n41045), .X(n45302) );
  inv_x4_sg U56886 ( .A(n41053), .X(n45304) );
  inv_x4_sg U56887 ( .A(n41089), .X(n45306) );
  inv_x4_sg U56888 ( .A(n41079), .X(n45308) );
  inv_x4_sg U56889 ( .A(n41113), .X(n45310) );
  inv_x4_sg U56890 ( .A(n41077), .X(n45312) );
  inv_x4_sg U56891 ( .A(n41125), .X(n45314) );
  inv_x4_sg U56892 ( .A(n41069), .X(n45316) );
  inv_x4_sg U56893 ( .A(n41097), .X(n45318) );
  inv_x4_sg U56894 ( .A(n41085), .X(n45320) );
  inv_x4_sg U56895 ( .A(n41065), .X(n45322) );
  inv_x4_sg U56896 ( .A(n41057), .X(n45324) );
  inv_x4_sg U56897 ( .A(n41049), .X(n45326) );
  inv_x8_sg U56898 ( .A(n29151), .X(n55460) );
  nand_x4_sg U56899 ( .A(n54935), .B(n20521), .X(n20538) );
  nand_x4_sg U56900 ( .A(n54367), .B(n18977), .X(n18994) );
  nand_x4_sg U56901 ( .A(n53802), .B(n17432), .X(n17449) );
  nand_x4_sg U56902 ( .A(n54084), .B(n46352), .X(n18215) );
  inv_x1_sg U56903 ( .A(n16836), .X(n53607) );
  inv_x1_sg U56904 ( .A(n16051), .X(n53328) );
  inv_x1_sg U56905 ( .A(n15270), .X(n53049) );
  inv_x1_sg U56906 ( .A(n13717), .X(n52492) );
  inv_x1_sg U56907 ( .A(n12937), .X(n52215) );
  inv_x1_sg U56908 ( .A(n12156), .X(n51940) );
  inv_x1_sg U56909 ( .A(n11376), .X(n51659) );
  nand_x4_sg U56910 ( .A(n18387), .B(n18386), .X(n18429) );
  inv_x4_sg U56911 ( .A(n16668), .X(n53527) );
  nand_x4_sg U56912 ( .A(n16662), .B(n16661), .X(n16668) );
  inv_x4_sg U56913 ( .A(n15102), .X(n52969) );
  nand_x4_sg U56914 ( .A(n15096), .B(n15095), .X(n15102) );
  inv_x4_sg U56915 ( .A(n12769), .X(n52135) );
  nand_x4_sg U56916 ( .A(n12763), .B(n12762), .X(n12769) );
  inv_x4_sg U56917 ( .A(n11208), .X(n51577) );
  nand_x4_sg U56918 ( .A(n11202), .B(n11201), .X(n11208) );
  inv_x4_sg U56919 ( .A(n21307), .X(n55217) );
  nand_x4_sg U56920 ( .A(n21300), .B(n21299), .X(n21307) );
  inv_x4_sg U56921 ( .A(n19762), .X(n54649) );
  nand_x4_sg U56922 ( .A(n19755), .B(n19754), .X(n19762) );
  nand_x4_sg U56923 ( .A(n15857), .B(n15856), .X(n15862) );
  nand_x4_sg U56924 ( .A(n54130), .B(n18304), .X(n18321) );
  inv_x4_sg U56925 ( .A(n18305), .X(n54130) );
  nand_x4_sg U56926 ( .A(n20707), .B(n20706), .X(n20749) );
  nand_x4_sg U56927 ( .A(n19163), .B(n19162), .X(n19205) );
  nand_x4_sg U56928 ( .A(n17618), .B(n17617), .X(n17660) );
  nand_x4_sg U56929 ( .A(n14497), .B(n14496), .X(n14539) );
  inv_x1_sg U56930 ( .A(n17075), .X(n53695) );
  inv_x1_sg U56931 ( .A(n15509), .X(n53137) );
  inv_x1_sg U56932 ( .A(n13956), .X(n52578) );
  inv_x1_sg U56933 ( .A(n13176), .X(n52303) );
  inv_x1_sg U56934 ( .A(n20937), .X(n55108) );
  inv_x1_sg U56935 ( .A(n19393), .X(n54540) );
  inv_x1_sg U56936 ( .A(n17848), .X(n53975) );
  inv_x1_sg U56937 ( .A(n14727), .X(n52855) );
  inv_x4_sg U56938 ( .A(n11009), .X(n51392) );
  nor_x4_sg U56939 ( .A(n10660), .B(n46565), .X(n11009) );
  nor_x4_sg U56940 ( .A(n10546), .B(n10545), .X(n10569) );
  inv_x2_sg U56941 ( .A(n10546), .X(n51307) );
  nand_x8_sg U56942 ( .A(n51306), .B(n46569), .X(n10546) );
  nand_x4_sg U56943 ( .A(n17095), .B(n53674), .X(n17054) );
  nand_x4_sg U56944 ( .A(n15529), .B(n53116), .X(n15488) );
  nand_x4_sg U56945 ( .A(n13976), .B(n52557), .X(n13935) );
  nand_x4_sg U56946 ( .A(n13196), .B(n52282), .X(n13155) );
  nand_x4_sg U56947 ( .A(n17200), .B(n17201), .X(n17116) );
  nand_x4_sg U56948 ( .A(n15634), .B(n15635), .X(n15550) );
  nand_x4_sg U56949 ( .A(n14081), .B(n14082), .X(n13997) );
  nand_x4_sg U56950 ( .A(n13301), .B(n13302), .X(n13217) );
  nand_x4_sg U56951 ( .A(n12520), .B(n12521), .X(n12436) );
  nand_x4_sg U56952 ( .A(n11740), .B(n11741), .X(n11656) );
  nand_x4_sg U56953 ( .A(n16414), .B(n16415), .X(n16331) );
  nor_x4_sg U56954 ( .A(n12344), .B(n46523), .X(n12416) );
  nand_x4_sg U56955 ( .A(n16980), .B(n16981), .X(n16978) );
  nand_x4_sg U56956 ( .A(n16195), .B(n16196), .X(n16193) );
  nand_x4_sg U56957 ( .A(n15414), .B(n15415), .X(n15412) );
  nand_x4_sg U56958 ( .A(n13861), .B(n13862), .X(n13859) );
  nand_x4_sg U56959 ( .A(n13081), .B(n13082), .X(n13079) );
  nand_x4_sg U56960 ( .A(n12300), .B(n12301), .X(n12298) );
  nand_x4_sg U56961 ( .A(n11520), .B(n11521), .X(n11518) );
  nand_x4_sg U56962 ( .A(n21611), .B(n21612), .X(n21609) );
  nand_x4_sg U56963 ( .A(n20842), .B(n20843), .X(n20840) );
  nand_x4_sg U56964 ( .A(n20066), .B(n20067), .X(n20064) );
  nand_x4_sg U56965 ( .A(n19298), .B(n19299), .X(n19296) );
  nand_x4_sg U56966 ( .A(n18521), .B(n18522), .X(n18519) );
  nand_x4_sg U56967 ( .A(n17753), .B(n17754), .X(n17751) );
  nand_x4_sg U56968 ( .A(n14632), .B(n14633), .X(n14630) );
  nor_x2_sg U56969 ( .A(n49696), .B(n49686), .X(n31799) );
  inv_x4_sg U56970 ( .A(n31801), .X(n49696) );
  inv_x4_sg U56971 ( .A(n18329), .X(n54105) );
  nor_x2_sg U56972 ( .A(n50555), .B(n50545), .X(n24133) );
  inv_x4_sg U56973 ( .A(n24135), .X(n50555) );
  nor_x2_sg U56974 ( .A(n40775), .B(n49738), .X(n31680) );
  inv_x4_sg U56975 ( .A(n31532), .X(n49738) );
  nor_x2_sg U56976 ( .A(n40776), .B(n49829), .X(n31356) );
  inv_x4_sg U56977 ( .A(n31171), .X(n49829) );
  nor_x2_sg U56978 ( .A(n40777), .B(n49965), .X(n30735) );
  inv_x4_sg U56979 ( .A(n30485), .X(n49965) );
  inv_x4_sg U56980 ( .A(n16803), .X(n53517) );
  inv_x4_sg U56981 ( .A(n16018), .X(n53233) );
  inv_x4_sg U56982 ( .A(n15237), .X(n52959) );
  inv_x4_sg U56983 ( .A(n13684), .X(n52399) );
  inv_x4_sg U56984 ( .A(n12904), .X(n52125) );
  inv_x4_sg U56985 ( .A(n12123), .X(n51847) );
  inv_x4_sg U56986 ( .A(n11343), .X(n51568) );
  inv_x4_sg U56987 ( .A(n17217), .X(n53716) );
  inv_x4_sg U56988 ( .A(n15651), .X(n53158) );
  inv_x4_sg U56989 ( .A(n14098), .X(n52599) );
  inv_x4_sg U56990 ( .A(n13318), .X(n52324) );
  nor_x2_sg U56991 ( .A(n40778), .B(n49647), .X(n31940) );
  inv_x4_sg U56992 ( .A(n31829), .X(n49647) );
  inv_x4_sg U56993 ( .A(n10956), .X(n51372) );
  inv_x4_sg U56994 ( .A(n10992), .X(n51453) );
  nor_x2_sg U56995 ( .A(n40779), .B(n50780), .X(n23295) );
  inv_x4_sg U56996 ( .A(n23074), .X(n50780) );
  inv_x4_sg U56997 ( .A(n16207), .X(n53310) );
  nor_x2_sg U56998 ( .A(n40780), .B(n50506), .X(n24274) );
  inv_x4_sg U56999 ( .A(n24163), .X(n50506) );
  nor_x2_sg U57000 ( .A(n40781), .B(n50597), .X(n24014) );
  inv_x4_sg U57001 ( .A(n23866), .X(n50597) );
  nor_x2_sg U57002 ( .A(n40782), .B(n50688), .X(n23690) );
  inv_x4_sg U57003 ( .A(n23505), .X(n50688) );
  inv_x4_sg U57004 ( .A(n21112), .X(n55001) );
  inv_x4_sg U57005 ( .A(n19568), .X(n54433) );
  nor_x4_sg U57006 ( .A(n18437), .B(n46346), .X(n18435) );
  inv_x4_sg U57007 ( .A(n18023), .X(n53868) );
  inv_x4_sg U57008 ( .A(n17242), .X(n53591) );
  inv_x4_sg U57009 ( .A(n16465), .X(n53311) );
  inv_x4_sg U57010 ( .A(n15676), .X(n53033) );
  inv_x4_sg U57011 ( .A(n14902), .X(n52748) );
  inv_x4_sg U57012 ( .A(n14123), .X(n52476) );
  inv_x4_sg U57013 ( .A(n13343), .X(n52199) );
  inv_x4_sg U57014 ( .A(n12561), .X(n51923) );
  nor_x4_sg U57015 ( .A(n12214), .B(n46523), .X(n12212) );
  inv_x4_sg U57016 ( .A(n11791), .X(n51643) );
  nor_x4_sg U57017 ( .A(n10655), .B(n46570), .X(n10653) );
  nand_x4_sg U57018 ( .A(n51377), .B(n51280), .X(n11036) );
  inv_x8_sg U57019 ( .A(n10660), .X(n51377) );
  nor_x2_sg U57020 ( .A(n50039), .B(n49995), .X(n29832) );
  inv_x4_sg U57021 ( .A(n29834), .X(n50039) );
  nor_x2_sg U57022 ( .A(n50898), .B(n50854), .X(n22167) );
  inv_x4_sg U57023 ( .A(n22169), .X(n50898) );
  inv_x4_sg U57024 ( .A(n16426), .X(n53440) );
  inv_x4_sg U57025 ( .A(n10968), .X(n51491) );
  nor_x4_sg U57026 ( .A(n46248), .B(n46254), .X(n21334) );
  nor_x4_sg U57027 ( .A(n46293), .B(n46299), .X(n19789) );
  nor_x4_sg U57028 ( .A(n46385), .B(n46396), .X(n16631) );
  nor_x4_sg U57029 ( .A(n46429), .B(n46440), .X(n15065) );
  nor_x4_sg U57030 ( .A(n46497), .B(n46508), .X(n12732) );
  nor_x4_sg U57031 ( .A(n46541), .B(n46552), .X(n11171) );
  inv_x4_sg U57032 ( .A(n45328), .X(n45329) );
  inv_x4_sg U57033 ( .A(n45330), .X(n45331) );
  inv_x4_sg U57034 ( .A(n45332), .X(n45333) );
  inv_x4_sg U57035 ( .A(n45334), .X(n45335) );
  nor_x2_sg U57036 ( .A(n21766), .B(n55445), .X(n21765) );
  inv_x4_sg U57037 ( .A(n21777), .X(n55445) );
  nor_x2_sg U57038 ( .A(n20996), .B(n55161), .X(n20995) );
  inv_x4_sg U57039 ( .A(n21006), .X(n55161) );
  nor_x2_sg U57040 ( .A(n20221), .B(n54877), .X(n20220) );
  inv_x4_sg U57041 ( .A(n20232), .X(n54877) );
  nor_x2_sg U57042 ( .A(n19452), .B(n54593), .X(n19451) );
  inv_x4_sg U57043 ( .A(n19462), .X(n54593) );
  nor_x2_sg U57044 ( .A(n18676), .B(n54309), .X(n18675) );
  inv_x4_sg U57045 ( .A(n18686), .X(n54309) );
  nor_x2_sg U57046 ( .A(n17907), .B(n54028), .X(n17906) );
  inv_x4_sg U57047 ( .A(n17917), .X(n54028) );
  nor_x2_sg U57048 ( .A(n17134), .B(n53744), .X(n17133) );
  inv_x4_sg U57049 ( .A(n17143), .X(n53744) );
  nor_x2_sg U57050 ( .A(n15568), .B(n53186), .X(n15567) );
  inv_x4_sg U57051 ( .A(n15577), .X(n53186) );
  nor_x2_sg U57052 ( .A(n14786), .B(n52908), .X(n14785) );
  inv_x4_sg U57053 ( .A(n14796), .X(n52908) );
  nor_x2_sg U57054 ( .A(n14015), .B(n52627), .X(n14014) );
  inv_x4_sg U57055 ( .A(n14024), .X(n52627) );
  nor_x2_sg U57056 ( .A(n13235), .B(n52352), .X(n13234) );
  inv_x4_sg U57057 ( .A(n13244), .X(n52352) );
  nor_x2_sg U57058 ( .A(n12454), .B(n52074), .X(n12453) );
  inv_x4_sg U57059 ( .A(n12463), .X(n52074) );
  nor_x2_sg U57060 ( .A(n11674), .B(n51798), .X(n11673) );
  inv_x4_sg U57061 ( .A(n11684), .X(n51798) );
  inv_x4_sg U57062 ( .A(n21278), .X(n55206) );
  inv_x4_sg U57063 ( .A(n19733), .X(n54638) );
  inv_x4_sg U57064 ( .A(n14298), .X(n52674) );
  inv_x4_sg U57065 ( .A(n10406), .X(n51284) );
  inv_x4_sg U57066 ( .A(n20394), .X(n54905) );
  inv_x4_sg U57067 ( .A(n18850), .X(n54337) );
  inv_x4_sg U57068 ( .A(n17305), .X(n53772) );
  nor_x2_sg U57069 ( .A(n46411), .B(n53216), .X(n15836) );
  inv_x4_sg U57070 ( .A(n15740), .X(n53216) );
  nor_x2_sg U57071 ( .A(n46523), .B(n51828), .X(n11941) );
  inv_x4_sg U57072 ( .A(n11845), .X(n51828) );
  nor_x2_sg U57073 ( .A(n46479), .B(n52380), .X(n13503) );
  inv_x4_sg U57074 ( .A(n13407), .X(n52380) );
  nor_x2_sg U57075 ( .A(n46299), .B(n54621), .X(n19718) );
  inv_x4_sg U57076 ( .A(n19622), .X(n54621) );
  nor_x2_sg U57077 ( .A(n46346), .B(n54054), .X(n18173) );
  inv_x4_sg U57078 ( .A(n18077), .X(n54054) );
  nor_x4_sg U57079 ( .A(n46402), .B(n46411), .X(n15994) );
  inv_x4_sg U57080 ( .A(n16745), .X(n53556) );
  inv_x4_sg U57081 ( .A(n15179), .X(n52998) );
  inv_x4_sg U57082 ( .A(n12846), .X(n52164) );
  inv_x4_sg U57083 ( .A(n10841), .X(n51406) );
  nor_x4_sg U57084 ( .A(n46555), .B(n46570), .X(n10841) );
  inv_x4_sg U57085 ( .A(n21342), .X(n55266) );
  inv_x4_sg U57086 ( .A(n20573), .X(n54987) );
  inv_x4_sg U57087 ( .A(n19797), .X(n54698) );
  inv_x4_sg U57088 ( .A(n19029), .X(n54419) );
  inv_x4_sg U57089 ( .A(n18252), .X(n54134) );
  inv_x4_sg U57090 ( .A(n17484), .X(n53854) );
  inv_x4_sg U57091 ( .A(n16706), .X(n53574) );
  inv_x4_sg U57092 ( .A(n15917), .X(n53290) );
  inv_x4_sg U57093 ( .A(n15140), .X(n53016) );
  inv_x4_sg U57094 ( .A(n14362), .X(n52734) );
  inv_x4_sg U57095 ( .A(n13583), .X(n52458) );
  inv_x4_sg U57096 ( .A(n12807), .X(n52182) );
  inv_x4_sg U57097 ( .A(n11246), .X(n51623) );
  inv_x4_sg U57098 ( .A(n10470), .X(n51344) );
  nor_x4_sg U57099 ( .A(n46561), .B(n46563), .X(n10694) );
  nor_x2_sg U57100 ( .A(n46254), .B(n55189), .X(n21263) );
  inv_x4_sg U57101 ( .A(n21167), .X(n55189) );
  nor_x2_sg U57102 ( .A(n46456), .B(n52656), .X(n14283) );
  inv_x4_sg U57103 ( .A(n14186), .X(n52656) );
  nor_x2_sg U57104 ( .A(n46570), .B(n51267), .X(n10391) );
  inv_x4_sg U57105 ( .A(n10294), .X(n51267) );
  inv_x4_sg U57106 ( .A(n21833), .X(n55294) );
  inv_x4_sg U57107 ( .A(n20288), .X(n54726) );
  inv_x4_sg U57108 ( .A(n18742), .X(n54160) );
  nand_x4_sg U57109 ( .A(n18209), .B(n18208), .X(n18216) );
  nor_x2_sg U57110 ( .A(n18208), .B(n18209), .X(n18207) );
  nor_x4_sg U57111 ( .A(n18205), .B(n41871), .X(n18209) );
  nand_x4_sg U57112 ( .A(n15875), .B(n15874), .X(n15882) );
  nor_x2_sg U57113 ( .A(n15874), .B(n15875), .X(n15873) );
  nor_x4_sg U57114 ( .A(n15890), .B(n15853), .X(n15875) );
  nand_x4_sg U57115 ( .A(n11980), .B(n11979), .X(n11987) );
  nor_x2_sg U57116 ( .A(n11979), .B(n11980), .X(n11978) );
  nor_x4_sg U57117 ( .A(n11995), .B(n11958), .X(n11980) );
  inv_x4_sg U57118 ( .A(n45336), .X(n45337) );
  inv_x4_sg U57119 ( .A(n45338), .X(n45339) );
  inv_x4_sg U57120 ( .A(n45340), .X(n45341) );
  inv_x4_sg U57121 ( .A(n45342), .X(n45343) );
  inv_x4_sg U57122 ( .A(n45344), .X(n45345) );
  inv_x4_sg U57123 ( .A(n45346), .X(n45347) );
  inv_x4_sg U57124 ( .A(n45348), .X(n45349) );
  inv_x4_sg U57125 ( .A(n45350), .X(n45351) );
  inv_x4_sg U57126 ( .A(n45352), .X(n45353) );
  inv_x4_sg U57127 ( .A(n45354), .X(n45355) );
  inv_x4_sg U57128 ( .A(n45356), .X(n45357) );
  inv_x4_sg U57129 ( .A(n45358), .X(n45359) );
  inv_x4_sg U57130 ( .A(n45360), .X(n45361) );
  inv_x4_sg U57131 ( .A(n45362), .X(n45363) );
  inv_x4_sg U57132 ( .A(n45364), .X(n45365) );
  inv_x4_sg U57133 ( .A(n45366), .X(n45367) );
  inv_x4_sg U57134 ( .A(n45368), .X(n45369) );
  inv_x4_sg U57135 ( .A(n45370), .X(n45371) );
  inv_x4_sg U57136 ( .A(n45372), .X(n45373) );
  inv_x4_sg U57137 ( .A(n45374), .X(n45375) );
  inv_x4_sg U57138 ( .A(n45376), .X(n45377) );
  inv_x4_sg U57139 ( .A(n45378), .X(n45379) );
  inv_x4_sg U57140 ( .A(n45380), .X(n45381) );
  inv_x4_sg U57141 ( .A(n45382), .X(n45383) );
  inv_x4_sg U57142 ( .A(n45384), .X(n45385) );
  inv_x4_sg U57143 ( .A(n45386), .X(n45387) );
  nand_x4_sg U57144 ( .A(n54056), .B(n46340), .X(n28215) );
  inv_x4_sg U57145 ( .A(n28208), .X(n54056) );
  nand_x4_sg U57146 ( .A(n54052), .B(n46344), .X(n28208) );
  inv_x4_sg U57147 ( .A(n28201), .X(n54052) );
  inv_x4_sg U57148 ( .A(n45388), .X(n45389) );
  nand_x4_sg U57149 ( .A(n21544), .B(n45389), .X(n21542) );
  inv_x4_sg U57150 ( .A(n45390), .X(n45391) );
  nand_x4_sg U57151 ( .A(n20774), .B(n45391), .X(n20772) );
  inv_x4_sg U57152 ( .A(n45392), .X(n45393) );
  nand_x4_sg U57153 ( .A(n19999), .B(n45393), .X(n19997) );
  inv_x4_sg U57154 ( .A(n45394), .X(n45395) );
  nand_x4_sg U57155 ( .A(n19230), .B(n45395), .X(n19228) );
  inv_x4_sg U57156 ( .A(n45396), .X(n45397) );
  nand_x4_sg U57157 ( .A(n18454), .B(n45397), .X(n18452) );
  inv_x4_sg U57158 ( .A(n45398), .X(n45399) );
  nand_x4_sg U57159 ( .A(n17685), .B(n45399), .X(n17683) );
  inv_x4_sg U57160 ( .A(n45400), .X(n45401) );
  nand_x4_sg U57161 ( .A(n14564), .B(n45401), .X(n14562) );
  inv_x4_sg U57162 ( .A(n45402), .X(n45403) );
  nand_x4_sg U57163 ( .A(n10672), .B(n45403), .X(n10670) );
  nor_x2_sg U57164 ( .A(n9406), .B(n40790), .X(n25372) );
  nor_x2_sg U57165 ( .A(n9406), .B(n40789), .X(n10265) );
  nand_x4_sg U57166 ( .A(n54044), .B(n46346), .X(n28201) );
  inv_x4_sg U57167 ( .A(n28194), .X(n54044) );
  nor_x2_sg U57168 ( .A(n40792), .B(n8475), .X(n32109) );
  nor_x2_sg U57169 ( .A(n40791), .B(n8775), .X(n24443) );
  nor_x4_sg U57170 ( .A(n46477), .B(n46479), .X(n13534) );
  nand_x4_sg U57171 ( .A(n51263), .B(n46568), .X(n25415) );
  inv_x4_sg U57172 ( .A(n25408), .X(n51263) );
  nor_x2_sg U57173 ( .A(n13540), .B(n13541), .X(n13539) );
  nand_x4_sg U57174 ( .A(n13541), .B(n13540), .X(n13548) );
  nor_x4_sg U57175 ( .A(n13556), .B(n13519), .X(n13541) );
  nand_x4_sg U57176 ( .A(n55192), .B(n46250), .X(n29334) );
  inv_x4_sg U57177 ( .A(n29327), .X(n55192) );
  nand_x4_sg U57178 ( .A(n55185), .B(n46252), .X(n29327) );
  inv_x4_sg U57179 ( .A(n29320), .X(n55185) );
  nand_x4_sg U57180 ( .A(n54908), .B(n46270), .X(n29053) );
  inv_x4_sg U57181 ( .A(n29046), .X(n54908) );
  nand_x4_sg U57182 ( .A(n54901), .B(n46272), .X(n29046) );
  inv_x4_sg U57183 ( .A(n29039), .X(n54901) );
  nand_x4_sg U57184 ( .A(n54624), .B(n46295), .X(n28773) );
  inv_x4_sg U57185 ( .A(n28766), .X(n54624) );
  nand_x4_sg U57186 ( .A(n54617), .B(n46297), .X(n28766) );
  inv_x4_sg U57187 ( .A(n28759), .X(n54617) );
  nand_x4_sg U57188 ( .A(n54340), .B(n46315), .X(n28494) );
  inv_x4_sg U57189 ( .A(n28487), .X(n54340) );
  nand_x4_sg U57190 ( .A(n54333), .B(n46317), .X(n28487) );
  inv_x4_sg U57191 ( .A(n28480), .X(n54333) );
  nand_x4_sg U57192 ( .A(n53775), .B(n46362), .X(n27936) );
  inv_x4_sg U57193 ( .A(n27929), .X(n53775) );
  nand_x4_sg U57194 ( .A(n53768), .B(n46364), .X(n27929) );
  inv_x4_sg U57195 ( .A(n27922), .X(n53768) );
  nand_x4_sg U57196 ( .A(n53497), .B(n46385), .X(n27656) );
  inv_x4_sg U57197 ( .A(n27649), .X(n53497) );
  nand_x4_sg U57198 ( .A(n53488), .B(n46387), .X(n27649) );
  inv_x4_sg U57199 ( .A(n27642), .X(n53488) );
  nand_x4_sg U57200 ( .A(n53218), .B(n46406), .X(n27376) );
  inv_x4_sg U57201 ( .A(n27369), .X(n53218) );
  nand_x4_sg U57202 ( .A(n53210), .B(n46409), .X(n27369) );
  inv_x4_sg U57203 ( .A(n27362), .X(n53210) );
  nand_x4_sg U57204 ( .A(n52939), .B(n46429), .X(n27096) );
  inv_x4_sg U57205 ( .A(n27089), .X(n52939) );
  nand_x4_sg U57206 ( .A(n52930), .B(n46431), .X(n27089) );
  inv_x4_sg U57207 ( .A(n27082), .X(n52930) );
  nand_x4_sg U57208 ( .A(n52659), .B(n46451), .X(n26817) );
  inv_x4_sg U57209 ( .A(n26810), .X(n52659) );
  nand_x4_sg U57210 ( .A(n52651), .B(n46454), .X(n26810) );
  inv_x4_sg U57211 ( .A(n26803), .X(n52651) );
  nand_x4_sg U57212 ( .A(n52382), .B(n46475), .X(n26539) );
  inv_x4_sg U57213 ( .A(n26532), .X(n52382) );
  nand_x4_sg U57214 ( .A(n52374), .B(n46477), .X(n26532) );
  inv_x4_sg U57215 ( .A(n26525), .X(n52374) );
  nand_x4_sg U57216 ( .A(n52105), .B(n46497), .X(n26260) );
  inv_x4_sg U57217 ( .A(n26253), .X(n52105) );
  nand_x4_sg U57218 ( .A(n52096), .B(n46499), .X(n26253) );
  inv_x4_sg U57219 ( .A(n26246), .X(n52096) );
  nand_x4_sg U57220 ( .A(n51830), .B(n46518), .X(n25979) );
  inv_x4_sg U57221 ( .A(n25972), .X(n51830) );
  nand_x4_sg U57222 ( .A(n51822), .B(n46521), .X(n25972) );
  inv_x4_sg U57223 ( .A(n25965), .X(n51822) );
  nand_x4_sg U57224 ( .A(n51548), .B(n46541), .X(n25701) );
  inv_x4_sg U57225 ( .A(n25694), .X(n51548) );
  nand_x4_sg U57226 ( .A(n51539), .B(n46543), .X(n25694) );
  inv_x4_sg U57227 ( .A(n25687), .X(n51539) );
  nand_x4_sg U57228 ( .A(n21729), .B(n55243), .X(n21686) );
  inv_x4_sg U57229 ( .A(n21417), .X(n55243) );
  nand_x4_sg U57230 ( .A(n20184), .B(n54675), .X(n20141) );
  inv_x4_sg U57231 ( .A(n19872), .X(n54675) );
  nand_x4_sg U57232 ( .A(n55177), .B(n46254), .X(n29320) );
  inv_x4_sg U57233 ( .A(n29313), .X(n55177) );
  nand_x4_sg U57234 ( .A(n54893), .B(n46274), .X(n29039) );
  inv_x4_sg U57235 ( .A(n29032), .X(n54893) );
  nand_x4_sg U57236 ( .A(n54609), .B(n46299), .X(n28759) );
  inv_x4_sg U57237 ( .A(n28752), .X(n54609) );
  nand_x4_sg U57238 ( .A(n54325), .B(n46319), .X(n28480) );
  inv_x4_sg U57239 ( .A(n28473), .X(n54325) );
  nand_x4_sg U57240 ( .A(n53760), .B(n46366), .X(n27922) );
  inv_x4_sg U57241 ( .A(n27915), .X(n53760) );
  nand_x4_sg U57242 ( .A(n53482), .B(n46389), .X(n27642) );
  inv_x4_sg U57243 ( .A(n27635), .X(n53482) );
  nand_x4_sg U57244 ( .A(n53202), .B(n46411), .X(n27362) );
  inv_x4_sg U57245 ( .A(n27355), .X(n53202) );
  nand_x4_sg U57246 ( .A(n52924), .B(n46433), .X(n27082) );
  inv_x4_sg U57247 ( .A(n27075), .X(n52924) );
  nand_x4_sg U57248 ( .A(n52643), .B(n46456), .X(n26803) );
  inv_x4_sg U57249 ( .A(n26796), .X(n52643) );
  nand_x4_sg U57250 ( .A(n52367), .B(n46479), .X(n26525) );
  inv_x4_sg U57251 ( .A(n26518), .X(n52367) );
  nand_x4_sg U57252 ( .A(n52090), .B(n46501), .X(n26246) );
  inv_x4_sg U57253 ( .A(n26239), .X(n52090) );
  nand_x4_sg U57254 ( .A(n51814), .B(n46523), .X(n25965) );
  inv_x4_sg U57255 ( .A(n25958), .X(n51814) );
  nand_x4_sg U57256 ( .A(n51532), .B(n46545), .X(n25687) );
  inv_x4_sg U57257 ( .A(n25680), .X(n51532) );
  nand_x4_sg U57258 ( .A(n51256), .B(n46570), .X(n25408) );
  inv_x4_sg U57259 ( .A(n25401), .X(n51256) );
  nor_x1_sg U57260 ( .A(n25081), .B(n25082), .X(n25079) );
  nor_x1_sg U57261 ( .A(n24794), .B(n24795), .X(n24792) );
  nor_x1_sg U57262 ( .A(n9973), .B(n9974), .X(n9971) );
  nor_x1_sg U57263 ( .A(n9686), .B(n9687), .X(n9684) );
  nor_x1_sg U57264 ( .A(n21969), .B(n21970), .X(n21966) );
  inv_x1_sg U57265 ( .A(n15878), .X(n53258) );
  nor_x2_sg U57266 ( .A(n53256), .B(n15892), .X(n15891) );
  inv_x4_sg U57267 ( .A(n15894), .X(n53256) );
  inv_x1_sg U57268 ( .A(n13544), .X(n52423) );
  nor_x2_sg U57269 ( .A(n52421), .B(n13558), .X(n13557) );
  inv_x4_sg U57270 ( .A(n13560), .X(n52421) );
  inv_x1_sg U57271 ( .A(n11983), .X(n51871) );
  nor_x2_sg U57272 ( .A(n51869), .B(n11997), .X(n11996) );
  inv_x4_sg U57273 ( .A(n11999), .X(n51869) );
  inv_x4_sg U57274 ( .A(n45404), .X(n45405) );
  nor_x2_sg U57275 ( .A(n16994), .B(n16995), .X(n16993) );
  inv_x4_sg U57276 ( .A(n45406), .X(n45407) );
  nor_x2_sg U57277 ( .A(n15428), .B(n15429), .X(n15427) );
  inv_x4_sg U57278 ( .A(n45408), .X(n45409) );
  nor_x2_sg U57279 ( .A(n13875), .B(n13876), .X(n13874) );
  nand_x4_sg U57280 ( .A(n13965), .B(n13966), .X(n13876) );
  inv_x4_sg U57281 ( .A(n45410), .X(n45411) );
  nor_x2_sg U57282 ( .A(n13095), .B(n13096), .X(n13094) );
  inv_x4_sg U57283 ( .A(n45412), .X(n45413) );
  nor_x2_sg U57284 ( .A(n11534), .B(n11535), .X(n11533) );
  inv_x4_sg U57285 ( .A(n45414), .X(n45415) );
  nor_x2_sg U57286 ( .A(n21746), .B(n21747), .X(n21745) );
  nand_x4_sg U57287 ( .A(n21835), .B(n55370), .X(n21747) );
  inv_x4_sg U57288 ( .A(n45416), .X(n45417) );
  nor_x2_sg U57289 ( .A(n20201), .B(n20202), .X(n20200) );
  nand_x4_sg U57290 ( .A(n20290), .B(n54802), .X(n20202) );
  nand_x4_sg U57291 ( .A(n16219), .B(n44439), .X(n16217) );
  inv_x4_sg U57292 ( .A(n55781), .X(n45421) );
  inv_x4_sg U57293 ( .A(n28739), .X(n55784) );
  inv_x4_sg U57294 ( .A(n27622), .X(n55785) );
  inv_x4_sg U57295 ( .A(n27342), .X(n55786) );
  inv_x4_sg U57296 ( .A(n18063), .X(n55789) );
  inv_x4_sg U57297 ( .A(n17290), .X(n55791) );
  inv_x4_sg U57298 ( .A(n14942), .X(n55793) );
  inv_x4_sg U57299 ( .A(n21916), .X(n55275) );
  inv_x4_sg U57300 ( .A(n20371), .X(n54707) );
  inv_x4_sg U57301 ( .A(n11039), .X(n51353) );
  inv_x4_sg U57302 ( .A(n15726), .X(n55469) );
  nor_x2_sg U57303 ( .A(n20558), .B(n20559), .X(n20557) );
  nor_x4_sg U57304 ( .A(n42337), .B(n20546), .X(n20559) );
  nor_x2_sg U57305 ( .A(n19014), .B(n19015), .X(n19013) );
  nor_x4_sg U57306 ( .A(n42338), .B(n19002), .X(n19015) );
  nor_x2_sg U57307 ( .A(n17469), .B(n17470), .X(n17468) );
  nor_x4_sg U57308 ( .A(n42339), .B(n17457), .X(n17470) );
  nor_x2_sg U57309 ( .A(n10994), .B(n51337), .X(n11012) );
  inv_x4_sg U57310 ( .A(n10993), .X(n51337) );
  inv_x4_sg U57311 ( .A(n20646), .X(n54971) );
  inv_x4_sg U57312 ( .A(n19102), .X(n54403) );
  inv_x4_sg U57313 ( .A(n17557), .X(n53838) );
  inv_x4_sg U57314 ( .A(n14438), .X(n52711) );
  inv_x4_sg U57315 ( .A(n45422), .X(n45423) );
  inv_x2_sg U57316 ( .A(n45424), .X(n45425) );
  nand_x4_sg U57317 ( .A(n21848), .B(n21849), .X(n21755) );
  inv_x4_sg U57318 ( .A(n45426), .X(n45427) );
  inv_x2_sg U57319 ( .A(n45428), .X(n45429) );
  nand_x4_sg U57320 ( .A(n21077), .B(n21078), .X(n20985) );
  inv_x4_sg U57321 ( .A(n45430), .X(n45431) );
  inv_x2_sg U57322 ( .A(n45432), .X(n45433) );
  nand_x4_sg U57323 ( .A(n20303), .B(n20304), .X(n20210) );
  inv_x4_sg U57324 ( .A(n45434), .X(n45435) );
  inv_x2_sg U57325 ( .A(n45436), .X(n45437) );
  nand_x4_sg U57326 ( .A(n19533), .B(n19534), .X(n19441) );
  inv_x4_sg U57327 ( .A(n45438), .X(n45439) );
  inv_x2_sg U57328 ( .A(n45440), .X(n45441) );
  nand_x4_sg U57329 ( .A(n18757), .B(n18758), .X(n18665) );
  inv_x4_sg U57330 ( .A(n45442), .X(n45443) );
  inv_x2_sg U57331 ( .A(n45444), .X(n45445) );
  nand_x4_sg U57332 ( .A(n17988), .B(n17989), .X(n17896) );
  inv_x4_sg U57333 ( .A(n45446), .X(n45447) );
  inv_x2_sg U57334 ( .A(n45448), .X(n45449) );
  nand_x4_sg U57335 ( .A(n14867), .B(n14868), .X(n14775) );
  inv_x4_sg U57336 ( .A(n45450), .X(n45451) );
  inv_x2_sg U57337 ( .A(n45452), .X(n45453) );
  nand_x4_sg U57338 ( .A(n11755), .B(n11756), .X(n11663) );
  inv_x4_sg U57339 ( .A(n45454), .X(n45455) );
  inv_x4_sg U57340 ( .A(n45456), .X(n45457) );
  inv_x4_sg U57341 ( .A(n45458), .X(n45459) );
  nand_x4_sg U57342 ( .A(n21344), .B(n45459), .X(n21343) );
  inv_x4_sg U57343 ( .A(n45460), .X(n45461) );
  nand_x4_sg U57344 ( .A(n20575), .B(n45461), .X(n20574) );
  inv_x4_sg U57345 ( .A(n45462), .X(n45463) );
  nand_x4_sg U57346 ( .A(n19799), .B(n45463), .X(n19798) );
  inv_x4_sg U57347 ( .A(n45464), .X(n45465) );
  nand_x4_sg U57348 ( .A(n19031), .B(n45465), .X(n19030) );
  nand_x4_sg U57349 ( .A(n44477), .B(n54104), .X(n18247) );
  inv_x4_sg U57350 ( .A(n18255), .X(n54104) );
  inv_x4_sg U57351 ( .A(n45466), .X(n45467) );
  nand_x4_sg U57352 ( .A(n17486), .B(n45467), .X(n17485) );
  inv_x4_sg U57353 ( .A(n45468), .X(n45469) );
  nand_x4_sg U57354 ( .A(n16708), .B(n45469), .X(n16707) );
  inv_x4_sg U57355 ( .A(n45470), .X(n45471) );
  nand_x4_sg U57356 ( .A(n15919), .B(n45471), .X(n15918) );
  inv_x4_sg U57357 ( .A(n45472), .X(n45473) );
  nand_x4_sg U57358 ( .A(n15142), .B(n45473), .X(n15141) );
  inv_x4_sg U57359 ( .A(n45474), .X(n45475) );
  nand_x4_sg U57360 ( .A(n14364), .B(n45475), .X(n14363) );
  inv_x4_sg U57361 ( .A(n45476), .X(n45477) );
  nand_x4_sg U57362 ( .A(n13585), .B(n45477), .X(n13584) );
  inv_x4_sg U57363 ( .A(n45478), .X(n45479) );
  nand_x4_sg U57364 ( .A(n12809), .B(n45479), .X(n12808) );
  inv_x4_sg U57365 ( .A(n45480), .X(n45481) );
  nand_x4_sg U57366 ( .A(n12024), .B(n45481), .X(n12023) );
  inv_x4_sg U57367 ( .A(n45482), .X(n45483) );
  nand_x4_sg U57368 ( .A(n11248), .B(n45483), .X(n11247) );
  inv_x4_sg U57369 ( .A(n45484), .X(n45485) );
  nand_x4_sg U57370 ( .A(n10472), .B(n45485), .X(n10471) );
  inv_x4_sg U57371 ( .A(n45486), .X(n45487) );
  inv_x4_sg U57372 ( .A(n45488), .X(n45489) );
  inv_x4_sg U57373 ( .A(n45490), .X(n45491) );
  inv_x4_sg U57374 ( .A(n45492), .X(n45493) );
  inv_x4_sg U57375 ( .A(n45494), .X(n45495) );
  nor_x4_sg U57376 ( .A(n12174), .B(n46521), .X(n12263) );
  inv_x4_sg U57377 ( .A(n12601), .X(n52057) );
  nor_x4_sg U57378 ( .A(n12482), .B(n46519), .X(n12601) );
  nand_x4_sg U57379 ( .A(n46569), .B(n46574), .X(n10286) );
  inv_x4_sg U57380 ( .A(n32101), .X(n49504) );
  inv_x4_sg U57381 ( .A(n24435), .X(n50363) );
  inv_x4_sg U57382 ( .A(n18776), .X(n54226) );
  nor_x4_sg U57383 ( .A(n18654), .B(n46344), .X(n18776) );
  inv_x4_sg U57384 ( .A(n11773), .X(n51714) );
  nor_x4_sg U57385 ( .A(n11638), .B(n46543), .X(n11773) );
  inv_x4_sg U57386 ( .A(n20803), .X(n54978) );
  inv_x4_sg U57387 ( .A(n19259), .X(n54410) );
  inv_x4_sg U57388 ( .A(n17714), .X(n53845) );
  inv_x4_sg U57389 ( .A(n14593), .X(n52725) );
  inv_x4_sg U57390 ( .A(n11482), .X(n51616) );
  inv_x4_sg U57391 ( .A(n29427), .X(n55451) );
  inv_x4_sg U57392 ( .A(n29145), .X(n55167) );
  inv_x4_sg U57393 ( .A(n28866), .X(n54883) );
  inv_x4_sg U57394 ( .A(n28586), .X(n54599) );
  inv_x4_sg U57395 ( .A(n28308), .X(n54315) );
  inv_x4_sg U57396 ( .A(n28028), .X(n54034) );
  inv_x4_sg U57397 ( .A(n27749), .X(n53750) );
  inv_x4_sg U57398 ( .A(n27468), .X(n53472) );
  inv_x4_sg U57399 ( .A(n27189), .X(n53192) );
  inv_x4_sg U57400 ( .A(n26909), .X(n52914) );
  inv_x4_sg U57401 ( .A(n26632), .X(n52633) );
  inv_x4_sg U57402 ( .A(n26353), .X(n52358) );
  inv_x4_sg U57403 ( .A(n26072), .X(n52080) );
  inv_x4_sg U57404 ( .A(n25793), .X(n51804) );
  nor_x2_sg U57405 ( .A(n55152), .B(n55139), .X(n20865) );
  nor_x2_sg U57406 ( .A(n20470), .B(n55139), .X(n20469) );
  inv_x4_sg U57407 ( .A(n20867), .X(n55139) );
  nor_x2_sg U57408 ( .A(n54584), .B(n54571), .X(n19321) );
  nor_x2_sg U57409 ( .A(n18926), .B(n54571), .X(n18925) );
  inv_x4_sg U57410 ( .A(n19323), .X(n54571) );
  nor_x2_sg U57411 ( .A(n54019), .B(n54006), .X(n17776) );
  nor_x2_sg U57412 ( .A(n17381), .B(n54006), .X(n17380) );
  inv_x4_sg U57413 ( .A(n17778), .X(n54006) );
  nor_x2_sg U57414 ( .A(n52899), .B(n52886), .X(n14655) );
  nor_x2_sg U57415 ( .A(n14262), .B(n52886), .X(n14261) );
  inv_x4_sg U57416 ( .A(n14657), .X(n52886) );
  nor_x2_sg U57417 ( .A(n16461), .B(n53411), .X(n16460) );
  nor_x2_sg U57418 ( .A(n53411), .B(n53394), .X(n16468) );
  inv_x4_sg U57419 ( .A(n16470), .X(n53411) );
  inv_x4_sg U57420 ( .A(n21888), .X(n55389) );
  inv_x4_sg U57421 ( .A(n21117), .X(n55104) );
  inv_x4_sg U57422 ( .A(n20343), .X(n54821) );
  inv_x4_sg U57423 ( .A(n19573), .X(n54536) );
  inv_x4_sg U57424 ( .A(n18028), .X(n53971) );
  inv_x4_sg U57425 ( .A(n14907), .X(n52851) );
  inv_x4_sg U57426 ( .A(n14317), .X(n52658) );
  nor_x4_sg U57427 ( .A(n46454), .B(n46456), .X(n14317) );
  inv_x4_sg U57428 ( .A(n21243), .X(n55423) );
  inv_x4_sg U57429 ( .A(n20471), .X(n55138) );
  inv_x4_sg U57430 ( .A(n19698), .X(n54855) );
  inv_x4_sg U57431 ( .A(n18927), .X(n54570) );
  inv_x4_sg U57432 ( .A(n18153), .X(n54287) );
  inv_x4_sg U57433 ( .A(n17382), .X(n54005) );
  inv_x4_sg U57434 ( .A(n16599), .X(n53724) );
  inv_x4_sg U57435 ( .A(n15033), .X(n53166) );
  inv_x4_sg U57436 ( .A(n14263), .X(n52885) );
  inv_x4_sg U57437 ( .A(n13484), .X(n52607) );
  inv_x4_sg U57438 ( .A(n12700), .X(n52332) );
  inv_x4_sg U57439 ( .A(n11922), .X(n52055) );
  inv_x4_sg U57440 ( .A(n11139), .X(n51775) );
  inv_x4_sg U57441 ( .A(n15959), .X(n53262) );
  inv_x4_sg U57442 ( .A(n11284), .X(n51587) );
  inv_x4_sg U57443 ( .A(n45528), .X(n45529) );
  nand_x4_sg U57444 ( .A(n53531), .B(n53568), .X(n16845) );
  inv_x4_sg U57445 ( .A(n16814), .X(n53568) );
  nand_x4_sg U57446 ( .A(n52973), .B(n53010), .X(n15279) );
  inv_x4_sg U57447 ( .A(n15248), .X(n53010) );
  nand_x4_sg U57448 ( .A(n52451), .B(n52414), .X(n13726) );
  inv_x4_sg U57449 ( .A(n13695), .X(n52451) );
  nand_x4_sg U57450 ( .A(n52139), .B(n52176), .X(n12946) );
  inv_x4_sg U57451 ( .A(n12915), .X(n52176) );
  nand_x4_sg U57452 ( .A(n51862), .B(n51899), .X(n12165) );
  inv_x4_sg U57453 ( .A(n12134), .X(n51899) );
  inv_x4_sg U57454 ( .A(n29589), .X(n55470) );
  inv_x4_sg U57455 ( .A(n45530), .X(n45531) );
  nand_x4_sg U57456 ( .A(n45531), .B(n17237), .X(n17216) );
  inv_x4_sg U57457 ( .A(n45532), .X(n45533) );
  nand_x4_sg U57458 ( .A(n45533), .B(n15671), .X(n15650) );
  inv_x4_sg U57459 ( .A(n45534), .X(n45535) );
  nand_x4_sg U57460 ( .A(n45535), .B(n14118), .X(n14097) );
  inv_x4_sg U57461 ( .A(n45536), .X(n45537) );
  nand_x4_sg U57462 ( .A(n45537), .B(n13338), .X(n13317) );
  inv_x4_sg U57463 ( .A(n21381), .X(n55253) );
  inv_x4_sg U57464 ( .A(n19836), .X(n54685) );
  inv_x4_sg U57465 ( .A(n14401), .X(n52721) );
  inv_x4_sg U57466 ( .A(n10509), .X(n51331) );
  inv_x4_sg U57467 ( .A(n45538), .X(n45539) );
  nor_x2_sg U57468 ( .A(n16841), .B(n16842), .X(n16840) );
  nand_x4_sg U57469 ( .A(n16899), .B(n16900), .X(n16842) );
  inv_x4_sg U57470 ( .A(n45540), .X(n45541) );
  nor_x2_sg U57471 ( .A(n16056), .B(n16057), .X(n16055) );
  inv_x4_sg U57472 ( .A(n45542), .X(n45543) );
  nor_x2_sg U57473 ( .A(n15275), .B(n15276), .X(n15274) );
  nand_x4_sg U57474 ( .A(n15333), .B(n15334), .X(n15276) );
  inv_x4_sg U57475 ( .A(n45544), .X(n45545) );
  nor_x2_sg U57476 ( .A(n13722), .B(n13723), .X(n13721) );
  nand_x4_sg U57477 ( .A(n13780), .B(n13781), .X(n13723) );
  inv_x4_sg U57478 ( .A(n45546), .X(n45547) );
  nor_x2_sg U57479 ( .A(n12942), .B(n12943), .X(n12941) );
  nand_x4_sg U57480 ( .A(n13000), .B(n13001), .X(n12943) );
  inv_x4_sg U57481 ( .A(n45548), .X(n45549) );
  nor_x2_sg U57482 ( .A(n12161), .B(n12162), .X(n12160) );
  inv_x4_sg U57483 ( .A(n45550), .X(n45551) );
  nor_x2_sg U57484 ( .A(n11381), .B(n11382), .X(n11380) );
  nand_x4_sg U57485 ( .A(n11439), .B(n11440), .X(n11382) );
  nor_x4_sg U57486 ( .A(n21398), .B(n21397), .X(n21399) );
  nor_x4_sg U57487 ( .A(n20627), .B(n20626), .X(n20628) );
  nor_x4_sg U57488 ( .A(n19853), .B(n19852), .X(n19854) );
  nor_x4_sg U57489 ( .A(n19083), .B(n19082), .X(n19084) );
  nor_x4_sg U57490 ( .A(n18308), .B(n18307), .X(n18309) );
  nor_x4_sg U57491 ( .A(n17538), .B(n17537), .X(n17539) );
  nor_x4_sg U57492 ( .A(n14418), .B(n14417), .X(n14419) );
  nor_x4_sg U57493 ( .A(n10526), .B(n10525), .X(n10527) );
  nor_x4_sg U57494 ( .A(n54142), .B(n18825), .X(n18397) );
  nor_x4_sg U57495 ( .A(n28346), .B(n28347), .X(n18825) );
  nor_x4_sg U57496 ( .A(n55275), .B(n21915), .X(n21487) );
  nor_x4_sg U57497 ( .A(n29464), .B(n29465), .X(n21915) );
  nor_x4_sg U57498 ( .A(n54707), .B(n20370), .X(n19942) );
  nor_x4_sg U57499 ( .A(n28903), .B(n28904), .X(n20370) );
  nor_x4_sg U57500 ( .A(n51353), .B(n11038), .X(n10615) );
  nor_x4_sg U57501 ( .A(n25551), .B(n25552), .X(n11038) );
  inv_x4_sg U57502 ( .A(n45552), .X(n45553) );
  inv_x4_sg U57503 ( .A(n45553), .X(n54040) );
  inv_x4_sg U57504 ( .A(n45554), .X(n45555) );
  inv_x4_sg U57505 ( .A(n45555), .X(n51810) );
  inv_x4_sg U57506 ( .A(n45556), .X(n45557) );
  inv_x4_sg U57507 ( .A(n45557), .X(n53198) );
  inv_x4_sg U57508 ( .A(n45558), .X(n45559) );
  inv_x4_sg U57509 ( .A(n45559), .X(n54889) );
  inv_x4_sg U57510 ( .A(n45560), .X(n45561) );
  inv_x4_sg U57511 ( .A(n45561), .X(n54321) );
  inv_x4_sg U57512 ( .A(n45562), .X(n45563) );
  inv_x4_sg U57513 ( .A(n45563), .X(n53756) );
  inv_x4_sg U57514 ( .A(n45564), .X(n45565) );
  inv_x4_sg U57515 ( .A(n45565), .X(n53478) );
  inv_x4_sg U57516 ( .A(n45566), .X(n45567) );
  inv_x4_sg U57517 ( .A(n45567), .X(n52920) );
  inv_x4_sg U57518 ( .A(n45568), .X(n45569) );
  inv_x4_sg U57519 ( .A(n45569), .X(n52086) );
  inv_x4_sg U57520 ( .A(n45570), .X(n45571) );
  inv_x4_sg U57521 ( .A(n45571), .X(n51528) );
  inv_x4_sg U57522 ( .A(n45572), .X(n45573) );
  inv_x4_sg U57523 ( .A(n45573), .X(n52639) );
  inv_x4_sg U57524 ( .A(n45574), .X(n45575) );
  inv_x4_sg U57525 ( .A(n45575), .X(n54605) );
  inv_x4_sg U57526 ( .A(n45576), .X(n45577) );
  inv_x4_sg U57527 ( .A(n45577), .X(n55173) );
  inv_x4_sg U57528 ( .A(n45578), .X(n45579) );
  inv_x4_sg U57529 ( .A(n45579), .X(n51252) );
  inv_x4_sg U57530 ( .A(n45580), .X(n45581) );
  nor_x2_sg U57531 ( .A(n46216), .B(n53706), .X(n27729) );
  inv_x4_sg U57532 ( .A(n27727), .X(n53706) );
  nor_x2_sg U57533 ( .A(n46220), .B(n53148), .X(n27169) );
  inv_x4_sg U57534 ( .A(n27167), .X(n53148) );
  nor_x2_sg U57535 ( .A(n46224), .B(n52589), .X(n26612) );
  inv_x4_sg U57536 ( .A(n26610), .X(n52589) );
  nor_x2_sg U57537 ( .A(n46226), .B(n52314), .X(n26333) );
  inv_x4_sg U57538 ( .A(n26331), .X(n52314) );
  nor_x2_sg U57539 ( .A(n46228), .B(n52038), .X(n26052) );
  inv_x4_sg U57540 ( .A(n26050), .X(n52038) );
  inv_x4_sg U57541 ( .A(n21671), .X(n55345) );
  inv_x4_sg U57542 ( .A(n20126), .X(n54777) );
  inv_x4_sg U57543 ( .A(n18580), .X(n54223) );
  inv_x4_sg U57544 ( .A(n14693), .X(n52807) );
  inv_x4_sg U57545 ( .A(n10800), .X(n51419) );
  inv_x4_sg U57546 ( .A(n21726), .X(n55374) );
  nor_x4_sg U57547 ( .A(n21714), .B(n46255), .X(n21726) );
  inv_x4_sg U57548 ( .A(n20957), .X(n55089) );
  nor_x4_sg U57549 ( .A(n20945), .B(n46275), .X(n20957) );
  inv_x4_sg U57550 ( .A(n20181), .X(n54806) );
  nor_x4_sg U57551 ( .A(n20169), .B(n46300), .X(n20181) );
  inv_x4_sg U57552 ( .A(n19413), .X(n54521) );
  nor_x4_sg U57553 ( .A(n19401), .B(n46320), .X(n19413) );
  inv_x4_sg U57554 ( .A(n17868), .X(n53956) );
  nor_x4_sg U57555 ( .A(n17856), .B(n46367), .X(n17868) );
  inv_x4_sg U57556 ( .A(n14747), .X(n52836) );
  nor_x4_sg U57557 ( .A(n14735), .B(n46452), .X(n14747) );
  inv_x4_sg U57558 ( .A(n20903), .X(n55060) );
  inv_x4_sg U57559 ( .A(n19359), .X(n54492) );
  inv_x4_sg U57560 ( .A(n17814), .X(n53927) );
  nor_x2_sg U57561 ( .A(n54257), .B(n54129), .X(n18626) );
  inv_x4_sg U57562 ( .A(n18628), .X(n54257) );
  nor_x2_sg U57563 ( .A(n51464), .B(n51338), .X(n10846) );
  inv_x4_sg U57564 ( .A(n10848), .X(n51464) );
  nor_x2_sg U57565 ( .A(n55392), .B(n55260), .X(n21717) );
  inv_x4_sg U57566 ( .A(n21719), .X(n55392) );
  nor_x2_sg U57567 ( .A(n54824), .B(n54692), .X(n20172) );
  inv_x4_sg U57568 ( .A(n20174), .X(n54824) );
  nor_x2_sg U57569 ( .A(n53590), .B(n16991), .X(n16990) );
  inv_x4_sg U57570 ( .A(n16992), .X(n53590) );
  nor_x2_sg U57571 ( .A(n53032), .B(n15425), .X(n15424) );
  inv_x4_sg U57572 ( .A(n15426), .X(n53032) );
  nor_x2_sg U57573 ( .A(n52475), .B(n13872), .X(n13871) );
  inv_x4_sg U57574 ( .A(n13873), .X(n52475) );
  nor_x2_sg U57575 ( .A(n52198), .B(n13092), .X(n13091) );
  inv_x4_sg U57576 ( .A(n13093), .X(n52198) );
  nor_x2_sg U57577 ( .A(n51642), .B(n11531), .X(n11530) );
  inv_x4_sg U57578 ( .A(n11532), .X(n51642) );
  nor_x2_sg U57579 ( .A(n52026), .B(n51901), .X(n12407) );
  inv_x4_sg U57580 ( .A(n12409), .X(n52026) );
  nor_x4_sg U57581 ( .A(n51354), .B(n46565), .X(n10803) );
  inv_x8_sg U57582 ( .A(n46557), .X(n51354) );
  nor_x4_sg U57583 ( .A(n55276), .B(n46250), .X(n21674) );
  inv_x8_sg U57584 ( .A(n46240), .X(n55276) );
  nor_x4_sg U57585 ( .A(n54708), .B(n46295), .X(n20129) );
  inv_x8_sg U57586 ( .A(n46285), .X(n54708) );
  inv_x4_sg U57587 ( .A(n16485), .X(n53277) );
  nand_x8_sg U57588 ( .A(n53266), .B(n53253), .X(n16485) );
  inv_x4_sg U57589 ( .A(n11810), .X(n51609) );
  nor_x2_sg U57590 ( .A(n49283), .B(n9373), .X(n25304) );
  inv_x4_sg U57591 ( .A(n31871), .X(n49283) );
  nor_x2_sg U57592 ( .A(n49293), .B(n9415), .X(n25329) );
  inv_x4_sg U57593 ( .A(n29912), .X(n49293) );
  nor_x2_sg U57594 ( .A(n50152), .B(n9415), .X(n10221) );
  inv_x4_sg U57595 ( .A(n22247), .X(n50152) );
  nor_x2_sg U57596 ( .A(n50142), .B(n9373), .X(n10198) );
  inv_x4_sg U57597 ( .A(n24205), .X(n50142) );
  inv_x4_sg U57598 ( .A(n32018), .X(n49554) );
  inv_x4_sg U57599 ( .A(n24352), .X(n50413) );
  nor_x2_sg U57600 ( .A(n49289), .B(n9385), .X(n25315) );
  inv_x4_sg U57601 ( .A(n30838), .X(n49289) );
  nor_x2_sg U57602 ( .A(n50148), .B(n9385), .X(n10207) );
  inv_x4_sg U57603 ( .A(n23172), .X(n50148) );
  nor_x4_sg U57604 ( .A(n11703), .B(n46552), .X(n11783) );
  nor_x4_sg U57605 ( .A(n46331), .B(n46340), .X(n18446) );
  nor_x4_sg U57606 ( .A(n46379), .B(n53509), .X(n17033) );
  nor_x4_sg U57607 ( .A(n46400), .B(n46404), .X(n16249) );
  nor_x4_sg U57608 ( .A(n46423), .B(n52951), .X(n15467) );
  nor_x4_sg U57609 ( .A(n46467), .B(n46473), .X(n13914) );
  nor_x4_sg U57610 ( .A(n46491), .B(n52117), .X(n13134) );
  nor_x4_sg U57611 ( .A(n46512), .B(n46516), .X(n12354) );
  nor_x4_sg U57612 ( .A(n50093), .B(n30197), .X(n29628) );
  inv_x4_sg U57613 ( .A(n30200), .X(n50093) );
  nor_x4_sg U57614 ( .A(n30198), .B(n30199), .X(n30197) );
  nor_x4_sg U57615 ( .A(n50952), .B(n22531), .X(n21965) );
  inv_x4_sg U57616 ( .A(n22534), .X(n50952) );
  nor_x4_sg U57617 ( .A(n22532), .B(n22533), .X(n22531) );
  nor_x4_sg U57618 ( .A(n55400), .B(n21545), .X(n21214) );
  inv_x4_sg U57619 ( .A(n21246), .X(n55400) );
  nor_x4_sg U57620 ( .A(n21546), .B(n21547), .X(n21545) );
  nor_x4_sg U57621 ( .A(n55355), .B(n21460), .X(n21206) );
  inv_x4_sg U57622 ( .A(n21250), .X(n55355) );
  nor_x4_sg U57623 ( .A(n21461), .B(n21462), .X(n21460) );
  nor_x4_sg U57624 ( .A(n55114), .B(n20775), .X(n20441) );
  inv_x4_sg U57625 ( .A(n20474), .X(n55114) );
  nor_x4_sg U57626 ( .A(n20776), .B(n20777), .X(n20775) );
  nor_x4_sg U57627 ( .A(n55071), .B(n20690), .X(n20433) );
  inv_x4_sg U57628 ( .A(n20478), .X(n55071) );
  nor_x4_sg U57629 ( .A(n20691), .B(n20692), .X(n20690) );
  nor_x4_sg U57630 ( .A(n54832), .B(n20000), .X(n19669) );
  inv_x4_sg U57631 ( .A(n19701), .X(n54832) );
  nor_x4_sg U57632 ( .A(n20001), .B(n20002), .X(n20000) );
  nor_x4_sg U57633 ( .A(n54787), .B(n19915), .X(n19661) );
  inv_x4_sg U57634 ( .A(n19705), .X(n54787) );
  nor_x4_sg U57635 ( .A(n19916), .B(n19917), .X(n19915) );
  nor_x4_sg U57636 ( .A(n54546), .B(n19231), .X(n18897) );
  inv_x4_sg U57637 ( .A(n18930), .X(n54546) );
  nor_x4_sg U57638 ( .A(n19232), .B(n19233), .X(n19231) );
  nor_x4_sg U57639 ( .A(n54503), .B(n19146), .X(n18889) );
  inv_x4_sg U57640 ( .A(n18934), .X(n54503) );
  nor_x4_sg U57641 ( .A(n19147), .B(n19148), .X(n19146) );
  nor_x4_sg U57642 ( .A(n54265), .B(n18455), .X(n18124) );
  inv_x4_sg U57643 ( .A(n18156), .X(n54265) );
  nor_x4_sg U57644 ( .A(n18456), .B(n18457), .X(n18455) );
  nor_x4_sg U57645 ( .A(n54218), .B(n18370), .X(n18116) );
  inv_x4_sg U57646 ( .A(n18160), .X(n54218) );
  nor_x4_sg U57647 ( .A(n18371), .B(n18372), .X(n18370) );
  nor_x4_sg U57648 ( .A(n53981), .B(n17686), .X(n17352) );
  inv_x4_sg U57649 ( .A(n17385), .X(n53981) );
  nor_x4_sg U57650 ( .A(n17687), .B(n17688), .X(n17686) );
  nor_x4_sg U57651 ( .A(n53938), .B(n17601), .X(n17344) );
  inv_x4_sg U57652 ( .A(n17389), .X(n53938) );
  nor_x4_sg U57653 ( .A(n17602), .B(n17603), .X(n17601) );
  nor_x4_sg U57654 ( .A(n53649), .B(n16825), .X(n16561) );
  inv_x4_sg U57655 ( .A(n16605), .X(n53649) );
  nor_x4_sg U57656 ( .A(n16826), .B(n16827), .X(n16825) );
  nor_x4_sg U57657 ( .A(n53371), .B(n16040), .X(n15779) );
  inv_x4_sg U57658 ( .A(n15823), .X(n53371) );
  nor_x4_sg U57659 ( .A(n16041), .B(n16042), .X(n16040) );
  nor_x4_sg U57660 ( .A(n53091), .B(n15259), .X(n14995) );
  inv_x4_sg U57661 ( .A(n15039), .X(n53091) );
  nor_x4_sg U57662 ( .A(n15260), .B(n15261), .X(n15259) );
  nor_x4_sg U57663 ( .A(n52861), .B(n14565), .X(n14233) );
  inv_x4_sg U57664 ( .A(n14266), .X(n52861) );
  nor_x4_sg U57665 ( .A(n14566), .B(n14567), .X(n14565) );
  nor_x4_sg U57666 ( .A(n52818), .B(n14480), .X(n14225) );
  inv_x4_sg U57667 ( .A(n14270), .X(n52818) );
  nor_x4_sg U57668 ( .A(n14481), .B(n14482), .X(n14480) );
  nor_x4_sg U57669 ( .A(n52533), .B(n13706), .X(n13446) );
  inv_x4_sg U57670 ( .A(n13490), .X(n52533) );
  nor_x4_sg U57671 ( .A(n13707), .B(n13708), .X(n13706) );
  nor_x4_sg U57672 ( .A(n52257), .B(n12926), .X(n12662) );
  inv_x4_sg U57673 ( .A(n12706), .X(n52257) );
  nor_x4_sg U57674 ( .A(n12927), .B(n12928), .X(n12926) );
  nor_x4_sg U57675 ( .A(n51982), .B(n12145), .X(n11884) );
  inv_x4_sg U57676 ( .A(n11928), .X(n51982) );
  nor_x4_sg U57677 ( .A(n12146), .B(n12147), .X(n12145) );
  nor_x4_sg U57678 ( .A(n51701), .B(n11365), .X(n11101) );
  inv_x4_sg U57679 ( .A(n11145), .X(n51701) );
  nor_x4_sg U57680 ( .A(n11366), .B(n11367), .X(n11365) );
  nor_x4_sg U57681 ( .A(n51472), .B(n10673), .X(n10341) );
  inv_x4_sg U57682 ( .A(n10374), .X(n51472) );
  nor_x4_sg U57683 ( .A(n10674), .B(n10675), .X(n10673) );
  nor_x4_sg U57684 ( .A(n51428), .B(n10588), .X(n10333) );
  inv_x4_sg U57685 ( .A(n10378), .X(n51428) );
  nor_x4_sg U57686 ( .A(n10589), .B(n10590), .X(n10588) );
  nor_x4_sg U57687 ( .A(n21796), .B(n46261), .X(n21877) );
  nor_x4_sg U57688 ( .A(n20251), .B(n46306), .X(n20332) );
  nor_x4_sg U57689 ( .A(n53654), .B(n16922), .X(n16910) );
  inv_x4_sg U57690 ( .A(n16916), .X(n53654) );
  nor_x4_sg U57691 ( .A(n16923), .B(n16924), .X(n16922) );
  nor_x4_sg U57692 ( .A(n53374), .B(n16137), .X(n16125) );
  inv_x4_sg U57693 ( .A(n16131), .X(n53374) );
  nor_x4_sg U57694 ( .A(n16138), .B(n16139), .X(n16137) );
  nor_x4_sg U57695 ( .A(n53096), .B(n15356), .X(n15344) );
  inv_x4_sg U57696 ( .A(n15350), .X(n53096) );
  nor_x4_sg U57697 ( .A(n15357), .B(n15358), .X(n15356) );
  nor_x4_sg U57698 ( .A(n52538), .B(n13803), .X(n13791) );
  inv_x4_sg U57699 ( .A(n13797), .X(n52538) );
  nor_x4_sg U57700 ( .A(n13804), .B(n13805), .X(n13803) );
  nor_x4_sg U57701 ( .A(n52262), .B(n13023), .X(n13011) );
  inv_x4_sg U57702 ( .A(n13017), .X(n52262) );
  nor_x4_sg U57703 ( .A(n13024), .B(n13025), .X(n13023) );
  nor_x4_sg U57704 ( .A(n51985), .B(n12242), .X(n12230) );
  inv_x4_sg U57705 ( .A(n12236), .X(n51985) );
  nor_x4_sg U57706 ( .A(n12243), .B(n12244), .X(n12242) );
  nor_x4_sg U57707 ( .A(n51706), .B(n11462), .X(n11450) );
  inv_x4_sg U57708 ( .A(n11456), .X(n51706) );
  nor_x4_sg U57709 ( .A(n11463), .B(n11464), .X(n11462) );
  nor_x4_sg U57710 ( .A(n20613), .B(n46270), .X(n20764) );
  nor_x4_sg U57711 ( .A(n19069), .B(n46315), .X(n19220) );
  nor_x4_sg U57712 ( .A(n17524), .B(n46362), .X(n17675) );
  nor_x4_sg U57713 ( .A(n14411), .B(n46451), .X(n14554) );
  nor_x4_sg U57714 ( .A(n46518), .B(n46512), .X(n12222) );
  nor_x4_sg U57715 ( .A(n46379), .B(n46385), .X(n16902) );
  nor_x4_sg U57716 ( .A(n46423), .B(n46429), .X(n15336) );
  nor_x4_sg U57717 ( .A(n46491), .B(n46497), .X(n13003) );
  nor_x4_sg U57718 ( .A(n46381), .B(n16854), .X(n17234) );
  nor_x4_sg U57719 ( .A(n46425), .B(n15288), .X(n15668) );
  nor_x4_sg U57720 ( .A(n46493), .B(n12955), .X(n13335) );
  nor_x4_sg U57721 ( .A(n18705), .B(n46353), .X(n18786) );
  nor_x4_sg U57722 ( .A(n46331), .B(n46346), .X(n18334) );
  nor_x4_sg U57723 ( .A(n10919), .B(n46573), .X(n10999) );
  nor_x4_sg U57724 ( .A(n46252), .B(n46244), .X(n21485) );
  nor_x4_sg U57725 ( .A(n46297), .B(n46289), .X(n19940) );
  nor_x4_sg U57726 ( .A(n55290), .B(n21437), .X(n21427) );
  inv_x4_sg U57727 ( .A(n21433), .X(n55290) );
  nor_x4_sg U57728 ( .A(n21438), .B(n21439), .X(n21437) );
  nor_x4_sg U57729 ( .A(n54998), .B(n20666), .X(n20656) );
  inv_x4_sg U57730 ( .A(n20662), .X(n54998) );
  nor_x4_sg U57731 ( .A(n20667), .B(n20668), .X(n20666) );
  nor_x4_sg U57732 ( .A(n54722), .B(n19892), .X(n19882) );
  inv_x4_sg U57733 ( .A(n19888), .X(n54722) );
  nor_x4_sg U57734 ( .A(n19893), .B(n19894), .X(n19892) );
  nor_x4_sg U57735 ( .A(n54430), .B(n19122), .X(n19112) );
  inv_x4_sg U57736 ( .A(n19118), .X(n54430) );
  nor_x4_sg U57737 ( .A(n19123), .B(n19124), .X(n19122) );
  nor_x4_sg U57738 ( .A(n54157), .B(n18347), .X(n18337) );
  inv_x4_sg U57739 ( .A(n18343), .X(n54157) );
  nor_x4_sg U57740 ( .A(n18348), .B(n18349), .X(n18347) );
  nor_x4_sg U57741 ( .A(n53865), .B(n17577), .X(n17567) );
  inv_x4_sg U57742 ( .A(n17573), .X(n53865) );
  nor_x4_sg U57743 ( .A(n17578), .B(n17579), .X(n17577) );
  nor_x4_sg U57744 ( .A(n53587), .B(n16795), .X(n16788) );
  inv_x4_sg U57745 ( .A(n16794), .X(n53587) );
  nor_x4_sg U57746 ( .A(n16796), .B(n16797), .X(n16795) );
  nor_x4_sg U57747 ( .A(n53307), .B(n16010), .X(n16003) );
  inv_x4_sg U57748 ( .A(n16009), .X(n53307) );
  nor_x4_sg U57749 ( .A(n16011), .B(n16012), .X(n16010) );
  nor_x4_sg U57750 ( .A(n53029), .B(n15229), .X(n15222) );
  inv_x4_sg U57751 ( .A(n15228), .X(n53029) );
  nor_x4_sg U57752 ( .A(n15230), .B(n15231), .X(n15229) );
  nor_x4_sg U57753 ( .A(n52745), .B(n14457), .X(n14447) );
  inv_x4_sg U57754 ( .A(n14453), .X(n52745) );
  nor_x4_sg U57755 ( .A(n14458), .B(n14459), .X(n14457) );
  nor_x4_sg U57756 ( .A(n52472), .B(n13676), .X(n13669) );
  inv_x4_sg U57757 ( .A(n13675), .X(n52472) );
  nor_x4_sg U57758 ( .A(n13677), .B(n13678), .X(n13676) );
  nor_x4_sg U57759 ( .A(n52195), .B(n12896), .X(n12889) );
  inv_x4_sg U57760 ( .A(n12895), .X(n52195) );
  nor_x4_sg U57761 ( .A(n12897), .B(n12898), .X(n12896) );
  nor_x4_sg U57762 ( .A(n51920), .B(n12115), .X(n12108) );
  inv_x4_sg U57763 ( .A(n12114), .X(n51920) );
  nor_x4_sg U57764 ( .A(n12116), .B(n12117), .X(n12115) );
  nor_x4_sg U57765 ( .A(n51639), .B(n11335), .X(n11328) );
  inv_x4_sg U57766 ( .A(n11334), .X(n51639) );
  nor_x4_sg U57767 ( .A(n11336), .B(n11337), .X(n11335) );
  nor_x4_sg U57768 ( .A(n51368), .B(n10565), .X(n10555) );
  inv_x4_sg U57769 ( .A(n10561), .X(n51368) );
  nor_x4_sg U57770 ( .A(n10566), .B(n10567), .X(n10565) );
  nor_x4_sg U57771 ( .A(n46381), .B(n46389), .X(n16749) );
  nor_x4_sg U57772 ( .A(n46425), .B(n46433), .X(n15183) );
  nor_x4_sg U57773 ( .A(n46493), .B(n46501), .X(n12850) );
  nor_x4_sg U57774 ( .A(n12030), .B(n46523), .X(n12069) );
  nor_x4_sg U57775 ( .A(n46471), .B(n46479), .X(n13630) );
  nor_x4_sg U57776 ( .A(n13735), .B(n46471), .X(n14115) );
  nor_x4_sg U57777 ( .A(n54947), .B(n46272), .X(n20714) );
  nor_x4_sg U57778 ( .A(n54379), .B(n46317), .X(n19170) );
  nor_x4_sg U57779 ( .A(n53814), .B(n46364), .X(n17625) );
  nor_x4_sg U57780 ( .A(n46445), .B(n46454), .X(n14504) );
  nand_x4_sg U57781 ( .A(n11590), .B(n11589), .X(n11595) );
  nor_x4_sg U57782 ( .A(n46535), .B(n46537), .X(n11590) );
  nand_x4_sg U57783 ( .A(n17050), .B(n17049), .X(n17055) );
  nor_x4_sg U57784 ( .A(n17099), .B(n46390), .X(n17049) );
  nand_x4_sg U57785 ( .A(n15484), .B(n15483), .X(n15489) );
  nor_x4_sg U57786 ( .A(n15533), .B(n46434), .X(n15483) );
  nand_x4_sg U57787 ( .A(n13931), .B(n13930), .X(n13936) );
  nor_x4_sg U57788 ( .A(n13980), .B(n46480), .X(n13930) );
  nand_x4_sg U57789 ( .A(n13151), .B(n13150), .X(n13156) );
  nor_x4_sg U57790 ( .A(n13200), .B(n46502), .X(n13150) );
  inv_x4_sg U57791 ( .A(n45582), .X(n45583) );
  nor_x4_sg U57792 ( .A(n49781), .B(n45583), .X(n31162) );
  inv_x4_sg U57793 ( .A(n31352), .X(n49781) );
  inv_x4_sg U57794 ( .A(n45584), .X(n45585) );
  nor_x4_sg U57795 ( .A(n50640), .B(n45585), .X(n23496) );
  inv_x4_sg U57796 ( .A(n23686), .X(n50640) );
  inv_x4_sg U57797 ( .A(n45586), .X(n45587) );
  nor_x4_sg U57798 ( .A(n49598), .B(n45587), .X(n31820) );
  inv_x4_sg U57799 ( .A(n31936), .X(n49598) );
  inv_x4_sg U57800 ( .A(n45588), .X(n45589) );
  nor_x4_sg U57801 ( .A(n50457), .B(n45589), .X(n24154) );
  inv_x4_sg U57802 ( .A(n24270), .X(n50457) );
  inv_x2_sg U57803 ( .A(n16288), .X(n53359) );
  nor_x4_sg U57804 ( .A(n16190), .B(n46409), .X(n16288) );
  nor_x2_sg U57805 ( .A(n49285), .B(n9367), .X(n25303) );
  inv_x4_sg U57806 ( .A(n31593), .X(n49285) );
  nor_x2_sg U57807 ( .A(n50144), .B(n9367), .X(n10195) );
  inv_x4_sg U57808 ( .A(n23927), .X(n50144) );
  nor_x2_sg U57809 ( .A(n49291), .B(n9394), .X(n25319) );
  inv_x4_sg U57810 ( .A(n30339), .X(n49291) );
  nor_x2_sg U57811 ( .A(n50150), .B(n9394), .X(n10211) );
  inv_x4_sg U57812 ( .A(n22673), .X(n50150) );
  nor_x2_sg U57813 ( .A(n50154), .B(n46603), .X(n10208) );
  inv_x4_sg U57814 ( .A(n10226), .X(n50154) );
  nand_x4_sg U57815 ( .A(n21274), .B(n21272), .X(n21279) );
  nor_x4_sg U57816 ( .A(n46250), .B(n46261), .X(n21272) );
  nand_x4_sg U57817 ( .A(n19729), .B(n19727), .X(n19734) );
  nor_x4_sg U57818 ( .A(n46295), .B(n46306), .X(n19727) );
  nand_x4_sg U57819 ( .A(n18183), .B(n18181), .X(n18188) );
  nor_x4_sg U57820 ( .A(n46340), .B(n46353), .X(n18181) );
  nand_x4_sg U57821 ( .A(n14294), .B(n14292), .X(n14299) );
  nor_x4_sg U57822 ( .A(n46451), .B(n46463), .X(n14292) );
  nand_x4_sg U57823 ( .A(n10402), .B(n10400), .X(n10407) );
  nor_x4_sg U57824 ( .A(n46565), .B(n46573), .X(n10400) );
  nor_x2_sg U57825 ( .A(n49295), .B(n46603), .X(n25316) );
  inv_x4_sg U57826 ( .A(n25334), .X(n49295) );
  nor_x4_sg U57827 ( .A(n46406), .B(n46416), .X(n15845) );
  nor_x4_sg U57828 ( .A(n46475), .B(n46485), .X(n13512) );
  nor_x4_sg U57829 ( .A(n46518), .B(n46528), .X(n11950) );
  nand_x4_sg U57830 ( .A(n12369), .B(n12368), .X(n12376) );
  nor_x4_sg U57831 ( .A(n12344), .B(n46519), .X(n12368) );
  nand_x4_sg U57832 ( .A(n16265), .B(n16266), .X(n16271) );
  nor_x4_sg U57833 ( .A(n46400), .B(n15925), .X(n16265) );
  inv_x4_sg U57834 ( .A(n21314), .X(n55210) );
  inv_x4_sg U57835 ( .A(n19769), .X(n54642) );
  inv_x4_sg U57836 ( .A(n14334), .X(n52678) );
  inv_x4_sg U57837 ( .A(n10442), .X(n51288) );
  inv_x4_sg U57838 ( .A(n45590), .X(n45591) );
  nor_x2_sg U57839 ( .A(n13523), .B(n52385), .X(n13520) );
  inv_x2_sg U57840 ( .A(n13523), .X(n52393) );
  nor_x4_sg U57841 ( .A(n45591), .B(n13537), .X(n13523) );
  nor_x4_sg U57842 ( .A(n13538), .B(n46477), .X(n13537) );
  inv_x4_sg U57843 ( .A(n45592), .X(n45593) );
  nor_x2_sg U57844 ( .A(n11962), .B(n51833), .X(n11959) );
  inv_x2_sg U57845 ( .A(n11962), .X(n51841) );
  nor_x4_sg U57846 ( .A(n45593), .B(n11976), .X(n11962) );
  nor_x4_sg U57847 ( .A(n11977), .B(n46521), .X(n11976) );
  inv_x4_sg U57848 ( .A(n45594), .X(n45595) );
  nor_x2_sg U57849 ( .A(n16644), .B(n53501), .X(n16641) );
  inv_x2_sg U57850 ( .A(n16644), .X(n53512) );
  nor_x4_sg U57851 ( .A(n45595), .B(n16657), .X(n16644) );
  nor_x4_sg U57852 ( .A(n16658), .B(n46387), .X(n16657) );
  inv_x4_sg U57853 ( .A(n45596), .X(n45597) );
  nor_x2_sg U57854 ( .A(n15078), .B(n52943), .X(n15075) );
  inv_x2_sg U57855 ( .A(n15078), .X(n52954) );
  nor_x4_sg U57856 ( .A(n45597), .B(n15091), .X(n15078) );
  nor_x4_sg U57857 ( .A(n15092), .B(n46431), .X(n15091) );
  inv_x4_sg U57858 ( .A(n45598), .X(n45599) );
  nor_x2_sg U57859 ( .A(n12745), .B(n52109), .X(n12742) );
  inv_x2_sg U57860 ( .A(n12745), .X(n52120) );
  nor_x4_sg U57861 ( .A(n45599), .B(n12758), .X(n12745) );
  nor_x4_sg U57862 ( .A(n12759), .B(n46499), .X(n12758) );
  inv_x4_sg U57863 ( .A(n45600), .X(n45601) );
  nor_x2_sg U57864 ( .A(n11184), .B(n51552), .X(n11181) );
  inv_x2_sg U57865 ( .A(n11184), .X(n51563) );
  nor_x4_sg U57866 ( .A(n45601), .B(n11197), .X(n11184) );
  nor_x4_sg U57867 ( .A(n11198), .B(n46543), .X(n11197) );
  nor_x2_sg U57868 ( .A(n15729), .B(n53208), .X(n15730) );
  inv_x4_sg U57869 ( .A(n15732), .X(n53208) );
  nor_x2_sg U57870 ( .A(n11834), .B(n51820), .X(n11835) );
  inv_x4_sg U57871 ( .A(n11837), .X(n51820) );
  nor_x2_sg U57872 ( .A(n13396), .B(n52372), .X(n13397) );
  inv_x4_sg U57873 ( .A(n13399), .X(n52372) );
  nor_x2_sg U57874 ( .A(n18066), .B(n43974), .X(n18067) );
  inv_x4_sg U57875 ( .A(n18069), .X(n54050) );
  nor_x2_sg U57876 ( .A(n19611), .B(n54615), .X(n19612) );
  inv_x4_sg U57877 ( .A(n19614), .X(n54615) );
  nor_x2_sg U57878 ( .A(n21156), .B(n55183), .X(n21157) );
  inv_x4_sg U57879 ( .A(n21159), .X(n55183) );
  nor_x2_sg U57880 ( .A(n14175), .B(n43975), .X(n14176) );
  inv_x4_sg U57881 ( .A(n14178), .X(n52649) );
  inv_x4_sg U57882 ( .A(n30343), .X(n49262) );
  nand_x2_sg U57883 ( .A(n49291), .B(n49262), .X(n30584) );
  inv_x4_sg U57884 ( .A(n22677), .X(n50121) );
  nand_x2_sg U57885 ( .A(n50150), .B(n50121), .X(n22918) );
  inv_x4_sg U57886 ( .A(n29916), .X(n49264) );
  nand_x2_sg U57887 ( .A(n49293), .B(n49264), .X(n30063) );
  inv_x4_sg U57888 ( .A(n22251), .X(n50123) );
  nand_x2_sg U57889 ( .A(n50152), .B(n50123), .X(n22398) );
  nand_x2_sg U57890 ( .A(n49283), .B(n49252), .X(n31972) );
  inv_x4_sg U57891 ( .A(n31875), .X(n49252) );
  nand_x2_sg U57892 ( .A(n50142), .B(n50111), .X(n24306) );
  inv_x4_sg U57893 ( .A(n24209), .X(n50111) );
  inv_x4_sg U57894 ( .A(n30842), .X(n49260) );
  nand_x2_sg U57895 ( .A(n49289), .B(n49260), .X(n31047) );
  inv_x4_sg U57896 ( .A(n23176), .X(n50119) );
  nand_x2_sg U57897 ( .A(n50148), .B(n50119), .X(n23381) );
  inv_x4_sg U57898 ( .A(n31597), .X(n49255) );
  nand_x2_sg U57899 ( .A(n49285), .B(n49255), .X(n31731) );
  inv_x4_sg U57900 ( .A(n23931), .X(n50114) );
  nand_x2_sg U57901 ( .A(n50144), .B(n50114), .X(n24065) );
  nand_x4_sg U57902 ( .A(n51671), .B(n51537), .X(n11619) );
  inv_x4_sg U57903 ( .A(n11515), .X(n51671) );
  nand_x4_sg U57904 ( .A(n55307), .B(n21434), .X(n21428) );
  inv_x4_sg U57905 ( .A(n21473), .X(n55307) );
  nand_x4_sg U57906 ( .A(n55025), .B(n20663), .X(n20657) );
  inv_x4_sg U57907 ( .A(n20703), .X(n55025) );
  nand_x4_sg U57908 ( .A(n54739), .B(n19889), .X(n19883) );
  inv_x4_sg U57909 ( .A(n19928), .X(n54739) );
  nand_x4_sg U57910 ( .A(n54457), .B(n19119), .X(n19113) );
  inv_x4_sg U57911 ( .A(n19159), .X(n54457) );
  nand_x4_sg U57912 ( .A(n54173), .B(n18344), .X(n18338) );
  inv_x4_sg U57913 ( .A(n18383), .X(n54173) );
  nand_x4_sg U57914 ( .A(n53892), .B(n17574), .X(n17568) );
  inv_x4_sg U57915 ( .A(n17614), .X(n53892) );
  nand_x4_sg U57916 ( .A(n52772), .B(n14454), .X(n14448) );
  inv_x4_sg U57917 ( .A(n14493), .X(n52772) );
  nand_x4_sg U57918 ( .A(n51385), .B(n10562), .X(n10556) );
  inv_x4_sg U57919 ( .A(n10601), .X(n51385) );
  nor_x4_sg U57920 ( .A(n46385), .B(n46389), .X(n16677) );
  nor_x4_sg U57921 ( .A(n46429), .B(n46433), .X(n15111) );
  nor_x4_sg U57922 ( .A(n46497), .B(n46501), .X(n12778) );
  nor_x4_sg U57923 ( .A(n46541), .B(n46545), .X(n11217) );
  inv_x4_sg U57924 ( .A(n29725), .X(n49265) );
  inv_x4_sg U57925 ( .A(n22060), .X(n50124) );
  inv_x4_sg U57926 ( .A(n30072), .X(n49263) );
  inv_x4_sg U57927 ( .A(n22407), .X(n50122) );
  inv_x4_sg U57928 ( .A(n31982), .X(n49251) );
  inv_x4_sg U57929 ( .A(n31741), .X(n49254) );
  inv_x4_sg U57930 ( .A(n24316), .X(n50110) );
  inv_x4_sg U57931 ( .A(n24075), .X(n50113) );
  inv_x4_sg U57932 ( .A(n30594), .X(n49261) );
  inv_x4_sg U57933 ( .A(n22928), .X(n50120) );
  inv_x4_sg U57934 ( .A(n32070), .X(n49249) );
  inv_x4_sg U57935 ( .A(n24404), .X(n50108) );
  inv_x4_sg U57936 ( .A(n23588), .X(n50117) );
  inv_x4_sg U57937 ( .A(n31254), .X(n49258) );
  inv_x4_sg U57938 ( .A(n31056), .X(n49259) );
  inv_x4_sg U57939 ( .A(n23390), .X(n50118) );
  inv_x4_sg U57940 ( .A(n31435), .X(n49256) );
  inv_x4_sg U57941 ( .A(n23769), .X(n50115) );
  nor_x4_sg U57942 ( .A(n46568), .B(n46570), .X(n10425) );
  inv_x4_sg U57943 ( .A(n10742), .X(n51408) );
  nor_x4_sg U57944 ( .A(n46555), .B(n46566), .X(n10742) );
  inv_x4_sg U57945 ( .A(n24495), .X(n50084) );
  inv_x4_sg U57946 ( .A(n9380), .X(n50943) );
  inv_x4_sg U57947 ( .A(n24511), .X(n50051) );
  inv_x4_sg U57948 ( .A(n24502), .X(n50074) );
  inv_x4_sg U57949 ( .A(n9388), .X(n50933) );
  inv_x4_sg U57950 ( .A(n9400), .X(n50910) );
  inv_x4_sg U57951 ( .A(n21350), .X(n55222) );
  nor_x4_sg U57952 ( .A(n46246), .B(n46254), .X(n21350) );
  inv_x4_sg U57953 ( .A(n19805), .X(n54654) );
  nor_x4_sg U57954 ( .A(n46291), .B(n46299), .X(n19805) );
  inv_x4_sg U57955 ( .A(n14370), .X(n52690) );
  nor_x4_sg U57956 ( .A(n46447), .B(n46456), .X(n14370) );
  inv_x4_sg U57957 ( .A(n10478), .X(n51300) );
  nor_x4_sg U57958 ( .A(n10518), .B(n46570), .X(n10478) );
  nor_x2_sg U57959 ( .A(n40783), .B(n49356), .X(n31266) );
  inv_x4_sg U57960 ( .A(n31267), .X(n49356) );
  inv_x4_sg U57961 ( .A(n31199), .X(n49916) );
  inv_x4_sg U57962 ( .A(n30768), .X(n50004) );
  inv_x4_sg U57963 ( .A(n16634), .X(n53496) );
  nand_x2_sg U57964 ( .A(n16635), .B(n53483), .X(n16634) );
  inv_x4_sg U57965 ( .A(n15068), .X(n52938) );
  nand_x2_sg U57966 ( .A(n15069), .B(n52925), .X(n15068) );
  nor_x2_sg U57967 ( .A(n40784), .B(n50215), .X(n23600) );
  inv_x4_sg U57968 ( .A(n23601), .X(n50215) );
  inv_x4_sg U57969 ( .A(n23533), .X(n50775) );
  inv_x4_sg U57970 ( .A(n23102), .X(n50863) );
  inv_x4_sg U57971 ( .A(n12735), .X(n52104) );
  nand_x2_sg U57972 ( .A(n12736), .B(n52091), .X(n12735) );
  inv_x4_sg U57973 ( .A(n11174), .X(n51547) );
  nand_x2_sg U57974 ( .A(n11175), .B(n51533), .X(n11174) );
  nor_x2_sg U57975 ( .A(n20383), .B(n20386), .X(n20384) );
  nor_x2_sg U57976 ( .A(n18839), .B(n18842), .X(n18840) );
  nor_x2_sg U57977 ( .A(n17294), .B(n17297), .X(n17295) );
  nand_x4_sg U57978 ( .A(n10857), .B(n51446), .X(n11002) );
  nor_x4_sg U57979 ( .A(n10782), .B(n46570), .X(n10857) );
  nor_x4_sg U57980 ( .A(n11638), .B(n46545), .X(n11636) );
  nand_x8_sg U57981 ( .A(n27683), .B(n16854), .X(n27690) );
  nor_x8_sg U57982 ( .A(n27676), .B(n46376), .X(n27683) );
  nand_x8_sg U57983 ( .A(n27123), .B(n15288), .X(n27130) );
  nor_x8_sg U57984 ( .A(n27116), .B(n46420), .X(n27123) );
  nand_x8_sg U57985 ( .A(n26566), .B(n13735), .X(n26573) );
  nor_x8_sg U57986 ( .A(n26559), .B(n52447), .X(n26566) );
  nand_x8_sg U57987 ( .A(n26287), .B(n12955), .X(n26294) );
  nor_x8_sg U57988 ( .A(n26280), .B(n46488), .X(n26287) );
  nand_x8_sg U57989 ( .A(n26006), .B(n12174), .X(n26013) );
  nor_x8_sg U57990 ( .A(n25999), .B(n51896), .X(n26006) );
  nand_x8_sg U57991 ( .A(n25728), .B(n11394), .X(n25735) );
  nor_x8_sg U57992 ( .A(n25721), .B(n46532), .X(n25728) );
  nor_x4_sg U57993 ( .A(n29335), .B(n55215), .X(n29340) );
  nor_x4_sg U57994 ( .A(n28774), .B(n54647), .X(n28779) );
  nor_x4_sg U57995 ( .A(n28216), .B(n54084), .X(n28221) );
  nor_x4_sg U57996 ( .A(n27657), .B(n53525), .X(n27662) );
  nor_x4_sg U57997 ( .A(n27377), .B(n53240), .X(n27382) );
  nor_x4_sg U57998 ( .A(n27097), .B(n52967), .X(n27102) );
  nor_x4_sg U57999 ( .A(n26540), .B(n52406), .X(n26545) );
  nor_x4_sg U58000 ( .A(n26261), .B(n52133), .X(n26266) );
  nor_x4_sg U58001 ( .A(n25980), .B(n51854), .X(n25985) );
  nor_x4_sg U58002 ( .A(n25702), .B(n46536), .X(n25707) );
  nor_x4_sg U58003 ( .A(n25423), .B(n51293), .X(n25428) );
  nor_x4_sg U58004 ( .A(n29054), .B(n54935), .X(n29059) );
  nor_x4_sg U58005 ( .A(n28495), .B(n54367), .X(n28500) );
  nor_x4_sg U58006 ( .A(n27937), .B(n53802), .X(n27942) );
  nor_x4_sg U58007 ( .A(n26818), .B(n52683), .X(n26823) );
  nand_x8_sg U58008 ( .A(n29361), .B(n29371), .X(n29368) );
  nor_x8_sg U58009 ( .A(n29354), .B(n55256), .X(n29361) );
  nand_x8_sg U58010 ( .A(n28800), .B(n28810), .X(n28807) );
  nor_x8_sg U58011 ( .A(n28793), .B(n54688), .X(n28800) );
  nand_x8_sg U58012 ( .A(n28242), .B(n28252), .X(n28249) );
  nor_x8_sg U58013 ( .A(n28235), .B(n54124), .X(n28242) );
  nor_x4_sg U58014 ( .A(n16239), .B(n46411), .X(n16313) );
  inv_x4_sg U58015 ( .A(n16501), .X(n53446) );
  nor_x4_sg U58016 ( .A(n16378), .B(n46407), .X(n16501) );
  inv_x4_sg U58017 ( .A(n45602), .X(n45603) );
  inv_x1_sg U58018 ( .A(n45603), .X(n55452) );
  inv_x4_sg U58019 ( .A(n45604), .X(n45605) );
  inv_x1_sg U58020 ( .A(n45605), .X(n55168) );
  inv_x4_sg U58021 ( .A(n45606), .X(n45607) );
  inv_x1_sg U58022 ( .A(n45607), .X(n54884) );
  inv_x4_sg U58023 ( .A(n45608), .X(n45609) );
  inv_x1_sg U58024 ( .A(n45609), .X(n54600) );
  inv_x4_sg U58025 ( .A(n45610), .X(n45611) );
  inv_x1_sg U58026 ( .A(n45611), .X(n54316) );
  inv_x4_sg U58027 ( .A(n45612), .X(n45613) );
  inv_x1_sg U58028 ( .A(n45613), .X(n54035) );
  inv_x4_sg U58029 ( .A(n45614), .X(n45615) );
  inv_x1_sg U58030 ( .A(n45615), .X(n53751) );
  inv_x4_sg U58031 ( .A(n45616), .X(n45617) );
  inv_x1_sg U58032 ( .A(n45617), .X(n53473) );
  inv_x4_sg U58033 ( .A(n45618), .X(n45619) );
  inv_x1_sg U58034 ( .A(n45619), .X(n53193) );
  inv_x4_sg U58035 ( .A(n45620), .X(n45621) );
  inv_x1_sg U58036 ( .A(n45621), .X(n52915) );
  inv_x4_sg U58037 ( .A(n45622), .X(n45623) );
  inv_x1_sg U58038 ( .A(n45623), .X(n52634) );
  inv_x4_sg U58039 ( .A(n45624), .X(n45625) );
  inv_x1_sg U58040 ( .A(n45625), .X(n52359) );
  inv_x4_sg U58041 ( .A(n45626), .X(n45627) );
  inv_x1_sg U58042 ( .A(n45627), .X(n52081) );
  inv_x4_sg U58043 ( .A(n45628), .X(n45629) );
  inv_x1_sg U58044 ( .A(n45629), .X(n51805) );
  inv_x4_sg U58045 ( .A(n45630), .X(n45631) );
  inv_x1_sg U58046 ( .A(n45631), .X(n51523) );
  inv_x4_sg U58047 ( .A(n45632), .X(n45633) );
  inv_x4_sg U58048 ( .A(n45633), .X(n51069) );
  inv_x4_sg U58049 ( .A(n45634), .X(n45635) );
  inv_x4_sg U58050 ( .A(n45635), .X(n50972) );
  inv_x4_sg U58051 ( .A(n45636), .X(n45637) );
  inv_x4_sg U58052 ( .A(n45637), .X(n51106) );
  inv_x4_sg U58053 ( .A(n45638), .X(n45639) );
  inv_x4_sg U58054 ( .A(n45639), .X(n51010) );
  inv_x4_sg U58055 ( .A(n45640), .X(n45641) );
  inv_x4_sg U58056 ( .A(n45641), .X(n51049) );
  inv_x4_sg U58057 ( .A(n45642), .X(n45643) );
  inv_x4_sg U58058 ( .A(n45643), .X(n51238) );
  inv_x4_sg U58059 ( .A(n45644), .X(n45645) );
  inv_x4_sg U58060 ( .A(n45645), .X(n51200) );
  nor_x4_sg U58061 ( .A(n16514), .B(n16511), .X(n16522) );
  nor_x4_sg U58062 ( .A(n14948), .B(n14945), .X(n14956) );
  nor_x4_sg U58063 ( .A(n12615), .B(n12612), .X(n12623) );
  nor_x4_sg U58064 ( .A(n11054), .B(n11051), .X(n11062) );
  nor_x4_sg U58065 ( .A(n53729), .B(n17288), .X(n17195) );
  nor_x4_sg U58066 ( .A(n27845), .B(n27846), .X(n17288) );
  inv_x4_sg U58067 ( .A(n17289), .X(n53729) );
  nor_x4_sg U58068 ( .A(n53171), .B(n15722), .X(n15629) );
  nor_x4_sg U58069 ( .A(n27287), .B(n27288), .X(n15722) );
  inv_x4_sg U58070 ( .A(n15723), .X(n53171) );
  nor_x4_sg U58071 ( .A(n52612), .B(n14169), .X(n14076) );
  nor_x4_sg U58072 ( .A(n26728), .B(n26729), .X(n14169) );
  inv_x4_sg U58073 ( .A(n14170), .X(n52612) );
  nor_x4_sg U58074 ( .A(n52337), .B(n13389), .X(n13296) );
  nor_x4_sg U58075 ( .A(n26450), .B(n26451), .X(n13389) );
  inv_x4_sg U58076 ( .A(n13390), .X(n52337) );
  nor_x4_sg U58077 ( .A(n52060), .B(n12607), .X(n12515) );
  nor_x4_sg U58078 ( .A(n26171), .B(n26172), .X(n12607) );
  inv_x4_sg U58079 ( .A(n12608), .X(n52060) );
  nor_x4_sg U58080 ( .A(n53449), .B(n16505), .X(n16409) );
  nor_x4_sg U58081 ( .A(n27566), .B(n27567), .X(n16505) );
  inv_x4_sg U58082 ( .A(n16506), .X(n53449) );
  nand_x4_sg U58083 ( .A(n55077), .B(n46280), .X(n20855) );
  inv_x4_sg U58084 ( .A(n20945), .X(n55077) );
  nand_x4_sg U58085 ( .A(n54509), .B(n46325), .X(n19311) );
  inv_x4_sg U58086 ( .A(n19401), .X(n54509) );
  nand_x4_sg U58087 ( .A(n53944), .B(n46372), .X(n17766) );
  inv_x4_sg U58088 ( .A(n17856), .X(n53944) );
  nand_x4_sg U58089 ( .A(n52824), .B(n46462), .X(n14645) );
  inv_x4_sg U58090 ( .A(n14735), .X(n52824) );
  inv_x4_sg U58091 ( .A(n45646), .X(n45647) );
  inv_x1_sg U58092 ( .A(n45647), .X(n55426) );
  inv_x4_sg U58093 ( .A(n45648), .X(n45649) );
  inv_x1_sg U58094 ( .A(n45649), .X(n55406) );
  inv_x4_sg U58095 ( .A(n45650), .X(n45651) );
  inv_x1_sg U58096 ( .A(n45651), .X(n55384) );
  inv_x4_sg U58097 ( .A(n45652), .X(n45653) );
  inv_x1_sg U58098 ( .A(n45653), .X(n55317) );
  inv_x4_sg U58099 ( .A(n45654), .X(n45655) );
  inv_x1_sg U58100 ( .A(n45655), .X(n55297) );
  inv_x4_sg U58101 ( .A(n45656), .X(n45657) );
  inv_x1_sg U58102 ( .A(n45657), .X(n55273) );
  inv_x4_sg U58103 ( .A(n45658), .X(n45659) );
  inv_x1_sg U58104 ( .A(n45659), .X(n55239) );
  inv_x4_sg U58105 ( .A(n45660), .X(n45661) );
  inv_x1_sg U58106 ( .A(n45661), .X(n55141) );
  inv_x4_sg U58107 ( .A(n45662), .X(n45663) );
  inv_x1_sg U58108 ( .A(n45663), .X(n55121) );
  inv_x4_sg U58109 ( .A(n45664), .X(n45665) );
  inv_x1_sg U58110 ( .A(n45665), .X(n55099) );
  inv_x4_sg U58111 ( .A(n45666), .X(n45667) );
  inv_x1_sg U58112 ( .A(n45667), .X(n55057) );
  inv_x4_sg U58113 ( .A(n45668), .X(n45669) );
  inv_x1_sg U58114 ( .A(n45669), .X(n55014) );
  inv_x4_sg U58115 ( .A(n45670), .X(n45671) );
  inv_x1_sg U58116 ( .A(n45671), .X(n54993) );
  inv_x4_sg U58117 ( .A(n45672), .X(n45673) );
  inv_x1_sg U58118 ( .A(n45673), .X(n54958) );
  inv_x4_sg U58119 ( .A(n45674), .X(n45675) );
  inv_x1_sg U58120 ( .A(n45675), .X(n54858) );
  inv_x4_sg U58121 ( .A(n45676), .X(n45677) );
  inv_x1_sg U58122 ( .A(n45677), .X(n54838) );
  inv_x4_sg U58123 ( .A(n45678), .X(n45679) );
  inv_x1_sg U58124 ( .A(n45679), .X(n54816) );
  inv_x4_sg U58125 ( .A(n45680), .X(n45681) );
  inv_x1_sg U58126 ( .A(n45681), .X(n54749) );
  inv_x4_sg U58127 ( .A(n45682), .X(n45683) );
  inv_x1_sg U58128 ( .A(n45683), .X(n54729) );
  inv_x4_sg U58129 ( .A(n45684), .X(n45685) );
  inv_x1_sg U58130 ( .A(n45685), .X(n54705) );
  inv_x4_sg U58131 ( .A(n45686), .X(n45687) );
  inv_x1_sg U58132 ( .A(n45687), .X(n54671) );
  inv_x4_sg U58133 ( .A(n45688), .X(n45689) );
  inv_x1_sg U58134 ( .A(n45689), .X(n54573) );
  inv_x4_sg U58135 ( .A(n45690), .X(n45691) );
  inv_x1_sg U58136 ( .A(n45691), .X(n54553) );
  inv_x4_sg U58137 ( .A(n45692), .X(n45693) );
  inv_x1_sg U58138 ( .A(n45693), .X(n54531) );
  inv_x4_sg U58139 ( .A(n45694), .X(n45695) );
  inv_x1_sg U58140 ( .A(n45695), .X(n54489) );
  inv_x4_sg U58141 ( .A(n45696), .X(n45697) );
  inv_x1_sg U58142 ( .A(n45697), .X(n54446) );
  inv_x4_sg U58143 ( .A(n45698), .X(n45699) );
  inv_x1_sg U58144 ( .A(n45699), .X(n54425) );
  inv_x4_sg U58145 ( .A(n45700), .X(n45701) );
  inv_x1_sg U58146 ( .A(n45701), .X(n54390) );
  inv_x4_sg U58147 ( .A(n45702), .X(n45703) );
  inv_x1_sg U58148 ( .A(n45703), .X(n54290) );
  inv_x4_sg U58149 ( .A(n45704), .X(n45705) );
  inv_x1_sg U58150 ( .A(n45705), .X(n54271) );
  inv_x4_sg U58151 ( .A(n45706), .X(n45707) );
  inv_x1_sg U58152 ( .A(n45707), .X(n54248) );
  inv_x4_sg U58153 ( .A(n45708), .X(n45709) );
  inv_x1_sg U58154 ( .A(n45709), .X(n54227) );
  inv_x4_sg U58155 ( .A(n45710), .X(n45711) );
  inv_x1_sg U58156 ( .A(n45711), .X(n54207) );
  inv_x4_sg U58157 ( .A(n45712), .X(n45713) );
  inv_x1_sg U58158 ( .A(n45713), .X(n54182) );
  inv_x4_sg U58159 ( .A(n45714), .X(n45715) );
  inv_x1_sg U58160 ( .A(n45715), .X(n54163) );
  inv_x4_sg U58161 ( .A(n45716), .X(n45717) );
  inv_x1_sg U58162 ( .A(n45717), .X(n54140) );
  inv_x4_sg U58163 ( .A(n45718), .X(n45719) );
  inv_x1_sg U58164 ( .A(n45719), .X(n54107) );
  inv_x4_sg U58165 ( .A(n45720), .X(n45721) );
  inv_x1_sg U58166 ( .A(n45721), .X(n54008) );
  inv_x4_sg U58167 ( .A(n45722), .X(n45723) );
  inv_x1_sg U58168 ( .A(n45723), .X(n53988) );
  inv_x4_sg U58169 ( .A(n45724), .X(n45725) );
  inv_x1_sg U58170 ( .A(n45725), .X(n53966) );
  inv_x4_sg U58171 ( .A(n45726), .X(n45727) );
  inv_x1_sg U58172 ( .A(n45727), .X(n53924) );
  inv_x4_sg U58173 ( .A(n45728), .X(n45729) );
  inv_x1_sg U58174 ( .A(n45729), .X(n53881) );
  inv_x4_sg U58175 ( .A(n45730), .X(n45731) );
  inv_x1_sg U58176 ( .A(n45731), .X(n53860) );
  inv_x4_sg U58177 ( .A(n45732), .X(n45733) );
  inv_x1_sg U58178 ( .A(n45733), .X(n53825) );
  inv_x4_sg U58179 ( .A(n45734), .X(n45735) );
  inv_x1_sg U58180 ( .A(n45735), .X(n53727) );
  inv_x4_sg U58181 ( .A(n45736), .X(n45737) );
  inv_x1_sg U58182 ( .A(n45737), .X(n53708) );
  inv_x4_sg U58183 ( .A(n45738), .X(n45739) );
  inv_x1_sg U58184 ( .A(n45739), .X(n53683) );
  inv_x4_sg U58185 ( .A(n45740), .X(n45741) );
  inv_x1_sg U58186 ( .A(n45741), .X(n53661) );
  inv_x4_sg U58187 ( .A(n45742), .X(n45743) );
  inv_x1_sg U58188 ( .A(n45743), .X(n53617) );
  inv_x4_sg U58189 ( .A(n45744), .X(n45745) );
  inv_x1_sg U58190 ( .A(n45745), .X(n53577) );
  inv_x4_sg U58191 ( .A(n45746), .X(n45747) );
  inv_x1_sg U58192 ( .A(n45747), .X(n53546) );
  inv_x4_sg U58193 ( .A(n45748), .X(n45749) );
  inv_x1_sg U58194 ( .A(n45749), .X(n53447) );
  inv_x4_sg U58195 ( .A(n45750), .X(n45751) );
  inv_x1_sg U58196 ( .A(n45751), .X(n53428) );
  inv_x4_sg U58197 ( .A(n45752), .X(n45753) );
  inv_x1_sg U58198 ( .A(n45753), .X(n53406) );
  inv_x4_sg U58199 ( .A(n45754), .X(n45755) );
  inv_x1_sg U58200 ( .A(n45755), .X(n53382) );
  inv_x4_sg U58201 ( .A(n45756), .X(n45757) );
  inv_x1_sg U58202 ( .A(n45757), .X(n53338) );
  inv_x4_sg U58203 ( .A(n45758), .X(n45759) );
  inv_x1_sg U58204 ( .A(n45759), .X(n53317) );
  inv_x4_sg U58205 ( .A(n45760), .X(n45761) );
  inv_x1_sg U58206 ( .A(n45761), .X(n53296) );
  inv_x4_sg U58207 ( .A(n45762), .X(n45763) );
  inv_x1_sg U58208 ( .A(n45763), .X(n53264) );
  inv_x4_sg U58209 ( .A(n45764), .X(n45765) );
  inv_x1_sg U58210 ( .A(n45765), .X(n53169) );
  inv_x4_sg U58211 ( .A(n45766), .X(n45767) );
  inv_x1_sg U58212 ( .A(n45767), .X(n53150) );
  inv_x4_sg U58213 ( .A(n45768), .X(n45769) );
  inv_x1_sg U58214 ( .A(n45769), .X(n53125) );
  inv_x4_sg U58215 ( .A(n45770), .X(n45771) );
  inv_x1_sg U58216 ( .A(n45771), .X(n53103) );
  inv_x4_sg U58217 ( .A(n45772), .X(n45773) );
  inv_x1_sg U58218 ( .A(n45773), .X(n53059) );
  inv_x4_sg U58219 ( .A(n45774), .X(n45775) );
  inv_x1_sg U58220 ( .A(n45775), .X(n53019) );
  inv_x4_sg U58221 ( .A(n45776), .X(n45777) );
  inv_x1_sg U58222 ( .A(n45777), .X(n52988) );
  inv_x4_sg U58223 ( .A(n45778), .X(n45779) );
  inv_x1_sg U58224 ( .A(n45779), .X(n52888) );
  inv_x4_sg U58225 ( .A(n45780), .X(n45781) );
  inv_x1_sg U58226 ( .A(n45781), .X(n52868) );
  inv_x4_sg U58227 ( .A(n45782), .X(n45783) );
  inv_x1_sg U58228 ( .A(n45783), .X(n52846) );
  inv_x4_sg U58229 ( .A(n45784), .X(n45785) );
  inv_x1_sg U58230 ( .A(n45785), .X(n52804) );
  inv_x4_sg U58231 ( .A(n45786), .X(n45787) );
  inv_x1_sg U58232 ( .A(n45787), .X(n52761) );
  inv_x4_sg U58233 ( .A(n45788), .X(n45789) );
  inv_x1_sg U58234 ( .A(n45789), .X(n52740) );
  inv_x4_sg U58235 ( .A(n45790), .X(n45791) );
  inv_x1_sg U58236 ( .A(n45791), .X(n52705) );
  inv_x4_sg U58237 ( .A(n45792), .X(n45793) );
  inv_x1_sg U58238 ( .A(n45793), .X(n52610) );
  inv_x4_sg U58239 ( .A(n45794), .X(n45795) );
  inv_x1_sg U58240 ( .A(n45795), .X(n52591) );
  inv_x4_sg U58241 ( .A(n45796), .X(n45797) );
  inv_x1_sg U58242 ( .A(n45797), .X(n52566) );
  inv_x4_sg U58243 ( .A(n45798), .X(n45799) );
  inv_x1_sg U58244 ( .A(n45799), .X(n52544) );
  inv_x4_sg U58245 ( .A(n45800), .X(n45801) );
  inv_x1_sg U58246 ( .A(n45801), .X(n52502) );
  inv_x4_sg U58247 ( .A(n45802), .X(n45803) );
  inv_x1_sg U58248 ( .A(n45803), .X(n52461) );
  inv_x4_sg U58249 ( .A(n45804), .X(n45805) );
  inv_x1_sg U58250 ( .A(n45805), .X(n52428) );
  inv_x4_sg U58251 ( .A(n45806), .X(n45807) );
  inv_x1_sg U58252 ( .A(n45807), .X(n52335) );
  inv_x4_sg U58253 ( .A(n45808), .X(n45809) );
  inv_x1_sg U58254 ( .A(n45809), .X(n52316) );
  inv_x4_sg U58255 ( .A(n45810), .X(n45811) );
  inv_x1_sg U58256 ( .A(n45811), .X(n52291) );
  inv_x4_sg U58257 ( .A(n45812), .X(n45813) );
  inv_x1_sg U58258 ( .A(n45813), .X(n52269) );
  inv_x4_sg U58259 ( .A(n45814), .X(n45815) );
  inv_x1_sg U58260 ( .A(n45815), .X(n52225) );
  inv_x4_sg U58261 ( .A(n45816), .X(n45817) );
  inv_x1_sg U58262 ( .A(n45817), .X(n52185) );
  inv_x4_sg U58263 ( .A(n45818), .X(n45819) );
  inv_x1_sg U58264 ( .A(n45819), .X(n52154) );
  inv_x4_sg U58265 ( .A(n45820), .X(n45821) );
  inv_x1_sg U58266 ( .A(n45821), .X(n52058) );
  inv_x4_sg U58267 ( .A(n45822), .X(n45823) );
  inv_x1_sg U58268 ( .A(n45823), .X(n52040) );
  inv_x4_sg U58269 ( .A(n45824), .X(n45825) );
  inv_x1_sg U58270 ( .A(n45825), .X(n52015) );
  inv_x4_sg U58271 ( .A(n45826), .X(n45827) );
  inv_x1_sg U58272 ( .A(n45827), .X(n51993) );
  inv_x4_sg U58273 ( .A(n45828), .X(n45829) );
  inv_x1_sg U58274 ( .A(n45829), .X(n51950) );
  inv_x4_sg U58275 ( .A(n45830), .X(n45831) );
  inv_x1_sg U58276 ( .A(n45831), .X(n51929) );
  inv_x4_sg U58277 ( .A(n45832), .X(n45833) );
  inv_x1_sg U58278 ( .A(n45833), .X(n51909) );
  inv_x4_sg U58279 ( .A(n45834), .X(n45835) );
  inv_x1_sg U58280 ( .A(n45835), .X(n51877) );
  inv_x4_sg U58281 ( .A(n45836), .X(n45837) );
  inv_x1_sg U58282 ( .A(n45837), .X(n51778) );
  inv_x4_sg U58283 ( .A(n45838), .X(n45839) );
  inv_x1_sg U58284 ( .A(n45839), .X(n51759) );
  inv_x4_sg U58285 ( .A(n45840), .X(n45841) );
  inv_x1_sg U58286 ( .A(n45841), .X(n51736) );
  inv_x4_sg U58287 ( .A(n45842), .X(n45843) );
  inv_x1_sg U58288 ( .A(n45843), .X(n51715) );
  inv_x4_sg U58289 ( .A(n45844), .X(n45845) );
  inv_x1_sg U58290 ( .A(n45845), .X(n51669) );
  inv_x4_sg U58291 ( .A(n45846), .X(n45847) );
  inv_x1_sg U58292 ( .A(n45847), .X(n51648) );
  inv_x4_sg U58293 ( .A(n45848), .X(n45849) );
  inv_x1_sg U58294 ( .A(n45849), .X(n51628) );
  inv_x4_sg U58295 ( .A(n45850), .X(n45851) );
  inv_x1_sg U58296 ( .A(n45851), .X(n51596) );
  inv_x4_sg U58297 ( .A(n45852), .X(n45853) );
  inv_x1_sg U58298 ( .A(n45853), .X(n51456) );
  inv_x4_sg U58299 ( .A(n45854), .X(n45855) );
  inv_x1_sg U58300 ( .A(n45855), .X(n51433) );
  inv_x4_sg U58301 ( .A(n45856), .X(n45857) );
  inv_x1_sg U58302 ( .A(n45857), .X(n51394) );
  inv_x4_sg U58303 ( .A(n45858), .X(n45859) );
  inv_x1_sg U58304 ( .A(n45859), .X(n51375) );
  inv_x4_sg U58305 ( .A(n45860), .X(n45861) );
  inv_x1_sg U58306 ( .A(n45861), .X(n51351) );
  inv_x4_sg U58307 ( .A(n45862), .X(n45863) );
  inv_x1_sg U58308 ( .A(n45863), .X(n51317) );
  inv_x4_sg U58309 ( .A(n45864), .X(n45865) );
  inv_x1_sg U58310 ( .A(n45865), .X(n51499) );
  inv_x4_sg U58311 ( .A(n45866), .X(n45867) );
  inv_x1_sg U58312 ( .A(n45867), .X(n52822) );
  inv_x4_sg U58313 ( .A(n45868), .X(n45869) );
  inv_x1_sg U58314 ( .A(n45869), .X(n55075) );
  inv_x4_sg U58315 ( .A(n45870), .X(n45871) );
  inv_x1_sg U58316 ( .A(n45871), .X(n54507) );
  inv_x4_sg U58317 ( .A(n45872), .X(n45873) );
  inv_x1_sg U58318 ( .A(n45873), .X(n53942) );
  inv_x4_sg U58319 ( .A(n45874), .X(n45875) );
  inv_x1_sg U58320 ( .A(n45875), .X(n52481) );
  inv_x4_sg U58321 ( .A(n45876), .X(n45877) );
  inv_x1_sg U58322 ( .A(n45877), .X(n53596) );
  inv_x4_sg U58323 ( .A(n45878), .X(n45879) );
  inv_x1_sg U58324 ( .A(n45879), .X(n53038) );
  inv_x4_sg U58325 ( .A(n45880), .X(n45881) );
  inv_x1_sg U58326 ( .A(n45881), .X(n52204) );
  inv_x4_sg U58327 ( .A(n45882), .X(n45883) );
  inv_x1_sg U58328 ( .A(n45883), .X(n51479) );
  inv_x4_sg U58329 ( .A(n45884), .X(n45885) );
  inv_x1_sg U58330 ( .A(n45885), .X(n51691) );
  inv_x4_sg U58331 ( .A(n45886), .X(n45887) );
  inv_x1_sg U58332 ( .A(n45887), .X(n55342) );
  inv_x4_sg U58333 ( .A(n45888), .X(n45889) );
  inv_x1_sg U58334 ( .A(n45889), .X(n54774) );
  inv_x4_sg U58335 ( .A(n45890), .X(n45891) );
  inv_x1_sg U58336 ( .A(n45891), .X(n51972) );
  inv_x4_sg U58337 ( .A(n45892), .X(n45893) );
  inv_x1_sg U58338 ( .A(n45893), .X(n55360) );
  inv_x4_sg U58339 ( .A(n45894), .X(n45895) );
  inv_x1_sg U58340 ( .A(n45895), .X(n54792) );
  inv_x4_sg U58341 ( .A(n45896), .X(n45897) );
  inv_x1_sg U58342 ( .A(n45897), .X(n51613) );
  inv_x4_sg U58343 ( .A(n45898), .X(n45899) );
  inv_x1_sg U58344 ( .A(n45899), .X(n53361) );
  inv_x4_sg U58345 ( .A(n45900), .X(n45901) );
  inv_x1_sg U58346 ( .A(n45901), .X(n52523) );
  inv_x4_sg U58347 ( .A(n45902), .X(n45903) );
  inv_x1_sg U58348 ( .A(n45903), .X(n53563) );
  inv_x4_sg U58349 ( .A(n45904), .X(n45905) );
  inv_x1_sg U58350 ( .A(n45905), .X(n53005) );
  inv_x4_sg U58351 ( .A(n45906), .X(n45907) );
  inv_x1_sg U58352 ( .A(n45907), .X(n52171) );
  inv_x4_sg U58353 ( .A(n45908), .X(n45909) );
  inv_x1_sg U58354 ( .A(n45909), .X(n52445) );
  inv_x4_sg U58355 ( .A(n45910), .X(n45911) );
  inv_x1_sg U58356 ( .A(n45911), .X(n51894) );
  inv_x4_sg U58357 ( .A(n45912), .X(n45913) );
  inv_x1_sg U58358 ( .A(n45913), .X(n53639) );
  inv_x4_sg U58359 ( .A(n45914), .X(n45915) );
  inv_x1_sg U58360 ( .A(n45915), .X(n53081) );
  inv_x4_sg U58361 ( .A(n45916), .X(n45917) );
  inv_x1_sg U58362 ( .A(n45917), .X(n52247) );
  inv_x4_sg U58363 ( .A(n45918), .X(n45919) );
  inv_x1_sg U58364 ( .A(n45919), .X(n53280) );
  inv_x4_sg U58365 ( .A(n45920), .X(n45921) );
  inv_x1_sg U58366 ( .A(n45921), .X(n51416) );
  inv_x4_sg U58367 ( .A(n45922), .X(n45923) );
  inv_x1_sg U58368 ( .A(n45923), .X(n52781) );
  inv_x4_sg U58369 ( .A(n45924), .X(n45925) );
  inv_x1_sg U58370 ( .A(n45925), .X(n55034) );
  inv_x4_sg U58371 ( .A(n45926), .X(n45927) );
  inv_x1_sg U58372 ( .A(n45927), .X(n54466) );
  inv_x4_sg U58373 ( .A(n45928), .X(n45929) );
  inv_x1_sg U58374 ( .A(n45929), .X(n53901) );
  inv_x4_sg U58375 ( .A(n45930), .X(n45931) );
  inv_x1_sg U58376 ( .A(n45931), .X(n54975) );
  inv_x4_sg U58377 ( .A(n45932), .X(n45933) );
  inv_x1_sg U58378 ( .A(n45933), .X(n54407) );
  inv_x4_sg U58379 ( .A(n45934), .X(n45935) );
  inv_x1_sg U58380 ( .A(n45935), .X(n53842) );
  inv_x4_sg U58381 ( .A(n45936), .X(n45937) );
  inv_x1_sg U58382 ( .A(n45937), .X(n52722) );
  inv_x4_sg U58383 ( .A(n45938), .X(n45939) );
  inv_x1_sg U58384 ( .A(n45939), .X(n54122) );
  inv_x4_sg U58385 ( .A(n45940), .X(n45941) );
  inv_x1_sg U58386 ( .A(n45941), .X(n55254) );
  inv_x4_sg U58387 ( .A(n45942), .X(n45943) );
  inv_x1_sg U58388 ( .A(n45943), .X(n54686) );
  inv_x4_sg U58389 ( .A(n45944), .X(n45945) );
  inv_x1_sg U58390 ( .A(n45945), .X(n51332) );
  inv_x4_sg U58391 ( .A(n45946), .X(n45947) );
  nor_x4_sg U58392 ( .A(n55428), .B(n21923), .X(n21828) );
  nor_x4_sg U58393 ( .A(n29523), .B(n29524), .X(n21923) );
  inv_x4_sg U58394 ( .A(n21924), .X(n55428) );
  nor_x4_sg U58395 ( .A(n55143), .B(n21150), .X(n21057) );
  nor_x4_sg U58396 ( .A(n29245), .B(n29246), .X(n21150) );
  inv_x4_sg U58397 ( .A(n21151), .X(n55143) );
  nor_x4_sg U58398 ( .A(n54860), .B(n20378), .X(n20283) );
  nor_x4_sg U58399 ( .A(n28962), .B(n28963), .X(n20378) );
  inv_x4_sg U58400 ( .A(n20379), .X(n54860) );
  nor_x4_sg U58401 ( .A(n54575), .B(n19606), .X(n19513) );
  nor_x4_sg U58402 ( .A(n28684), .B(n28685), .X(n19606) );
  inv_x4_sg U58403 ( .A(n19607), .X(n54575) );
  nor_x4_sg U58404 ( .A(n54292), .B(n18833), .X(n18737) );
  nor_x4_sg U58405 ( .A(n28405), .B(n28406), .X(n18833) );
  inv_x4_sg U58406 ( .A(n18834), .X(n54292) );
  nor_x4_sg U58407 ( .A(n54010), .B(n18061), .X(n17968) );
  nor_x4_sg U58408 ( .A(n28126), .B(n28127), .X(n18061) );
  inv_x4_sg U58409 ( .A(n18062), .X(n54010) );
  nor_x4_sg U58410 ( .A(n52890), .B(n14940), .X(n14847) );
  nor_x4_sg U58411 ( .A(n27007), .B(n27008), .X(n14940) );
  inv_x4_sg U58412 ( .A(n14941), .X(n52890) );
  nor_x4_sg U58413 ( .A(n51780), .B(n11828), .X(n11735) );
  nor_x4_sg U58414 ( .A(n25891), .B(n25892), .X(n11828) );
  inv_x4_sg U58415 ( .A(n11829), .X(n51780) );
  nor_x4_sg U58416 ( .A(n51501), .B(n11044), .X(n10951) );
  nor_x4_sg U58417 ( .A(n25610), .B(n25611), .X(n11044) );
  inv_x4_sg U58418 ( .A(n11045), .X(n51501) );
  inv_x4_sg U58419 ( .A(n40999), .X(n45948) );
  inv_x4_sg U58420 ( .A(n40929), .X(n45950) );
  inv_x4_sg U58421 ( .A(n41027), .X(n45952) );
  inv_x4_sg U58422 ( .A(n41009), .X(n45954) );
  inv_x4_sg U58423 ( .A(n40993), .X(n45956) );
  inv_x4_sg U58424 ( .A(n40975), .X(n45958) );
  inv_x4_sg U58425 ( .A(n40987), .X(n45960) );
  inv_x4_sg U58426 ( .A(n40969), .X(n45962) );
  inv_x4_sg U58427 ( .A(n40941), .X(n45964) );
  inv_x4_sg U58428 ( .A(n40923), .X(n45966) );
  inv_x4_sg U58429 ( .A(n41015), .X(n45968) );
  inv_x4_sg U58430 ( .A(n40957), .X(n45970) );
  inv_x4_sg U58431 ( .A(n41033), .X(n45972) );
  inv_x4_sg U58432 ( .A(n40911), .X(n45974) );
  nor_x8_sg U58433 ( .A(n46252), .B(n46248), .X(n21290) );
  nor_x8_sg U58434 ( .A(n46297), .B(n46293), .X(n19745) );
  nor_x8_sg U58435 ( .A(n54921), .B(n46272), .X(n20520) );
  nor_x8_sg U58436 ( .A(n54353), .B(n46317), .X(n18976) );
  nor_x8_sg U58437 ( .A(n53788), .B(n46364), .X(n17431) );
  nor_x8_sg U58438 ( .A(n46568), .B(n46563), .X(n10418) );
  nand_x4_sg U58439 ( .A(n11321), .B(n11191), .X(n11284) );
  nor_x8_sg U58440 ( .A(n51560), .B(n46543), .X(n11191) );
  nor_x8_sg U58441 ( .A(n46337), .B(n46344), .X(n18198) );
  nand_x4_sg U58442 ( .A(n15996), .B(n15864), .X(n15959) );
  nor_x8_sg U58443 ( .A(n46409), .B(n46404), .X(n15864) );
  nor_x8_sg U58444 ( .A(n46449), .B(n46454), .X(n14310) );
  nand_x4_sg U58445 ( .A(n51952), .B(n51819), .X(n12400) );
  nand_x4_sg U58446 ( .A(n53619), .B(n46388), .X(n17079) );
  nand_x4_sg U58447 ( .A(n53061), .B(n46432), .X(n15513) );
  nand_x4_sg U58448 ( .A(n52227), .B(n46500), .X(n13180) );
  nand_x4_sg U58449 ( .A(n52504), .B(n46478), .X(n13960) );
  nand_x4_sg U58450 ( .A(n55036), .B(n54898), .X(n20941) );
  nand_x4_sg U58451 ( .A(n55036), .B(n46269), .X(n21125) );
  inv_x8_sg U58452 ( .A(n20837), .X(n55036) );
  nand_x4_sg U58453 ( .A(n54468), .B(n54330), .X(n19397) );
  nand_x4_sg U58454 ( .A(n54468), .B(n46314), .X(n19581) );
  inv_x8_sg U58455 ( .A(n19293), .X(n54468) );
  nand_x4_sg U58456 ( .A(n53903), .B(n53765), .X(n17852) );
  nand_x4_sg U58457 ( .A(n53903), .B(n46361), .X(n18036) );
  inv_x8_sg U58458 ( .A(n17748), .X(n53903) );
  nand_x4_sg U58459 ( .A(n52783), .B(n52648), .X(n14731) );
  nand_x4_sg U58460 ( .A(n52783), .B(n46450), .X(n14915) );
  inv_x8_sg U58461 ( .A(n14627), .X(n52783) );
  inv_x4_sg U58462 ( .A(n45976), .X(n45977) );
  inv_x1_sg U58463 ( .A(n45977), .X(n54945) );
  inv_x4_sg U58464 ( .A(n45978), .X(n45979) );
  inv_x1_sg U58465 ( .A(n45979), .X(n54377) );
  inv_x4_sg U58466 ( .A(n45980), .X(n45981) );
  inv_x1_sg U58467 ( .A(n45981), .X(n53812) );
  inv_x4_sg U58468 ( .A(n45982), .X(n45983) );
  inv_x4_sg U58469 ( .A(n45984), .X(n45985) );
  inv_x4_sg U58470 ( .A(n45986), .X(n45987) );
  inv_x4_sg U58471 ( .A(n45988), .X(n45989) );
  inv_x1_sg U58472 ( .A(n45989), .X(n54919) );
  inv_x4_sg U58473 ( .A(n45990), .X(n45991) );
  inv_x1_sg U58474 ( .A(n45991), .X(n54351) );
  inv_x4_sg U58475 ( .A(n45992), .X(n45993) );
  inv_x1_sg U58476 ( .A(n45993), .X(n53786) );
  inv_x4_sg U58477 ( .A(n45994), .X(n45995) );
  inv_x1_sg U58478 ( .A(n45995), .X(n53507) );
  inv_x4_sg U58479 ( .A(n45996), .X(n45997) );
  inv_x1_sg U58480 ( .A(n45997), .X(n52949) );
  inv_x4_sg U58481 ( .A(n45998), .X(n45999) );
  inv_x1_sg U58482 ( .A(n45999), .X(n52115) );
  inv_x4_sg U58483 ( .A(n46000), .X(n46001) );
  inv_x4_sg U58484 ( .A(n46002), .X(n46003) );
  inv_x4_sg U58485 ( .A(n46004), .X(n46005) );
  inv_x4_sg U58486 ( .A(n46006), .X(n46007) );
  inv_x4_sg U58487 ( .A(n46008), .X(n46009) );
  inv_x4_sg U58488 ( .A(n46010), .X(n46011) );
  inv_x4_sg U58489 ( .A(n46012), .X(n46013) );
  inv_x4_sg U58490 ( .A(n46014), .X(n46015) );
  inv_x4_sg U58491 ( .A(n46016), .X(n46017) );
  inv_x4_sg U58492 ( .A(n46018), .X(n46019) );
  inv_x4_sg U58493 ( .A(n46020), .X(n46021) );
  inv_x4_sg U58494 ( .A(n46022), .X(n46023) );
  inv_x4_sg U58495 ( .A(n46024), .X(n46025) );
  inv_x4_sg U58496 ( .A(n46026), .X(n46027) );
  inv_x4_sg U58497 ( .A(n46028), .X(n46029) );
  inv_x1_sg U58498 ( .A(n46029), .X(n51586) );
  inv_x4_sg U58499 ( .A(n46030), .X(n46031) );
  inv_x1_sg U58500 ( .A(n46031), .X(n51558) );
  inv_x4_sg U58501 ( .A(n46032), .X(n46033) );
  inv_x4_sg U58502 ( .A(n46034), .X(n46035) );
  inv_x4_sg U58503 ( .A(n46036), .X(n46037) );
  inv_x4_sg U58504 ( .A(n46038), .X(n46039) );
  inv_x4_sg U58505 ( .A(n46040), .X(n46041) );
  inv_x4_sg U58506 ( .A(n46042), .X(n46043) );
  inv_x4_sg U58507 ( .A(n46044), .X(n46045) );
  inv_x4_sg U58508 ( .A(n46046), .X(n46047) );
  inv_x4_sg U58509 ( .A(n46048), .X(n46049) );
  inv_x4_sg U58510 ( .A(n46050), .X(n46051) );
  inv_x4_sg U58511 ( .A(n46052), .X(n46053) );
  inv_x4_sg U58512 ( .A(n46054), .X(n46055) );
  inv_x4_sg U58513 ( .A(n46056), .X(n46057) );
  inv_x4_sg U58514 ( .A(n46058), .X(n46059) );
  inv_x4_sg U58515 ( .A(n46060), .X(n46061) );
  inv_x4_sg U58516 ( .A(n46062), .X(n46063) );
  inv_x4_sg U58517 ( .A(n46064), .X(n46065) );
  inv_x4_sg U58518 ( .A(n46066), .X(n46067) );
  inv_x4_sg U58519 ( .A(n46068), .X(n46069) );
  inv_x4_sg U58520 ( .A(n46070), .X(n46071) );
  inv_x4_sg U58521 ( .A(n46072), .X(n46073) );
  inv_x4_sg U58522 ( .A(n46074), .X(n46075) );
  inv_x4_sg U58523 ( .A(n46076), .X(n46077) );
  inv_x4_sg U58524 ( .A(n46078), .X(n46079) );
  inv_x4_sg U58525 ( .A(n46080), .X(n46081) );
  inv_x4_sg U58526 ( .A(n46082), .X(n46083) );
  inv_x4_sg U58527 ( .A(n46084), .X(n46085) );
  inv_x4_sg U58528 ( .A(n40921), .X(n46086) );
  inv_x8_sg U58529 ( .A(n46086), .X(n46087) );
  inv_x4_sg U58530 ( .A(n41043), .X(n46088) );
  inv_x8_sg U58531 ( .A(n46088), .X(n46089) );
  inv_x4_sg U58532 ( .A(n41025), .X(n46090) );
  inv_x8_sg U58533 ( .A(n46090), .X(n46091) );
  inv_x4_sg U58534 ( .A(n41007), .X(n46092) );
  inv_x8_sg U58535 ( .A(n46092), .X(n46093) );
  inv_x4_sg U58536 ( .A(n40967), .X(n46094) );
  inv_x8_sg U58537 ( .A(n46094), .X(n46095) );
  inv_x4_sg U58538 ( .A(n41031), .X(n46096) );
  inv_x8_sg U58539 ( .A(n46096), .X(n46097) );
  inv_x4_sg U58540 ( .A(n41013), .X(n46098) );
  inv_x8_sg U58541 ( .A(n46098), .X(n46099) );
  inv_x4_sg U58542 ( .A(n40997), .X(n46100) );
  inv_x8_sg U58543 ( .A(n46100), .X(n46101) );
  inv_x4_sg U58544 ( .A(n40985), .X(n46102) );
  inv_x8_sg U58545 ( .A(n46102), .X(n46103) );
  inv_x4_sg U58546 ( .A(n40927), .X(n46104) );
  inv_x8_sg U58547 ( .A(n46104), .X(n46105) );
  inv_x4_sg U58548 ( .A(n40955), .X(n46106) );
  inv_x8_sg U58549 ( .A(n46106), .X(n46107) );
  inv_x4_sg U58550 ( .A(n40939), .X(n46108) );
  inv_x8_sg U58551 ( .A(n46108), .X(n46109) );
  inv_x4_sg U58552 ( .A(n40991), .X(n46110) );
  inv_x8_sg U58553 ( .A(n46110), .X(n46111) );
  inv_x4_sg U58554 ( .A(n40973), .X(n46112) );
  inv_x8_sg U58555 ( .A(n46112), .X(n46113) );
  inv_x4_sg U58556 ( .A(n40945), .X(n46114) );
  inv_x8_sg U58557 ( .A(n46114), .X(n46115) );
  inv_x4_sg U58558 ( .A(n41005), .X(n46116) );
  inv_x8_sg U58559 ( .A(n46116), .X(n46117) );
  inv_x4_sg U58560 ( .A(n40953), .X(n46118) );
  inv_x8_sg U58561 ( .A(n46118), .X(n46119) );
  inv_x4_sg U58562 ( .A(n41041), .X(n46120) );
  inv_x8_sg U58563 ( .A(n46120), .X(n46121) );
  inv_x4_sg U58564 ( .A(n41023), .X(n46122) );
  inv_x8_sg U58565 ( .A(n46122), .X(n46123) );
  inv_x4_sg U58566 ( .A(n40983), .X(n46124) );
  inv_x8_sg U58567 ( .A(n46124), .X(n46125) );
  inv_x4_sg U58568 ( .A(n40937), .X(n46126) );
  inv_x8_sg U58569 ( .A(n46126), .X(n46127) );
  inv_x4_sg U58570 ( .A(n40951), .X(n46128) );
  inv_x8_sg U58571 ( .A(n46128), .X(n46129) );
  inv_x4_sg U58572 ( .A(n40919), .X(n46130) );
  inv_x8_sg U58573 ( .A(n46130), .X(n46131) );
  inv_x4_sg U58574 ( .A(n40915), .X(n46132) );
  inv_x8_sg U58575 ( .A(n46132), .X(n46133) );
  inv_x4_sg U58576 ( .A(n41039), .X(n46134) );
  inv_x8_sg U58577 ( .A(n46134), .X(n46135) );
  inv_x4_sg U58578 ( .A(n41021), .X(n46136) );
  inv_x8_sg U58579 ( .A(n46136), .X(n46137) );
  inv_x4_sg U58580 ( .A(n40933), .X(n46138) );
  inv_x8_sg U58581 ( .A(n46138), .X(n46139) );
  inv_x4_sg U58582 ( .A(n40963), .X(n46140) );
  inv_x8_sg U58583 ( .A(n46140), .X(n46141) );
  inv_x4_sg U58584 ( .A(n40979), .X(n46142) );
  inv_x8_sg U58585 ( .A(n46142), .X(n46143) );
  inv_x4_sg U58586 ( .A(n41037), .X(n46144) );
  inv_x8_sg U58587 ( .A(n46144), .X(n46145) );
  inv_x4_sg U58588 ( .A(n41019), .X(n46146) );
  inv_x8_sg U58589 ( .A(n46146), .X(n46147) );
  inv_x4_sg U58590 ( .A(n40965), .X(n46148) );
  inv_x8_sg U58591 ( .A(n46148), .X(n46149) );
  inv_x4_sg U58592 ( .A(n40949), .X(n46150) );
  inv_x8_sg U58593 ( .A(n46150), .X(n46151) );
  inv_x4_sg U58594 ( .A(n40935), .X(n46152) );
  inv_x8_sg U58595 ( .A(n46152), .X(n46153) );
  inv_x4_sg U58596 ( .A(n41029), .X(n46154) );
  inv_x8_sg U58597 ( .A(n46154), .X(n46155) );
  inv_x4_sg U58598 ( .A(n41011), .X(n46156) );
  inv_x8_sg U58599 ( .A(n46156), .X(n46157) );
  inv_x4_sg U58600 ( .A(n40995), .X(n46158) );
  inv_x8_sg U58601 ( .A(n46158), .X(n46159) );
  inv_x4_sg U58602 ( .A(n40981), .X(n46160) );
  inv_x8_sg U58603 ( .A(n46160), .X(n46161) );
  inv_x4_sg U58604 ( .A(n40913), .X(n46162) );
  inv_x8_sg U58605 ( .A(n46162), .X(n46163) );
  inv_x4_sg U58606 ( .A(n40925), .X(n46164) );
  inv_x8_sg U58607 ( .A(n46164), .X(n46165) );
  inv_x4_sg U58608 ( .A(n40977), .X(n46166) );
  inv_x8_sg U58609 ( .A(n46166), .X(n46167) );
  inv_x4_sg U58610 ( .A(n40961), .X(n46168) );
  inv_x8_sg U58611 ( .A(n46168), .X(n46169) );
  inv_x4_sg U58612 ( .A(n41017), .X(n46170) );
  inv_x8_sg U58613 ( .A(n46170), .X(n46171) );
  inv_x4_sg U58614 ( .A(n40959), .X(n46172) );
  inv_x8_sg U58615 ( .A(n46172), .X(n46173) );
  inv_x4_sg U58616 ( .A(n41035), .X(n46174) );
  inv_x8_sg U58617 ( .A(n46174), .X(n46175) );
  inv_x4_sg U58618 ( .A(n40947), .X(n46176) );
  inv_x8_sg U58619 ( .A(n46176), .X(n46177) );
  inv_x4_sg U58620 ( .A(n40989), .X(n46178) );
  inv_x8_sg U58621 ( .A(n46178), .X(n46179) );
  inv_x4_sg U58622 ( .A(n40971), .X(n46180) );
  inv_x8_sg U58623 ( .A(n46180), .X(n46181) );
  inv_x4_sg U58624 ( .A(n40943), .X(n46182) );
  inv_x8_sg U58625 ( .A(n46182), .X(n46183) );
  inv_x4_sg U58626 ( .A(n40931), .X(n46184) );
  inv_x8_sg U58627 ( .A(n46184), .X(n46185) );
  inv_x4_sg U58628 ( .A(n40917), .X(n46186) );
  inv_x8_sg U58629 ( .A(n46186), .X(n46187) );
  nand_x2_sg U58630 ( .A(n55458), .B(n46583), .X(n29633) );
  nand_x4_sg U58631 ( .A(n54184), .B(n46343), .X(n18612) );
  inv_x8_sg U58632 ( .A(n18574), .X(n54184) );
  inv_x8_sg U58633 ( .A(n21714), .X(n55362) );
  nand_x4_sg U58634 ( .A(n55362), .B(n46260), .X(n21624) );
  inv_x8_sg U58635 ( .A(n20169), .X(n54794) );
  nand_x4_sg U58636 ( .A(n54794), .B(n46305), .X(n20079) );
  nand_x4_sg U58637 ( .A(n51995), .B(n46529), .X(n12315) );
  nand_x4_sg U58638 ( .A(n51995), .B(n46525), .X(n12417) );
  nand_x4_sg U58639 ( .A(n51995), .B(n51819), .X(n12580) );
  inv_x8_sg U58640 ( .A(n12404), .X(n51995) );
  nand_x4_sg U58641 ( .A(n53663), .B(n46395), .X(n16994) );
  nand_x4_sg U58642 ( .A(n53663), .B(n46388), .X(n17261) );
  inv_x8_sg U58643 ( .A(n17083), .X(n53663) );
  nand_x4_sg U58644 ( .A(n53105), .B(n46439), .X(n15428) );
  nand_x4_sg U58645 ( .A(n53105), .B(n46432), .X(n15695) );
  inv_x8_sg U58646 ( .A(n15517), .X(n53105) );
  nand_x4_sg U58647 ( .A(n52546), .B(n46478), .X(n14142) );
  nand_x4_sg U58648 ( .A(n52546), .B(n46484), .X(n13875) );
  inv_x8_sg U58649 ( .A(n13964), .X(n52546) );
  nand_x4_sg U58650 ( .A(n52271), .B(n46507), .X(n13095) );
  nand_x4_sg U58651 ( .A(n52271), .B(n46500), .X(n13362) );
  inv_x8_sg U58652 ( .A(n13184), .X(n52271) );
  inv_x4_sg U58653 ( .A(n41137), .X(n46188) );
  inv_x8_sg U58654 ( .A(n46188), .X(state[0]) );
  inv_x4_sg U58655 ( .A(n41001), .X(n46190) );
  inv_x8_sg U58656 ( .A(n46190), .X(n46191) );
  nand_x4_sg U58657 ( .A(n51717), .B(n46551), .X(n11534) );
  nand_x4_sg U58658 ( .A(n51717), .B(n51537), .X(n11805) );
  inv_x8_sg U58659 ( .A(n11623), .X(n51717) );
  inv_x4_sg U58660 ( .A(n41003), .X(n46192) );
  inv_x8_sg U58661 ( .A(n46192), .X(n46193) );
  inv_x8_sg U58662 ( .A(n10923), .X(n51458) );
  nor_x2_sg U58663 ( .A(n46232), .B(n51458), .X(n25495) );
  nand_x4_sg U58664 ( .A(n55319), .B(n46251), .X(n21703) );
  nand_x4_sg U58665 ( .A(n55319), .B(n46249), .X(n21896) );
  inv_x8_sg U58666 ( .A(n21774), .X(n55319) );
  nand_x4_sg U58667 ( .A(n54751), .B(n46296), .X(n20158) );
  nand_x4_sg U58668 ( .A(n54751), .B(n46294), .X(n20351) );
  inv_x8_sg U58669 ( .A(n20229), .X(n54751) );
  inv_x8_sg U58670 ( .A(n16299), .X(n53384) );
  nand_x4_sg U58671 ( .A(n53384), .B(n46417), .X(n16210) );
  nand_x4_sg U58672 ( .A(n53384), .B(n53207), .X(n16479) );
  inv_x4_sg U58673 ( .A(n41135), .X(n46194) );
  inv_x8_sg U58674 ( .A(n46194), .X(n46195) );
  nor_x2_sg U58675 ( .A(n46204), .B(n55299), .X(n29379) );
  nand_x4_sg U58676 ( .A(n55299), .B(n55202), .X(n21913) );
  inv_x8_sg U58677 ( .A(n21532), .X(n55299) );
  nor_x2_sg U58678 ( .A(n46208), .B(n54731), .X(n28818) );
  nand_x4_sg U58679 ( .A(n54731), .B(n54634), .X(n20368) );
  inv_x8_sg U58680 ( .A(n19987), .X(n54731) );
  nor_x2_sg U58681 ( .A(n46212), .B(n54165), .X(n28260) );
  nand_x4_sg U58682 ( .A(n54165), .B(n54070), .X(n18823) );
  inv_x8_sg U58683 ( .A(n18442), .X(n54165) );
  nand_x4_sg U58684 ( .A(n46268), .B(n54995), .X(n21112) );
  inv_x8_sg U58685 ( .A(n20717), .X(n54995) );
  nand_x4_sg U58686 ( .A(n46313), .B(n54427), .X(n19568) );
  inv_x8_sg U58687 ( .A(n19173), .X(n54427) );
  nand_x4_sg U58688 ( .A(n46360), .B(n53862), .X(n18023) );
  inv_x8_sg U58689 ( .A(n17628), .X(n53862) );
  nand_x4_sg U58690 ( .A(n52742), .B(n52670), .X(n14902) );
  inv_x8_sg U58691 ( .A(n14507), .X(n52742) );
  nor_x2_sg U58692 ( .A(n46204), .B(n55344), .X(n29393) );
  inv_x8_sg U58693 ( .A(n21653), .X(n55344) );
  nor_x2_sg U58694 ( .A(n46208), .B(n54776), .X(n28832) );
  inv_x8_sg U58695 ( .A(n20108), .X(n54776) );
  inv_x8_sg U58696 ( .A(n18623), .X(n54229) );
  nand_x4_sg U58697 ( .A(n54229), .B(n46345), .X(n18808) );
  nand_x4_sg U58698 ( .A(n54229), .B(n46352), .X(n18534) );
  nand_x4_sg U58699 ( .A(n46558), .B(n51334), .X(n10875) );
  nand_x4_sg U58700 ( .A(n46567), .B(n51435), .X(n10955) );
  inv_x8_sg U58701 ( .A(n10843), .X(n51435) );
  nand_x4_sg U58702 ( .A(n51435), .B(n46574), .X(n10753) );
  nor_x2_sg U58703 ( .A(n46212), .B(n54209), .X(n28274) );
  nand_x4_sg U58704 ( .A(n18638), .B(n54209), .X(n18595) );
  nand_x4_sg U58705 ( .A(n54209), .B(n46352), .X(n18561) );
  inv_x8_sg U58706 ( .A(n18654), .X(n54209) );
  nor_x2_sg U58707 ( .A(n46222), .B(n52806), .X(n26875) );
  inv_x8_sg U58708 ( .A(n14674), .X(n52806) );
  nor_x2_sg U58709 ( .A(n46206), .B(n55059), .X(n29111) );
  inv_x8_sg U58710 ( .A(n20884), .X(n55059) );
  nor_x2_sg U58711 ( .A(n46210), .B(n54491), .X(n28552) );
  inv_x8_sg U58712 ( .A(n19340), .X(n54491) );
  nor_x2_sg U58713 ( .A(n46214), .B(n53926), .X(n27994) );
  inv_x8_sg U58714 ( .A(n17795), .X(n53926) );
  nand_x4_sg U58715 ( .A(n53227), .B(n53298), .X(n16465) );
  inv_x8_sg U58716 ( .A(n16069), .X(n53298) );
  nor_x2_sg U58717 ( .A(n46206), .B(n55016), .X(n29097) );
  nand_x4_sg U58718 ( .A(n55016), .B(n46268), .X(n21143) );
  inv_x8_sg U58719 ( .A(n20762), .X(n55016) );
  nor_x2_sg U58720 ( .A(n46210), .B(n54448), .X(n28538) );
  nand_x4_sg U58721 ( .A(n54448), .B(n46313), .X(n19599) );
  inv_x8_sg U58722 ( .A(n19218), .X(n54448) );
  nor_x2_sg U58723 ( .A(n46214), .B(n53883), .X(n27980) );
  nand_x4_sg U58724 ( .A(n53883), .B(n46360), .X(n18054) );
  inv_x8_sg U58725 ( .A(n17673), .X(n53883) );
  inv_x8_sg U58726 ( .A(n16442), .X(n53408) );
  nor_x2_sg U58727 ( .A(n46218), .B(n53408), .X(n27448) );
  inv_x8_sg U58728 ( .A(n11768), .X(n51738) );
  nor_x2_sg U58729 ( .A(n46230), .B(n51738), .X(n25773) );
  inv_x8_sg U58730 ( .A(n21091), .X(n55101) );
  nor_x2_sg U58731 ( .A(n46206), .B(n55101), .X(n29125) );
  inv_x8_sg U58732 ( .A(n19547), .X(n54533) );
  nor_x2_sg U58733 ( .A(n46210), .B(n54533), .X(n28566) );
  inv_x8_sg U58734 ( .A(n18002), .X(n53968) );
  nor_x2_sg U58735 ( .A(n46214), .B(n53968), .X(n28008) );
  inv_x8_sg U58736 ( .A(n18771), .X(n54250) );
  nor_x2_sg U58737 ( .A(n46212), .B(n54250), .X(n28288) );
  inv_x8_sg U58738 ( .A(n14881), .X(n52848) );
  nor_x2_sg U58739 ( .A(n46222), .B(n52848), .X(n26889) );
  inv_x8_sg U58740 ( .A(n21862), .X(n55386) );
  nor_x2_sg U58741 ( .A(n46204), .B(n55386), .X(n29407) );
  inv_x8_sg U58742 ( .A(n20317), .X(n54818) );
  nor_x2_sg U58743 ( .A(n46208), .B(n54818), .X(n28846) );
  nor_x2_sg U58744 ( .A(n46222), .B(n52763), .X(n26861) );
  nand_x4_sg U58745 ( .A(n52763), .B(n52670), .X(n14933) );
  inv_x8_sg U58746 ( .A(n14552), .X(n52763) );
  nand_x8_sg U58747 ( .A(n46241), .B(n46256), .X(n21417) );
  nand_x4_sg U58748 ( .A(n55256), .B(n46241), .X(n21746) );
  nand_x8_sg U58749 ( .A(n46286), .B(n46301), .X(n19872) );
  nand_x4_sg U58750 ( .A(n54688), .B(n46286), .X(n20201) );
  nand_x4_sg U58751 ( .A(n46513), .B(n51854), .X(n12339) );
  nor_x2_sg U58752 ( .A(n46228), .B(n51931), .X(n26023) );
  nand_x4_sg U58753 ( .A(n51931), .B(n51839), .X(n12596) );
  nand_x4_sg U58754 ( .A(n51931), .B(n46529), .X(n12161) );
  inv_x8_sg U58755 ( .A(n12218), .X(n51931) );
  nor_x2_sg U58756 ( .A(n46230), .B(n51650), .X(n25745) );
  nand_x4_sg U58757 ( .A(n51650), .B(n46539), .X(n11821) );
  nand_x4_sg U58758 ( .A(n51650), .B(n46551), .X(n11381) );
  inv_x8_sg U58759 ( .A(n11438), .X(n51650) );
  nor_x2_sg U58760 ( .A(n46218), .B(n53319), .X(n27420) );
  nand_x4_sg U58761 ( .A(n53319), .B(n53227), .X(n16496) );
  nand_x4_sg U58762 ( .A(n53319), .B(n46417), .X(n16056) );
  inv_x8_sg U58763 ( .A(n16113), .X(n53319) );
  nor_x2_sg U58764 ( .A(n46216), .B(n53598), .X(n27700) );
  nand_x4_sg U58765 ( .A(n53598), .B(n46383), .X(n17277) );
  nand_x4_sg U58766 ( .A(n53598), .B(n46395), .X(n16841) );
  inv_x8_sg U58767 ( .A(n16898), .X(n53598) );
  nor_x2_sg U58768 ( .A(n46220), .B(n53040), .X(n27140) );
  nand_x4_sg U58769 ( .A(n53040), .B(n46427), .X(n15711) );
  nand_x4_sg U58770 ( .A(n53040), .B(n46439), .X(n15275) );
  inv_x8_sg U58771 ( .A(n15332), .X(n53040) );
  nor_x2_sg U58772 ( .A(n46224), .B(n52483), .X(n26583) );
  nand_x4_sg U58773 ( .A(n52483), .B(n46484), .X(n13722) );
  nand_x4_sg U58774 ( .A(n52483), .B(n52391), .X(n14158) );
  inv_x8_sg U58775 ( .A(n13779), .X(n52483) );
  nor_x2_sg U58776 ( .A(n46226), .B(n52206), .X(n26304) );
  nand_x4_sg U58777 ( .A(n52206), .B(n46495), .X(n13378) );
  nand_x4_sg U58778 ( .A(n52206), .B(n46507), .X(n12942) );
  inv_x8_sg U58779 ( .A(n12999), .X(n52206) );
  inv_x4_sg U58780 ( .A(n41133), .X(n46199) );
  inv_x8_sg U58781 ( .A(n46199), .X(n46200) );
  inv_x4_sg U58782 ( .A(n46200), .X(n55458) );
  nand_x1_sg U58783 ( .A(n46510), .B(n8842), .X(n8841) );
  nand_x1_sg U58784 ( .A(n46487), .B(n8797), .X(n8796) );
  nand_x1_sg U58785 ( .A(n46263), .B(n9111), .X(n9110) );
  nand_x1_sg U58786 ( .A(n46375), .B(n9260), .X(n9259) );
  nand_x1_sg U58787 ( .A(n46553), .B(n8880), .X(n8879) );
  nand_x1_sg U58788 ( .A(n10359), .B(n10360), .X(n10358) );
  nand_x1_sg U58789 ( .A(n11126), .B(n11127), .X(n11125) );
  nand_x1_sg U58790 ( .A(n11909), .B(n11910), .X(n11908) );
  nand_x1_sg U58791 ( .A(n12687), .B(n12688), .X(n12686) );
  nand_x1_sg U58792 ( .A(n13471), .B(n13472), .X(n13470) );
  nand_x1_sg U58793 ( .A(n15020), .B(n15021), .X(n15019) );
  nand_x1_sg U58794 ( .A(n15805), .B(n15806), .X(n15804) );
  nand_x1_sg U58795 ( .A(n16586), .B(n16587), .X(n16585) );
  nand_x1_sg U58796 ( .A(n18141), .B(n18142), .X(n18140) );
  nand_x1_sg U58797 ( .A(n19686), .B(n19687), .X(n19685) );
  nand_x1_sg U58798 ( .A(n21231), .B(n21232), .X(n21230) );
  nand_x1_sg U58799 ( .A(n13314), .B(n13225), .X(n13313) );
  nand_x1_sg U58800 ( .A(n14094), .B(n14005), .X(n14093) );
  nand_x1_sg U58801 ( .A(n15647), .B(n15558), .X(n15646) );
  nand_x1_sg U58802 ( .A(n17213), .B(n17124), .X(n17212) );
  nand_x1_sg U58803 ( .A(n12533), .B(n12444), .X(n12532) );
  nand_x1_sg U58804 ( .A(n46419), .B(n9341), .X(n9340) );
  nand_x1_sg U58805 ( .A(n46398), .B(n9292), .X(n9291) );
  nand_x1_sg U58806 ( .A(n46398), .B(n9298), .X(n9297) );
  nand_x1_sg U58807 ( .A(n46327), .B(n9222), .X(n9221) );
  nand_x1_sg U58808 ( .A(n46531), .B(n8917), .X(n8916) );
  nand_x1_sg U58809 ( .A(n46465), .B(n8956), .X(n8955) );
  nand_x1_sg U58810 ( .A(n14250), .B(n14251), .X(n14249) );
  nand_x1_sg U58811 ( .A(n17369), .B(n17370), .X(n17368) );
  nand_x1_sg U58812 ( .A(n18914), .B(n18915), .X(n18913) );
  nand_x1_sg U58813 ( .A(n20458), .B(n20459), .X(n20457) );
  nand_x1_sg U58814 ( .A(n12499), .B(n12501), .X(n12500) );
  nand_x1_sg U58815 ( .A(n13280), .B(n13282), .X(n13281) );
  nand_x1_sg U58816 ( .A(n14060), .B(n14062), .X(n14061) );
  nand_x1_sg U58817 ( .A(n15613), .B(n15615), .X(n15614) );
  nand_x1_sg U58818 ( .A(n17179), .B(n17181), .X(n17180) );
  nand_x1_sg U58819 ( .A(n46442), .B(n8975), .X(n8974) );
  nand_x1_sg U58820 ( .A(n46442), .B(n8981), .X(n8980) );
  nand_x1_sg U58821 ( .A(n51890), .B(n52025), .X(n12589) );
  nand_x1_sg U58822 ( .A(n17868), .B(n17869), .X(n17867) );
  nand_x1_sg U58823 ( .A(n19413), .B(n19414), .X(n19412) );
  nand_x1_sg U58824 ( .A(n20957), .B(n20958), .X(n20956) );
  nand_x1_sg U58825 ( .A(n14747), .B(n14748), .X(n14746) );
  nand_x1_sg U58826 ( .A(n13199), .B(n13198), .X(n13196) );
  nand_x1_sg U58827 ( .A(n13979), .B(n13978), .X(n13976) );
  nand_x1_sg U58828 ( .A(n15532), .B(n15531), .X(n15529) );
  nand_x1_sg U58829 ( .A(n17098), .B(n17097), .X(n17095) );
  nand_x1_sg U58830 ( .A(n20181), .B(n20182), .X(n20180) );
  nand_x1_sg U58831 ( .A(n21726), .B(n21727), .X(n21725) );
  inv_x1_sg U58832 ( .A(n18333), .X(n54147) );
  inv_x1_sg U58833 ( .A(n10551), .X(n51358) );
  inv_x1_sg U58834 ( .A(n19878), .X(n54712) );
  inv_x1_sg U58835 ( .A(n21423), .X(n55280) );
  nand_x1_sg U58836 ( .A(n9039), .B(n46577), .X(n9038) );
  nand_x1_sg U58837 ( .A(n46283), .B(n9140), .X(n9139) );
  nand_x1_sg U58838 ( .A(n46283), .B(n9146), .X(n9145) );
  nand_x1_sg U58839 ( .A(n46355), .B(n42629), .X(n9082) );
  nand_x1_sg U58840 ( .A(n46355), .B(n9067), .X(n9066) );
  nand_x1_sg U58841 ( .A(n46308), .B(n41354), .X(n9196) );
  nand_x1_sg U58842 ( .A(n46308), .B(n9201), .X(n9200) );
  nand_x1_sg U58843 ( .A(n24502), .B(n46607), .X(n24501) );
  nand_x1_sg U58844 ( .A(n21974), .B(n21951), .X(n21972) );
  nand_x1_sg U58845 ( .A(n29639), .B(n29606), .X(n29637) );
  inv_x1_sg U58846 ( .A(n26984), .X(n52661) );
  inv_x1_sg U58847 ( .A(n25581), .X(n51279) );
  inv_x1_sg U58848 ( .A(n26705), .X(n52384) );
  inv_x1_sg U58849 ( .A(n28939), .X(n54626) );
  inv_x1_sg U58850 ( .A(n29500), .X(n55194) );
  inv_x1_sg U58851 ( .A(n27543), .X(n53220) );
  inv_x1_sg U58852 ( .A(n26148), .X(n51832) );
  inv_x1_sg U58853 ( .A(n25587), .X(n51272) );
  inv_x1_sg U58854 ( .A(n26978), .X(n52669) );
  inv_x1_sg U58855 ( .A(n28933), .X(n54633) );
  inv_x1_sg U58856 ( .A(n29494), .X(n55201) );
  inv_x1_sg U58857 ( .A(n26699), .X(n52390) );
  inv_x1_sg U58858 ( .A(n26142), .X(n51838) );
  inv_x1_sg U58859 ( .A(n27537), .X(n53226) );
  inv_x1_sg U58860 ( .A(n28370), .X(n54083) );
  nand_x2_sg U58861 ( .A(n50146), .B(n50117), .X(n23760) );
  nand_x2_sg U58862 ( .A(n49287), .B(n49258), .X(n31426) );
  inv_x1_sg U58863 ( .A(n44787), .X(n50985) );
  inv_x1_sg U58864 ( .A(n44785), .X(n51004) );
  inv_x1_sg U58865 ( .A(n44783), .X(n51023) );
  inv_x1_sg U58866 ( .A(n44781), .X(n51042) );
  inv_x1_sg U58867 ( .A(n44779), .X(n51062) );
  inv_x1_sg U58868 ( .A(n44777), .X(n51081) );
  inv_x1_sg U58869 ( .A(n44775), .X(n51100) );
  inv_x1_sg U58870 ( .A(n44773), .X(n51119) );
  inv_x1_sg U58871 ( .A(n44771), .X(n51138) );
  inv_x1_sg U58872 ( .A(n44769), .X(n51157) );
  inv_x1_sg U58873 ( .A(n44767), .X(n51175) );
  inv_x1_sg U58874 ( .A(n44765), .X(n51194) );
  inv_x1_sg U58875 ( .A(n44763), .X(n51213) );
  inv_x1_sg U58876 ( .A(n44761), .X(n51232) );
  inv_x1_sg U58877 ( .A(n44759), .X(n51251) );
  nand_x1_sg U58878 ( .A(n16222), .B(n15817), .X(n16220) );
  nand_x1_sg U58879 ( .A(n10765), .B(n10371), .X(n10763) );
  nand_x1_sg U58880 ( .A(n13548), .B(n13550), .X(n13549) );
  nand_x1_sg U58881 ( .A(n17466), .B(n17465), .X(n17463) );
  nand_x1_sg U58882 ( .A(n19011), .B(n19010), .X(n19008) );
  nand_x1_sg U58883 ( .A(n20555), .B(n20554), .X(n20552) );
  nand_x1_sg U58884 ( .A(n10451), .B(n10450), .X(n10448) );
  nand_x1_sg U58885 ( .A(n14343), .B(n14342), .X(n14340) );
  nand_x1_sg U58886 ( .A(n19778), .B(n19777), .X(n19775) );
  nand_x1_sg U58887 ( .A(n21323), .B(n21322), .X(n21320) );
  nand_x1_sg U58888 ( .A(n11375), .B(n11376), .X(n11374) );
  nand_x1_sg U58889 ( .A(n12155), .B(n12156), .X(n12154) );
  nand_x1_sg U58890 ( .A(n12936), .B(n12937), .X(n12935) );
  nand_x1_sg U58891 ( .A(n15269), .B(n15270), .X(n15268) );
  nand_x1_sg U58892 ( .A(n16050), .B(n16051), .X(n16049) );
  nand_x1_sg U58893 ( .A(n16835), .B(n16836), .X(n16834) );
  nand_x1_sg U58894 ( .A(n18232), .B(n18231), .X(n18229) );
  inv_x1_sg U58895 ( .A(n17420), .X(n53783) );
  inv_x1_sg U58896 ( .A(n18965), .X(n54348) );
  inv_x1_sg U58897 ( .A(n20509), .X(n54916) );
  nand_x1_sg U58898 ( .A(n14880), .B(n14915), .X(n14913) );
  nand_x1_sg U58899 ( .A(n18001), .B(n18036), .X(n18034) );
  nand_x1_sg U58900 ( .A(n19546), .B(n19581), .X(n19579) );
  nand_x1_sg U58901 ( .A(n21090), .B(n21125), .X(n21123) );
  nand_x1_sg U58902 ( .A(n12003), .B(n12002), .X(n12000) );
  nand_x1_sg U58903 ( .A(n15898), .B(n15897), .X(n15895) );
  nand_x1_sg U58904 ( .A(n11226), .B(n11225), .X(n11223) );
  nand_x1_sg U58905 ( .A(n12787), .B(n12786), .X(n12784) );
  nand_x1_sg U58906 ( .A(n15120), .B(n15119), .X(n15117) );
  nand_x1_sg U58907 ( .A(n16686), .B(n16685), .X(n16683) );
  nand_x1_sg U58908 ( .A(n51622), .B(n11272), .X(n11271) );
  nand_x1_sg U58909 ( .A(n52181), .B(n12833), .X(n12832) );
  nand_x1_sg U58910 ( .A(n53015), .B(n15166), .X(n15165) );
  nand_x1_sg U58911 ( .A(n53573), .B(n16732), .X(n16731) );
  nand_x1_sg U58912 ( .A(n51904), .B(n12051), .X(n12050) );
  nand_x1_sg U58913 ( .A(n53289), .B(n15946), .X(n15945) );
  nand_x1_sg U58914 ( .A(n14539), .B(n14549), .X(n14548) );
  nand_x1_sg U58915 ( .A(n17660), .B(n17670), .X(n17669) );
  nand_x1_sg U58916 ( .A(n19205), .B(n19215), .X(n19214) );
  nand_x1_sg U58917 ( .A(n20749), .B(n20759), .X(n20758) );
  nand_x2_sg U58918 ( .A(n13530), .B(n46484), .X(n13526) );
  nand_x1_sg U58919 ( .A(n17450), .B(n17452), .X(n17451) );
  nand_x1_sg U58920 ( .A(n18995), .B(n18997), .X(n18996) );
  nand_x1_sg U58921 ( .A(n20539), .B(n20541), .X(n20540) );
  nand_x1_sg U58922 ( .A(n13716), .B(n13717), .X(n13715) );
  nand_x2_sg U58923 ( .A(n53844), .B(n17703), .X(n17701) );
  nand_x2_sg U58924 ( .A(n54409), .B(n19248), .X(n19246) );
  nand_x2_sg U58925 ( .A(n54977), .B(n20792), .X(n20790) );
  nand_x2_sg U58926 ( .A(n54125), .B(n18472), .X(n18470) );
  nand_x2_sg U58927 ( .A(n51335), .B(n10690), .X(n10688) );
  nand_x2_sg U58928 ( .A(n52448), .B(n13812), .X(n13810) );
  nand_x2_sg U58929 ( .A(n53283), .B(n16146), .X(n16144) );
  nand_x2_sg U58930 ( .A(n51897), .B(n12251), .X(n12249) );
  nand_x2_sg U58931 ( .A(n51615), .B(n11471), .X(n11469) );
  nand_x2_sg U58932 ( .A(n52173), .B(n13032), .X(n13030) );
  nand_x2_sg U58933 ( .A(n53007), .B(n15365), .X(n15363) );
  nand_x2_sg U58934 ( .A(n53565), .B(n16931), .X(n16929) );
  nand_x1_sg U58935 ( .A(n11208), .B(n11210), .X(n11209) );
  nand_x1_sg U58936 ( .A(n12769), .B(n12771), .X(n12770) );
  nand_x1_sg U58937 ( .A(n15102), .B(n15104), .X(n15103) );
  nand_x1_sg U58938 ( .A(n16668), .B(n16670), .X(n16669) );
  nand_x1_sg U58939 ( .A(n10435), .B(n10437), .X(n10436) );
  nand_x1_sg U58940 ( .A(n14327), .B(n14329), .X(n14328) );
  nand_x1_sg U58941 ( .A(n19762), .B(n19764), .X(n19763) );
  nand_x1_sg U58942 ( .A(n21307), .B(n21309), .X(n21308) );
  nand_x2_sg U58943 ( .A(n54689), .B(n20017), .X(n20015) );
  nand_x2_sg U58944 ( .A(n55257), .B(n21562), .X(n21560) );
  nand_x1_sg U58945 ( .A(n11987), .B(n11989), .X(n11988) );
  nand_x1_sg U58946 ( .A(n15882), .B(n15884), .X(n15883) );
  nand_x1_sg U58947 ( .A(n18216), .B(n18218), .X(n18217) );
  nand_x2_sg U58948 ( .A(n52724), .B(n14582), .X(n14580) );
  nand_x1_sg U58949 ( .A(n43938), .B(n11965), .X(n11968) );
  nand_x1_sg U58950 ( .A(n15862), .B(n15860), .X(n15863) );
  nand_x1_sg U58951 ( .A(n43843), .B(n11187), .X(n11190) );
  nand_x1_sg U58952 ( .A(n43841), .B(n12748), .X(n12751) );
  nand_x1_sg U58953 ( .A(n43839), .B(n15081), .X(n15084) );
  nand_x1_sg U58954 ( .A(n43837), .B(n16647), .X(n16650) );
  nand_x1_sg U58955 ( .A(n13775), .B(n14168), .X(n14166) );
  nand_x1_sg U58956 ( .A(n14646), .B(n14645), .X(n14643) );
  nand_x1_sg U58957 ( .A(n17767), .B(n17766), .X(n17764) );
  nand_x1_sg U58958 ( .A(n19312), .B(n19311), .X(n19309) );
  nand_x1_sg U58959 ( .A(n20856), .B(n20855), .X(n20853) );
  nand_x1_sg U58960 ( .A(n20080), .B(n20079), .X(n20077) );
  nand_x1_sg U58961 ( .A(n21625), .B(n21624), .X(n21622) );
  nand_x2_sg U58962 ( .A(n17431), .B(n46372), .X(n17428) );
  nand_x2_sg U58963 ( .A(n18976), .B(n46325), .X(n18973) );
  nand_x2_sg U58964 ( .A(n20520), .B(n46280), .X(n20517) );
  nand_x2_sg U58965 ( .A(n11191), .B(n46551), .X(n11187) );
  nand_x2_sg U58966 ( .A(n12752), .B(n46507), .X(n12748) );
  nand_x2_sg U58967 ( .A(n15085), .B(n46439), .X(n15081) );
  nand_x2_sg U58968 ( .A(n16651), .B(n46395), .X(n16647) );
  nand_x2_sg U58969 ( .A(n18198), .B(n18184), .X(n18195) );
  nand_x2_sg U58970 ( .A(n14310), .B(n46462), .X(n14307) );
  nand_x2_sg U58971 ( .A(n10418), .B(n46574), .X(n10415) );
  nand_x2_sg U58972 ( .A(n19745), .B(n19730), .X(n19742) );
  nand_x2_sg U58973 ( .A(n21290), .B(n21275), .X(n21287) );
  nand_x2_sg U58974 ( .A(n11969), .B(n11952), .X(n11965) );
  nand_x2_sg U58975 ( .A(n15864), .B(n15847), .X(n15860) );
  nor_x1_sg U58976 ( .A(n26721), .B(n52364), .X(n8785) );
  nand_x4_sg U58977 ( .A(n13456), .B(n52606), .X(n8813) );
  nor_x1_sg U58978 ( .A(n13458), .B(n13459), .X(n13457) );
  nand_x4_sg U58979 ( .A(n13459), .B(n13458), .X(n13456) );
  nand_x1_sg U58980 ( .A(n52003), .B(n11892), .X(n11891) );
  nand_x1_sg U58981 ( .A(n52535), .B(n13450), .X(n13449) );
  nand_x1_sg U58982 ( .A(n52554), .B(n13454), .X(n13453) );
  nand_x1_sg U58983 ( .A(n53392), .B(n15787), .X(n15786) );
  nand_x1_sg U58984 ( .A(n51442), .B(n10341), .X(n10340) );
  nand_x1_sg U58985 ( .A(n52831), .B(n14233), .X(n14232) );
  nand_x1_sg U58986 ( .A(n53951), .B(n17352), .X(n17351) );
  nand_x1_sg U58987 ( .A(n54236), .B(n18124), .X(n18123) );
  nand_x1_sg U58988 ( .A(n54516), .B(n18897), .X(n18896) );
  nand_x1_sg U58989 ( .A(n54801), .B(n19669), .X(n19668) );
  nand_x1_sg U58990 ( .A(n55084), .B(n20441), .X(n20440) );
  nand_x1_sg U58991 ( .A(n55369), .B(n21214), .X(n21213) );
  nand_x2_sg U58992 ( .A(n13485), .B(n13456), .X(n13484) );
  nand_x1_sg U58993 ( .A(n43273), .B(n13839), .X(n13485) );
  nand_x4_sg U58994 ( .A(n11115), .B(n51790), .X(n8882) );
  nand_x1_sg U58995 ( .A(n51775), .B(n43203), .X(n11115) );
  nand_x4_sg U58996 ( .A(n11898), .B(n43230), .X(n8900) );
  nand_x1_sg U58997 ( .A(n52055), .B(n42347), .X(n11898) );
  nand_x4_sg U58998 ( .A(n12676), .B(n52346), .X(n8848) );
  nand_x1_sg U58999 ( .A(n52332), .B(n43201), .X(n12676) );
  nand_x4_sg U59000 ( .A(n13460), .B(n52621), .X(n8799) );
  nand_x1_sg U59001 ( .A(n52607), .B(n43199), .X(n13460) );
  nand_x4_sg U59002 ( .A(n14239), .B(n52900), .X(n9002) );
  nand_x1_sg U59003 ( .A(n52885), .B(n44693), .X(n14239) );
  nand_x4_sg U59004 ( .A(n15009), .B(n53180), .X(n8992) );
  nand_x1_sg U59005 ( .A(n53166), .B(n43197), .X(n15009) );
  nand_x4_sg U59006 ( .A(n16575), .B(n53738), .X(n9300) );
  nand_x1_sg U59007 ( .A(n53724), .B(n43195), .X(n16575) );
  nand_x4_sg U59008 ( .A(n17358), .B(n54020), .X(n9262) );
  nand_x1_sg U59009 ( .A(n54005), .B(n44691), .X(n17358) );
  nand_x4_sg U59010 ( .A(n18130), .B(n43228), .X(n9054) );
  nand_x1_sg U59011 ( .A(n54287), .B(n42345), .X(n18130) );
  nand_x4_sg U59012 ( .A(n18903), .B(n54585), .X(n9224) );
  nand_x1_sg U59013 ( .A(n54570), .B(n44689), .X(n18903) );
  nand_x4_sg U59014 ( .A(n19675), .B(n43226), .X(n9166) );
  nand_x1_sg U59015 ( .A(n54855), .B(n42343), .X(n19675) );
  nand_x4_sg U59016 ( .A(n20447), .B(n55153), .X(n9148) );
  nand_x1_sg U59017 ( .A(n55138), .B(n44687), .X(n20447) );
  nand_x4_sg U59018 ( .A(n21220), .B(n43224), .X(n9090) );
  nand_x1_sg U59019 ( .A(n55423), .B(n42341), .X(n21220) );
  nand_x4_sg U59020 ( .A(n11924), .B(n11925), .X(n11896) );
  nand_x1_sg U59021 ( .A(n11892), .B(n11893), .X(n11924) );
  nand_x4_sg U59022 ( .A(n13486), .B(n13487), .X(n13458) );
  nand_x1_sg U59023 ( .A(n13454), .B(n13455), .X(n13486) );
  nand_x4_sg U59024 ( .A(n15819), .B(n15820), .X(n15791) );
  nand_x1_sg U59025 ( .A(n15787), .B(n15788), .X(n15819) );
  nand_x4_sg U59026 ( .A(n10373), .B(n10374), .X(n10345) );
  nand_x1_sg U59027 ( .A(n10341), .B(n10342), .X(n10373) );
  nand_x4_sg U59028 ( .A(n14265), .B(n14266), .X(n14237) );
  nand_x1_sg U59029 ( .A(n14233), .B(n14234), .X(n14265) );
  nand_x4_sg U59030 ( .A(n17384), .B(n17385), .X(n17356) );
  nand_x1_sg U59031 ( .A(n17352), .B(n17353), .X(n17384) );
  nand_x4_sg U59032 ( .A(n18155), .B(n18156), .X(n18128) );
  nand_x1_sg U59033 ( .A(n18124), .B(n18125), .X(n18155) );
  nand_x4_sg U59034 ( .A(n18929), .B(n18930), .X(n18901) );
  nand_x1_sg U59035 ( .A(n18897), .B(n18898), .X(n18929) );
  nand_x4_sg U59036 ( .A(n19700), .B(n19701), .X(n19673) );
  nand_x1_sg U59037 ( .A(n19669), .B(n19670), .X(n19700) );
  nand_x4_sg U59038 ( .A(n20473), .B(n20474), .X(n20445) );
  nand_x1_sg U59039 ( .A(n20441), .B(n20442), .X(n20473) );
  nand_x4_sg U59040 ( .A(n21245), .B(n21246), .X(n21218) );
  nand_x1_sg U59041 ( .A(n21214), .B(n21215), .X(n21245) );
  nand_x4_sg U59042 ( .A(n13836), .B(n13837), .X(n13459) );
  nand_x1_sg U59043 ( .A(n52584), .B(n43273), .X(n13837) );
  nand_x4_sg U59044 ( .A(n13488), .B(n13489), .X(n13455) );
  nand_x1_sg U59045 ( .A(n13450), .B(n13451), .X(n13488) );
  nand_x4_sg U59046 ( .A(n10335), .B(n51441), .X(n9020) );
  nor_x1_sg U59047 ( .A(n10337), .B(n10338), .X(n10336) );
  nand_x4_sg U59048 ( .A(n10343), .B(n51496), .X(n9018) );
  nor_x1_sg U59049 ( .A(n10345), .B(n10346), .X(n10344) );
  nand_x4_sg U59050 ( .A(n11111), .B(n51774), .X(n8868) );
  nor_x1_sg U59051 ( .A(n11113), .B(n11114), .X(n11112) );
  nand_x4_sg U59052 ( .A(n11894), .B(n52054), .X(n8911) );
  nor_x1_sg U59053 ( .A(n11896), .B(n11897), .X(n11895) );
  nand_x4_sg U59054 ( .A(n12672), .B(n52331), .X(n8830) );
  nor_x1_sg U59055 ( .A(n12674), .B(n12675), .X(n12673) );
  nand_x4_sg U59056 ( .A(n14227), .B(n52830), .X(n8954) );
  nor_x1_sg U59057 ( .A(n14229), .B(n14230), .X(n14228) );
  nand_x4_sg U59058 ( .A(n14235), .B(n52884), .X(n8946) );
  nor_x1_sg U59059 ( .A(n14237), .B(n14238), .X(n14236) );
  nand_x4_sg U59060 ( .A(n15005), .B(n53165), .X(n8969) );
  nor_x1_sg U59061 ( .A(n15007), .B(n15008), .X(n15006) );
  nand_x4_sg U59062 ( .A(n15789), .B(n53444), .X(n9349) );
  nor_x1_sg U59063 ( .A(n15791), .B(n15792), .X(n15790) );
  nand_x4_sg U59064 ( .A(n16571), .B(n53723), .X(n9286) );
  nor_x1_sg U59065 ( .A(n16573), .B(n16574), .X(n16572) );
  nand_x4_sg U59066 ( .A(n17346), .B(n53950), .X(n9258) );
  nor_x1_sg U59067 ( .A(n17348), .B(n17349), .X(n17347) );
  nand_x4_sg U59068 ( .A(n17354), .B(n54004), .X(n9248) );
  nor_x1_sg U59069 ( .A(n17356), .B(n17357), .X(n17355) );
  nand_x4_sg U59070 ( .A(n18118), .B(n54235), .X(n9065) );
  nor_x1_sg U59071 ( .A(n18120), .B(n18121), .X(n18119) );
  nand_x4_sg U59072 ( .A(n18126), .B(n54286), .X(n9081) );
  nor_x1_sg U59073 ( .A(n18128), .B(n18129), .X(n18127) );
  nand_x4_sg U59074 ( .A(n18891), .B(n54515), .X(n9220) );
  nor_x1_sg U59075 ( .A(n18893), .B(n18894), .X(n18892) );
  nand_x4_sg U59076 ( .A(n18899), .B(n54569), .X(n9210) );
  nor_x1_sg U59077 ( .A(n18901), .B(n18902), .X(n18900) );
  nand_x4_sg U59078 ( .A(n19663), .B(n54800), .X(n9199) );
  nor_x1_sg U59079 ( .A(n19665), .B(n19666), .X(n19664) );
  nand_x4_sg U59080 ( .A(n19671), .B(n54854), .X(n9171) );
  nor_x1_sg U59081 ( .A(n19673), .B(n19674), .X(n19672) );
  nand_x4_sg U59082 ( .A(n20435), .B(n55083), .X(n9144) );
  nor_x1_sg U59083 ( .A(n20437), .B(n20438), .X(n20436) );
  nand_x4_sg U59084 ( .A(n20443), .B(n55137), .X(n9134) );
  nor_x1_sg U59085 ( .A(n20445), .B(n20446), .X(n20444) );
  nand_x4_sg U59086 ( .A(n21208), .B(n55368), .X(n9109) );
  nor_x1_sg U59087 ( .A(n21210), .B(n21211), .X(n21209) );
  nand_x4_sg U59088 ( .A(n21216), .B(n55422), .X(n9115) );
  nor_x1_sg U59089 ( .A(n21218), .B(n21219), .X(n21217) );
  nand_x4_sg U59090 ( .A(n51510), .B(n10347), .X(n9016) );
  nor_x1_sg U59091 ( .A(n10349), .B(n10350), .X(n10348) );
  nand_x4_sg U59092 ( .A(n53460), .B(n15793), .X(n9336) );
  nor_x1_sg U59093 ( .A(n15795), .B(n15796), .X(n15794) );
  nand_x4_sg U59094 ( .A(n10347), .B(n10370), .X(n10368) );
  nand_x4_sg U59095 ( .A(n15793), .B(n15816), .X(n15814) );
  nand_x4_sg U59096 ( .A(n10338), .B(n10337), .X(n10335) );
  nand_x4_sg U59097 ( .A(n14230), .B(n14229), .X(n14227) );
  nand_x4_sg U59098 ( .A(n17349), .B(n17348), .X(n17346) );
  nand_x4_sg U59099 ( .A(n18121), .B(n18120), .X(n18118) );
  nand_x4_sg U59100 ( .A(n18894), .B(n18893), .X(n18891) );
  nand_x4_sg U59101 ( .A(n19666), .B(n19665), .X(n19663) );
  nand_x4_sg U59102 ( .A(n20438), .B(n20437), .X(n20435) );
  nand_x4_sg U59103 ( .A(n21211), .B(n21210), .X(n21208) );
  nand_x4_sg U59104 ( .A(n10346), .B(n10345), .X(n10343) );
  nand_x4_sg U59105 ( .A(n11114), .B(n11113), .X(n11111) );
  nand_x4_sg U59106 ( .A(n11897), .B(n11896), .X(n11894) );
  nand_x4_sg U59107 ( .A(n12675), .B(n12674), .X(n12672) );
  nand_x4_sg U59108 ( .A(n14238), .B(n14237), .X(n14235) );
  nand_x4_sg U59109 ( .A(n15008), .B(n15007), .X(n15005) );
  nand_x4_sg U59110 ( .A(n15792), .B(n15791), .X(n15789) );
  nand_x4_sg U59111 ( .A(n16574), .B(n16573), .X(n16571) );
  nand_x4_sg U59112 ( .A(n17357), .B(n17356), .X(n17354) );
  nand_x4_sg U59113 ( .A(n18129), .B(n18128), .X(n18126) );
  nand_x4_sg U59114 ( .A(n18902), .B(n18901), .X(n18899) );
  nand_x4_sg U59115 ( .A(n19674), .B(n19673), .X(n19671) );
  nand_x4_sg U59116 ( .A(n20446), .B(n20445), .X(n20443) );
  nand_x4_sg U59117 ( .A(n21219), .B(n21218), .X(n21216) );
  nand_x4_sg U59118 ( .A(n10350), .B(n10349), .X(n10347) );
  nand_x4_sg U59119 ( .A(n15796), .B(n15795), .X(n15793) );
  nand_x1_sg U59120 ( .A(n51329), .B(n10316), .X(n10315) );
  nand_x1_sg U59121 ( .A(n54683), .B(n19644), .X(n19643) );
  nand_x1_sg U59122 ( .A(n55251), .B(n21189), .X(n21188) );
  nand_x1_sg U59123 ( .A(n51703), .B(n11105), .X(n11104) );
  nand_x1_sg U59124 ( .A(n51725), .B(n11109), .X(n11108) );
  nand_x1_sg U59125 ( .A(n51984), .B(n11888), .X(n11887) );
  nand_x1_sg U59126 ( .A(n52259), .B(n12666), .X(n12665) );
  nand_x1_sg U59127 ( .A(n52279), .B(n12670), .X(n12669) );
  nand_x1_sg U59128 ( .A(n53093), .B(n14999), .X(n14998) );
  nand_x1_sg U59129 ( .A(n53113), .B(n15003), .X(n15002) );
  nand_x1_sg U59130 ( .A(n53373), .B(n15783), .X(n15782) );
  nand_x1_sg U59131 ( .A(n53651), .B(n16565), .X(n16564) );
  nand_x1_sg U59132 ( .A(n53671), .B(n16569), .X(n16568) );
  nand_x1_sg U59133 ( .A(n51405), .B(n10333), .X(n10332) );
  nand_x1_sg U59134 ( .A(n51682), .B(n11101), .X(n11100) );
  nand_x1_sg U59135 ( .A(n51963), .B(n11884), .X(n11883) );
  nand_x1_sg U59136 ( .A(n52238), .B(n12662), .X(n12661) );
  nand_x1_sg U59137 ( .A(n52515), .B(n13446), .X(n13445) );
  nand_x1_sg U59138 ( .A(n52794), .B(n14225), .X(n14224) );
  nand_x1_sg U59139 ( .A(n53072), .B(n14995), .X(n14994) );
  nand_x1_sg U59140 ( .A(n53351), .B(n15779), .X(n15778) );
  nand_x1_sg U59141 ( .A(n53630), .B(n16561), .X(n16560) );
  nand_x1_sg U59142 ( .A(n53914), .B(n17344), .X(n17343) );
  nand_x1_sg U59143 ( .A(n54194), .B(n18116), .X(n18115) );
  nand_x1_sg U59144 ( .A(n54479), .B(n18889), .X(n18888) );
  nand_x1_sg U59145 ( .A(n54761), .B(n19661), .X(n19660) );
  nand_x1_sg U59146 ( .A(n55047), .B(n20433), .X(n20432) );
  nand_x1_sg U59147 ( .A(n55329), .B(n21206), .X(n21205) );
  nor_x1_sg U59148 ( .A(n10357), .B(n41400), .X(n10355) );
  nand_x1_sg U59149 ( .A(n41400), .B(n10357), .X(n10356) );
  nor_x1_sg U59150 ( .A(n11124), .B(n41398), .X(n11122) );
  nand_x1_sg U59151 ( .A(n41398), .B(n11124), .X(n11123) );
  nor_x1_sg U59152 ( .A(n11907), .B(n41396), .X(n11905) );
  nand_x1_sg U59153 ( .A(n41396), .B(n11907), .X(n11906) );
  nor_x1_sg U59154 ( .A(n12685), .B(n41394), .X(n12683) );
  nand_x1_sg U59155 ( .A(n41394), .B(n12685), .X(n12684) );
  nor_x1_sg U59156 ( .A(n13469), .B(n41390), .X(n13467) );
  nand_x1_sg U59157 ( .A(n41390), .B(n13469), .X(n13468) );
  nor_x1_sg U59158 ( .A(n15018), .B(n41386), .X(n15016) );
  nand_x1_sg U59159 ( .A(n41386), .B(n15018), .X(n15017) );
  nor_x1_sg U59160 ( .A(n15803), .B(n41382), .X(n15801) );
  nand_x1_sg U59161 ( .A(n41382), .B(n15803), .X(n15802) );
  nor_x1_sg U59162 ( .A(n16584), .B(n41380), .X(n16582) );
  nand_x1_sg U59163 ( .A(n41380), .B(n16584), .X(n16583) );
  nor_x1_sg U59164 ( .A(n18139), .B(n41191), .X(n18137) );
  nand_x1_sg U59165 ( .A(n41191), .B(n18139), .X(n18138) );
  nor_x1_sg U59166 ( .A(n19684), .B(n41372), .X(n19682) );
  nand_x1_sg U59167 ( .A(n41372), .B(n19684), .X(n19683) );
  nor_x1_sg U59168 ( .A(n21229), .B(n41368), .X(n21227) );
  nand_x1_sg U59169 ( .A(n41368), .B(n21229), .X(n21228) );
  nand_x2_sg U59170 ( .A(n11140), .B(n11111), .X(n11139) );
  nand_x1_sg U59171 ( .A(n43277), .B(n11498), .X(n11140) );
  nand_x2_sg U59172 ( .A(n11923), .B(n11894), .X(n11922) );
  nand_x1_sg U59173 ( .A(n42379), .B(n12278), .X(n11923) );
  nand_x2_sg U59174 ( .A(n12701), .B(n12672), .X(n12700) );
  nand_x1_sg U59175 ( .A(n43275), .B(n13059), .X(n12701) );
  nand_x2_sg U59176 ( .A(n14264), .B(n14235), .X(n14263) );
  nand_x1_sg U59177 ( .A(n43295), .B(n14609), .X(n14264) );
  nand_x2_sg U59178 ( .A(n15034), .B(n15005), .X(n15033) );
  nand_x1_sg U59179 ( .A(n43271), .B(n15392), .X(n15034) );
  nand_x2_sg U59180 ( .A(n16600), .B(n16571), .X(n16599) );
  nand_x1_sg U59181 ( .A(n43269), .B(n16958), .X(n16600) );
  nand_x2_sg U59182 ( .A(n17383), .B(n17354), .X(n17382) );
  nand_x1_sg U59183 ( .A(n43293), .B(n17730), .X(n17383) );
  nand_x2_sg U59184 ( .A(n18154), .B(n18126), .X(n18153) );
  nand_x1_sg U59185 ( .A(n42377), .B(n18499), .X(n18154) );
  nand_x2_sg U59186 ( .A(n18928), .B(n18899), .X(n18927) );
  nand_x1_sg U59187 ( .A(n43291), .B(n19275), .X(n18928) );
  nand_x2_sg U59188 ( .A(n19699), .B(n19671), .X(n19698) );
  nand_x1_sg U59189 ( .A(n42375), .B(n20044), .X(n19699) );
  nand_x2_sg U59190 ( .A(n20472), .B(n20443), .X(n20471) );
  nand_x1_sg U59191 ( .A(n43289), .B(n20819), .X(n20472) );
  nand_x2_sg U59192 ( .A(n21244), .B(n21216), .X(n21243) );
  nand_x1_sg U59193 ( .A(n42373), .B(n21589), .X(n21244) );
  nand_x1_sg U59194 ( .A(n41740), .B(n10324), .X(n10322) );
  nand_x1_sg U59195 ( .A(n41760), .B(n11092), .X(n11090) );
  nand_x1_sg U59196 ( .A(n41758), .B(n11875), .X(n11873) );
  nand_x1_sg U59197 ( .A(n41756), .B(n12653), .X(n12651) );
  nand_x1_sg U59198 ( .A(n41754), .B(n13437), .X(n13435) );
  nand_x1_sg U59199 ( .A(n41778), .B(n14216), .X(n14214) );
  nand_x1_sg U59200 ( .A(n41752), .B(n14986), .X(n14984) );
  nand_x1_sg U59201 ( .A(n41736), .B(n15770), .X(n15768) );
  nand_x1_sg U59202 ( .A(n41750), .B(n16552), .X(n16550) );
  nand_x1_sg U59203 ( .A(n41776), .B(n17335), .X(n17333) );
  nand_x1_sg U59204 ( .A(n41748), .B(n18107), .X(n18105) );
  nand_x1_sg U59205 ( .A(n41774), .B(n18880), .X(n18878) );
  nand_x1_sg U59206 ( .A(n41746), .B(n19652), .X(n19650) );
  nand_x1_sg U59207 ( .A(n41772), .B(n20424), .X(n20422) );
  nand_x1_sg U59208 ( .A(n41744), .B(n21197), .X(n21195) );
  nand_x4_sg U59209 ( .A(n41725), .B(n13163), .X(n12690) );
  nand_x4_sg U59210 ( .A(n41717), .B(n15496), .X(n15023) );
  nand_x4_sg U59211 ( .A(n41713), .B(n17062), .X(n16589) );
  nand_x4_sg U59212 ( .A(n45451), .B(n11602), .X(n11129) );
  nand_x4_sg U59213 ( .A(n45447), .B(n14714), .X(n14253) );
  nor_x1_sg U59214 ( .A(n41725), .B(n13163), .X(n13161) );
  nor_x1_sg U59215 ( .A(n41717), .B(n15496), .X(n15494) );
  nor_x1_sg U59216 ( .A(n41713), .B(n17062), .X(n17060) );
  nor_x1_sg U59217 ( .A(n45451), .B(n11602), .X(n11600) );
  nor_x1_sg U59218 ( .A(n45447), .B(n14714), .X(n14712) );
  nand_x1_sg U59219 ( .A(n41728), .B(n42302), .X(n10381) );
  nand_x1_sg U59220 ( .A(n51655), .B(n51656), .X(n11148) );
  nand_x1_sg U59221 ( .A(n51936), .B(n51937), .X(n11931) );
  nand_x1_sg U59222 ( .A(n52211), .B(n52212), .X(n12709) );
  nand_x1_sg U59223 ( .A(n52488), .B(n52489), .X(n13493) );
  nand_x1_sg U59224 ( .A(n42320), .B(n52775), .X(n14273) );
  nand_x1_sg U59225 ( .A(n53045), .B(n53046), .X(n15042) );
  nand_x1_sg U59226 ( .A(n53324), .B(n53325), .X(n15826) );
  nand_x1_sg U59227 ( .A(n53603), .B(n53604), .X(n16608) );
  nand_x1_sg U59228 ( .A(n42318), .B(n53895), .X(n17392) );
  nand_x1_sg U59229 ( .A(n41730), .B(n42304), .X(n18163) );
  nand_x1_sg U59230 ( .A(n42316), .B(n54460), .X(n18937) );
  nand_x1_sg U59231 ( .A(n42308), .B(n54742), .X(n19708) );
  nand_x1_sg U59232 ( .A(n42314), .B(n55028), .X(n20481) );
  nand_x1_sg U59233 ( .A(n42306), .B(n55310), .X(n21253) );
  nand_x4_sg U59234 ( .A(n16223), .B(n16217), .X(n15817) );
  nand_x4_sg U59235 ( .A(n10766), .B(n10760), .X(n10371) );
  nand_x4_sg U59236 ( .A(n11141), .B(n11142), .X(n11113) );
  nand_x1_sg U59237 ( .A(n11109), .B(n11110), .X(n11141) );
  nand_x4_sg U59238 ( .A(n12702), .B(n12703), .X(n12674) );
  nand_x1_sg U59239 ( .A(n12670), .B(n12671), .X(n12702) );
  nand_x4_sg U59240 ( .A(n15035), .B(n15036), .X(n15007) );
  nand_x1_sg U59241 ( .A(n15003), .B(n15004), .X(n15035) );
  nand_x4_sg U59242 ( .A(n16601), .B(n16602), .X(n16573) );
  nand_x1_sg U59243 ( .A(n16569), .B(n16570), .X(n16601) );
  nand_x4_sg U59244 ( .A(n10378), .B(n10379), .X(n10337) );
  nand_x1_sg U59245 ( .A(n10333), .B(n10334), .X(n10379) );
  nand_x4_sg U59246 ( .A(n14270), .B(n14271), .X(n14229) );
  nand_x1_sg U59247 ( .A(n14225), .B(n14226), .X(n14271) );
  nand_x4_sg U59248 ( .A(n17389), .B(n17390), .X(n17348) );
  nand_x1_sg U59249 ( .A(n17344), .B(n17345), .X(n17390) );
  nand_x4_sg U59250 ( .A(n18160), .B(n18161), .X(n18120) );
  nand_x1_sg U59251 ( .A(n18116), .B(n18117), .X(n18161) );
  nand_x4_sg U59252 ( .A(n18934), .B(n18935), .X(n18893) );
  nand_x1_sg U59253 ( .A(n18889), .B(n18890), .X(n18935) );
  nand_x4_sg U59254 ( .A(n19705), .B(n19706), .X(n19665) );
  nand_x1_sg U59255 ( .A(n19661), .B(n19662), .X(n19706) );
  nand_x4_sg U59256 ( .A(n20478), .B(n20479), .X(n20437) );
  nand_x1_sg U59257 ( .A(n20433), .B(n20434), .X(n20479) );
  nand_x4_sg U59258 ( .A(n21250), .B(n21251), .X(n21210) );
  nand_x1_sg U59259 ( .A(n21206), .B(n21207), .X(n21251) );
  nor_x1_sg U59260 ( .A(n10320), .B(n41451), .X(n10319) );
  nor_x1_sg U59261 ( .A(n11871), .B(n41465), .X(n11870) );
  nor_x1_sg U59262 ( .A(n15766), .B(n41449), .X(n15765) );
  nor_x1_sg U59263 ( .A(n19648), .B(n41455), .X(n19647) );
  nor_x1_sg U59264 ( .A(n21193), .B(n41453), .X(n21192) );
  nand_x4_sg U59265 ( .A(n10624), .B(n10625), .X(n10338) );
  nand_x1_sg U59266 ( .A(n51426), .B(n10376), .X(n10625) );
  nand_x4_sg U59267 ( .A(n14516), .B(n14517), .X(n14230) );
  nand_x1_sg U59268 ( .A(n52816), .B(n14268), .X(n14517) );
  nand_x4_sg U59269 ( .A(n17637), .B(n17638), .X(n17349) );
  nand_x1_sg U59270 ( .A(n53936), .B(n17387), .X(n17638) );
  nand_x4_sg U59271 ( .A(n18406), .B(n18407), .X(n18121) );
  nand_x1_sg U59272 ( .A(n54216), .B(n18158), .X(n18407) );
  nand_x4_sg U59273 ( .A(n19182), .B(n19183), .X(n18894) );
  nand_x1_sg U59274 ( .A(n54501), .B(n18932), .X(n19183) );
  nand_x4_sg U59275 ( .A(n19951), .B(n19952), .X(n19666) );
  nand_x1_sg U59276 ( .A(n54785), .B(n19703), .X(n19952) );
  nand_x4_sg U59277 ( .A(n20726), .B(n20727), .X(n20438) );
  nand_x1_sg U59278 ( .A(n55069), .B(n20476), .X(n20727) );
  nand_x4_sg U59279 ( .A(n21496), .B(n21497), .X(n21211) );
  nand_x1_sg U59280 ( .A(n55353), .B(n21248), .X(n21497) );
  nand_x4_sg U59281 ( .A(n10714), .B(n10715), .X(n10346) );
  nand_x1_sg U59282 ( .A(n51471), .B(n10716), .X(n10715) );
  nand_x4_sg U59283 ( .A(n11495), .B(n11496), .X(n11114) );
  nand_x1_sg U59284 ( .A(n51751), .B(n43277), .X(n11496) );
  nand_x4_sg U59285 ( .A(n12275), .B(n12276), .X(n11897) );
  nand_x1_sg U59286 ( .A(n52034), .B(n42379), .X(n12276) );
  nand_x4_sg U59287 ( .A(n13056), .B(n13057), .X(n12675) );
  nand_x1_sg U59288 ( .A(n52309), .B(n43275), .X(n13057) );
  nand_x4_sg U59289 ( .A(n14606), .B(n14607), .X(n14238) );
  nand_x1_sg U59290 ( .A(n52860), .B(n43295), .X(n14607) );
  nand_x4_sg U59291 ( .A(n15389), .B(n15390), .X(n15008) );
  nand_x1_sg U59292 ( .A(n53143), .B(n43271), .X(n15390) );
  nand_x4_sg U59293 ( .A(n16170), .B(n16171), .X(n15792) );
  nand_x1_sg U59294 ( .A(n53420), .B(n43267), .X(n16171) );
  nand_x4_sg U59295 ( .A(n16955), .B(n16956), .X(n16574) );
  nand_x1_sg U59296 ( .A(n53701), .B(n43269), .X(n16956) );
  nand_x4_sg U59297 ( .A(n17727), .B(n17728), .X(n17357) );
  nand_x1_sg U59298 ( .A(n53980), .B(n43293), .X(n17728) );
  nand_x4_sg U59299 ( .A(n18496), .B(n18497), .X(n18129) );
  nand_x1_sg U59300 ( .A(n54264), .B(n42377), .X(n18497) );
  nand_x4_sg U59301 ( .A(n19272), .B(n19273), .X(n18902) );
  nand_x1_sg U59302 ( .A(n54545), .B(n43291), .X(n19273) );
  nand_x4_sg U59303 ( .A(n20041), .B(n20042), .X(n19674) );
  nand_x1_sg U59304 ( .A(n54831), .B(n42375), .X(n20042) );
  nand_x4_sg U59305 ( .A(n20816), .B(n20817), .X(n20446) );
  nand_x1_sg U59306 ( .A(n55113), .B(n43289), .X(n20817) );
  nand_x4_sg U59307 ( .A(n21586), .B(n21587), .X(n21219) );
  nand_x1_sg U59308 ( .A(n55399), .B(n42373), .X(n21587) );
  nand_x4_sg U59309 ( .A(n10372), .B(n10343), .X(n10349) );
  nand_x1_sg U59310 ( .A(n10716), .B(n10717), .X(n10372) );
  nand_x4_sg U59311 ( .A(n15818), .B(n15789), .X(n15795) );
  nand_x1_sg U59312 ( .A(n43267), .B(n16173), .X(n15818) );
  nand_x4_sg U59313 ( .A(n16279), .B(n53457), .X(n16277) );
  nand_x1_sg U59314 ( .A(n42765), .B(n15811), .X(n16279) );
  nor_x1_sg U59315 ( .A(n15811), .B(n42765), .X(n16280) );
  nand_x4_sg U59316 ( .A(n11603), .B(n51787), .X(n11602) );
  nand_x1_sg U59317 ( .A(n41919), .B(n11132), .X(n11603) );
  nor_x1_sg U59318 ( .A(n11132), .B(n41919), .X(n11604) );
  nand_x4_sg U59319 ( .A(n18603), .B(n54299), .X(n18602) );
  nand_x1_sg U59320 ( .A(n41903), .B(n18146), .X(n18603) );
  nor_x1_sg U59321 ( .A(n18146), .B(n41903), .X(n18604) );
  nand_x4_sg U59322 ( .A(n20149), .B(n54867), .X(n20148) );
  nand_x1_sg U59323 ( .A(n41897), .B(n19691), .X(n20149) );
  nor_x1_sg U59324 ( .A(n19691), .B(n41897), .X(n20150) );
  nand_x4_sg U59325 ( .A(n21694), .B(n55435), .X(n21693) );
  nand_x1_sg U59326 ( .A(n41891), .B(n21236), .X(n21694) );
  nor_x1_sg U59327 ( .A(n21236), .B(n41891), .X(n21695) );
  nand_x4_sg U59328 ( .A(n13890), .B(n52580), .X(n13885) );
  nand_x1_sg U59329 ( .A(n52575), .B(n13892), .X(n13890) );
  nor_x1_sg U59330 ( .A(n13892), .B(n52575), .X(n13891) );
  nand_x4_sg U59331 ( .A(n10325), .B(n10326), .X(n9024) );
  nor_x1_sg U59332 ( .A(n41729), .B(n42303), .X(n10327) );
  nand_x4_sg U59333 ( .A(n11093), .B(n11094), .X(n8866) );
  nor_x1_sg U59334 ( .A(n11097), .B(n11098), .X(n11095) );
  nand_x4_sg U59335 ( .A(n11876), .B(n11877), .X(n8905) );
  nor_x1_sg U59336 ( .A(n11880), .B(n11881), .X(n11878) );
  nand_x4_sg U59337 ( .A(n12654), .B(n12655), .X(n8828) );
  nor_x1_sg U59338 ( .A(n12658), .B(n12659), .X(n12656) );
  nand_x4_sg U59339 ( .A(n13438), .B(n13439), .X(n8807) );
  nor_x1_sg U59340 ( .A(n13442), .B(n13443), .X(n13440) );
  nand_x4_sg U59341 ( .A(n14217), .B(n14218), .X(n8944) );
  nor_x1_sg U59342 ( .A(n42321), .B(n14222), .X(n14219) );
  nand_x4_sg U59343 ( .A(n14987), .B(n14988), .X(n8967) );
  nor_x1_sg U59344 ( .A(n14991), .B(n14992), .X(n14989) );
  nand_x4_sg U59345 ( .A(n15771), .B(n15772), .X(n9330) );
  nor_x1_sg U59346 ( .A(n15775), .B(n15776), .X(n15773) );
  nand_x4_sg U59347 ( .A(n16553), .B(n16554), .X(n9284) );
  nor_x1_sg U59348 ( .A(n16557), .B(n16558), .X(n16555) );
  nand_x4_sg U59349 ( .A(n17336), .B(n17337), .X(n9246) );
  nor_x1_sg U59350 ( .A(n42319), .B(n17341), .X(n17338) );
  nand_x4_sg U59351 ( .A(n18108), .B(n18109), .X(n9073) );
  nor_x1_sg U59352 ( .A(n41731), .B(n42305), .X(n18110) );
  nand_x4_sg U59353 ( .A(n18881), .B(n18882), .X(n9208) );
  nor_x1_sg U59354 ( .A(n42317), .B(n18886), .X(n18883) );
  nand_x4_sg U59355 ( .A(n19653), .B(n19654), .X(n9187) );
  nor_x1_sg U59356 ( .A(n42309), .B(n19658), .X(n19655) );
  nand_x4_sg U59357 ( .A(n20425), .B(n20426), .X(n9132) );
  nor_x1_sg U59358 ( .A(n42315), .B(n20430), .X(n20427) );
  nand_x4_sg U59359 ( .A(n21198), .B(n21199), .X(n9113) );
  nor_x1_sg U59360 ( .A(n42307), .B(n21203), .X(n21200) );
  nand_x4_sg U59361 ( .A(n10351), .B(n51522), .X(n9014) );
  nand_x1_sg U59362 ( .A(n10354), .B(n42931), .X(n10351) );
  nor_x1_sg U59363 ( .A(n42931), .B(n10354), .X(n10352) );
  nand_x4_sg U59364 ( .A(n11118), .B(n51803), .X(n8895) );
  nand_x1_sg U59365 ( .A(n11121), .B(n42927), .X(n11118) );
  nor_x1_sg U59366 ( .A(n42927), .B(n11121), .X(n11119) );
  nand_x4_sg U59367 ( .A(n11901), .B(n52079), .X(n8929) );
  nand_x1_sg U59368 ( .A(n11904), .B(n42024), .X(n11901) );
  nor_x1_sg U59369 ( .A(n42024), .B(n11904), .X(n11902) );
  nand_x4_sg U59370 ( .A(n12679), .B(n52357), .X(n8859) );
  nand_x1_sg U59371 ( .A(n12682), .B(n42020), .X(n12679) );
  nor_x1_sg U59372 ( .A(n42020), .B(n12682), .X(n12680) );
  nand_x4_sg U59373 ( .A(n13463), .B(n52632), .X(n8821) );
  nand_x1_sg U59374 ( .A(n13466), .B(n42016), .X(n13463) );
  nor_x1_sg U59375 ( .A(n42016), .B(n13466), .X(n13464) );
  nand_x4_sg U59376 ( .A(n14242), .B(n52913), .X(n9009) );
  nand_x1_sg U59377 ( .A(n14245), .B(n42923), .X(n14242) );
  nor_x1_sg U59378 ( .A(n42923), .B(n14245), .X(n14243) );
  nand_x4_sg U59379 ( .A(n15012), .B(n53191), .X(n8998) );
  nand_x1_sg U59380 ( .A(n15015), .B(n42012), .X(n15012) );
  nor_x1_sg U59381 ( .A(n42012), .B(n15015), .X(n15013) );
  nand_x4_sg U59382 ( .A(n15797), .B(n53471), .X(n9324) );
  nand_x1_sg U59383 ( .A(n15800), .B(n42919), .X(n15797) );
  nor_x1_sg U59384 ( .A(n42919), .B(n15800), .X(n15798) );
  nand_x4_sg U59385 ( .A(n16578), .B(n53749), .X(n9315) );
  nand_x1_sg U59386 ( .A(n16581), .B(n42008), .X(n16578) );
  nor_x1_sg U59387 ( .A(n42008), .B(n16581), .X(n16579) );
  nand_x4_sg U59388 ( .A(n17361), .B(n54033), .X(n9275) );
  nand_x1_sg U59389 ( .A(n17364), .B(n42915), .X(n17361) );
  nor_x1_sg U59390 ( .A(n42915), .B(n17364), .X(n17362) );
  nand_x4_sg U59391 ( .A(n18133), .B(n54314), .X(n9087) );
  nand_x1_sg U59392 ( .A(n18136), .B(n42911), .X(n18133) );
  nor_x1_sg U59393 ( .A(n42911), .B(n18136), .X(n18134) );
  nand_x4_sg U59394 ( .A(n18906), .B(n54598), .X(n9237) );
  nand_x1_sg U59395 ( .A(n18909), .B(n42907), .X(n18906) );
  nor_x1_sg U59396 ( .A(n42907), .B(n18909), .X(n18907) );
  nand_x4_sg U59397 ( .A(n19678), .B(n54882), .X(n9179) );
  nand_x1_sg U59398 ( .A(n19681), .B(n42903), .X(n19678) );
  nor_x1_sg U59399 ( .A(n42903), .B(n19681), .X(n19679) );
  nand_x4_sg U59400 ( .A(n20450), .B(n55166), .X(n9161) );
  nand_x1_sg U59401 ( .A(n20453), .B(n42899), .X(n20450) );
  nor_x1_sg U59402 ( .A(n42899), .B(n20453), .X(n20451) );
  nand_x4_sg U59403 ( .A(n21223), .B(n55450), .X(n9099) );
  nand_x1_sg U59404 ( .A(n21226), .B(n42895), .X(n21223) );
  nor_x1_sg U59405 ( .A(n42895), .B(n21226), .X(n21224) );
  nand_x4_sg U59406 ( .A(n11143), .B(n11144), .X(n11110) );
  nand_x1_sg U59407 ( .A(n11105), .B(n11106), .X(n11143) );
  nand_x4_sg U59408 ( .A(n11926), .B(n11927), .X(n11893) );
  nand_x1_sg U59409 ( .A(n11888), .B(n11889), .X(n11926) );
  nand_x4_sg U59410 ( .A(n12704), .B(n12705), .X(n12671) );
  nand_x1_sg U59411 ( .A(n12666), .B(n12667), .X(n12704) );
  nand_x4_sg U59412 ( .A(n15037), .B(n15038), .X(n15004) );
  nand_x1_sg U59413 ( .A(n14999), .B(n15000), .X(n15037) );
  nand_x4_sg U59414 ( .A(n15821), .B(n15822), .X(n15788) );
  nand_x1_sg U59415 ( .A(n15783), .B(n15784), .X(n15821) );
  nand_x4_sg U59416 ( .A(n16603), .B(n16604), .X(n16570) );
  nand_x1_sg U59417 ( .A(n16565), .B(n16566), .X(n16603) );
  nand_x4_sg U59418 ( .A(n11145), .B(n11146), .X(n11106) );
  nand_x1_sg U59419 ( .A(n11101), .B(n11102), .X(n11146) );
  nand_x4_sg U59420 ( .A(n11928), .B(n11929), .X(n11889) );
  nand_x1_sg U59421 ( .A(n11884), .B(n11885), .X(n11929) );
  nand_x4_sg U59422 ( .A(n12706), .B(n12707), .X(n12667) );
  nand_x1_sg U59423 ( .A(n12662), .B(n12663), .X(n12707) );
  nand_x4_sg U59424 ( .A(n13490), .B(n13491), .X(n13451) );
  nand_x1_sg U59425 ( .A(n13446), .B(n13447), .X(n13491) );
  nand_x4_sg U59426 ( .A(n15039), .B(n15040), .X(n15000) );
  nand_x1_sg U59427 ( .A(n14995), .B(n14996), .X(n15040) );
  nand_x4_sg U59428 ( .A(n15823), .B(n15824), .X(n15784) );
  nand_x1_sg U59429 ( .A(n15779), .B(n15780), .X(n15824) );
  nand_x4_sg U59430 ( .A(n16605), .B(n16606), .X(n16566) );
  nand_x1_sg U59431 ( .A(n16561), .B(n16562), .X(n16606) );
  nand_x4_sg U59432 ( .A(n11548), .B(n11542), .X(n11547) );
  nand_x4_sg U59433 ( .A(n13109), .B(n13103), .X(n13108) );
  nand_x4_sg U59434 ( .A(n13889), .B(n13883), .X(n13888) );
  nand_x4_sg U59435 ( .A(n14658), .B(n14652), .X(n14657) );
  nand_x4_sg U59436 ( .A(n15442), .B(n15436), .X(n15441) );
  nand_x4_sg U59437 ( .A(n17008), .B(n17002), .X(n17007) );
  nand_x4_sg U59438 ( .A(n17779), .B(n17773), .X(n17778) );
  nand_x4_sg U59439 ( .A(n18547), .B(n18541), .X(n18546) );
  nand_x4_sg U59440 ( .A(n19324), .B(n19318), .X(n19323) );
  nand_x4_sg U59441 ( .A(n20092), .B(n20086), .X(n20091) );
  nand_x4_sg U59442 ( .A(n20868), .B(n20862), .X(n20867) );
  nand_x4_sg U59443 ( .A(n21637), .B(n21631), .X(n21636) );
  nand_x4_sg U59444 ( .A(n13849), .B(n13802), .X(n13847) );
  nand_x4_sg U59445 ( .A(n10763), .B(n10764), .X(n10350) );
  nand_x1_sg U59446 ( .A(n51497), .B(n51509), .X(n10764) );
  nand_x4_sg U59447 ( .A(n16220), .B(n16221), .X(n15796) );
  nand_x1_sg U59448 ( .A(n53445), .B(n53459), .X(n16221) );
  nand_x4_sg U59449 ( .A(n13498), .B(n13419), .X(n13425) );
  nand_x4_sg U59450 ( .A(n10335), .B(n10375), .X(n10342) );
  nand_x1_sg U59451 ( .A(n10376), .B(n10377), .X(n10375) );
  nand_x4_sg U59452 ( .A(n14227), .B(n14267), .X(n14234) );
  nand_x1_sg U59453 ( .A(n14268), .B(n14269), .X(n14267) );
  nand_x4_sg U59454 ( .A(n17346), .B(n17386), .X(n17353) );
  nand_x1_sg U59455 ( .A(n17387), .B(n17388), .X(n17386) );
  nand_x4_sg U59456 ( .A(n18118), .B(n18157), .X(n18125) );
  nand_x1_sg U59457 ( .A(n18158), .B(n18159), .X(n18157) );
  nand_x4_sg U59458 ( .A(n18891), .B(n18931), .X(n18898) );
  nand_x1_sg U59459 ( .A(n18932), .B(n18933), .X(n18931) );
  nand_x4_sg U59460 ( .A(n19663), .B(n19702), .X(n19670) );
  nand_x1_sg U59461 ( .A(n19703), .B(n19704), .X(n19702) );
  nand_x4_sg U59462 ( .A(n20435), .B(n20475), .X(n20442) );
  nand_x1_sg U59463 ( .A(n20476), .B(n20477), .X(n20475) );
  nand_x4_sg U59464 ( .A(n21208), .B(n21247), .X(n21215) );
  nand_x1_sg U59465 ( .A(n21248), .B(n21249), .X(n21247) );
  nand_x4_sg U59466 ( .A(n12336), .B(n12281), .X(n12334) );
  nand_x4_sg U59467 ( .A(n13745), .B(n13744), .X(n13489) );
  nand_x4_sg U59468 ( .A(n12235), .B(n12234), .X(n11925) );
  nand_x4_sg U59469 ( .A(n13796), .B(n13795), .X(n13487) );
  nand_x4_sg U59470 ( .A(n16130), .B(n16129), .X(n15820) );
  nand_x4_sg U59471 ( .A(n18457), .B(n18456), .X(n18156) );
  nand_x4_sg U59472 ( .A(n10675), .B(n10674), .X(n10374) );
  nand_x4_sg U59473 ( .A(n14567), .B(n14566), .X(n14266) );
  nand_x4_sg U59474 ( .A(n17688), .B(n17687), .X(n17385) );
  nand_x4_sg U59475 ( .A(n19233), .B(n19232), .X(n18930) );
  nand_x4_sg U59476 ( .A(n20002), .B(n20001), .X(n19701) );
  nand_x4_sg U59477 ( .A(n20777), .B(n20776), .X(n20474) );
  nand_x4_sg U59478 ( .A(n21547), .B(n21546), .X(n21246) );
  nand_x1_sg U59479 ( .A(n41994), .B(n46510), .X(n8854) );
  nand_x1_sg U59480 ( .A(n42883), .B(n46510), .X(n8850) );
  nand_x1_sg U59481 ( .A(n44128), .B(n46510), .X(n8839) );
  nand_x1_sg U59482 ( .A(n44126), .B(n46510), .X(n8825) );
  nand_x1_sg U59483 ( .A(n41990), .B(n46487), .X(n8816) );
  nand_x1_sg U59484 ( .A(n42881), .B(n46487), .X(n8810) );
  nand_x1_sg U59485 ( .A(n44124), .B(n46487), .X(n8794) );
  nand_x1_sg U59486 ( .A(n44122), .B(n46487), .X(n8790) );
  nand_x1_sg U59487 ( .A(n41966), .B(n46263), .X(n9120) );
  nand_x1_sg U59488 ( .A(n42857), .B(n46263), .X(n9104) );
  nand_x1_sg U59489 ( .A(n44387), .B(n46263), .X(n9124) );
  nand_x1_sg U59490 ( .A(n41974), .B(n46375), .X(n9270) );
  nand_x1_sg U59491 ( .A(n42867), .B(n46375), .X(n9266) );
  nand_x1_sg U59492 ( .A(n44397), .B(n46375), .X(n9243) );
  nand_x1_sg U59493 ( .A(n42002), .B(n46553), .X(n8890) );
  nand_x1_sg U59494 ( .A(n42889), .B(n46553), .X(n8883) );
  nand_x1_sg U59495 ( .A(n44136), .B(n46553), .X(n8877) );
  nand_x1_sg U59496 ( .A(n44134), .B(n46553), .X(n8863) );
  nand_x1_sg U59497 ( .A(n11276), .B(n11277), .X(n11275) );
  nand_x1_sg U59498 ( .A(n12055), .B(n12056), .X(n12054) );
  nand_x1_sg U59499 ( .A(n12837), .B(n12838), .X(n12836) );
  nand_x1_sg U59500 ( .A(n15170), .B(n15171), .X(n15169) );
  nand_x1_sg U59501 ( .A(n15950), .B(n15951), .X(n15949) );
  nand_x1_sg U59502 ( .A(n16736), .B(n16737), .X(n16735) );
  nand_x1_sg U59503 ( .A(n10502), .B(n10503), .X(n10501) );
  nand_x1_sg U59504 ( .A(n14393), .B(n14394), .X(n14392) );
  nand_x1_sg U59505 ( .A(n18283), .B(n18284), .X(n18282) );
  nand_x1_sg U59506 ( .A(n19829), .B(n19830), .X(n19828) );
  nand_x1_sg U59507 ( .A(n21374), .B(n21375), .X(n21373) );
  nand_x1_sg U59508 ( .A(n41764), .B(n41530), .X(n20186) );
  nand_x1_sg U59509 ( .A(n41762), .B(n41528), .X(n21731) );
  nand_x1_sg U59510 ( .A(n41742), .B(n41526), .X(n10860) );
  nor_x1_sg U59511 ( .A(n11084), .B(n51604), .X(n11082) );
  nand_x1_sg U59512 ( .A(n51604), .B(n11084), .X(n11083) );
  nor_x1_sg U59513 ( .A(n11867), .B(n51885), .X(n11865) );
  nand_x1_sg U59514 ( .A(n51885), .B(n11867), .X(n11866) );
  nor_x1_sg U59515 ( .A(n12645), .B(n52162), .X(n12643) );
  nand_x1_sg U59516 ( .A(n52162), .B(n12645), .X(n12644) );
  nor_x1_sg U59517 ( .A(n13429), .B(n52436), .X(n13427) );
  nand_x1_sg U59518 ( .A(n52436), .B(n13429), .X(n13428) );
  nand_x1_sg U59519 ( .A(n52719), .B(n14208), .X(n14207) );
  nor_x1_sg U59520 ( .A(n14978), .B(n52996), .X(n14976) );
  nand_x1_sg U59521 ( .A(n52996), .B(n14978), .X(n14977) );
  nor_x1_sg U59522 ( .A(n15762), .B(n53272), .X(n15760) );
  nand_x1_sg U59523 ( .A(n53272), .B(n15762), .X(n15761) );
  nor_x1_sg U59524 ( .A(n16544), .B(n53554), .X(n16542) );
  nand_x1_sg U59525 ( .A(n53554), .B(n16544), .X(n16543) );
  nand_x1_sg U59526 ( .A(n53833), .B(n17327), .X(n17326) );
  nand_x1_sg U59527 ( .A(n54120), .B(n18099), .X(n18098) );
  nand_x1_sg U59528 ( .A(n54398), .B(n18872), .X(n18871) );
  nand_x1_sg U59529 ( .A(n54966), .B(n20416), .X(n20415) );
  nand_x1_sg U59530 ( .A(n14447), .B(n14448), .X(n14446) );
  nand_x1_sg U59531 ( .A(n18337), .B(n18338), .X(n18336) );
  nand_x1_sg U59532 ( .A(n19882), .B(n19883), .X(n19881) );
  nand_x1_sg U59533 ( .A(n21427), .B(n21428), .X(n21426) );
  nor_x1_sg U59534 ( .A(n41494), .B(n13224), .X(n13222) );
  nor_x1_sg U59535 ( .A(n41492), .B(n15557), .X(n15555) );
  nor_x1_sg U59536 ( .A(n41490), .B(n17123), .X(n17121) );
  nor_x1_sg U59537 ( .A(n41426), .B(n11711), .X(n11709) );
  nand_x1_sg U59538 ( .A(n11711), .B(n41426), .X(n11710) );
  nor_x1_sg U59539 ( .A(n41424), .B(n12491), .X(n12489) );
  nand_x1_sg U59540 ( .A(n12491), .B(n41424), .X(n12490) );
  nor_x1_sg U59541 ( .A(n41422), .B(n13272), .X(n13270) );
  nand_x1_sg U59542 ( .A(n13272), .B(n41422), .X(n13271) );
  nor_x1_sg U59543 ( .A(n41420), .B(n14052), .X(n14050) );
  nand_x1_sg U59544 ( .A(n14052), .B(n41420), .X(n14051) );
  nor_x1_sg U59545 ( .A(n41416), .B(n15605), .X(n15603) );
  nand_x1_sg U59546 ( .A(n15605), .B(n41416), .X(n15604) );
  nor_x1_sg U59547 ( .A(n41414), .B(n17171), .X(n17169) );
  nand_x1_sg U59548 ( .A(n17171), .B(n41414), .X(n17170) );
  nor_x1_sg U59549 ( .A(n14248), .B(n41388), .X(n14246) );
  nand_x1_sg U59550 ( .A(n41388), .B(n14248), .X(n14247) );
  nor_x1_sg U59551 ( .A(n17367), .B(n41376), .X(n17365) );
  nand_x1_sg U59552 ( .A(n41376), .B(n17367), .X(n17366) );
  nor_x1_sg U59553 ( .A(n18912), .B(n41374), .X(n18910) );
  nand_x1_sg U59554 ( .A(n41374), .B(n18912), .X(n18911) );
  nor_x1_sg U59555 ( .A(n20456), .B(n41370), .X(n20454) );
  nand_x1_sg U59556 ( .A(n41370), .B(n20456), .X(n20455) );
  nor_x1_sg U59557 ( .A(n51764), .B(n11663), .X(n11662) );
  nor_x1_sg U59558 ( .A(n52873), .B(n14775), .X(n14774) );
  nand_x2_sg U59559 ( .A(n10969), .B(n10970), .X(n10968) );
  nand_x1_sg U59560 ( .A(n51485), .B(n10883), .X(n10970) );
  nand_x2_sg U59561 ( .A(n16427), .B(n16428), .X(n16426) );
  nand_x1_sg U59562 ( .A(n53434), .B(n16338), .X(n16428) );
  nand_x2_sg U59563 ( .A(n14865), .B(n14866), .X(n14864) );
  nand_x1_sg U59564 ( .A(n52873), .B(n14775), .X(n14866) );
  nand_x2_sg U59565 ( .A(n17986), .B(n17987), .X(n17985) );
  nand_x1_sg U59566 ( .A(n53993), .B(n17896), .X(n17987) );
  nand_x2_sg U59567 ( .A(n19531), .B(n19532), .X(n19530) );
  nand_x1_sg U59568 ( .A(n54558), .B(n19441), .X(n19532) );
  nand_x2_sg U59569 ( .A(n21075), .B(n21076), .X(n21074) );
  nand_x1_sg U59570 ( .A(n55126), .B(n20985), .X(n21076) );
  nand_x2_sg U59571 ( .A(n11753), .B(n11754), .X(n11752) );
  nand_x1_sg U59572 ( .A(n51764), .B(n11663), .X(n11754) );
  nand_x2_sg U59573 ( .A(n18755), .B(n18756), .X(n18754) );
  nand_x1_sg U59574 ( .A(n54276), .B(n18665), .X(n18756) );
  nand_x2_sg U59575 ( .A(n20301), .B(n20302), .X(n20300) );
  nand_x1_sg U59576 ( .A(n54843), .B(n20210), .X(n20302) );
  nand_x2_sg U59577 ( .A(n21846), .B(n21847), .X(n21845) );
  nand_x1_sg U59578 ( .A(n55411), .B(n21755), .X(n21847) );
  nor_x1_sg U59579 ( .A(n43129), .B(n41830), .X(n11156) );
  nor_x1_sg U59580 ( .A(n43127), .B(n41828), .X(n12717) );
  nand_x4_sg U59581 ( .A(n52488), .B(n13646), .X(n13437) );
  nand_x1_sg U59582 ( .A(n13647), .B(n44703), .X(n13646) );
  nand_x4_sg U59583 ( .A(n41730), .B(n18310), .X(n18107) );
  nand_x1_sg U59584 ( .A(n18311), .B(n43211), .X(n18310) );
  nand_x4_sg U59585 ( .A(n42320), .B(n14420), .X(n14216) );
  nand_x1_sg U59586 ( .A(n14421), .B(n43219), .X(n14420) );
  nand_x4_sg U59587 ( .A(n42318), .B(n17540), .X(n17335) );
  nand_x1_sg U59588 ( .A(n17541), .B(n43217), .X(n17540) );
  nand_x4_sg U59589 ( .A(n42316), .B(n19085), .X(n18880) );
  nand_x1_sg U59590 ( .A(n19086), .B(n43215), .X(n19085) );
  nand_x4_sg U59591 ( .A(n42314), .B(n20629), .X(n20424) );
  nand_x1_sg U59592 ( .A(n20630), .B(n43213), .X(n20629) );
  nand_x4_sg U59593 ( .A(n41728), .B(n10528), .X(n10324) );
  nand_x1_sg U59594 ( .A(n10529), .B(n43205), .X(n10528) );
  nand_x4_sg U59595 ( .A(n51655), .B(n11305), .X(n11092) );
  nand_x1_sg U59596 ( .A(n11306), .B(n44709), .X(n11305) );
  nand_x4_sg U59597 ( .A(n51936), .B(n12085), .X(n11875) );
  nand_x1_sg U59598 ( .A(n12086), .B(n44707), .X(n12085) );
  nand_x4_sg U59599 ( .A(n52211), .B(n12866), .X(n12653) );
  nand_x1_sg U59600 ( .A(n12867), .B(n44705), .X(n12866) );
  nand_x4_sg U59601 ( .A(n53045), .B(n15199), .X(n14986) );
  nand_x1_sg U59602 ( .A(n15200), .B(n44701), .X(n15199) );
  nand_x4_sg U59603 ( .A(n53324), .B(n15980), .X(n15770) );
  nand_x1_sg U59604 ( .A(n15981), .B(n44699), .X(n15980) );
  nand_x4_sg U59605 ( .A(n53603), .B(n16765), .X(n16552) );
  nand_x1_sg U59606 ( .A(n16766), .B(n44697), .X(n16765) );
  nand_x4_sg U59607 ( .A(n42308), .B(n19855), .X(n19652) );
  nand_x1_sg U59608 ( .A(n19856), .B(n43209), .X(n19855) );
  nand_x4_sg U59609 ( .A(n42306), .B(n21400), .X(n21197) );
  nand_x1_sg U59610 ( .A(n21401), .B(n43207), .X(n21400) );
  nand_x4_sg U59611 ( .A(n43167), .B(n12383), .X(n11912) );
  nand_x4_sg U59612 ( .A(n41721), .B(n13943), .X(n13474) );
  nand_x4_sg U59613 ( .A(n45443), .B(n17835), .X(n17372) );
  nand_x4_sg U59614 ( .A(n45439), .B(n18602), .X(n18143) );
  nand_x4_sg U59615 ( .A(n45435), .B(n19380), .X(n18917) );
  nand_x4_sg U59616 ( .A(n45431), .B(n20148), .X(n19688) );
  nand_x4_sg U59617 ( .A(n45427), .B(n20924), .X(n20461) );
  nand_x4_sg U59618 ( .A(n45423), .B(n21693), .X(n21233) );
  nand_x4_sg U59619 ( .A(n41883), .B(n11067), .X(n8874) );
  nand_x1_sg U59620 ( .A(n41830), .B(n43129), .X(n11067) );
  nand_x4_sg U59621 ( .A(n41881), .B(n12628), .X(n8836) );
  nand_x1_sg U59622 ( .A(n41828), .B(n43127), .X(n12628) );
  nand_x1_sg U59623 ( .A(n41826), .B(n43125), .X(n14961) );
  nand_x1_sg U59624 ( .A(n41824), .B(n43123), .X(n16527) );
  nand_x1_sg U59625 ( .A(n51385), .B(n51360), .X(n10600) );
  nand_x1_sg U59626 ( .A(n54173), .B(n54149), .X(n18382) );
  nand_x1_sg U59627 ( .A(n54739), .B(n54714), .X(n19927) );
  nand_x1_sg U59628 ( .A(n55307), .B(n55282), .X(n21472) );
  nand_x1_sg U59629 ( .A(n52772), .B(n52757), .X(n14492) );
  nand_x1_sg U59630 ( .A(n53892), .B(n53877), .X(n17613) );
  nand_x1_sg U59631 ( .A(n54457), .B(n54442), .X(n19158) );
  nand_x1_sg U59632 ( .A(n55025), .B(n55010), .X(n20702) );
  nand_x4_sg U59633 ( .A(n44449), .B(n20864), .X(n20862) );
  nand_x4_sg U59634 ( .A(n10762), .B(n45455), .X(n10760) );
  nand_x4_sg U59635 ( .A(n44455), .B(n14654), .X(n14652) );
  nand_x4_sg U59636 ( .A(n44453), .B(n17775), .X(n17773) );
  nand_x4_sg U59637 ( .A(n44451), .B(n19320), .X(n19318) );
  nor_x1_sg U59638 ( .A(n43167), .B(n12383), .X(n12381) );
  nor_x1_sg U59639 ( .A(n41721), .B(n13943), .X(n13941) );
  nor_x1_sg U59640 ( .A(n45443), .B(n17835), .X(n17833) );
  nor_x1_sg U59641 ( .A(n45439), .B(n18602), .X(n18600) );
  nor_x1_sg U59642 ( .A(n45435), .B(n19380), .X(n19378) );
  nor_x1_sg U59643 ( .A(n45431), .B(n20148), .X(n20146) );
  nor_x1_sg U59644 ( .A(n45427), .B(n20924), .X(n20922) );
  nor_x1_sg U59645 ( .A(n45423), .B(n21693), .X(n21691) );
  nand_x1_sg U59646 ( .A(n51555), .B(n51564), .X(n11155) );
  nand_x1_sg U59647 ( .A(n52112), .B(n52121), .X(n12716) );
  nand_x1_sg U59648 ( .A(n52946), .B(n52955), .X(n15049) );
  nand_x1_sg U59649 ( .A(n53504), .B(n53513), .X(n16615) );
  nand_x4_sg U59650 ( .A(n10628), .B(n51411), .X(n10622) );
  nor_x1_sg U59651 ( .A(n10630), .B(n10631), .X(n10629) );
  nand_x4_sg U59652 ( .A(n18410), .B(n54204), .X(n18404) );
  nor_x1_sg U59653 ( .A(n18412), .B(n18413), .X(n18411) );
  nand_x4_sg U59654 ( .A(n19955), .B(n54772), .X(n19949) );
  nor_x1_sg U59655 ( .A(n19957), .B(n19958), .X(n19956) );
  nand_x4_sg U59656 ( .A(n21500), .B(n55340), .X(n21494) );
  nor_x1_sg U59657 ( .A(n21502), .B(n21503), .X(n21501) );
  nor_x1_sg U59658 ( .A(n9355), .B(n9032), .X(\L2_0/n4120 ) );
  nor_x1_sg U59659 ( .A(n9355), .B(n9028), .X(\L2_0/n4108 ) );
  nor_x1_sg U59660 ( .A(n42006), .B(n9355), .X(\L2_0/n4104 ) );
  nor_x1_sg U59661 ( .A(n9355), .B(n9041), .X(\L2_0/n4100 ) );
  nor_x1_sg U59662 ( .A(n9355), .B(n9039), .X(\L2_0/n4096 ) );
  nor_x1_sg U59663 ( .A(n9355), .B(n9024), .X(\L2_0/n4092 ) );
  nor_x1_sg U59664 ( .A(n42893), .B(n9355), .X(\L2_0/n4088 ) );
  nor_x1_sg U59665 ( .A(n9355), .B(n9020), .X(\L2_0/n4084 ) );
  nor_x1_sg U59666 ( .A(n44401), .B(n9355), .X(\L2_0/n4080 ) );
  nor_x1_sg U59667 ( .A(n9355), .B(n9018), .X(\L2_0/n4076 ) );
  nand_x4_sg U59668 ( .A(n12386), .B(n12387), .X(n11915) );
  nand_x1_sg U59669 ( .A(n43303), .B(n12332), .X(n12387) );
  nand_x4_sg U59670 ( .A(n10729), .B(n10665), .X(n10682) );
  nand_x4_sg U59671 ( .A(n53872), .B(n17536), .X(n17515) );
  nand_x4_sg U59672 ( .A(n54437), .B(n19081), .X(n19060) );
  nand_x4_sg U59673 ( .A(n55005), .B(n20625), .X(n20604) );
  nand_x4_sg U59674 ( .A(n10383), .B(n10384), .X(n10320) );
  nand_x1_sg U59675 ( .A(n51344), .B(n10471), .X(n10383) );
  nand_x1_sg U59676 ( .A(n10316), .B(n10317), .X(n10384) );
  nand_x4_sg U59677 ( .A(n11933), .B(n11934), .X(n11871) );
  nand_x1_sg U59678 ( .A(n51905), .B(n12023), .X(n11933) );
  nand_x1_sg U59679 ( .A(n11867), .B(n11868), .X(n11934) );
  nand_x4_sg U59680 ( .A(n13495), .B(n13496), .X(n13433) );
  nand_x1_sg U59681 ( .A(n52458), .B(n13584), .X(n13495) );
  nand_x1_sg U59682 ( .A(n13429), .B(n13430), .X(n13496) );
  nand_x4_sg U59683 ( .A(n15828), .B(n15829), .X(n15766) );
  nand_x1_sg U59684 ( .A(n53290), .B(n15918), .X(n15828) );
  nand_x1_sg U59685 ( .A(n15762), .B(n15763), .X(n15829) );
  nand_x4_sg U59686 ( .A(n17394), .B(n17395), .X(n17331) );
  nand_x1_sg U59687 ( .A(n53854), .B(n17485), .X(n17394) );
  nand_x1_sg U59688 ( .A(n17327), .B(n17328), .X(n17395) );
  nand_x4_sg U59689 ( .A(n18939), .B(n18940), .X(n18876) );
  nand_x1_sg U59690 ( .A(n54419), .B(n19030), .X(n18939) );
  nand_x1_sg U59691 ( .A(n18872), .B(n18873), .X(n18940) );
  nand_x4_sg U59692 ( .A(n19710), .B(n19711), .X(n19648) );
  nand_x1_sg U59693 ( .A(n54698), .B(n19798), .X(n19710) );
  nand_x1_sg U59694 ( .A(n19644), .B(n19645), .X(n19711) );
  nand_x4_sg U59695 ( .A(n20483), .B(n20484), .X(n20420) );
  nand_x1_sg U59696 ( .A(n54987), .B(n20574), .X(n20483) );
  nand_x1_sg U59697 ( .A(n20416), .B(n20417), .X(n20484) );
  nand_x4_sg U59698 ( .A(n21255), .B(n21256), .X(n21193) );
  nand_x1_sg U59699 ( .A(n55266), .B(n21343), .X(n21255) );
  nand_x1_sg U59700 ( .A(n21189), .B(n21190), .X(n21256) );
  nand_x4_sg U59701 ( .A(n19887), .B(n19888), .X(n19885) );
  nand_x1_sg U59702 ( .A(n19882), .B(n54740), .X(n19887) );
  nand_x4_sg U59703 ( .A(n21432), .B(n21433), .X(n21430) );
  nand_x1_sg U59704 ( .A(n21427), .B(n55308), .X(n21432) );
  nand_x4_sg U59705 ( .A(n52551), .B(n13790), .X(n13745) );
  nand_x1_sg U59706 ( .A(n42795), .B(n13791), .X(n13790) );
  nor_x1_sg U59707 ( .A(n13791), .B(n42795), .X(n13792) );
  nand_x4_sg U59708 ( .A(n13797), .B(n13798), .X(n13795) );
  nand_x1_sg U59709 ( .A(n13791), .B(n42794), .X(n13798) );
  nand_x4_sg U59710 ( .A(n14452), .B(n14453), .X(n14450) );
  nand_x1_sg U59711 ( .A(n14447), .B(n52773), .X(n14452) );
  nand_x4_sg U59712 ( .A(n18342), .B(n18343), .X(n18340) );
  nand_x1_sg U59713 ( .A(n18337), .B(n54174), .X(n18342) );
  nand_x4_sg U59714 ( .A(n52000), .B(n12229), .X(n12184) );
  nand_x1_sg U59715 ( .A(n42799), .B(n12230), .X(n12229) );
  nor_x1_sg U59716 ( .A(n12230), .B(n42799), .X(n12231) );
  nand_x4_sg U59717 ( .A(n12236), .B(n12237), .X(n12234) );
  nand_x1_sg U59718 ( .A(n12230), .B(n42798), .X(n12237) );
  nand_x4_sg U59719 ( .A(n53389), .B(n16124), .X(n16079) );
  nand_x1_sg U59720 ( .A(n42781), .B(n16125), .X(n16124) );
  nor_x1_sg U59721 ( .A(n16125), .B(n42781), .X(n16126) );
  nand_x4_sg U59722 ( .A(n16131), .B(n16132), .X(n16129) );
  nand_x1_sg U59723 ( .A(n16125), .B(n42780), .X(n16132) );
  nor_x1_sg U59724 ( .A(n11088), .B(n41467), .X(n11087) );
  nor_x1_sg U59725 ( .A(n12649), .B(n41463), .X(n12648) );
  nor_x1_sg U59726 ( .A(n13433), .B(n41217), .X(n13432) );
  nor_x1_sg U59727 ( .A(n14212), .B(n41475), .X(n14211) );
  nor_x1_sg U59728 ( .A(n14982), .B(n41461), .X(n14981) );
  nor_x1_sg U59729 ( .A(n16548), .B(n41459), .X(n16547) );
  nor_x1_sg U59730 ( .A(n17331), .B(n41473), .X(n17330) );
  nor_x1_sg U59731 ( .A(n18103), .B(n41457), .X(n18102) );
  nor_x1_sg U59732 ( .A(n18876), .B(n41471), .X(n18875) );
  nor_x1_sg U59733 ( .A(n20420), .B(n41469), .X(n20419) );
  nand_x4_sg U59734 ( .A(n11912), .B(n11913), .X(n11907) );
  nand_x1_sg U59735 ( .A(n43286), .B(n11915), .X(n11913) );
  nand_x4_sg U59736 ( .A(n12690), .B(n12691), .X(n12685) );
  nand_x1_sg U59737 ( .A(n43284), .B(n12693), .X(n12691) );
  nand_x4_sg U59738 ( .A(n13474), .B(n13475), .X(n13469) );
  nand_x1_sg U59739 ( .A(n43282), .B(n13477), .X(n13475) );
  nand_x4_sg U59740 ( .A(n15023), .B(n15024), .X(n15018) );
  nand_x1_sg U59741 ( .A(n43280), .B(n15026), .X(n15024) );
  nand_x4_sg U59742 ( .A(n16589), .B(n16590), .X(n16584) );
  nand_x1_sg U59743 ( .A(n43278), .B(n16592), .X(n16590) );
  nand_x4_sg U59744 ( .A(n18081), .B(n54075), .X(n9063) );
  nor_x1_sg U59745 ( .A(n18083), .B(n43998), .X(n18082) );
  nor_x1_sg U59746 ( .A(n10300), .B(n43111), .X(n10299) );
  nor_x1_sg U59747 ( .A(n14192), .B(n43147), .X(n14191) );
  nor_x1_sg U59748 ( .A(n19628), .B(n43119), .X(n19627) );
  nor_x1_sg U59749 ( .A(n21173), .B(n43115), .X(n21172) );
  nand_x4_sg U59750 ( .A(n10362), .B(n10363), .X(n10357) );
  nand_x1_sg U59751 ( .A(n41920), .B(n10365), .X(n10363) );
  nand_x4_sg U59752 ( .A(n11129), .B(n11130), .X(n11124) );
  nand_x1_sg U59753 ( .A(n41918), .B(n11132), .X(n11130) );
  nand_x4_sg U59754 ( .A(n14253), .B(n14254), .X(n14248) );
  nand_x1_sg U59755 ( .A(n41911), .B(n14256), .X(n14254) );
  nand_x4_sg U59756 ( .A(n15808), .B(n15809), .X(n15803) );
  nand_x1_sg U59757 ( .A(n42764), .B(n15811), .X(n15809) );
  nand_x4_sg U59758 ( .A(n17372), .B(n17373), .X(n17367) );
  nand_x1_sg U59759 ( .A(n41906), .B(n17375), .X(n17373) );
  nand_x4_sg U59760 ( .A(n18143), .B(n18144), .X(n18139) );
  nand_x1_sg U59761 ( .A(n41902), .B(n18146), .X(n18144) );
  nand_x4_sg U59762 ( .A(n18917), .B(n18918), .X(n18912) );
  nand_x1_sg U59763 ( .A(n41898), .B(n18920), .X(n18918) );
  nand_x4_sg U59764 ( .A(n19688), .B(n19689), .X(n19684) );
  nand_x1_sg U59765 ( .A(n41896), .B(n19691), .X(n19689) );
  nand_x4_sg U59766 ( .A(n20461), .B(n20462), .X(n20456) );
  nand_x1_sg U59767 ( .A(n41892), .B(n20464), .X(n20462) );
  nand_x4_sg U59768 ( .A(n21233), .B(n21234), .X(n21229) );
  nand_x1_sg U59769 ( .A(n41890), .B(n21236), .X(n21234) );
  nand_x4_sg U59770 ( .A(n11549), .B(n11550), .X(n11544) );
  nand_x1_sg U59771 ( .A(n51748), .B(n42384), .X(n11550) );
  nand_x4_sg U59772 ( .A(n16227), .B(n16228), .X(n16219) );
  nand_x1_sg U59773 ( .A(n53417), .B(n42380), .X(n16228) );
  nand_x4_sg U59774 ( .A(n18548), .B(n18549), .X(n18543) );
  nand_x1_sg U59775 ( .A(n54261), .B(n43300), .X(n18549) );
  nand_x4_sg U59776 ( .A(n20093), .B(n20094), .X(n20088) );
  nand_x1_sg U59777 ( .A(n54828), .B(n43298), .X(n20094) );
  nand_x4_sg U59778 ( .A(n21638), .B(n21639), .X(n21633) );
  nand_x1_sg U59779 ( .A(n55396), .B(n43296), .X(n21639) );
  nand_x4_sg U59780 ( .A(n12329), .B(n12330), .X(n12324) );
  nand_x1_sg U59781 ( .A(n52030), .B(n43303), .X(n12330) );
  nand_x4_sg U59782 ( .A(n12384), .B(n12385), .X(n12383) );
  nand_x1_sg U59783 ( .A(n52031), .B(n43286), .X(n12385) );
  nand_x4_sg U59784 ( .A(n13164), .B(n13165), .X(n13163) );
  nand_x1_sg U59785 ( .A(n52306), .B(n43284), .X(n13165) );
  nand_x4_sg U59786 ( .A(n13944), .B(n13945), .X(n13943) );
  nand_x1_sg U59787 ( .A(n52581), .B(n43282), .X(n13945) );
  nand_x4_sg U59788 ( .A(n15497), .B(n15498), .X(n15496) );
  nand_x1_sg U59789 ( .A(n53140), .B(n43280), .X(n15498) );
  nand_x4_sg U59790 ( .A(n17063), .B(n17064), .X(n17062) );
  nand_x1_sg U59791 ( .A(n53698), .B(n43278), .X(n17064) );
  nand_x4_sg U59792 ( .A(n52423), .B(n13549), .X(n13498) );
  nand_x4_sg U59793 ( .A(n18458), .B(n18452), .X(n18456) );
  nand_x4_sg U59794 ( .A(n10676), .B(n10670), .X(n10674) );
  nand_x4_sg U59795 ( .A(n14568), .B(n14562), .X(n14566) );
  nand_x4_sg U59796 ( .A(n20003), .B(n19997), .X(n20001) );
  nand_x4_sg U59797 ( .A(n21548), .B(n21542), .X(n21546) );
  nand_x4_sg U59798 ( .A(n17689), .B(n17683), .X(n17687) );
  nand_x4_sg U59799 ( .A(n19234), .B(n19228), .X(n19232) );
  nand_x4_sg U59800 ( .A(n20778), .B(n20772), .X(n20776) );
  nand_x4_sg U59801 ( .A(n51802), .B(n11133), .X(n11121) );
  nand_x1_sg U59802 ( .A(n41661), .B(n42052), .X(n11133) );
  nor_x1_sg U59803 ( .A(n42052), .B(n41661), .X(n11136) );
  nand_x4_sg U59804 ( .A(n52078), .B(n11916), .X(n11904) );
  nand_x1_sg U59805 ( .A(n41659), .B(n42050), .X(n11916) );
  nor_x1_sg U59806 ( .A(n42050), .B(n41659), .X(n11919) );
  nand_x4_sg U59807 ( .A(n52356), .B(n12694), .X(n12682) );
  nand_x1_sg U59808 ( .A(n41392), .B(n42048), .X(n12694) );
  nor_x1_sg U59809 ( .A(n42048), .B(n41392), .X(n12697) );
  nand_x4_sg U59810 ( .A(n52631), .B(n13478), .X(n13466) );
  nand_x1_sg U59811 ( .A(n41193), .B(n42046), .X(n13478) );
  nor_x1_sg U59812 ( .A(n42046), .B(n41193), .X(n13481) );
  nand_x4_sg U59813 ( .A(n52912), .B(n14257), .X(n14245) );
  nand_x1_sg U59814 ( .A(n43951), .B(n42044), .X(n14257) );
  nor_x1_sg U59815 ( .A(n42044), .B(n43951), .X(n14260) );
  nand_x4_sg U59816 ( .A(n53190), .B(n15027), .X(n15015) );
  nand_x1_sg U59817 ( .A(n41384), .B(n42042), .X(n15027) );
  nor_x1_sg U59818 ( .A(n42042), .B(n41384), .X(n15030) );
  nand_x4_sg U59819 ( .A(n53748), .B(n16593), .X(n16581) );
  nand_x1_sg U59820 ( .A(n41378), .B(n42040), .X(n16593) );
  nor_x1_sg U59821 ( .A(n42040), .B(n41378), .X(n16596) );
  nand_x4_sg U59822 ( .A(n54032), .B(n17376), .X(n17364) );
  nand_x1_sg U59823 ( .A(n43949), .B(n42038), .X(n17376) );
  nor_x1_sg U59824 ( .A(n42038), .B(n43949), .X(n17379) );
  nand_x4_sg U59825 ( .A(n54313), .B(n18147), .X(n18136) );
  nand_x1_sg U59826 ( .A(n41657), .B(n42036), .X(n18147) );
  nor_x1_sg U59827 ( .A(n42036), .B(n41657), .X(n18150) );
  nand_x4_sg U59828 ( .A(n54597), .B(n18921), .X(n18909) );
  nand_x1_sg U59829 ( .A(n43947), .B(n42034), .X(n18921) );
  nor_x1_sg U59830 ( .A(n42034), .B(n43947), .X(n18924) );
  nand_x4_sg U59831 ( .A(n54881), .B(n19692), .X(n19681) );
  nand_x1_sg U59832 ( .A(n41655), .B(n42032), .X(n19692) );
  nor_x1_sg U59833 ( .A(n42032), .B(n41655), .X(n19695) );
  nand_x4_sg U59834 ( .A(n55165), .B(n20465), .X(n20453) );
  nand_x1_sg U59835 ( .A(n43945), .B(n42030), .X(n20465) );
  nor_x1_sg U59836 ( .A(n42030), .B(n43945), .X(n20468) );
  nand_x4_sg U59837 ( .A(n55449), .B(n21237), .X(n21226) );
  nand_x1_sg U59838 ( .A(n41653), .B(n42028), .X(n21237) );
  nor_x1_sg U59839 ( .A(n42028), .B(n41653), .X(n21240) );
  nand_x4_sg U59840 ( .A(n10823), .B(n51507), .X(n10821) );
  nand_x1_sg U59841 ( .A(n41921), .B(n10365), .X(n10823) );
  nor_x1_sg U59842 ( .A(n10365), .B(n41921), .X(n10824) );
  nand_x4_sg U59843 ( .A(n14715), .B(n52897), .X(n14714) );
  nand_x1_sg U59844 ( .A(n41912), .B(n14256), .X(n14715) );
  nor_x1_sg U59845 ( .A(n14256), .B(n41912), .X(n14716) );
  nand_x4_sg U59846 ( .A(n17836), .B(n54017), .X(n17835) );
  nand_x1_sg U59847 ( .A(n41907), .B(n17375), .X(n17836) );
  nor_x1_sg U59848 ( .A(n17375), .B(n41907), .X(n17837) );
  nand_x4_sg U59849 ( .A(n19381), .B(n54582), .X(n19380) );
  nand_x1_sg U59850 ( .A(n41899), .B(n18920), .X(n19381) );
  nor_x1_sg U59851 ( .A(n18920), .B(n41899), .X(n19382) );
  nand_x4_sg U59852 ( .A(n20925), .B(n55150), .X(n20924) );
  nand_x1_sg U59853 ( .A(n41893), .B(n20464), .X(n20925) );
  nor_x1_sg U59854 ( .A(n20464), .B(n41893), .X(n20926) );
  nand_x4_sg U59855 ( .A(n13110), .B(n52305), .X(n13105) );
  nand_x1_sg U59856 ( .A(n52300), .B(n13112), .X(n13110) );
  nor_x1_sg U59857 ( .A(n13112), .B(n52300), .X(n13111) );
  nand_x4_sg U59858 ( .A(n15443), .B(n53139), .X(n15438) );
  nand_x1_sg U59859 ( .A(n53134), .B(n15445), .X(n15443) );
  nor_x1_sg U59860 ( .A(n15445), .B(n53134), .X(n15444) );
  nand_x4_sg U59861 ( .A(n17009), .B(n53697), .X(n17004) );
  nand_x1_sg U59862 ( .A(n53692), .B(n17011), .X(n17009) );
  nor_x1_sg U59863 ( .A(n17011), .B(n53692), .X(n17010) );
  nand_x4_sg U59864 ( .A(n13315), .B(n52325), .X(n13224) );
  nand_x1_sg U59865 ( .A(n52324), .B(n13317), .X(n13315) );
  nor_x1_sg U59866 ( .A(n13317), .B(n52324), .X(n13316) );
  nand_x4_sg U59867 ( .A(n14095), .B(n52600), .X(n14004) );
  nand_x1_sg U59868 ( .A(n52599), .B(n14097), .X(n14095) );
  nor_x1_sg U59869 ( .A(n14097), .B(n52599), .X(n14096) );
  nand_x4_sg U59870 ( .A(n15648), .B(n53159), .X(n15557) );
  nand_x1_sg U59871 ( .A(n53158), .B(n15650), .X(n15648) );
  nor_x1_sg U59872 ( .A(n15650), .B(n53158), .X(n15649) );
  nand_x4_sg U59873 ( .A(n17214), .B(n53717), .X(n17123) );
  nand_x1_sg U59874 ( .A(n53716), .B(n17216), .X(n17214) );
  nor_x1_sg U59875 ( .A(n17216), .B(n53716), .X(n17215) );
  nand_x4_sg U59876 ( .A(n11849), .B(n51843), .X(n8909) );
  nor_x1_sg U59877 ( .A(n11851), .B(n11852), .X(n11850) );
  nand_x4_sg U59878 ( .A(n15744), .B(n53229), .X(n9334) );
  nor_x1_sg U59879 ( .A(n15746), .B(n15747), .X(n15745) );
  nand_x4_sg U59880 ( .A(n10620), .B(n51427), .X(n10590) );
  nor_x1_sg U59881 ( .A(n10622), .B(n10623), .X(n10621) );
  nand_x4_sg U59882 ( .A(n12178), .B(n51981), .X(n12147) );
  nor_x1_sg U59883 ( .A(n12180), .B(n12181), .X(n12179) );
  nand_x4_sg U59884 ( .A(n13739), .B(n52532), .X(n13708) );
  nor_x1_sg U59885 ( .A(n13741), .B(n13742), .X(n13740) );
  nand_x4_sg U59886 ( .A(n14512), .B(n52817), .X(n14482) );
  nor_x1_sg U59887 ( .A(n14514), .B(n14515), .X(n14513) );
  nand_x4_sg U59888 ( .A(n16073), .B(n53370), .X(n16042) );
  nor_x1_sg U59889 ( .A(n16075), .B(n16076), .X(n16074) );
  nand_x4_sg U59890 ( .A(n17633), .B(n53937), .X(n17603) );
  nor_x1_sg U59891 ( .A(n17635), .B(n17636), .X(n17634) );
  nand_x4_sg U59892 ( .A(n18402), .B(n54217), .X(n18372) );
  nor_x1_sg U59893 ( .A(n18404), .B(n18405), .X(n18403) );
  nand_x4_sg U59894 ( .A(n19178), .B(n54502), .X(n19148) );
  nor_x1_sg U59895 ( .A(n19180), .B(n19181), .X(n19179) );
  nand_x4_sg U59896 ( .A(n19947), .B(n54786), .X(n19917) );
  nor_x1_sg U59897 ( .A(n19949), .B(n19950), .X(n19948) );
  nand_x4_sg U59898 ( .A(n20722), .B(n55070), .X(n20692) );
  nor_x1_sg U59899 ( .A(n20724), .B(n20725), .X(n20723) );
  nand_x4_sg U59900 ( .A(n21492), .B(n55354), .X(n21462) );
  nor_x1_sg U59901 ( .A(n21494), .B(n21495), .X(n21493) );
  nand_x4_sg U59902 ( .A(n13499), .B(n13415), .X(n13422) );
  nand_x4_sg U59903 ( .A(n12328), .B(n12322), .X(n12327) );
  nand_x4_sg U59904 ( .A(n17321), .B(n53832), .X(n9252) );
  nor_x1_sg U59905 ( .A(n17323), .B(n17324), .X(n17322) );
  nand_x4_sg U59906 ( .A(n18866), .B(n54397), .X(n9214) );
  nor_x1_sg U59907 ( .A(n18868), .B(n18869), .X(n18867) );
  nand_x4_sg U59908 ( .A(n20410), .B(n54965), .X(n9138) );
  nor_x1_sg U59909 ( .A(n20412), .B(n20413), .X(n20411) );
  nand_x4_sg U59910 ( .A(n10366), .B(n51521), .X(n10354) );
  nor_x1_sg U59911 ( .A(n10368), .B(n10369), .X(n10367) );
  nand_x4_sg U59912 ( .A(n15812), .B(n53470), .X(n15800) );
  nor_x1_sg U59913 ( .A(n15814), .B(n15815), .X(n15813) );
  nand_x4_sg U59914 ( .A(n13866), .B(n13867), .X(n13801) );
  nand_x1_sg U59915 ( .A(n52543), .B(n45409), .X(n13867) );
  nand_x1_sg U59916 ( .A(n52548), .B(n44146), .X(n13866) );
  nand_x4_sg U59917 ( .A(n11852), .B(n11851), .X(n11849) );
  nand_x4_sg U59918 ( .A(n15747), .B(n15746), .X(n15744) );
  nand_x4_sg U59919 ( .A(n11078), .B(n51603), .X(n8872) );
  nor_x1_sg U59920 ( .A(n11080), .B(n11081), .X(n11079) );
  nand_x4_sg U59921 ( .A(n11861), .B(n51884), .X(n8907) );
  nor_x1_sg U59922 ( .A(n11863), .B(n11864), .X(n11862) );
  nand_x4_sg U59923 ( .A(n12639), .B(n52161), .X(n8834) );
  nor_x1_sg U59924 ( .A(n12641), .B(n12642), .X(n12640) );
  nand_x4_sg U59925 ( .A(n13423), .B(n52435), .X(n8787) );
  nor_x1_sg U59926 ( .A(n13425), .B(n13426), .X(n13424) );
  nand_x4_sg U59927 ( .A(n14972), .B(n52995), .X(n8973) );
  nor_x1_sg U59928 ( .A(n14974), .B(n14975), .X(n14973) );
  nand_x4_sg U59929 ( .A(n16538), .B(n53553), .X(n9290) );
  nor_x1_sg U59930 ( .A(n16540), .B(n16541), .X(n16539) );
  nand_x4_sg U59931 ( .A(n10310), .B(n51328), .X(n9028) );
  nor_x1_sg U59932 ( .A(n10312), .B(n10313), .X(n10311) );
  nand_x4_sg U59933 ( .A(n14202), .B(n52718), .X(n8948) );
  nor_x1_sg U59934 ( .A(n14204), .B(n14205), .X(n14203) );
  nand_x4_sg U59935 ( .A(n15756), .B(n53271), .X(n9332) );
  nor_x1_sg U59936 ( .A(n15758), .B(n15759), .X(n15757) );
  nand_x4_sg U59937 ( .A(n18093), .B(n54119), .X(n9061) );
  nor_x1_sg U59938 ( .A(n18095), .B(n18096), .X(n18094) );
  nand_x4_sg U59939 ( .A(n19638), .B(n54682), .X(n9193) );
  nor_x1_sg U59940 ( .A(n19640), .B(n19641), .X(n19639) );
  nand_x4_sg U59941 ( .A(n21183), .B(n55250), .X(n9095) );
  nor_x1_sg U59942 ( .A(n21185), .B(n21186), .X(n21184) );
  nand_x4_sg U59943 ( .A(n53328), .B(n16054), .X(n16043) );
  nand_x1_sg U59944 ( .A(n53321), .B(n53313), .X(n16054) );
  nand_x4_sg U59945 ( .A(n51659), .B(n11379), .X(n11368) );
  nand_x1_sg U59946 ( .A(n51652), .B(n51645), .X(n11379) );
  nand_x4_sg U59947 ( .A(n51940), .B(n12159), .X(n12148) );
  nand_x1_sg U59948 ( .A(n51933), .B(n51925), .X(n12159) );
  nand_x4_sg U59949 ( .A(n52215), .B(n12940), .X(n12929) );
  nand_x1_sg U59950 ( .A(n52208), .B(n52201), .X(n12940) );
  nand_x4_sg U59951 ( .A(n53049), .B(n15273), .X(n15262) );
  nand_x1_sg U59952 ( .A(n53042), .B(n53035), .X(n15273) );
  nand_x4_sg U59953 ( .A(n53607), .B(n16839), .X(n16828) );
  nand_x1_sg U59954 ( .A(n53600), .B(n53593), .X(n16839) );
  nand_x1_sg U59955 ( .A(n52665), .B(n52674), .X(n14280) );
  nand_x4_sg U59956 ( .A(n18081), .B(n18170), .X(n18088) );
  nand_x1_sg U59957 ( .A(n54062), .B(n54074), .X(n18170) );
  nand_x1_sg U59958 ( .A(n51276), .B(n51284), .X(n10388) );
  nand_x1_sg U59959 ( .A(n54630), .B(n54638), .X(n19715) );
  nand_x1_sg U59960 ( .A(n55198), .B(n55206), .X(n21260) );
  nand_x4_sg U59961 ( .A(n10710), .B(n10711), .X(n10675) );
  nand_x1_sg U59962 ( .A(n10712), .B(n51451), .X(n10711) );
  nand_x1_sg U59963 ( .A(n10713), .B(n51470), .X(n10710) );
  nand_x4_sg U59964 ( .A(n11491), .B(n11492), .X(n11455) );
  nand_x1_sg U59965 ( .A(n11493), .B(n51730), .X(n11492) );
  nand_x1_sg U59966 ( .A(n11494), .B(n51750), .X(n11491) );
  nand_x4_sg U59967 ( .A(n12271), .B(n12272), .X(n12235) );
  nand_x1_sg U59968 ( .A(n12273), .B(n52008), .X(n12272) );
  nand_x1_sg U59969 ( .A(n12274), .B(n52033), .X(n12271) );
  nand_x4_sg U59970 ( .A(n13052), .B(n13053), .X(n13016) );
  nand_x1_sg U59971 ( .A(n13054), .B(n52286), .X(n13053) );
  nand_x1_sg U59972 ( .A(n13055), .B(n52308), .X(n13052) );
  nand_x4_sg U59973 ( .A(n13832), .B(n13833), .X(n13796) );
  nand_x1_sg U59974 ( .A(n13834), .B(n52561), .X(n13833) );
  nand_x1_sg U59975 ( .A(n13835), .B(n52583), .X(n13832) );
  nand_x4_sg U59976 ( .A(n14602), .B(n14603), .X(n14567) );
  nand_x1_sg U59977 ( .A(n14604), .B(n52842), .X(n14603) );
  nand_x1_sg U59978 ( .A(n14605), .B(n52859), .X(n14602) );
  nand_x4_sg U59979 ( .A(n15385), .B(n15386), .X(n15349) );
  nand_x1_sg U59980 ( .A(n15387), .B(n53120), .X(n15386) );
  nand_x1_sg U59981 ( .A(n15388), .B(n53142), .X(n15385) );
  nand_x4_sg U59982 ( .A(n16166), .B(n16167), .X(n16130) );
  nand_x1_sg U59983 ( .A(n16168), .B(n53399), .X(n16167) );
  nand_x1_sg U59984 ( .A(n16169), .B(n53419), .X(n16166) );
  nand_x4_sg U59985 ( .A(n16951), .B(n16952), .X(n16915) );
  nand_x1_sg U59986 ( .A(n16953), .B(n53678), .X(n16952) );
  nand_x1_sg U59987 ( .A(n16954), .B(n53700), .X(n16951) );
  nand_x4_sg U59988 ( .A(n17723), .B(n17724), .X(n17688) );
  nand_x1_sg U59989 ( .A(n17725), .B(n53962), .X(n17724) );
  nand_x1_sg U59990 ( .A(n17726), .B(n53979), .X(n17723) );
  nand_x4_sg U59991 ( .A(n18492), .B(n18493), .X(n18457) );
  nand_x1_sg U59992 ( .A(n18494), .B(n54244), .X(n18493) );
  nand_x1_sg U59993 ( .A(n18495), .B(n54263), .X(n18492) );
  nand_x4_sg U59994 ( .A(n19268), .B(n19269), .X(n19233) );
  nand_x1_sg U59995 ( .A(n19270), .B(n54527), .X(n19269) );
  nand_x1_sg U59996 ( .A(n19271), .B(n54544), .X(n19268) );
  nand_x4_sg U59997 ( .A(n20037), .B(n20038), .X(n20002) );
  nand_x1_sg U59998 ( .A(n20039), .B(n54812), .X(n20038) );
  nand_x1_sg U59999 ( .A(n20040), .B(n54830), .X(n20037) );
  nand_x4_sg U60000 ( .A(n20812), .B(n20813), .X(n20777) );
  nand_x1_sg U60001 ( .A(n20814), .B(n55095), .X(n20813) );
  nand_x1_sg U60002 ( .A(n20815), .B(n55112), .X(n20812) );
  nand_x4_sg U60003 ( .A(n21582), .B(n21583), .X(n21547) );
  nand_x1_sg U60004 ( .A(n21584), .B(n55380), .X(n21583) );
  nand_x1_sg U60005 ( .A(n21585), .B(n55398), .X(n21582) );
  nor_x1_sg U60006 ( .A(n42851), .B(n10821), .X(n10822) );
  nor_x1_sg U60007 ( .A(n42849), .B(n16277), .X(n16278) );
  nand_x4_sg U60008 ( .A(n10448), .B(n10449), .X(n10313) );
  nand_x4_sg U60009 ( .A(n14340), .B(n14341), .X(n14205) );
  nand_x4_sg U60010 ( .A(n17463), .B(n17464), .X(n17324) );
  nand_x4_sg U60011 ( .A(n19008), .B(n19009), .X(n18869) );
  nand_x4_sg U60012 ( .A(n19775), .B(n19776), .X(n19641) );
  nand_x4_sg U60013 ( .A(n20552), .B(n20553), .X(n20413) );
  nand_x4_sg U60014 ( .A(n21320), .B(n21321), .X(n21186) );
  nand_x4_sg U60015 ( .A(n17787), .B(n17733), .X(n17785) );
  nand_x4_sg U60016 ( .A(n19332), .B(n19278), .X(n19330) );
  nand_x4_sg U60017 ( .A(n20876), .B(n20822), .X(n20874) );
  nand_x4_sg U60018 ( .A(n16231), .B(n16176), .X(n16225) );
  nand_x4_sg U60019 ( .A(n14666), .B(n14612), .X(n14664) );
  nand_x4_sg U60020 ( .A(n52409), .B(n13418), .X(n13415) );
  nand_x4_sg U60021 ( .A(n19859), .B(n19860), .X(n19852) );
  nor_x1_sg U60022 ( .A(n54694), .B(n19863), .X(n19861) );
  nand_x4_sg U60023 ( .A(n21404), .B(n21405), .X(n21397) );
  nor_x1_sg U60024 ( .A(n55262), .B(n21408), .X(n21406) );
  nand_x4_sg U60025 ( .A(n11556), .B(n11501), .X(n11554) );
  nand_x4_sg U60026 ( .A(n14424), .B(n14425), .X(n14417) );
  nor_x1_sg U60027 ( .A(n52730), .B(n14428), .X(n14426) );
  nand_x4_sg U60028 ( .A(n13117), .B(n13062), .X(n13115) );
  nand_x4_sg U60029 ( .A(n13897), .B(n13842), .X(n13895) );
  nand_x4_sg U60030 ( .A(n15450), .B(n15395), .X(n15448) );
  nand_x4_sg U60031 ( .A(n17016), .B(n16961), .X(n17014) );
  nand_x4_sg U60032 ( .A(n18555), .B(n18502), .X(n18553) );
  nand_x4_sg U60033 ( .A(n54811), .B(n20050), .X(n20047) );
  nand_x4_sg U60034 ( .A(n55379), .B(n21595), .X(n21592) );
  nand_x4_sg U60035 ( .A(n52424), .B(n13422), .X(n13419) );
  nand_x4_sg U60036 ( .A(n53398), .B(n16179), .X(n16176) );
  nand_x4_sg U60037 ( .A(n52841), .B(n14615), .X(n14612) );
  nand_x4_sg U60038 ( .A(n13419), .B(n13420), .X(n8801) );
  nand_x4_sg U60039 ( .A(n13415), .B(n13416), .X(n8819) );
  nand_x4_sg U60040 ( .A(n51450), .B(n10723), .X(n10720) );
  nand_x4_sg U60041 ( .A(n51729), .B(n11504), .X(n11501) );
  nand_x4_sg U60042 ( .A(n52007), .B(n12284), .X(n12281) );
  nand_x4_sg U60043 ( .A(n52285), .B(n13065), .X(n13062) );
  nand_x4_sg U60044 ( .A(n53119), .B(n15398), .X(n15395) );
  nand_x4_sg U60045 ( .A(n53677), .B(n16964), .X(n16961) );
  nand_x4_sg U60046 ( .A(n54243), .B(n18505), .X(n18502) );
  nand_x1_sg U60047 ( .A(n14490), .B(n52772), .X(n14489) );
  nor_x1_sg U60048 ( .A(n14491), .B(n52766), .X(n14490) );
  nand_x1_sg U60049 ( .A(n18380), .B(n54173), .X(n18379) );
  nor_x1_sg U60050 ( .A(n18381), .B(n54168), .X(n18380) );
  nand_x1_sg U60051 ( .A(n19925), .B(n54739), .X(n19924) );
  nor_x1_sg U60052 ( .A(n19926), .B(n54734), .X(n19925) );
  nand_x1_sg U60053 ( .A(n21470), .B(n55307), .X(n21469) );
  nor_x1_sg U60054 ( .A(n21471), .B(n55302), .X(n21470) );
  nand_x4_sg U60055 ( .A(n17324), .B(n17323), .X(n17321) );
  nand_x4_sg U60056 ( .A(n18869), .B(n18868), .X(n18866) );
  nand_x4_sg U60057 ( .A(n20413), .B(n20412), .X(n20410) );
  nand_x4_sg U60058 ( .A(n13848), .B(n13847), .X(n13840) );
  nand_x4_sg U60059 ( .A(n11081), .B(n11080), .X(n11078) );
  nand_x4_sg U60060 ( .A(n12642), .B(n12641), .X(n12639) );
  nand_x4_sg U60061 ( .A(n14975), .B(n14974), .X(n14972) );
  nand_x4_sg U60062 ( .A(n16541), .B(n16540), .X(n16538) );
  nand_x4_sg U60063 ( .A(n11864), .B(n11863), .X(n11861) );
  nand_x4_sg U60064 ( .A(n13426), .B(n13425), .X(n13423) );
  nand_x4_sg U60065 ( .A(n15759), .B(n15758), .X(n15756) );
  nand_x4_sg U60066 ( .A(n10313), .B(n10312), .X(n10310) );
  nand_x4_sg U60067 ( .A(n14205), .B(n14204), .X(n14202) );
  nand_x4_sg U60068 ( .A(n18096), .B(n18095), .X(n18093) );
  nand_x4_sg U60069 ( .A(n19641), .B(n19640), .X(n19638) );
  nand_x4_sg U60070 ( .A(n21186), .B(n21185), .X(n21183) );
  nand_x4_sg U60071 ( .A(n12534), .B(n12535), .X(n12443) );
  nand_x4_sg U60072 ( .A(n13746), .B(n13747), .X(n13744) );
  nand_x4_sg U60073 ( .A(n11849), .B(n11938), .X(n11856) );
  nand_x4_sg U60074 ( .A(n15744), .B(n15833), .X(n15751) );
  nand_x4_sg U60075 ( .A(n13840), .B(n52582), .X(n13834) );
  nor_x1_sg U60076 ( .A(n13847), .B(n13848), .X(n13846) );
  nand_x4_sg U60077 ( .A(n12359), .B(n12364), .X(n12336) );
  nand_x4_sg U60078 ( .A(n13919), .B(n13924), .X(n13897) );
  nand_x4_sg U60079 ( .A(n11332), .B(n11331), .X(n11147) );
  nand_x4_sg U60080 ( .A(n12112), .B(n12111), .X(n11930) );
  nand_x4_sg U60081 ( .A(n12893), .B(n12892), .X(n12708) );
  nand_x4_sg U60082 ( .A(n13673), .B(n13672), .X(n13492) );
  nand_x4_sg U60083 ( .A(n15226), .B(n15225), .X(n15041) );
  nand_x4_sg U60084 ( .A(n16007), .B(n16006), .X(n15825) );
  nand_x4_sg U60085 ( .A(n16792), .B(n16791), .X(n16607) );
  nand_x4_sg U60086 ( .A(n10559), .B(n10558), .X(n10380) );
  nand_x4_sg U60087 ( .A(n14451), .B(n14450), .X(n14272) );
  nand_x4_sg U60088 ( .A(n17571), .B(n17570), .X(n17391) );
  nand_x4_sg U60089 ( .A(n18341), .B(n18340), .X(n18162) );
  nand_x4_sg U60090 ( .A(n19116), .B(n19115), .X(n18936) );
  nand_x4_sg U60091 ( .A(n19886), .B(n19885), .X(n19707) );
  nand_x4_sg U60092 ( .A(n20660), .B(n20659), .X(n20480) );
  nand_x4_sg U60093 ( .A(n21431), .B(n21430), .X(n21252) );
  nand_x4_sg U60094 ( .A(n11404), .B(n11403), .X(n11144) );
  nand_x4_sg U60095 ( .A(n12184), .B(n12183), .X(n11927) );
  nand_x4_sg U60096 ( .A(n12965), .B(n12964), .X(n12705) );
  nand_x4_sg U60097 ( .A(n15298), .B(n15297), .X(n15038) );
  nand_x4_sg U60098 ( .A(n16864), .B(n16863), .X(n16604) );
  nand_x4_sg U60099 ( .A(n11455), .B(n11454), .X(n11142) );
  nand_x4_sg U60100 ( .A(n13016), .B(n13015), .X(n12703) );
  nand_x4_sg U60101 ( .A(n15349), .B(n15348), .X(n15036) );
  nand_x4_sg U60102 ( .A(n16915), .B(n16914), .X(n16602) );
  nand_x4_sg U60103 ( .A(n16079), .B(n16078), .X(n15822) );
  nand_x4_sg U60104 ( .A(n10590), .B(n10589), .X(n10378) );
  nand_x4_sg U60105 ( .A(n14482), .B(n14481), .X(n14270) );
  nand_x4_sg U60106 ( .A(n17603), .B(n17602), .X(n17389) );
  nand_x4_sg U60107 ( .A(n18372), .B(n18371), .X(n18160) );
  nand_x4_sg U60108 ( .A(n19148), .B(n19147), .X(n18934) );
  nand_x4_sg U60109 ( .A(n19917), .B(n19916), .X(n19705) );
  nand_x4_sg U60110 ( .A(n20692), .B(n20691), .X(n20478) );
  nand_x4_sg U60111 ( .A(n21462), .B(n21461), .X(n21250) );
  nand_x4_sg U60112 ( .A(n10385), .B(n10310), .X(n10317) );
  nand_x1_sg U60113 ( .A(n51327), .B(n10450), .X(n10385) );
  nand_x4_sg U60114 ( .A(n14277), .B(n14202), .X(n14209) );
  nand_x1_sg U60115 ( .A(n52717), .B(n14342), .X(n14277) );
  nand_x4_sg U60116 ( .A(n17396), .B(n17321), .X(n17328) );
  nand_x1_sg U60117 ( .A(n53831), .B(n17465), .X(n17396) );
  nand_x4_sg U60118 ( .A(n18167), .B(n18093), .X(n18100) );
  nand_x4_sg U60119 ( .A(n18941), .B(n18866), .X(n18873) );
  nand_x1_sg U60120 ( .A(n54396), .B(n19010), .X(n18941) );
  nand_x4_sg U60121 ( .A(n19712), .B(n19638), .X(n19645) );
  nand_x1_sg U60122 ( .A(n54681), .B(n19777), .X(n19712) );
  nand_x4_sg U60123 ( .A(n20485), .B(n20410), .X(n20417) );
  nand_x1_sg U60124 ( .A(n54964), .B(n20554), .X(n20485) );
  nand_x4_sg U60125 ( .A(n21257), .B(n21183), .X(n21190) );
  nand_x1_sg U60126 ( .A(n55249), .B(n21322), .X(n21257) );
  nand_x4_sg U60127 ( .A(n18554), .B(n18553), .X(n18547) );
  nand_x4_sg U60128 ( .A(n11555), .B(n11554), .X(n11548) );
  nand_x4_sg U60129 ( .A(n13116), .B(n13115), .X(n13109) );
  nand_x4_sg U60130 ( .A(n13896), .B(n13895), .X(n13889) );
  nand_x4_sg U60131 ( .A(n15449), .B(n15448), .X(n15442) );
  nand_x4_sg U60132 ( .A(n17015), .B(n17014), .X(n17008) );
  nand_x4_sg U60133 ( .A(n16226), .B(n16225), .X(n16223) );
  nand_x4_sg U60134 ( .A(n13801), .B(n13800), .X(n13802) );
  nand_x4_sg U60135 ( .A(n20099), .B(n20098), .X(n20092) );
  nand_x4_sg U60136 ( .A(n21644), .B(n21643), .X(n21637) );
  nand_x4_sg U60137 ( .A(n17786), .B(n17785), .X(n17779) );
  nand_x4_sg U60138 ( .A(n19331), .B(n19330), .X(n19324) );
  nand_x4_sg U60139 ( .A(n20875), .B(n20874), .X(n20868) );
  nand_x4_sg U60140 ( .A(n14665), .B(n14664), .X(n14658) );
  nand_x4_sg U60141 ( .A(n11367), .B(n11366), .X(n11145) );
  nand_x4_sg U60142 ( .A(n12147), .B(n12146), .X(n11928) );
  nand_x4_sg U60143 ( .A(n12928), .B(n12927), .X(n12706) );
  nand_x4_sg U60144 ( .A(n13708), .B(n13707), .X(n13490) );
  nand_x4_sg U60145 ( .A(n15261), .B(n15260), .X(n15039) );
  nand_x4_sg U60146 ( .A(n16042), .B(n16041), .X(n15823) );
  nand_x4_sg U60147 ( .A(n16827), .B(n16826), .X(n16605) );
  nand_x4_sg U60148 ( .A(n10769), .B(n10768), .X(n10766) );
  nand_x4_sg U60149 ( .A(n11501), .B(n11502), .X(n11494) );
  nand_x4_sg U60150 ( .A(n16176), .B(n16177), .X(n16169) );
  nand_x4_sg U60151 ( .A(n20047), .B(n20048), .X(n20040) );
  nand_x4_sg U60152 ( .A(n21592), .B(n21593), .X(n21585) );
  nand_x4_sg U60153 ( .A(n13062), .B(n13063), .X(n13055) );
  nand_x4_sg U60154 ( .A(n15395), .B(n15396), .X(n15388) );
  nand_x4_sg U60155 ( .A(n16961), .B(n16962), .X(n16954) );
  nand_x4_sg U60156 ( .A(n18502), .B(n18503), .X(n18495) );
  nand_x4_sg U60157 ( .A(n10720), .B(n10721), .X(n10713) );
  nand_x4_sg U60158 ( .A(n14612), .B(n14613), .X(n14605) );
  nand_x4_sg U60159 ( .A(n12281), .B(n12282), .X(n12274) );
  nor_x1_sg U60160 ( .A(n51988), .B(n12360), .X(n12358) );
  nor_x1_sg U60161 ( .A(n44660), .B(n13921), .X(n13918) );
  nor_x1_sg U60162 ( .A(n54223), .B(n18578), .X(n18576) );
  nor_x1_sg U60163 ( .A(n9355), .B(n9016), .X(\L2_0/n4072 ) );
  nor_x1_sg U60164 ( .A(n9355), .B(n9014), .X(\L2_0/n4068 ) );
  nand_x1_sg U60165 ( .A(n44094), .B(n46487), .X(n8792) );
  nand_x1_sg U60166 ( .A(n41980), .B(n46419), .X(n9319) );
  nand_x1_sg U60167 ( .A(n42873), .B(n46419), .X(n9344) );
  nand_x1_sg U60168 ( .A(n44116), .B(n46419), .X(n9327) );
  nand_x1_sg U60169 ( .A(n46419), .B(n44114), .X(n9317) );
  nand_x1_sg U60170 ( .A(n41976), .B(n46398), .X(n9308) );
  nand_x1_sg U60171 ( .A(n42869), .B(n46398), .X(n9304) );
  nand_x1_sg U60172 ( .A(n44112), .B(n46398), .X(n9295) );
  nand_x1_sg U60173 ( .A(n44110), .B(n46398), .X(n9281) );
  nand_x1_sg U60174 ( .A(n41988), .B(n46465), .X(n8957) );
  nand_x1_sg U60175 ( .A(n42879), .B(n46465), .X(n8999) );
  nand_x1_sg U60176 ( .A(n44399), .B(n46465), .X(n8941) );
  nand_x1_sg U60177 ( .A(n41972), .B(n46327), .X(n9232) );
  nand_x1_sg U60178 ( .A(n42863), .B(n46327), .X(n9228) );
  nand_x1_sg U60179 ( .A(n44393), .B(n46327), .X(n9205) );
  nand_x1_sg U60180 ( .A(n41998), .B(n46531), .X(n8924) );
  nand_x1_sg U60181 ( .A(n42887), .B(n46531), .X(n8920) );
  nand_x1_sg U60182 ( .A(n44132), .B(n46531), .X(n8934) );
  nand_x1_sg U60183 ( .A(n44130), .B(n46531), .X(n8926) );
  nor_x1_sg U60184 ( .A(n11233), .B(n11234), .X(n11232) );
  nand_x2_sg U60185 ( .A(n11233), .B(n11234), .X(n11235) );
  nor_x1_sg U60186 ( .A(n12794), .B(n12795), .X(n12793) );
  nand_x2_sg U60187 ( .A(n12794), .B(n12795), .X(n12796) );
  nor_x1_sg U60188 ( .A(n15127), .B(n15128), .X(n15126) );
  nand_x2_sg U60189 ( .A(n15127), .B(n15128), .X(n15129) );
  nor_x1_sg U60190 ( .A(n16693), .B(n16694), .X(n16692) );
  nand_x2_sg U60191 ( .A(n16693), .B(n16694), .X(n16695) );
  nor_x1_sg U60192 ( .A(n11631), .B(n41251), .X(n11630) );
  nor_x1_sg U60193 ( .A(n16307), .B(n41237), .X(n16306) );
  nor_x1_sg U60194 ( .A(n18631), .B(n41249), .X(n18630) );
  nor_x1_sg U60195 ( .A(n20177), .B(n41247), .X(n20176) );
  nor_x1_sg U60196 ( .A(n21722), .B(n41245), .X(n21721) );
  nor_x1_sg U60197 ( .A(n41699), .B(n12425), .X(n12423) );
  nor_x1_sg U60198 ( .A(n41695), .B(n13206), .X(n13204) );
  nor_x1_sg U60199 ( .A(n41691), .B(n13986), .X(n13984) );
  nor_x1_sg U60200 ( .A(n41687), .B(n15539), .X(n15537) );
  nor_x1_sg U60201 ( .A(n41683), .B(n17105), .X(n17103) );
  nor_x1_sg U60202 ( .A(n53898), .B(n53916), .X(n17798) );
  nor_x1_sg U60203 ( .A(n54463), .B(n54481), .X(n19343) );
  nor_x1_sg U60204 ( .A(n55031), .B(n55049), .X(n20887) );
  nor_x1_sg U60205 ( .A(n51547), .B(n11066), .X(n11068) );
  nor_x1_sg U60206 ( .A(n52104), .B(n12627), .X(n12629) );
  nor_x1_sg U60207 ( .A(n52938), .B(n14960), .X(n14962) );
  nor_x1_sg U60208 ( .A(n53496), .B(n16526), .X(n16528) );
  nand_x1_sg U60209 ( .A(n42449), .B(n13617), .X(n13615) );
  nand_x1_sg U60210 ( .A(n17514), .B(n17515), .X(n17513) );
  nand_x1_sg U60211 ( .A(n19059), .B(n19060), .X(n19058) );
  nand_x1_sg U60212 ( .A(n20603), .B(n20604), .X(n20602) );
  nand_x1_sg U60213 ( .A(n41770), .B(n41534), .X(n11640) );
  nand_x1_sg U60214 ( .A(n41786), .B(n41542), .X(n14752) );
  nand_x1_sg U60215 ( .A(n41738), .B(n41524), .X(n16315) );
  nand_x1_sg U60216 ( .A(n41784), .B(n41540), .X(n17873) );
  nand_x1_sg U60217 ( .A(n41782), .B(n41538), .X(n19418) );
  nand_x1_sg U60218 ( .A(n41780), .B(n41536), .X(n20962) );
  nand_x1_sg U60219 ( .A(n41766), .B(n41532), .X(n18640) );
  nor_x1_sg U60220 ( .A(n41187), .B(n42699), .X(n17517) );
  nor_x1_sg U60221 ( .A(n41185), .B(n42697), .X(n19062) );
  nor_x1_sg U60222 ( .A(n41183), .B(n42693), .X(n20606) );
  nor_x1_sg U60223 ( .A(n13686), .B(n13641), .X(n13682) );
  nand_x1_sg U60224 ( .A(n18181), .B(n18182), .X(n18180) );
  nand_x1_sg U60225 ( .A(n11328), .B(n11327), .X(n11329) );
  nand_x1_sg U60226 ( .A(n12108), .B(n12107), .X(n12109) );
  nand_x1_sg U60227 ( .A(n12889), .B(n12888), .X(n12890) );
  nand_x1_sg U60228 ( .A(n13669), .B(n13668), .X(n13670) );
  nand_x1_sg U60229 ( .A(n15222), .B(n15221), .X(n15223) );
  nand_x1_sg U60230 ( .A(n16003), .B(n16002), .X(n16004) );
  nand_x1_sg U60231 ( .A(n16788), .B(n16787), .X(n16789) );
  nand_x1_sg U60232 ( .A(n10555), .B(n10556), .X(n10554) );
  nand_x1_sg U60233 ( .A(n17567), .B(n17568), .X(n17566) );
  nand_x1_sg U60234 ( .A(n19112), .B(n19113), .X(n19111) );
  nand_x1_sg U60235 ( .A(n20656), .B(n20657), .X(n20655) );
  nand_x1_sg U60236 ( .A(n13723), .B(n13722), .X(n13724) );
  nand_x1_sg U60237 ( .A(n51460), .B(n11002), .X(n11011) );
  nor_x1_sg U60238 ( .A(n41496), .B(n12443), .X(n12441) );
  nor_x1_sg U60239 ( .A(n41219), .B(n14004), .X(n14002) );
  nand_x1_sg U60240 ( .A(n11667), .B(n43005), .X(n11666) );
  nand_x1_sg U60241 ( .A(n12447), .B(n43001), .X(n12446) );
  nand_x1_sg U60242 ( .A(n13228), .B(n42997), .X(n13227) );
  nand_x1_sg U60243 ( .A(n14008), .B(n42993), .X(n14007) );
  nand_x1_sg U60244 ( .A(n14779), .B(n42989), .X(n14778) );
  nand_x1_sg U60245 ( .A(n15561), .B(n42985), .X(n15560) );
  nand_x1_sg U60246 ( .A(n17127), .B(n42977), .X(n17126) );
  nand_x1_sg U60247 ( .A(n17900), .B(n42973), .X(n17899) );
  nand_x1_sg U60248 ( .A(n18669), .B(n42969), .X(n18668) );
  nand_x1_sg U60249 ( .A(n19445), .B(n42965), .X(n19444) );
  nand_x1_sg U60250 ( .A(n20214), .B(n42961), .X(n20213) );
  nand_x1_sg U60251 ( .A(n20989), .B(n42957), .X(n20988) );
  nand_x1_sg U60252 ( .A(n21759), .B(n42953), .X(n21758) );
  nor_x1_sg U60253 ( .A(n41418), .B(n14823), .X(n14821) );
  nand_x1_sg U60254 ( .A(n14823), .B(n41418), .X(n14822) );
  nor_x1_sg U60255 ( .A(n41412), .B(n17944), .X(n17942) );
  nand_x1_sg U60256 ( .A(n17944), .B(n41412), .X(n17943) );
  nor_x1_sg U60257 ( .A(n41410), .B(n18713), .X(n18711) );
  nand_x1_sg U60258 ( .A(n18713), .B(n41410), .X(n18712) );
  nor_x1_sg U60259 ( .A(n41408), .B(n19489), .X(n19487) );
  nand_x1_sg U60260 ( .A(n19489), .B(n41408), .X(n19488) );
  nor_x1_sg U60261 ( .A(n41406), .B(n20259), .X(n20257) );
  nand_x1_sg U60262 ( .A(n20259), .B(n41406), .X(n20258) );
  nor_x1_sg U60263 ( .A(n41404), .B(n21033), .X(n21031) );
  nand_x1_sg U60264 ( .A(n21033), .B(n41404), .X(n21032) );
  nor_x1_sg U60265 ( .A(n41402), .B(n21804), .X(n21802) );
  nand_x1_sg U60266 ( .A(n21804), .B(n41402), .X(n21803) );
  nor_x1_sg U60267 ( .A(n54638), .B(n54630), .X(n19731) );
  nor_x1_sg U60268 ( .A(n55206), .B(n55198), .X(n21276) );
  nor_x1_sg U60269 ( .A(n51284), .B(n51276), .X(n10404) );
  nor_x1_sg U60270 ( .A(n53993), .B(n17896), .X(n17895) );
  nor_x1_sg U60271 ( .A(n54276), .B(n18665), .X(n18664) );
  nor_x1_sg U60272 ( .A(n54558), .B(n19441), .X(n19440) );
  nor_x1_sg U60273 ( .A(n54843), .B(n20210), .X(n20209) );
  nor_x1_sg U60274 ( .A(n55126), .B(n20985), .X(n20984) );
  nor_x1_sg U60275 ( .A(n55411), .B(n21755), .X(n21754) );
  nor_x1_sg U60276 ( .A(n11002), .B(n44503), .X(n11001) );
  nand_x1_sg U60277 ( .A(n10618), .B(n10619), .X(n10617) );
  nand_x1_sg U60278 ( .A(n18400), .B(n18401), .X(n18399) );
  nand_x1_sg U60279 ( .A(n19945), .B(n19946), .X(n19944) );
  nand_x1_sg U60280 ( .A(n21490), .B(n21491), .X(n21489) );
  nand_x1_sg U60281 ( .A(n14510), .B(n14511), .X(n14509) );
  nand_x1_sg U60282 ( .A(n17631), .B(n17632), .X(n17630) );
  nand_x1_sg U60283 ( .A(n19176), .B(n19177), .X(n19175) );
  nand_x1_sg U60284 ( .A(n20720), .B(n20721), .X(n20719) );
  nor_x1_sg U60285 ( .A(n17312), .B(n42441), .X(n17400) );
  nor_x1_sg U60286 ( .A(n18857), .B(n42439), .X(n18945) );
  nor_x1_sg U60287 ( .A(n20401), .B(n42437), .X(n20489) );
  nor_x1_sg U60288 ( .A(n10743), .B(n10742), .X(n10740) );
  nand_x1_sg U60289 ( .A(n10742), .B(n10743), .X(n10741) );
  nor_x1_sg U60290 ( .A(n20138), .B(n20139), .X(n20137) );
  nand_x1_sg U60291 ( .A(n20139), .B(n20138), .X(n20140) );
  nor_x1_sg U60292 ( .A(n21683), .B(n21684), .X(n21682) );
  nand_x1_sg U60293 ( .A(n21684), .B(n21683), .X(n21685) );
  nand_x1_sg U60294 ( .A(n20202), .B(n20201), .X(n20203) );
  nand_x1_sg U60295 ( .A(n21747), .B(n21746), .X(n21748) );
  nor_x1_sg U60296 ( .A(n13203), .B(n43109), .X(n13339) );
  nor_x1_sg U60297 ( .A(n13983), .B(n43107), .X(n14119) );
  nor_x1_sg U60298 ( .A(n15536), .B(n43105), .X(n15672) );
  nor_x1_sg U60299 ( .A(n17102), .B(n43103), .X(n17238) );
  nor_x1_sg U60300 ( .A(n42811), .B(n41502), .X(n13681) );
  nand_x1_sg U60301 ( .A(n13876), .B(n13875), .X(n13877) );
  nor_x1_sg U60302 ( .A(n18770), .B(n54064), .X(n18769) );
  nand_x1_sg U60303 ( .A(n15892), .B(n53256), .X(n15893) );
  nand_x1_sg U60304 ( .A(n13558), .B(n52421), .X(n13559) );
  nand_x1_sg U60305 ( .A(n11997), .B(n51869), .X(n11998) );
  nor_x1_sg U60306 ( .A(n18653), .B(n46340), .X(n18727) );
  nor_x1_sg U60307 ( .A(n17707), .B(n46367), .X(n17706) );
  nor_x1_sg U60308 ( .A(n19252), .B(n46320), .X(n19251) );
  nor_x1_sg U60309 ( .A(n20796), .B(n46275), .X(n20795) );
  nor_x1_sg U60310 ( .A(n11475), .B(n46546), .X(n11474) );
  nor_x1_sg U60311 ( .A(n13036), .B(n46502), .X(n13035) );
  nor_x1_sg U60312 ( .A(n15369), .B(n46434), .X(n15368) );
  nor_x1_sg U60313 ( .A(n16935), .B(n46390), .X(n16934) );
  nor_x1_sg U60314 ( .A(n52836), .B(n14883), .X(n14882) );
  nor_x1_sg U60315 ( .A(n53956), .B(n18004), .X(n18003) );
  nor_x1_sg U60316 ( .A(n54521), .B(n19549), .X(n19548) );
  nor_x1_sg U60317 ( .A(n54806), .B(n20319), .X(n20318) );
  nor_x1_sg U60318 ( .A(n55089), .B(n21093), .X(n21092) );
  nor_x1_sg U60319 ( .A(n55374), .B(n21864), .X(n21863) );
  nand_x4_sg U60320 ( .A(n42272), .B(n13321), .X(n13280) );
  nand_x4_sg U60321 ( .A(n42264), .B(n15654), .X(n15613) );
  nand_x4_sg U60322 ( .A(n42260), .B(n17220), .X(n17179) );
  nand_x4_sg U60323 ( .A(n46356), .B(n46363), .X(n17651) );
  nand_x4_sg U60324 ( .A(n46309), .B(n46316), .X(n19196) );
  nand_x4_sg U60325 ( .A(n46264), .B(n46271), .X(n20740) );
  nand_x4_sg U60326 ( .A(n54149), .B(n18388), .X(n18346) );
  nand_x1_sg U60327 ( .A(n54148), .B(n18389), .X(n18388) );
  nand_x4_sg U60328 ( .A(n52757), .B(n14498), .X(n14456) );
  nand_x1_sg U60329 ( .A(n52756), .B(n14499), .X(n14498) );
  nand_x4_sg U60330 ( .A(n54714), .B(n19933), .X(n19891) );
  nand_x1_sg U60331 ( .A(n54713), .B(n19934), .X(n19933) );
  nand_x4_sg U60332 ( .A(n55282), .B(n21478), .X(n21436) );
  nand_x1_sg U60333 ( .A(n55281), .B(n21479), .X(n21478) );
  nand_x4_sg U60334 ( .A(n44201), .B(n13529), .X(n13499) );
  nand_x1_sg U60335 ( .A(n43936), .B(n13526), .X(n13529) );
  nand_x4_sg U60336 ( .A(n41251), .B(n11631), .X(n11605) );
  nand_x4_sg U60337 ( .A(n41237), .B(n16307), .X(n16281) );
  nand_x4_sg U60338 ( .A(n41249), .B(n18631), .X(n18605) );
  nand_x4_sg U60339 ( .A(n41247), .B(n20177), .X(n20151) );
  nand_x4_sg U60340 ( .A(n41245), .B(n21722), .X(n21696) );
  nand_x4_sg U60341 ( .A(n12413), .B(n12412), .X(n12386) );
  nand_x4_sg U60342 ( .A(n53794), .B(n17310), .X(n9254) );
  nand_x1_sg U60343 ( .A(n42441), .B(n17312), .X(n17310) );
  nand_x4_sg U60344 ( .A(n54359), .B(n18855), .X(n9216) );
  nand_x1_sg U60345 ( .A(n42439), .B(n18857), .X(n18855) );
  nand_x1_sg U60346 ( .A(n42437), .B(n20401), .X(n20399) );
  nand_x4_sg U60347 ( .A(n41346), .B(n41175), .X(n11851) );
  nand_x4_sg U60348 ( .A(n41342), .B(n41173), .X(n15746) );
  nand_x4_sg U60349 ( .A(n41177), .B(n54629), .X(n19628) );
  nand_x4_sg U60350 ( .A(n18171), .B(n54061), .X(n18083) );
  nand_x4_sg U60351 ( .A(n42192), .B(n11338), .X(n11337) );
  nand_x1_sg U60352 ( .A(n51610), .B(n11339), .X(n11338) );
  nand_x4_sg U60353 ( .A(n42190), .B(n12118), .X(n12117) );
  nand_x1_sg U60354 ( .A(n51891), .B(n12119), .X(n12118) );
  nand_x4_sg U60355 ( .A(n41709), .B(n12899), .X(n12898) );
  nand_x1_sg U60356 ( .A(n52168), .B(n12900), .X(n12899) );
  nand_x4_sg U60357 ( .A(n41707), .B(n13679), .X(n13678) );
  nand_x1_sg U60358 ( .A(n52442), .B(n13680), .X(n13679) );
  nand_x4_sg U60359 ( .A(n41705), .B(n15232), .X(n15231) );
  nand_x1_sg U60360 ( .A(n53002), .B(n15233), .X(n15232) );
  nand_x4_sg U60361 ( .A(n42188), .B(n16013), .X(n16012) );
  nand_x1_sg U60362 ( .A(n53278), .B(n16014), .X(n16013) );
  nand_x4_sg U60363 ( .A(n41703), .B(n16798), .X(n16797) );
  nand_x1_sg U60364 ( .A(n53560), .B(n16799), .X(n16798) );
  nand_x4_sg U60365 ( .A(n41707), .B(n13650), .X(n13643) );
  nand_x1_sg U60366 ( .A(n41502), .B(n42811), .X(n13650) );
  nand_x2_sg U60367 ( .A(n53327), .B(n16070), .X(n16051) );
  nand_x1_sg U60368 ( .A(n16071), .B(n16072), .X(n16070) );
  nand_x2_sg U60369 ( .A(n51658), .B(n11395), .X(n11376) );
  nand_x1_sg U60370 ( .A(n11396), .B(n11397), .X(n11395) );
  nand_x2_sg U60371 ( .A(n52214), .B(n12956), .X(n12937) );
  nand_x1_sg U60372 ( .A(n12957), .B(n12958), .X(n12956) );
  nand_x2_sg U60373 ( .A(n53048), .B(n15289), .X(n15270) );
  nand_x1_sg U60374 ( .A(n15290), .B(n15291), .X(n15289) );
  nand_x2_sg U60375 ( .A(n53606), .B(n16855), .X(n16836) );
  nand_x1_sg U60376 ( .A(n16856), .B(n16857), .X(n16855) );
  nand_x2_sg U60377 ( .A(n51939), .B(n12175), .X(n12156) );
  nand_x1_sg U60378 ( .A(n12176), .B(n12177), .X(n12175) );
  nand_x2_sg U60379 ( .A(n52491), .B(n13736), .X(n13717) );
  nand_x1_sg U60380 ( .A(n13737), .B(n13738), .X(n13736) );
  nand_x4_sg U60381 ( .A(n11624), .B(n11625), .X(n11535) );
  nand_x4_sg U60382 ( .A(n13185), .B(n13186), .X(n13096) );
  nand_x4_sg U60383 ( .A(n15518), .B(n15519), .X(n15429) );
  nand_x4_sg U60384 ( .A(n16300), .B(n16301), .X(n16211) );
  nand_x4_sg U60385 ( .A(n17084), .B(n17085), .X(n16995) );
  nand_x4_sg U60386 ( .A(n12405), .B(n12406), .X(n12316) );
  nand_x4_sg U60387 ( .A(n12219), .B(n12220), .X(n12162) );
  nand_x4_sg U60388 ( .A(n46285), .B(n46296), .X(n20029) );
  nand_x4_sg U60389 ( .A(n46240), .B(n46251), .X(n21574) );
  nand_x4_sg U60390 ( .A(n14736), .B(n14737), .X(n14646) );
  nand_x4_sg U60391 ( .A(n17857), .B(n17858), .X(n17767) );
  nand_x4_sg U60392 ( .A(n19402), .B(n19403), .X(n19312) );
  nand_x4_sg U60393 ( .A(n20946), .B(n20947), .X(n20856) );
  nand_x4_sg U60394 ( .A(n45537), .B(n13201), .X(n13194) );
  nand_x1_sg U60395 ( .A(n43109), .B(n13203), .X(n13201) );
  nand_x4_sg U60396 ( .A(n45535), .B(n13981), .X(n13974) );
  nand_x1_sg U60397 ( .A(n43107), .B(n13983), .X(n13981) );
  nand_x4_sg U60398 ( .A(n45533), .B(n15534), .X(n15527) );
  nand_x1_sg U60399 ( .A(n43105), .B(n15536), .X(n15534) );
  nand_x4_sg U60400 ( .A(n45531), .B(n17100), .X(n17093) );
  nand_x1_sg U60401 ( .A(n43103), .B(n17102), .X(n17100) );
  nand_x4_sg U60402 ( .A(n10958), .B(n51443), .X(n10876) );
  nand_x1_sg U60403 ( .A(n51372), .B(n10955), .X(n10958) );
  nor_x1_sg U60404 ( .A(n10955), .B(n51372), .X(n10959) );
  nand_x4_sg U60405 ( .A(n18233), .B(n18225), .X(n18231) );
  nand_x4_sg U60406 ( .A(n46557), .B(n46567), .X(n10702) );
  nand_x4_sg U60407 ( .A(n20170), .B(n20171), .X(n20080) );
  nand_x4_sg U60408 ( .A(n21715), .B(n21716), .X(n21625) );
  nand_x4_sg U60409 ( .A(n19985), .B(n19986), .X(n19931) );
  nand_x4_sg U60410 ( .A(n21530), .B(n21531), .X(n21476) );
  nor_x1_sg U60411 ( .A(n20287), .B(n54726), .X(n20291) );
  nor_x1_sg U60412 ( .A(n21832), .B(n55294), .X(n21836) );
  nand_x4_sg U60413 ( .A(n20349), .B(n54815), .X(n20144) );
  nand_x1_sg U60414 ( .A(n20316), .B(n20351), .X(n20349) );
  nor_x1_sg U60415 ( .A(n20351), .B(n20316), .X(n20350) );
  nand_x4_sg U60416 ( .A(n21894), .B(n55383), .X(n21689) );
  nand_x1_sg U60417 ( .A(n21861), .B(n21896), .X(n21894) );
  nor_x1_sg U60418 ( .A(n21896), .B(n21861), .X(n21895) );
  nor_x1_sg U60419 ( .A(n12011), .B(n12012), .X(n12010) );
  nor_x1_sg U60420 ( .A(n13572), .B(n13573), .X(n13571) );
  nor_x1_sg U60421 ( .A(n15906), .B(n15907), .X(n15905) );
  nand_x4_sg U60422 ( .A(n14913), .B(n52845), .X(n14710) );
  nor_x1_sg U60423 ( .A(n14915), .B(n14880), .X(n14914) );
  nand_x4_sg U60424 ( .A(n18034), .B(n53965), .X(n17831) );
  nor_x1_sg U60425 ( .A(n18036), .B(n18001), .X(n18035) );
  nand_x4_sg U60426 ( .A(n19579), .B(n54530), .X(n19376) );
  nor_x1_sg U60427 ( .A(n19581), .B(n19546), .X(n19580) );
  nand_x4_sg U60428 ( .A(n21123), .B(n55098), .X(n20920) );
  nor_x1_sg U60429 ( .A(n21125), .B(n21090), .X(n21124) );
  nand_x4_sg U60430 ( .A(n54197), .B(n18609), .X(n18538) );
  nand_x1_sg U60431 ( .A(n18610), .B(n54196), .X(n18609) );
  nor_x1_sg U60432 ( .A(n18610), .B(n54196), .X(n18611) );
  nand_x4_sg U60433 ( .A(n54764), .B(n20155), .X(n20083) );
  nand_x1_sg U60434 ( .A(n20156), .B(n54763), .X(n20155) );
  nor_x1_sg U60435 ( .A(n20156), .B(n54763), .X(n20157) );
  nand_x4_sg U60436 ( .A(n55332), .B(n21700), .X(n21628) );
  nand_x1_sg U60437 ( .A(n21701), .B(n55331), .X(n21700) );
  nor_x1_sg U60438 ( .A(n21701), .B(n55331), .X(n21702) );
  nand_x4_sg U60439 ( .A(n10658), .B(n10659), .X(n10604) );
  nand_x4_sg U60440 ( .A(n16114), .B(n16115), .X(n16057) );
  nor_x1_sg U60441 ( .A(n46585), .B(n26234), .X(\L1_0/n4499 ) );
  nor_x1_sg U60442 ( .A(n55661), .B(n46585), .X(\L1_0/n4498 ) );
  nor_x1_sg U60443 ( .A(n46585), .B(n26241), .X(\L1_0/n4495 ) );
  nor_x1_sg U60444 ( .A(n55662), .B(n46585), .X(\L1_0/n4494 ) );
  nor_x1_sg U60445 ( .A(n46585), .B(n26248), .X(\L1_0/n4491 ) );
  nor_x1_sg U60446 ( .A(n55663), .B(n46585), .X(\L1_0/n4490 ) );
  nor_x1_sg U60447 ( .A(n46585), .B(n26255), .X(\L1_0/n4487 ) );
  nor_x1_sg U60448 ( .A(n55664), .B(n46585), .X(\L1_0/n4486 ) );
  nor_x1_sg U60449 ( .A(n55670), .B(n46587), .X(\L1_0/n4422 ) );
  nor_x1_sg U60450 ( .A(n46587), .B(n26513), .X(\L1_0/n4419 ) );
  nor_x1_sg U60451 ( .A(n55671), .B(n46587), .X(\L1_0/n4418 ) );
  nor_x1_sg U60452 ( .A(n46587), .B(n26520), .X(\L1_0/n4415 ) );
  nor_x1_sg U60453 ( .A(n55672), .B(n46587), .X(\L1_0/n4414 ) );
  nor_x1_sg U60454 ( .A(n46587), .B(n26527), .X(\L1_0/n4411 ) );
  nor_x1_sg U60455 ( .A(n55673), .B(n46587), .X(\L1_0/n4410 ) );
  nor_x1_sg U60456 ( .A(n46587), .B(n26534), .X(\L1_0/n4407 ) );
  nor_x1_sg U60457 ( .A(n55674), .B(n46587), .X(\L1_0/n4406 ) );
  nor_x1_sg U60458 ( .A(n46591), .B(n27910), .X(\L1_0/n4019 ) );
  nor_x1_sg U60459 ( .A(n55721), .B(n46591), .X(\L1_0/n4018 ) );
  nor_x1_sg U60460 ( .A(n46591), .B(n27917), .X(\L1_0/n4015 ) );
  nor_x1_sg U60461 ( .A(n55722), .B(n46591), .X(\L1_0/n4014 ) );
  nor_x1_sg U60462 ( .A(n46591), .B(n27924), .X(\L1_0/n4011 ) );
  nor_x1_sg U60463 ( .A(n55723), .B(n46591), .X(\L1_0/n4010 ) );
  nor_x1_sg U60464 ( .A(n46591), .B(n27931), .X(\L1_0/n4007 ) );
  nor_x1_sg U60465 ( .A(n55724), .B(n46591), .X(\L1_0/n4006 ) );
  nor_x1_sg U60466 ( .A(n46591), .B(n55582), .X(\L1_0/n3999 ) );
  nor_x1_sg U60467 ( .A(n44048), .B(n46591), .X(\L1_0/n3998 ) );
  nor_x1_sg U60468 ( .A(n28459), .B(n28468), .X(\L1_0/n3859 ) );
  nor_x1_sg U60469 ( .A(n55741), .B(n28459), .X(\L1_0/n3858 ) );
  nor_x1_sg U60470 ( .A(n28459), .B(n28475), .X(\L1_0/n3855 ) );
  nor_x1_sg U60471 ( .A(n55742), .B(n28459), .X(\L1_0/n3854 ) );
  nor_x1_sg U60472 ( .A(n28459), .B(n28482), .X(\L1_0/n3851 ) );
  nor_x1_sg U60473 ( .A(n55743), .B(n28459), .X(\L1_0/n3850 ) );
  nor_x1_sg U60474 ( .A(n28459), .B(n28489), .X(\L1_0/n3847 ) );
  nor_x1_sg U60475 ( .A(n55744), .B(n28459), .X(\L1_0/n3846 ) );
  nor_x1_sg U60476 ( .A(n46596), .B(n29308), .X(\L1_0/n3619 ) );
  nor_x1_sg U60477 ( .A(n55771), .B(n46596), .X(\L1_0/n3618 ) );
  nor_x1_sg U60478 ( .A(n46596), .B(n29315), .X(\L1_0/n3615 ) );
  nor_x1_sg U60479 ( .A(n55772), .B(n46596), .X(\L1_0/n3614 ) );
  nor_x1_sg U60480 ( .A(n46596), .B(n29322), .X(\L1_0/n3611 ) );
  nor_x1_sg U60481 ( .A(n55773), .B(n46596), .X(\L1_0/n3610 ) );
  nor_x1_sg U60482 ( .A(n46596), .B(n29329), .X(\L1_0/n3607 ) );
  nor_x1_sg U60483 ( .A(n55774), .B(n46596), .X(\L1_0/n3606 ) );
  nor_x1_sg U60484 ( .A(n17643), .B(n17644), .X(n17642) );
  nor_x1_sg U60485 ( .A(n19188), .B(n19189), .X(n19187) );
  nor_x1_sg U60486 ( .A(n20732), .B(n20733), .X(n20731) );
  nor_x1_sg U60487 ( .A(n14522), .B(n14523), .X(n14521) );
  nor_x1_sg U60488 ( .A(n12189), .B(n12190), .X(n12188) );
  nor_x1_sg U60489 ( .A(n16084), .B(n16085), .X(n16083) );
  nand_x4_sg U60490 ( .A(n11407), .B(n51689), .X(n11400) );
  nor_x1_sg U60491 ( .A(n11409), .B(n11410), .X(n11408) );
  nand_x4_sg U60492 ( .A(n12968), .B(n52244), .X(n12961) );
  nor_x1_sg U60493 ( .A(n12970), .B(n12971), .X(n12969) );
  nor_x1_sg U60494 ( .A(n13750), .B(n13751), .X(n13749) );
  nand_x4_sg U60495 ( .A(n15301), .B(n53078), .X(n15294) );
  nor_x1_sg U60496 ( .A(n15303), .B(n15304), .X(n15302) );
  nand_x4_sg U60497 ( .A(n16867), .B(n53636), .X(n16860) );
  nor_x1_sg U60498 ( .A(n16869), .B(n16870), .X(n16868) );
  nand_x4_sg U60499 ( .A(n12370), .B(n12371), .X(n12312) );
  nand_x1_sg U60500 ( .A(n51922), .B(n12362), .X(n12371) );
  nand_x1_sg U60501 ( .A(n51898), .B(n12361), .X(n12370) );
  nand_x4_sg U60502 ( .A(n14465), .B(n14466), .X(n14413) );
  nor_x1_sg U60503 ( .A(n46585), .B(n55535), .X(\L1_0/n4479 ) );
  nor_x1_sg U60504 ( .A(n44058), .B(n46585), .X(\L1_0/n4478 ) );
  nor_x1_sg U60505 ( .A(n46585), .B(n55536), .X(\L1_0/n4475 ) );
  nor_x1_sg U60506 ( .A(n44495), .B(n46585), .X(\L1_0/n4474 ) );
  nor_x1_sg U60507 ( .A(n46587), .B(n55544), .X(\L1_0/n4395 ) );
  nor_x1_sg U60508 ( .A(n44493), .B(n46587), .X(\L1_0/n4394 ) );
  nor_x1_sg U60509 ( .A(n46589), .B(n27070), .X(\L1_0/n4259 ) );
  nor_x1_sg U60510 ( .A(n55691), .B(n46589), .X(\L1_0/n4258 ) );
  nor_x1_sg U60511 ( .A(n46589), .B(n27077), .X(\L1_0/n4255 ) );
  nor_x1_sg U60512 ( .A(n55692), .B(n46589), .X(\L1_0/n4254 ) );
  nor_x1_sg U60513 ( .A(n46589), .B(n27084), .X(\L1_0/n4251 ) );
  nor_x1_sg U60514 ( .A(n55693), .B(n46589), .X(\L1_0/n4250 ) );
  nor_x1_sg U60515 ( .A(n46589), .B(n27091), .X(\L1_0/n4247 ) );
  nor_x1_sg U60516 ( .A(n55694), .B(n46589), .X(\L1_0/n4246 ) );
  nor_x1_sg U60517 ( .A(n28459), .B(n55598), .X(\L1_0/n3839 ) );
  nor_x1_sg U60518 ( .A(n44046), .B(n28459), .X(\L1_0/n3838 ) );
  nor_x1_sg U60519 ( .A(n46596), .B(n55623), .X(\L1_0/n3595 ) );
  nor_x1_sg U60520 ( .A(n44217), .B(n46596), .X(\L1_0/n3594 ) );
  nor_x1_sg U60521 ( .A(n46596), .B(n55624), .X(\L1_0/n3587 ) );
  nor_x1_sg U60522 ( .A(n44040), .B(n46596), .X(\L1_0/n3586 ) );
  nand_x4_sg U60523 ( .A(n19900), .B(n19901), .X(n19848) );
  nand_x4_sg U60524 ( .A(n21445), .B(n21446), .X(n21393) );
  nor_x1_sg U60525 ( .A(n9355), .B(n9034), .X(\L2_0/n4124 ) );
  nor_x1_sg U60526 ( .A(n9355), .B(n9030), .X(\L2_0/n4116 ) );
  nor_x1_sg U60527 ( .A(n9355), .B(n9047), .X(\L2_0/n4112 ) );
  nor_x1_sg U60528 ( .A(n46589), .B(n55559), .X(\L1_0/n4239 ) );
  nor_x1_sg U60529 ( .A(n44052), .B(n46589), .X(\L1_0/n4238 ) );
  nor_x1_sg U60530 ( .A(n46589), .B(n55560), .X(\L1_0/n4235 ) );
  nor_x1_sg U60531 ( .A(n44491), .B(n46589), .X(\L1_0/n4234 ) );
  nor_x1_sg U60532 ( .A(n55763), .B(n46616), .X(\L1_0/n3690 ) );
  nor_x1_sg U60533 ( .A(n46616), .B(n29048), .X(\L1_0/n3687 ) );
  nor_x1_sg U60534 ( .A(n55764), .B(n46616), .X(\L1_0/n3686 ) );
  nor_x1_sg U60535 ( .A(n46616), .B(n55614), .X(\L1_0/n3679 ) );
  nor_x1_sg U60536 ( .A(n44042), .B(n46616), .X(\L1_0/n3678 ) );
  nor_x1_sg U60537 ( .A(n46615), .B(n25396), .X(\L1_0/n4739 ) );
  nor_x1_sg U60538 ( .A(n46615), .B(n55631), .X(\L1_0/n4738 ) );
  nor_x1_sg U60539 ( .A(n46615), .B(n25403), .X(\L1_0/n4735 ) );
  nor_x1_sg U60540 ( .A(n46615), .B(n55632), .X(\L1_0/n4734 ) );
  nor_x1_sg U60541 ( .A(n46615), .B(n25410), .X(\L1_0/n4731 ) );
  nor_x1_sg U60542 ( .A(n46615), .B(n55633), .X(\L1_0/n4730 ) );
  nor_x1_sg U60543 ( .A(n46615), .B(n25417), .X(\L1_0/n4727 ) );
  nor_x1_sg U60544 ( .A(n46615), .B(n55634), .X(\L1_0/n4726 ) );
  nor_x1_sg U60545 ( .A(n46615), .B(n55514), .X(\L1_0/n4715 ) );
  nor_x1_sg U60546 ( .A(n46615), .B(n44243), .X(\L1_0/n4714 ) );
  nor_x1_sg U60547 ( .A(n46615), .B(n55515), .X(\L1_0/n4707 ) );
  nor_x1_sg U60548 ( .A(n46615), .B(n44064), .X(\L1_0/n4706 ) );
  nor_x1_sg U60549 ( .A(n46615), .B(n55516), .X(\L1_0/n4699 ) );
  nor_x1_sg U60550 ( .A(n46615), .B(n43934), .X(\L1_0/n4698 ) );
  nor_x1_sg U60551 ( .A(n55653), .B(n46612), .X(\L1_0/n4570 ) );
  nor_x1_sg U60552 ( .A(n46612), .B(n25974), .X(\L1_0/n4567 ) );
  nor_x1_sg U60553 ( .A(n55654), .B(n46612), .X(\L1_0/n4566 ) );
  nor_x1_sg U60554 ( .A(n46612), .B(n55529), .X(\L1_0/n4555 ) );
  nor_x1_sg U60555 ( .A(n44241), .B(n46612), .X(\L1_0/n4554 ) );
  nor_x1_sg U60556 ( .A(n46625), .B(n26812), .X(\L1_0/n4327 ) );
  nor_x1_sg U60557 ( .A(n46625), .B(n55684), .X(\L1_0/n4326 ) );
  nor_x1_sg U60558 ( .A(n46611), .B(n25696), .X(\L1_0/n4647 ) );
  nor_x1_sg U60559 ( .A(n46611), .B(n55644), .X(\L1_0/n4646 ) );
  nor_x1_sg U60560 ( .A(n46611), .B(n55521), .X(\L1_0/n4639 ) );
  nor_x1_sg U60561 ( .A(n46611), .B(n44062), .X(\L1_0/n4638 ) );
  nor_x1_sg U60562 ( .A(n46611), .B(n55522), .X(\L1_0/n4635 ) );
  nor_x1_sg U60563 ( .A(n46611), .B(n44499), .X(\L1_0/n4634 ) );
  nor_x1_sg U60564 ( .A(n46623), .B(n27371), .X(\L1_0/n4167 ) );
  nor_x1_sg U60565 ( .A(n46623), .B(n55704), .X(\L1_0/n4166 ) );
  nor_x1_sg U60566 ( .A(n46623), .B(n55568), .X(\L1_0/n4155 ) );
  nor_x1_sg U60567 ( .A(n46623), .B(n45487), .X(\L1_0/n4154 ) );
  nor_x1_sg U60568 ( .A(n46621), .B(n27651), .X(\L1_0/n4087 ) );
  nor_x1_sg U60569 ( .A(n46621), .B(n55714), .X(\L1_0/n4086 ) );
  nor_x1_sg U60570 ( .A(n46621), .B(n55574), .X(\L1_0/n4079 ) );
  nor_x1_sg U60571 ( .A(n46621), .B(n44050), .X(\L1_0/n4078 ) );
  nor_x1_sg U60572 ( .A(n46621), .B(n55575), .X(\L1_0/n4075 ) );
  nor_x1_sg U60573 ( .A(n46621), .B(n44487), .X(\L1_0/n4074 ) );
  nor_x1_sg U60574 ( .A(n46619), .B(n28768), .X(\L1_0/n3767 ) );
  nor_x1_sg U60575 ( .A(n46619), .B(n55754), .X(\L1_0/n3766 ) );
  nor_x1_sg U60576 ( .A(n46619), .B(n55607), .X(\L1_0/n3755 ) );
  nor_x1_sg U60577 ( .A(n46619), .B(n44225), .X(\L1_0/n3754 ) );
  nor_x1_sg U60578 ( .A(n46619), .B(n55608), .X(\L1_0/n3747 ) );
  nor_x1_sg U60579 ( .A(n46619), .B(n44223), .X(\L1_0/n3746 ) );
  nand_x4_sg U60580 ( .A(n12309), .B(n51989), .X(n12307) );
  nand_x1_sg U60581 ( .A(n12312), .B(n12311), .X(n12309) );
  nor_x1_sg U60582 ( .A(n12311), .B(n12312), .X(n12310) );
  nor_x1_sg U60583 ( .A(n46585), .B(n26326), .X(\L1_0/n4447 ) );
  nor_x1_sg U60584 ( .A(n55669), .B(n46585), .X(\L1_0/n4446 ) );
  nor_x1_sg U60585 ( .A(n46587), .B(n26605), .X(\L1_0/n4367 ) );
  nor_x1_sg U60586 ( .A(n55679), .B(n46587), .X(\L1_0/n4366 ) );
  nor_x1_sg U60587 ( .A(n46612), .B(n26045), .X(\L1_0/n4527 ) );
  nor_x1_sg U60588 ( .A(n55659), .B(n46612), .X(\L1_0/n4526 ) );
  nor_x1_sg U60589 ( .A(n46621), .B(n27722), .X(\L1_0/n4047 ) );
  nor_x1_sg U60590 ( .A(n46621), .B(n55719), .X(\L1_0/n4046 ) );
  nor_x1_sg U60591 ( .A(n46616), .B(n29027), .X(\L1_0/n3699 ) );
  nor_x1_sg U60592 ( .A(n55761), .B(n46616), .X(\L1_0/n3698 ) );
  nor_x1_sg U60593 ( .A(n46616), .B(n29034), .X(\L1_0/n3695 ) );
  nor_x1_sg U60594 ( .A(n55762), .B(n46616), .X(\L1_0/n3694 ) );
  nor_x1_sg U60595 ( .A(n46616), .B(n29041), .X(\L1_0/n3691 ) );
  nor_x1_sg U60596 ( .A(n46612), .B(n25953), .X(\L1_0/n4579 ) );
  nor_x1_sg U60597 ( .A(n55651), .B(n46612), .X(\L1_0/n4578 ) );
  nor_x1_sg U60598 ( .A(n46612), .B(n25960), .X(\L1_0/n4575 ) );
  nor_x1_sg U60599 ( .A(n55652), .B(n46612), .X(\L1_0/n4574 ) );
  nor_x1_sg U60600 ( .A(n46612), .B(n25967), .X(\L1_0/n4571 ) );
  nor_x1_sg U60601 ( .A(n46611), .B(n25675), .X(\L1_0/n4659 ) );
  nor_x1_sg U60602 ( .A(n46611), .B(n55641), .X(\L1_0/n4658 ) );
  nor_x1_sg U60603 ( .A(n46611), .B(n25682), .X(\L1_0/n4655 ) );
  nor_x1_sg U60604 ( .A(n46611), .B(n55642), .X(\L1_0/n4654 ) );
  nor_x1_sg U60605 ( .A(n46611), .B(n25689), .X(\L1_0/n4651 ) );
  nor_x1_sg U60606 ( .A(n46611), .B(n55643), .X(\L1_0/n4650 ) );
  nor_x1_sg U60607 ( .A(n46625), .B(n26791), .X(\L1_0/n4339 ) );
  nor_x1_sg U60608 ( .A(n46625), .B(n55681), .X(\L1_0/n4338 ) );
  nor_x1_sg U60609 ( .A(n46625), .B(n26798), .X(\L1_0/n4335 ) );
  nor_x1_sg U60610 ( .A(n46625), .B(n55682), .X(\L1_0/n4334 ) );
  nor_x1_sg U60611 ( .A(n46625), .B(n26805), .X(\L1_0/n4331 ) );
  nor_x1_sg U60612 ( .A(n46625), .B(n55683), .X(\L1_0/n4330 ) );
  nor_x1_sg U60613 ( .A(n46623), .B(n27350), .X(\L1_0/n4179 ) );
  nor_x1_sg U60614 ( .A(n46623), .B(n55701), .X(\L1_0/n4178 ) );
  nor_x1_sg U60615 ( .A(n46623), .B(n27357), .X(\L1_0/n4175 ) );
  nor_x1_sg U60616 ( .A(n46623), .B(n55702), .X(\L1_0/n4174 ) );
  nor_x1_sg U60617 ( .A(n46623), .B(n27364), .X(\L1_0/n4171 ) );
  nor_x1_sg U60618 ( .A(n46623), .B(n55703), .X(\L1_0/n4170 ) );
  nor_x1_sg U60619 ( .A(n46621), .B(n27630), .X(\L1_0/n4099 ) );
  nor_x1_sg U60620 ( .A(n46621), .B(n55711), .X(\L1_0/n4098 ) );
  nor_x1_sg U60621 ( .A(n46621), .B(n27637), .X(\L1_0/n4095 ) );
  nor_x1_sg U60622 ( .A(n46621), .B(n55712), .X(\L1_0/n4094 ) );
  nor_x1_sg U60623 ( .A(n46621), .B(n27644), .X(\L1_0/n4091 ) );
  nor_x1_sg U60624 ( .A(n46621), .B(n55713), .X(\L1_0/n4090 ) );
  nor_x1_sg U60625 ( .A(n46619), .B(n28747), .X(\L1_0/n3779 ) );
  nor_x1_sg U60626 ( .A(n46619), .B(n55751), .X(\L1_0/n3778 ) );
  nor_x1_sg U60627 ( .A(n46619), .B(n28754), .X(\L1_0/n3775 ) );
  nor_x1_sg U60628 ( .A(n46619), .B(n55752), .X(\L1_0/n3774 ) );
  nor_x1_sg U60629 ( .A(n46619), .B(n28761), .X(\L1_0/n3771 ) );
  nor_x1_sg U60630 ( .A(n46619), .B(n55753), .X(\L1_0/n3770 ) );
  nand_x4_sg U60631 ( .A(n52867), .B(n14872), .X(n14831) );
  nand_x4_sg U60632 ( .A(n51758), .B(n11760), .X(n11719) );
  nand_x4_sg U60633 ( .A(n10873), .B(n51444), .X(n10361) );
  nand_x1_sg U60634 ( .A(n10876), .B(n10875), .X(n10873) );
  nor_x1_sg U60635 ( .A(n10875), .B(n10876), .X(n10874) );
  nor_x1_sg U60636 ( .A(n16122), .B(n16123), .X(n16121) );
  nor_x1_sg U60637 ( .A(n10667), .B(n10668), .X(n10666) );
  nor_x1_sg U60638 ( .A(n18449), .B(n18450), .X(n18448) );
  nor_x1_sg U60639 ( .A(n19994), .B(n19995), .X(n19993) );
  nor_x1_sg U60640 ( .A(n21539), .B(n21540), .X(n21538) );
  nor_x1_sg U60641 ( .A(n11447), .B(n11448), .X(n11446) );
  nor_x1_sg U60642 ( .A(n13008), .B(n13009), .X(n13007) );
  nor_x1_sg U60643 ( .A(n15341), .B(n15342), .X(n15340) );
  nor_x1_sg U60644 ( .A(n16907), .B(n16908), .X(n16906) );
  nor_x1_sg U60645 ( .A(n12227), .B(n12228), .X(n12226) );
  inv_x4_sg U60646 ( .A(n45421), .X(n46614) );
  nor_x1_sg U60647 ( .A(n13756), .B(n13757), .X(n13754) );
  nand_x4_sg U60648 ( .A(n16328), .B(n53404), .X(n15807) );
  nor_x1_sg U60649 ( .A(n16330), .B(n16331), .X(n16329) );
  nand_x4_sg U60650 ( .A(n13994), .B(n52564), .X(n13473) );
  nor_x1_sg U60651 ( .A(n13996), .B(n13997), .X(n13995) );
  nor_x1_sg U60652 ( .A(n10636), .B(n10637), .X(n10634) );
  nor_x1_sg U60653 ( .A(n18418), .B(n18419), .X(n18416) );
  nor_x1_sg U60654 ( .A(n19963), .B(n19964), .X(n19961) );
  nor_x1_sg U60655 ( .A(n21508), .B(n21509), .X(n21506) );
  nor_x1_sg U60656 ( .A(n16090), .B(n16091), .X(n16088) );
  nor_x1_sg U60657 ( .A(n14528), .B(n14529), .X(n14526) );
  nor_x1_sg U60658 ( .A(n17649), .B(n17650), .X(n17647) );
  nor_x1_sg U60659 ( .A(n19194), .B(n19195), .X(n19192) );
  nor_x1_sg U60660 ( .A(n20738), .B(n20739), .X(n20736) );
  nor_x1_sg U60661 ( .A(n12195), .B(n12196), .X(n12193) );
  nand_x4_sg U60662 ( .A(n12433), .B(n52012), .X(n11911) );
  nor_x1_sg U60663 ( .A(n12435), .B(n12436), .X(n12434) );
  nand_x4_sg U60664 ( .A(n11653), .B(n51734), .X(n11128) );
  nor_x1_sg U60665 ( .A(n11655), .B(n11656), .X(n11654) );
  nand_x4_sg U60666 ( .A(n13214), .B(n52289), .X(n12689) );
  nor_x1_sg U60667 ( .A(n13216), .B(n13217), .X(n13215) );
  nand_x4_sg U60668 ( .A(n15547), .B(n53123), .X(n15022) );
  nor_x1_sg U60669 ( .A(n15549), .B(n15550), .X(n15548) );
  nand_x4_sg U60670 ( .A(n17113), .B(n53681), .X(n16588) );
  nor_x1_sg U60671 ( .A(n17115), .B(n17116), .X(n17114) );
  nand_x4_sg U60672 ( .A(n14719), .B(n14720), .X(n14662) );
  nand_x4_sg U60673 ( .A(n17840), .B(n17841), .X(n17783) );
  nand_x4_sg U60674 ( .A(n19385), .B(n19386), .X(n19328) );
  nand_x4_sg U60675 ( .A(n20929), .B(n20930), .X(n20872) );
  nand_x4_sg U60676 ( .A(n18511), .B(n18447), .X(n18464) );
  nand_x4_sg U60677 ( .A(n17742), .B(n17678), .X(n17695) );
  nand_x4_sg U60678 ( .A(n19287), .B(n19223), .X(n19240) );
  nand_x4_sg U60679 ( .A(n20831), .B(n20767), .X(n20784) );
  nand_x4_sg U60680 ( .A(n20056), .B(n19992), .X(n20009) );
  nand_x4_sg U60681 ( .A(n21601), .B(n21537), .X(n21554) );
  nand_x4_sg U60682 ( .A(n14621), .B(n14557), .X(n14574) );
  nand_x4_sg U60683 ( .A(n51554), .B(n11063), .X(n8862) );
  nand_x1_sg U60684 ( .A(n44685), .B(n11065), .X(n11063) );
  nand_x4_sg U60685 ( .A(n52111), .B(n12624), .X(n8824) );
  nand_x1_sg U60686 ( .A(n44683), .B(n12626), .X(n12624) );
  nand_x4_sg U60687 ( .A(n52945), .B(n14957), .X(n8963) );
  nand_x1_sg U60688 ( .A(n44681), .B(n14959), .X(n14957) );
  nand_x4_sg U60689 ( .A(n53503), .B(n16523), .X(n9280) );
  nand_x1_sg U60690 ( .A(n44679), .B(n16525), .X(n16523) );
  nand_x4_sg U60691 ( .A(n54221), .B(n18488), .X(n18461) );
  nand_x1_sg U60692 ( .A(n43472), .B(n18490), .X(n18488) );
  nor_x1_sg U60693 ( .A(n18490), .B(n43472), .X(n18491) );
  nor_x1_sg U60694 ( .A(n46278), .B(n9159), .X(\L2_0/n3076 ) );
  nor_x1_sg U60695 ( .A(n41968), .B(n46278), .X(\L2_0/n3064 ) );
  nor_x1_sg U60696 ( .A(n46278), .B(n9132), .X(\L2_0/n3052 ) );
  nor_x1_sg U60697 ( .A(n44389), .B(n46278), .X(\L2_0/n3040 ) );
  nor_x1_sg U60698 ( .A(n46278), .B(n9161), .X(\L2_0/n3028 ) );
  nor_x1_sg U60699 ( .A(n46549), .B(n8886), .X(\L2_0/n4036 ) );
  nor_x1_sg U60700 ( .A(n42002), .B(n46549), .X(\L2_0/n4024 ) );
  nor_x1_sg U60701 ( .A(n46549), .B(n8866), .X(\L2_0/n4012 ) );
  nor_x1_sg U60702 ( .A(n44134), .B(n46549), .X(\L2_0/n4000 ) );
  nor_x1_sg U60703 ( .A(n46549), .B(n8895), .X(\L2_0/n3988 ) );
  nor_x1_sg U60704 ( .A(n46505), .B(n8857), .X(\L2_0/n3876 ) );
  nor_x1_sg U60705 ( .A(n41994), .B(n46505), .X(\L2_0/n3864 ) );
  nor_x1_sg U60706 ( .A(n46505), .B(n8828), .X(\L2_0/n3852 ) );
  nor_x1_sg U60707 ( .A(n44126), .B(n46505), .X(\L2_0/n3840 ) );
  nor_x1_sg U60708 ( .A(n46505), .B(n8859), .X(\L2_0/n3828 ) );
  nor_x1_sg U60709 ( .A(n46460), .B(n8960), .X(\L2_0/n3716 ) );
  nor_x1_sg U60710 ( .A(n41988), .B(n46460), .X(\L2_0/n3704 ) );
  nor_x1_sg U60711 ( .A(n46460), .B(n8944), .X(\L2_0/n3692 ) );
  nor_x1_sg U60712 ( .A(n44399), .B(n46460), .X(\L2_0/n3680 ) );
  nor_x1_sg U60713 ( .A(n46460), .B(n9009), .X(\L2_0/n3668 ) );
  nor_x1_sg U60714 ( .A(n46415), .B(n9322), .X(\L2_0/n3556 ) );
  nor_x1_sg U60715 ( .A(n41980), .B(n46415), .X(\L2_0/n3544 ) );
  nor_x1_sg U60716 ( .A(n46415), .B(n9330), .X(\L2_0/n3532 ) );
  nor_x1_sg U60717 ( .A(n44114), .B(n46415), .X(\L2_0/n3520 ) );
  nor_x1_sg U60718 ( .A(n46415), .B(n9324), .X(\L2_0/n3508 ) );
  nor_x1_sg U60719 ( .A(n46370), .B(n9273), .X(\L2_0/n3396 ) );
  nor_x1_sg U60720 ( .A(n41974), .B(n46370), .X(\L2_0/n3384 ) );
  nor_x1_sg U60721 ( .A(n46370), .B(n9246), .X(\L2_0/n3372 ) );
  nor_x1_sg U60722 ( .A(n44397), .B(n46370), .X(\L2_0/n3360 ) );
  nor_x1_sg U60723 ( .A(n46370), .B(n9275), .X(\L2_0/n3348 ) );
  nor_x1_sg U60724 ( .A(n46323), .B(n9235), .X(\L2_0/n3236 ) );
  nor_x1_sg U60725 ( .A(n41972), .B(n46323), .X(\L2_0/n3224 ) );
  nor_x1_sg U60726 ( .A(n46323), .B(n9208), .X(\L2_0/n3212 ) );
  nor_x1_sg U60727 ( .A(n44393), .B(n46323), .X(\L2_0/n3200 ) );
  nor_x1_sg U60728 ( .A(n46323), .B(n9237), .X(\L2_0/n3188 ) );
  nor_x1_sg U60729 ( .A(n46527), .B(n8933), .X(\L2_0/n3956 ) );
  nor_x1_sg U60730 ( .A(n41998), .B(n46527), .X(\L2_0/n3944 ) );
  nor_x1_sg U60731 ( .A(n46527), .B(n8905), .X(\L2_0/n3932 ) );
  nor_x1_sg U60732 ( .A(n44130), .B(n46527), .X(\L2_0/n3920 ) );
  nor_x1_sg U60733 ( .A(n46527), .B(n8929), .X(\L2_0/n3908 ) );
  nor_x1_sg U60734 ( .A(n46437), .B(n8990), .X(\L2_0/n3636 ) );
  nor_x1_sg U60735 ( .A(n41984), .B(n46437), .X(\L2_0/n3624 ) );
  nor_x1_sg U60736 ( .A(n46437), .B(n8967), .X(\L2_0/n3612 ) );
  nor_x1_sg U60737 ( .A(n44118), .B(n46437), .X(\L2_0/n3600 ) );
  nor_x1_sg U60738 ( .A(n46437), .B(n8998), .X(\L2_0/n3588 ) );
  nor_x1_sg U60739 ( .A(n46483), .B(n8819), .X(\L2_0/n3796 ) );
  nor_x1_sg U60740 ( .A(n41990), .B(n46483), .X(\L2_0/n3784 ) );
  nor_x1_sg U60741 ( .A(n46483), .B(n8807), .X(\L2_0/n3772 ) );
  nor_x1_sg U60742 ( .A(n44122), .B(n46483), .X(\L2_0/n3760 ) );
  nor_x1_sg U60743 ( .A(n46483), .B(n8821), .X(\L2_0/n3748 ) );
  nor_x1_sg U60744 ( .A(n46393), .B(n9311), .X(\L2_0/n3476 ) );
  nor_x1_sg U60745 ( .A(n41976), .B(n46393), .X(\L2_0/n3464 ) );
  nor_x1_sg U60746 ( .A(n46393), .B(n9284), .X(\L2_0/n3452 ) );
  nor_x1_sg U60747 ( .A(n44110), .B(n46393), .X(\L2_0/n3440 ) );
  nor_x1_sg U60748 ( .A(n46393), .B(n9315), .X(\L2_0/n3428 ) );
  nor_x1_sg U60749 ( .A(n46258), .B(n9123), .X(\L2_0/n2996 ) );
  nor_x1_sg U60750 ( .A(n41966), .B(n46258), .X(\L2_0/n2984 ) );
  nor_x1_sg U60751 ( .A(n46258), .B(n9113), .X(\L2_0/n2972 ) );
  nor_x1_sg U60752 ( .A(n44387), .B(n46258), .X(\L2_0/n2960 ) );
  nor_x1_sg U60753 ( .A(n46258), .B(n9099), .X(\L2_0/n2948 ) );
  nand_x4_sg U60754 ( .A(n43246), .B(n17551), .X(n17538) );
  nand_x1_sg U60755 ( .A(n42363), .B(n41800), .X(n17551) );
  nand_x4_sg U60756 ( .A(n43244), .B(n19096), .X(n19083) );
  nand_x1_sg U60757 ( .A(n42361), .B(n41798), .X(n19096) );
  nand_x4_sg U60758 ( .A(n43242), .B(n20640), .X(n20627) );
  nand_x1_sg U60759 ( .A(n42359), .B(n41796), .X(n20640) );
  nand_x4_sg U60760 ( .A(n51632), .B(n11312), .X(n11303) );
  nand_x1_sg U60761 ( .A(n11313), .B(n11314), .X(n11312) );
  nand_x4_sg U60762 ( .A(n43240), .B(n12873), .X(n12864) );
  nand_x1_sg U60763 ( .A(n12874), .B(n12875), .X(n12873) );
  nand_x4_sg U60764 ( .A(n43238), .B(n15206), .X(n15197) );
  nand_x1_sg U60765 ( .A(n15207), .B(n15208), .X(n15206) );
  nand_x4_sg U60766 ( .A(n43236), .B(n16772), .X(n16763) );
  nand_x1_sg U60767 ( .A(n16773), .B(n16774), .X(n16772) );
  nand_x4_sg U60768 ( .A(n52261), .B(n13048), .X(n13025) );
  nand_x1_sg U60769 ( .A(n42455), .B(n13050), .X(n13048) );
  nor_x1_sg U60770 ( .A(n13050), .B(n42455), .X(n13051) );
  nand_x4_sg U60771 ( .A(n53095), .B(n15381), .X(n15358) );
  nand_x1_sg U60772 ( .A(n42453), .B(n15383), .X(n15381) );
  nor_x1_sg U60773 ( .A(n15383), .B(n42453), .X(n15384) );
  nand_x4_sg U60774 ( .A(n53653), .B(n16947), .X(n16924) );
  nand_x1_sg U60775 ( .A(n42451), .B(n16949), .X(n16947) );
  nor_x1_sg U60776 ( .A(n16949), .B(n42451), .X(n16950) );
  nand_x4_sg U60777 ( .A(n51705), .B(n11487), .X(n11464) );
  nand_x1_sg U60778 ( .A(n42457), .B(n11489), .X(n11487) );
  nor_x1_sg U60779 ( .A(n11489), .B(n42457), .X(n11490) );
  nand_x4_sg U60780 ( .A(n19859), .B(n19895), .X(n19894) );
  nand_x1_sg U60781 ( .A(n19896), .B(n19897), .X(n19895) );
  nand_x4_sg U60782 ( .A(n21404), .B(n21440), .X(n21439) );
  nand_x1_sg U60783 ( .A(n21441), .B(n21442), .X(n21440) );
  nor_x1_sg U60784 ( .A(n44136), .B(n46549), .X(\L2_0/n4004 ) );
  nor_x1_sg U60785 ( .A(n44132), .B(n46527), .X(\L2_0/n3924 ) );
  nor_x1_sg U60786 ( .A(n44128), .B(n46505), .X(\L2_0/n3844 ) );
  nor_x1_sg U60787 ( .A(n44124), .B(n46483), .X(\L2_0/n3764 ) );
  nor_x1_sg U60788 ( .A(n42879), .B(n46460), .X(\L2_0/n3688 ) );
  nor_x1_sg U60789 ( .A(n44120), .B(n46437), .X(\L2_0/n3604 ) );
  nor_x1_sg U60790 ( .A(n44116), .B(n46415), .X(\L2_0/n3524 ) );
  nor_x1_sg U60791 ( .A(n44112), .B(n46393), .X(\L2_0/n3444 ) );
  nor_x1_sg U60792 ( .A(n42889), .B(n46549), .X(\L2_0/n4008 ) );
  nor_x1_sg U60793 ( .A(n42887), .B(n46527), .X(\L2_0/n3928 ) );
  nor_x1_sg U60794 ( .A(n42883), .B(n46505), .X(\L2_0/n3848 ) );
  nor_x1_sg U60795 ( .A(n42881), .B(n46483), .X(\L2_0/n3768 ) );
  nor_x1_sg U60796 ( .A(n42875), .B(n46437), .X(\L2_0/n3608 ) );
  nor_x1_sg U60797 ( .A(n42873), .B(n46415), .X(\L2_0/n3528 ) );
  nor_x1_sg U60798 ( .A(n42869), .B(n46393), .X(\L2_0/n3448 ) );
  nor_x1_sg U60799 ( .A(n42867), .B(n46370), .X(\L2_0/n3368 ) );
  nor_x1_sg U60800 ( .A(n42863), .B(n46323), .X(\L2_0/n3208 ) );
  nor_x1_sg U60801 ( .A(n42859), .B(n46278), .X(\L2_0/n3048 ) );
  nor_x1_sg U60802 ( .A(n42857), .B(n46258), .X(\L2_0/n2968 ) );
  nor_x1_sg U60803 ( .A(n44094), .B(n46483), .X(\L2_0/n3812 ) );
  nand_x4_sg U60804 ( .A(n18589), .B(n18590), .X(n18531) );
  nand_x1_sg U60805 ( .A(n54127), .B(n54144), .X(n18589) );
  nand_x1_sg U60806 ( .A(n18583), .B(n18579), .X(n18590) );
  nand_x4_sg U60807 ( .A(n14424), .B(n14460), .X(n14459) );
  nand_x1_sg U60808 ( .A(n14461), .B(n14462), .X(n14460) );
  nand_x4_sg U60809 ( .A(n12312), .B(n51987), .X(n12363) );
  nand_x4_sg U60810 ( .A(n18314), .B(n18350), .X(n18349) );
  nand_x1_sg U60811 ( .A(n18351), .B(n18352), .X(n18350) );
  nand_x4_sg U60812 ( .A(n51633), .B(n11301), .X(n11277) );
  nand_x4_sg U60813 ( .A(n51914), .B(n12081), .X(n12056) );
  nand_x4_sg U60814 ( .A(n52189), .B(n12862), .X(n12838) );
  nand_x4_sg U60815 ( .A(n52466), .B(n13642), .X(n13617) );
  nand_x4_sg U60816 ( .A(n53023), .B(n15195), .X(n15171) );
  nand_x4_sg U60817 ( .A(n53301), .B(n15976), .X(n15951) );
  nand_x4_sg U60818 ( .A(n53581), .B(n16761), .X(n16737) );
  nand_x4_sg U60819 ( .A(n51362), .B(n10524), .X(n10503) );
  nand_x4_sg U60820 ( .A(n52752), .B(n14416), .X(n14394) );
  nand_x4_sg U60821 ( .A(n54151), .B(n18306), .X(n18284) );
  nand_x4_sg U60822 ( .A(n54716), .B(n19851), .X(n19830) );
  nand_x4_sg U60823 ( .A(n55284), .B(n21396), .X(n21375) );
  nand_x4_sg U60824 ( .A(n11150), .B(n11151), .X(n11088) );
  nand_x1_sg U60825 ( .A(n51623), .B(n11247), .X(n11150) );
  nand_x1_sg U60826 ( .A(n11084), .B(n11085), .X(n11151) );
  nand_x4_sg U60827 ( .A(n12711), .B(n12712), .X(n12649) );
  nand_x1_sg U60828 ( .A(n52182), .B(n12808), .X(n12711) );
  nand_x1_sg U60829 ( .A(n12645), .B(n12646), .X(n12712) );
  nand_x4_sg U60830 ( .A(n14275), .B(n14276), .X(n14212) );
  nand_x1_sg U60831 ( .A(n52734), .B(n14363), .X(n14275) );
  nand_x1_sg U60832 ( .A(n14208), .B(n14209), .X(n14276) );
  nand_x4_sg U60833 ( .A(n15044), .B(n15045), .X(n14982) );
  nand_x1_sg U60834 ( .A(n53016), .B(n15141), .X(n15044) );
  nand_x1_sg U60835 ( .A(n14978), .B(n14979), .X(n15045) );
  nand_x4_sg U60836 ( .A(n16610), .B(n16611), .X(n16548) );
  nand_x1_sg U60837 ( .A(n53574), .B(n16707), .X(n16610) );
  nand_x1_sg U60838 ( .A(n16544), .B(n16545), .X(n16611) );
  nand_x4_sg U60839 ( .A(n18165), .B(n18166), .X(n18103) );
  nand_x1_sg U60840 ( .A(n54134), .B(n18253), .X(n18165) );
  nand_x1_sg U60841 ( .A(n18099), .B(n18100), .X(n18166) );
  nand_x4_sg U60842 ( .A(n11333), .B(n11334), .X(n11331) );
  nand_x1_sg U60843 ( .A(n51653), .B(n11328), .X(n11333) );
  nand_x4_sg U60844 ( .A(n12113), .B(n12114), .X(n12111) );
  nand_x1_sg U60845 ( .A(n51934), .B(n12108), .X(n12113) );
  nand_x4_sg U60846 ( .A(n12894), .B(n12895), .X(n12892) );
  nand_x1_sg U60847 ( .A(n52209), .B(n12889), .X(n12894) );
  nand_x4_sg U60848 ( .A(n13674), .B(n13675), .X(n13672) );
  nand_x1_sg U60849 ( .A(n52486), .B(n13669), .X(n13674) );
  nand_x4_sg U60850 ( .A(n15227), .B(n15228), .X(n15225) );
  nand_x1_sg U60851 ( .A(n53043), .B(n15222), .X(n15227) );
  nand_x4_sg U60852 ( .A(n16008), .B(n16009), .X(n16006) );
  nand_x1_sg U60853 ( .A(n53322), .B(n16003), .X(n16008) );
  nand_x4_sg U60854 ( .A(n16793), .B(n16794), .X(n16791) );
  nand_x1_sg U60855 ( .A(n53601), .B(n16788), .X(n16793) );
  nand_x4_sg U60856 ( .A(n10560), .B(n10561), .X(n10558) );
  nand_x1_sg U60857 ( .A(n10555), .B(n51386), .X(n10560) );
  nand_x4_sg U60858 ( .A(n51722), .B(n11449), .X(n11404) );
  nand_x1_sg U60859 ( .A(n42801), .B(n11450), .X(n11449) );
  nor_x1_sg U60860 ( .A(n11450), .B(n42801), .X(n11451) );
  nand_x4_sg U60861 ( .A(n52276), .B(n13010), .X(n12965) );
  nand_x1_sg U60862 ( .A(n42797), .B(n13011), .X(n13010) );
  nor_x1_sg U60863 ( .A(n13011), .B(n42797), .X(n13012) );
  nand_x4_sg U60864 ( .A(n53110), .B(n15343), .X(n15298) );
  nand_x1_sg U60865 ( .A(n42793), .B(n15344), .X(n15343) );
  nor_x1_sg U60866 ( .A(n15344), .B(n42793), .X(n15345) );
  nand_x4_sg U60867 ( .A(n53668), .B(n16909), .X(n16864) );
  nand_x1_sg U60868 ( .A(n42791), .B(n16910), .X(n16909) );
  nor_x1_sg U60869 ( .A(n16910), .B(n42791), .X(n16911) );
  nand_x4_sg U60870 ( .A(n11456), .B(n11457), .X(n11454) );
  nand_x1_sg U60871 ( .A(n11450), .B(n42800), .X(n11457) );
  nand_x4_sg U60872 ( .A(n13017), .B(n13018), .X(n13015) );
  nand_x1_sg U60873 ( .A(n13011), .B(n42796), .X(n13018) );
  nand_x4_sg U60874 ( .A(n15350), .B(n15351), .X(n15348) );
  nand_x1_sg U60875 ( .A(n15344), .B(n42792), .X(n15351) );
  nand_x4_sg U60876 ( .A(n16916), .B(n16917), .X(n16914) );
  nand_x1_sg U60877 ( .A(n16910), .B(n42790), .X(n16917) );
  nand_x4_sg U60878 ( .A(n17572), .B(n17573), .X(n17570) );
  nand_x1_sg U60879 ( .A(n17567), .B(n53893), .X(n17572) );
  nand_x4_sg U60880 ( .A(n19117), .B(n19118), .X(n19115) );
  nand_x1_sg U60881 ( .A(n19112), .B(n54458), .X(n19117) );
  nand_x4_sg U60882 ( .A(n20661), .B(n20662), .X(n20659) );
  nand_x1_sg U60883 ( .A(n20656), .B(n55026), .X(n20661) );
  nand_x4_sg U60884 ( .A(n14619), .B(n14620), .X(n14617) );
  nand_x4_sg U60885 ( .A(n17740), .B(n17741), .X(n17738) );
  nand_x4_sg U60886 ( .A(n18509), .B(n18510), .X(n18507) );
  nand_x4_sg U60887 ( .A(n19285), .B(n19286), .X(n19283) );
  nand_x4_sg U60888 ( .A(n20829), .B(n20830), .X(n20827) );
  nand_x4_sg U60889 ( .A(n20054), .B(n20055), .X(n20052) );
  nand_x4_sg U60890 ( .A(n21599), .B(n21600), .X(n21597) );
  nand_x4_sg U60891 ( .A(n10727), .B(n10728), .X(n10725) );
  nand_x4_sg U60892 ( .A(n13551), .B(n13552), .X(n13540) );
  nand_x1_sg U60893 ( .A(n52401), .B(n13547), .X(n13551) );
  nand_x1_sg U60894 ( .A(n13546), .B(n52407), .X(n13552) );
  nand_x4_sg U60895 ( .A(n14701), .B(n14702), .X(n14642) );
  nand_x4_sg U60896 ( .A(n16162), .B(n16163), .X(n16139) );
  nand_x1_sg U60897 ( .A(n53366), .B(n42399), .X(n16163) );
  nand_x4_sg U60898 ( .A(n20033), .B(n20034), .X(n20006) );
  nand_x1_sg U60899 ( .A(n54781), .B(n42429), .X(n20034) );
  nand_x4_sg U60900 ( .A(n21578), .B(n21579), .X(n21551) );
  nand_x1_sg U60901 ( .A(n55349), .B(n42427), .X(n21579) );
  nand_x4_sg U60902 ( .A(n10706), .B(n10707), .X(n10679) );
  nand_x1_sg U60903 ( .A(n51422), .B(n43342), .X(n10707) );
  nand_x4_sg U60904 ( .A(n10770), .B(n10771), .X(n10762) );
  nand_x1_sg U60905 ( .A(n51468), .B(n42382), .X(n10771) );
  nand_x4_sg U60906 ( .A(n14659), .B(n14660), .X(n14654) );
  nand_x1_sg U60907 ( .A(n52857), .B(n42392), .X(n14660) );
  nand_x4_sg U60908 ( .A(n17780), .B(n17781), .X(n17775) );
  nand_x1_sg U60909 ( .A(n53977), .B(n42390), .X(n17781) );
  nand_x4_sg U60910 ( .A(n19325), .B(n19326), .X(n19320) );
  nand_x1_sg U60911 ( .A(n54542), .B(n42388), .X(n19326) );
  nand_x4_sg U60912 ( .A(n20869), .B(n20870), .X(n20864) );
  nand_x1_sg U60913 ( .A(n55110), .B(n42386), .X(n20870) );
  nand_x4_sg U60914 ( .A(n14598), .B(n14599), .X(n14571) );
  nand_x1_sg U60915 ( .A(n52812), .B(n43345), .X(n14599) );
  nand_x4_sg U60916 ( .A(n12267), .B(n12268), .X(n12244) );
  nand_x1_sg U60917 ( .A(n51977), .B(n43309), .X(n12268) );
  nor_x1_sg U60918 ( .A(n46278), .B(n9128), .X(\L2_0/n3084 ) );
  nor_x1_sg U60919 ( .A(n46278), .B(n9140), .X(\L2_0/n3080 ) );
  nor_x1_sg U60920 ( .A(n46278), .B(n9136), .X(\L2_0/n3072 ) );
  nor_x1_sg U60921 ( .A(n46278), .B(n9138), .X(\L2_0/n3068 ) );
  nor_x1_sg U60922 ( .A(n46278), .B(n9142), .X(\L2_0/n3060 ) );
  nor_x1_sg U60923 ( .A(n46278), .B(n9146), .X(\L2_0/n3056 ) );
  nor_x1_sg U60924 ( .A(n46278), .B(n9144), .X(\L2_0/n3044 ) );
  nor_x1_sg U60925 ( .A(n46278), .B(n9134), .X(\L2_0/n3036 ) );
  nor_x1_sg U60926 ( .A(n46278), .B(n9148), .X(\L2_0/n3032 ) );
  nor_x1_sg U60927 ( .A(n46549), .B(n8862), .X(\L2_0/n4044 ) );
  nor_x1_sg U60928 ( .A(n46549), .B(n8874), .X(\L2_0/n4040 ) );
  nor_x1_sg U60929 ( .A(n46549), .B(n8870), .X(\L2_0/n4032 ) );
  nor_x1_sg U60930 ( .A(n46549), .B(n8872), .X(\L2_0/n4028 ) );
  nor_x1_sg U60931 ( .A(n46549), .B(n8876), .X(\L2_0/n4020 ) );
  nor_x1_sg U60932 ( .A(n46549), .B(n8880), .X(\L2_0/n4016 ) );
  nor_x1_sg U60933 ( .A(n46549), .B(n8868), .X(\L2_0/n3996 ) );
  nor_x1_sg U60934 ( .A(n46549), .B(n8882), .X(\L2_0/n3992 ) );
  nor_x1_sg U60935 ( .A(n46505), .B(n8824), .X(\L2_0/n3884 ) );
  nor_x1_sg U60936 ( .A(n46505), .B(n8836), .X(\L2_0/n3880 ) );
  nor_x1_sg U60937 ( .A(n46505), .B(n8832), .X(\L2_0/n3872 ) );
  nor_x1_sg U60938 ( .A(n46505), .B(n8834), .X(\L2_0/n3868 ) );
  nor_x1_sg U60939 ( .A(n46505), .B(n8838), .X(\L2_0/n3860 ) );
  nor_x1_sg U60940 ( .A(n46505), .B(n8842), .X(\L2_0/n3856 ) );
  nor_x1_sg U60941 ( .A(n46505), .B(n8830), .X(\L2_0/n3836 ) );
  nor_x1_sg U60942 ( .A(n46505), .B(n8848), .X(\L2_0/n3832 ) );
  nor_x1_sg U60943 ( .A(n46460), .B(n8940), .X(\L2_0/n3724 ) );
  nor_x1_sg U60944 ( .A(n46460), .B(n8950), .X(\L2_0/n3720 ) );
  nor_x1_sg U60945 ( .A(n46460), .B(n8938), .X(\L2_0/n3712 ) );
  nor_x1_sg U60946 ( .A(n46460), .B(n8948), .X(\L2_0/n3708 ) );
  nor_x1_sg U60947 ( .A(n46460), .B(n8952), .X(\L2_0/n3700 ) );
  nor_x1_sg U60948 ( .A(n46460), .B(n8956), .X(\L2_0/n3696 ) );
  nor_x1_sg U60949 ( .A(n46460), .B(n8954), .X(\L2_0/n3684 ) );
  nor_x1_sg U60950 ( .A(n46460), .B(n8946), .X(\L2_0/n3676 ) );
  nor_x1_sg U60951 ( .A(n46460), .B(n9002), .X(\L2_0/n3672 ) );
  nor_x1_sg U60952 ( .A(n46415), .B(n41360), .X(\L2_0/n3564 ) );
  nor_x1_sg U60953 ( .A(n46415), .B(n9334), .X(\L2_0/n3560 ) );
  nor_x1_sg U60954 ( .A(n46415), .B(n9347), .X(\L2_0/n3552 ) );
  nor_x1_sg U60955 ( .A(n46415), .B(n9332), .X(\L2_0/n3548 ) );
  nor_x1_sg U60956 ( .A(n46415), .B(n9351), .X(\L2_0/n3540 ) );
  nor_x1_sg U60957 ( .A(n46415), .B(n9341), .X(\L2_0/n3536 ) );
  nor_x1_sg U60958 ( .A(n46415), .B(n9349), .X(\L2_0/n3516 ) );
  nor_x1_sg U60959 ( .A(n46415), .B(n9336), .X(\L2_0/n3512 ) );
  nor_x1_sg U60960 ( .A(n46370), .B(n9242), .X(\L2_0/n3404 ) );
  nor_x1_sg U60961 ( .A(n46370), .B(n9254), .X(\L2_0/n3400 ) );
  nor_x1_sg U60962 ( .A(n46370), .B(n9250), .X(\L2_0/n3392 ) );
  nor_x1_sg U60963 ( .A(n46370), .B(n9252), .X(\L2_0/n3388 ) );
  nor_x1_sg U60964 ( .A(n46370), .B(n9256), .X(\L2_0/n3380 ) );
  nor_x1_sg U60965 ( .A(n46370), .B(n9260), .X(\L2_0/n3376 ) );
  nor_x1_sg U60966 ( .A(n46370), .B(n9258), .X(\L2_0/n3364 ) );
  nor_x1_sg U60967 ( .A(n46370), .B(n9248), .X(\L2_0/n3356 ) );
  nor_x1_sg U60968 ( .A(n46370), .B(n9262), .X(\L2_0/n3352 ) );
  nor_x1_sg U60969 ( .A(n46323), .B(n9204), .X(\L2_0/n3244 ) );
  nor_x1_sg U60970 ( .A(n46323), .B(n9216), .X(\L2_0/n3240 ) );
  nor_x1_sg U60971 ( .A(n46323), .B(n9212), .X(\L2_0/n3232 ) );
  nor_x1_sg U60972 ( .A(n46323), .B(n9214), .X(\L2_0/n3228 ) );
  nor_x1_sg U60973 ( .A(n46323), .B(n9218), .X(\L2_0/n3220 ) );
  nor_x1_sg U60974 ( .A(n46323), .B(n9222), .X(\L2_0/n3216 ) );
  nor_x1_sg U60975 ( .A(n46323), .B(n9220), .X(\L2_0/n3204 ) );
  nor_x1_sg U60976 ( .A(n46323), .B(n9210), .X(\L2_0/n3196 ) );
  nor_x1_sg U60977 ( .A(n46323), .B(n9224), .X(\L2_0/n3192 ) );
  nor_x1_sg U60978 ( .A(n46527), .B(n41366), .X(\L2_0/n3964 ) );
  nor_x1_sg U60979 ( .A(n46527), .B(n8909), .X(\L2_0/n3960 ) );
  nor_x1_sg U60980 ( .A(n46527), .B(n8923), .X(\L2_0/n3952 ) );
  nor_x1_sg U60981 ( .A(n46527), .B(n8907), .X(\L2_0/n3948 ) );
  nor_x1_sg U60982 ( .A(n46527), .B(n8913), .X(\L2_0/n3940 ) );
  nor_x1_sg U60983 ( .A(n46527), .B(n8917), .X(\L2_0/n3936 ) );
  nor_x1_sg U60984 ( .A(n46527), .B(n8911), .X(\L2_0/n3916 ) );
  nor_x1_sg U60985 ( .A(n46527), .B(n8900), .X(\L2_0/n3912 ) );
  nor_x1_sg U60986 ( .A(n46437), .B(n8963), .X(\L2_0/n3644 ) );
  nor_x1_sg U60987 ( .A(n46437), .B(n8975), .X(\L2_0/n3640 ) );
  nor_x1_sg U60988 ( .A(n46437), .B(n8971), .X(\L2_0/n3632 ) );
  nor_x1_sg U60989 ( .A(n46437), .B(n8973), .X(\L2_0/n3628 ) );
  nor_x1_sg U60990 ( .A(n46437), .B(n8977), .X(\L2_0/n3620 ) );
  nor_x1_sg U60991 ( .A(n46437), .B(n8981), .X(\L2_0/n3616 ) );
  nor_x1_sg U60992 ( .A(n46437), .B(n8969), .X(\L2_0/n3596 ) );
  nor_x1_sg U60993 ( .A(n46437), .B(n8992), .X(\L2_0/n3592 ) );
  nor_x1_sg U60994 ( .A(n46483), .B(n41364), .X(\L2_0/n3804 ) );
  nor_x1_sg U60995 ( .A(n46483), .B(n8789), .X(\L2_0/n3800 ) );
  nor_x1_sg U60996 ( .A(n46483), .B(n8801), .X(\L2_0/n3792 ) );
  nor_x1_sg U60997 ( .A(n46483), .B(n8787), .X(\L2_0/n3788 ) );
  nor_x1_sg U60998 ( .A(n46483), .B(n41362), .X(\L2_0/n3780 ) );
  nor_x1_sg U60999 ( .A(n46483), .B(n8797), .X(\L2_0/n3776 ) );
  nor_x1_sg U61000 ( .A(n46483), .B(n8813), .X(\L2_0/n3756 ) );
  nor_x1_sg U61001 ( .A(n46483), .B(n8799), .X(\L2_0/n3752 ) );
  nor_x1_sg U61002 ( .A(n46393), .B(n9280), .X(\L2_0/n3484 ) );
  nor_x1_sg U61003 ( .A(n46393), .B(n9292), .X(\L2_0/n3480 ) );
  nor_x1_sg U61004 ( .A(n46393), .B(n9288), .X(\L2_0/n3472 ) );
  nor_x1_sg U61005 ( .A(n46393), .B(n9290), .X(\L2_0/n3468 ) );
  nor_x1_sg U61006 ( .A(n46393), .B(n9294), .X(\L2_0/n3460 ) );
  nor_x1_sg U61007 ( .A(n46393), .B(n9298), .X(\L2_0/n3456 ) );
  nor_x1_sg U61008 ( .A(n46393), .B(n9286), .X(\L2_0/n3436 ) );
  nor_x1_sg U61009 ( .A(n46393), .B(n9300), .X(\L2_0/n3432 ) );
  nor_x1_sg U61010 ( .A(n46258), .B(n9119), .X(\L2_0/n3004 ) );
  nor_x1_sg U61011 ( .A(n46258), .B(n9097), .X(\L2_0/n3000 ) );
  nor_x1_sg U61012 ( .A(n46258), .B(n9107), .X(\L2_0/n2992 ) );
  nor_x1_sg U61013 ( .A(n46258), .B(n9095), .X(\L2_0/n2988 ) );
  nor_x1_sg U61014 ( .A(n46258), .B(n9117), .X(\L2_0/n2980 ) );
  nor_x1_sg U61015 ( .A(n46258), .B(n9111), .X(\L2_0/n2976 ) );
  nor_x1_sg U61016 ( .A(n46258), .B(n9109), .X(\L2_0/n2964 ) );
  nor_x1_sg U61017 ( .A(n46258), .B(n9115), .X(\L2_0/n2956 ) );
  nor_x1_sg U61018 ( .A(n46258), .B(n9090), .X(\L2_0/n2952 ) );
  nand_x4_sg U61019 ( .A(n54189), .B(n18438), .X(n18421) );
  nand_x1_sg U61020 ( .A(n18429), .B(n18439), .X(n18438) );
  nand_x4_sg U61021 ( .A(n51400), .B(n10656), .X(n10639) );
  nand_x1_sg U61022 ( .A(n44082), .B(n10657), .X(n10656) );
  nand_x1_sg U61023 ( .A(n51308), .B(n51319), .X(n10657) );
  nand_x4_sg U61024 ( .A(n52046), .B(n12588), .X(n12573) );
  nand_x4_sg U61025 ( .A(n54756), .B(n19983), .X(n19966) );
  nand_x1_sg U61026 ( .A(n44080), .B(n19984), .X(n19983) );
  nand_x1_sg U61027 ( .A(n54662), .B(n54673), .X(n19984) );
  nand_x4_sg U61028 ( .A(n55324), .B(n21528), .X(n21511) );
  nand_x1_sg U61029 ( .A(n44078), .B(n21529), .X(n21528) );
  nand_x1_sg U61030 ( .A(n55230), .B(n55241), .X(n21529) );
  nand_x4_sg U61031 ( .A(n52530), .B(n13809), .X(n13752) );
  nand_x1_sg U61032 ( .A(n52491), .B(n13810), .X(n13809) );
  nand_x4_sg U61033 ( .A(n52578), .B(n13961), .X(n13948) );
  nand_x1_sg U61034 ( .A(n52505), .B(n52494), .X(n13962) );
  nand_x4_sg U61035 ( .A(n53960), .B(n17815), .X(n17787) );
  nand_x4_sg U61036 ( .A(n54525), .B(n19360), .X(n19332) );
  nand_x4_sg U61037 ( .A(n55093), .B(n20904), .X(n20876) );
  nand_x4_sg U61038 ( .A(n53397), .B(n16259), .X(n16231) );
  nand_x4_sg U61039 ( .A(n52840), .B(n14694), .X(n14666) );
  nand_x1_sg U61040 ( .A(n52726), .B(n52747), .X(n14695) );
  nand_x4_sg U61041 ( .A(n51348), .B(n10575), .X(n10535) );
  nand_x1_sg U61042 ( .A(n51347), .B(n10569), .X(n10575) );
  nor_x1_sg U61043 ( .A(n51347), .B(n10569), .X(n10576) );
  nand_x4_sg U61044 ( .A(n41875), .B(n10592), .X(n10589) );
  nand_x4_sg U61045 ( .A(n14483), .B(n14484), .X(n14481) );
  nand_x4_sg U61046 ( .A(n17604), .B(n17605), .X(n17602) );
  nand_x4_sg U61047 ( .A(n18373), .B(n18374), .X(n18371) );
  nand_x4_sg U61048 ( .A(n19149), .B(n19150), .X(n19147) );
  nand_x4_sg U61049 ( .A(n41879), .B(n19919), .X(n19916) );
  nand_x4_sg U61050 ( .A(n20693), .B(n20694), .X(n20691) );
  nand_x4_sg U61051 ( .A(n41877), .B(n21464), .X(n21461) );
  nand_x4_sg U61052 ( .A(n17397), .B(n17317), .X(n17323) );
  nand_x4_sg U61053 ( .A(n18942), .B(n18862), .X(n18868) );
  nand_x4_sg U61054 ( .A(n20486), .B(n20406), .X(n20412) );
  nand_x4_sg U61055 ( .A(n52453), .B(n13968), .X(n14149) );
  nand_x2_sg U61056 ( .A(n46500), .B(n26239), .X(n26238) );
  nand_x2_sg U61057 ( .A(n46432), .B(n27075), .X(n27074) );
  nand_x2_sg U61058 ( .A(n46388), .B(n27635), .X(n27634) );
  nand_x2_sg U61059 ( .A(n46345), .B(n28194), .X(n28193) );
  nand_x4_sg U61060 ( .A(n54702), .B(n19902), .X(n19862) );
  nand_x1_sg U61061 ( .A(n54701), .B(n19896), .X(n19902) );
  nor_x1_sg U61062 ( .A(n54701), .B(n19896), .X(n19903) );
  nand_x4_sg U61063 ( .A(n55270), .B(n21447), .X(n21407) );
  nand_x1_sg U61064 ( .A(n55269), .B(n21441), .X(n21447) );
  nor_x1_sg U61065 ( .A(n55269), .B(n21441), .X(n21448) );
  nand_x4_sg U61066 ( .A(n10885), .B(n51520), .X(n10369) );
  nand_x1_sg U61067 ( .A(n10888), .B(n43009), .X(n10885) );
  nor_x1_sg U61068 ( .A(n43009), .B(n10888), .X(n10886) );
  nand_x4_sg U61069 ( .A(n16340), .B(n53469), .X(n15815) );
  nand_x1_sg U61070 ( .A(n16343), .B(n42981), .X(n16340) );
  nor_x1_sg U61071 ( .A(n42981), .B(n16343), .X(n16341) );
  nand_x4_sg U61072 ( .A(n10925), .B(n51514), .X(n10888) );
  nand_x1_sg U61073 ( .A(n10928), .B(n44333), .X(n10925) );
  nor_x1_sg U61074 ( .A(n44333), .B(n10928), .X(n10926) );
  nand_x4_sg U61075 ( .A(n16383), .B(n53454), .X(n16343) );
  nand_x1_sg U61076 ( .A(n16386), .B(n44331), .X(n16383) );
  nor_x1_sg U61077 ( .A(n44331), .B(n16386), .X(n16384) );
  nand_x4_sg U61078 ( .A(n12474), .B(n52043), .X(n12452) );
  nand_x1_sg U61079 ( .A(n41431), .B(n12476), .X(n12474) );
  nor_x1_sg U61080 ( .A(n12476), .B(n52018), .X(n12475) );
  nand_x4_sg U61081 ( .A(n13255), .B(n52319), .X(n13233) );
  nand_x1_sg U61082 ( .A(n41430), .B(n13257), .X(n13255) );
  nor_x1_sg U61083 ( .A(n13257), .B(n52294), .X(n13256) );
  nand_x4_sg U61084 ( .A(n14035), .B(n52594), .X(n14013) );
  nand_x1_sg U61085 ( .A(n41585), .B(n14037), .X(n14035) );
  nor_x1_sg U61086 ( .A(n14037), .B(n52569), .X(n14036) );
  nand_x4_sg U61087 ( .A(n15588), .B(n53153), .X(n15566) );
  nand_x1_sg U61088 ( .A(n41429), .B(n15590), .X(n15588) );
  nor_x1_sg U61089 ( .A(n15590), .B(n53128), .X(n15589) );
  nand_x4_sg U61090 ( .A(n17154), .B(n53711), .X(n17132) );
  nand_x1_sg U61091 ( .A(n41427), .B(n17156), .X(n17154) );
  nor_x1_sg U61092 ( .A(n17156), .B(n53686), .X(n17155) );
  nand_x4_sg U61093 ( .A(n11695), .B(n51762), .X(n11672) );
  nand_x1_sg U61094 ( .A(n51739), .B(n11697), .X(n11695) );
  nor_x1_sg U61095 ( .A(n11697), .B(n51739), .X(n11696) );
  nand_x4_sg U61096 ( .A(n14807), .B(n52871), .X(n14784) );
  nand_x1_sg U61097 ( .A(n52849), .B(n14809), .X(n14807) );
  nor_x1_sg U61098 ( .A(n14809), .B(n52849), .X(n14808) );
  nand_x4_sg U61099 ( .A(n17928), .B(n53991), .X(n17905) );
  nand_x1_sg U61100 ( .A(n53969), .B(n17930), .X(n17928) );
  nor_x1_sg U61101 ( .A(n17930), .B(n53969), .X(n17929) );
  nand_x4_sg U61102 ( .A(n19473), .B(n54556), .X(n19450) );
  nand_x1_sg U61103 ( .A(n54534), .B(n19475), .X(n19473) );
  nor_x1_sg U61104 ( .A(n19475), .B(n54534), .X(n19474) );
  nand_x4_sg U61105 ( .A(n20243), .B(n54841), .X(n20219) );
  nand_x1_sg U61106 ( .A(n54819), .B(n20245), .X(n20243) );
  nor_x1_sg U61107 ( .A(n20245), .B(n54819), .X(n20244) );
  nand_x4_sg U61108 ( .A(n21017), .B(n55124), .X(n20994) );
  nand_x1_sg U61109 ( .A(n55102), .B(n21019), .X(n21017) );
  nor_x1_sg U61110 ( .A(n21019), .B(n55102), .X(n21018) );
  nand_x4_sg U61111 ( .A(n21788), .B(n55409), .X(n21764) );
  nand_x1_sg U61112 ( .A(n55387), .B(n21790), .X(n21788) );
  nor_x1_sg U61113 ( .A(n21790), .B(n55387), .X(n21789) );
  nand_x4_sg U61114 ( .A(n11713), .B(n51782), .X(n11711) );
  nand_x1_sg U61115 ( .A(n51781), .B(n11715), .X(n11713) );
  nor_x1_sg U61116 ( .A(n11715), .B(n51781), .X(n11714) );
  nand_x4_sg U61117 ( .A(n12493), .B(n52062), .X(n12491) );
  nand_x1_sg U61118 ( .A(n52061), .B(n12495), .X(n12493) );
  nor_x1_sg U61119 ( .A(n12495), .B(n52061), .X(n12494) );
  nand_x4_sg U61120 ( .A(n13274), .B(n52339), .X(n13272) );
  nand_x1_sg U61121 ( .A(n52338), .B(n13276), .X(n13274) );
  nor_x1_sg U61122 ( .A(n13276), .B(n52338), .X(n13275) );
  nand_x4_sg U61123 ( .A(n14054), .B(n52614), .X(n14052) );
  nand_x1_sg U61124 ( .A(n52613), .B(n14056), .X(n14054) );
  nor_x1_sg U61125 ( .A(n14056), .B(n52613), .X(n14055) );
  nand_x4_sg U61126 ( .A(n15607), .B(n53173), .X(n15605) );
  nand_x1_sg U61127 ( .A(n53172), .B(n15609), .X(n15607) );
  nor_x1_sg U61128 ( .A(n15609), .B(n53172), .X(n15608) );
  nand_x4_sg U61129 ( .A(n17173), .B(n53731), .X(n17171) );
  nand_x1_sg U61130 ( .A(n53730), .B(n17175), .X(n17173) );
  nor_x1_sg U61131 ( .A(n17175), .B(n53730), .X(n17174) );
  nand_x4_sg U61132 ( .A(n18715), .B(n54294), .X(n18713) );
  nand_x1_sg U61133 ( .A(n54293), .B(n18717), .X(n18715) );
  nor_x1_sg U61134 ( .A(n18717), .B(n54293), .X(n18716) );
  nand_x4_sg U61135 ( .A(n20261), .B(n54862), .X(n20259) );
  nand_x1_sg U61136 ( .A(n54861), .B(n20263), .X(n20261) );
  nor_x1_sg U61137 ( .A(n20263), .B(n54861), .X(n20262) );
  nand_x4_sg U61138 ( .A(n21806), .B(n55430), .X(n21804) );
  nand_x1_sg U61139 ( .A(n55429), .B(n21808), .X(n21806) );
  nor_x1_sg U61140 ( .A(n21808), .B(n55429), .X(n21807) );
  nand_x4_sg U61141 ( .A(n53453), .B(n16418), .X(n16386) );
  nand_x1_sg U61142 ( .A(n53441), .B(n16419), .X(n16418) );
  nor_x1_sg U61143 ( .A(n16419), .B(n53441), .X(n16420) );
  nand_x4_sg U61144 ( .A(n51513), .B(n10960), .X(n10928) );
  nand_x1_sg U61145 ( .A(n51492), .B(n10961), .X(n10960) );
  nor_x1_sg U61146 ( .A(n10961), .B(n51492), .X(n10962) );
  nand_x4_sg U61147 ( .A(n11557), .B(n11558), .X(n11504) );
  nand_x1_sg U61148 ( .A(n11489), .B(n42456), .X(n11557) );
  nand_x4_sg U61149 ( .A(n16232), .B(n16233), .X(n16179) );
  nand_x1_sg U61150 ( .A(n42399), .B(n16165), .X(n16232) );
  nand_x4_sg U61151 ( .A(n53858), .B(n17587), .X(n17547) );
  nand_x1_sg U61152 ( .A(n53857), .B(n17581), .X(n17587) );
  nor_x1_sg U61153 ( .A(n53857), .B(n17581), .X(n17588) );
  nand_x4_sg U61154 ( .A(n54423), .B(n19132), .X(n19092) );
  nand_x1_sg U61155 ( .A(n54422), .B(n19126), .X(n19132) );
  nor_x1_sg U61156 ( .A(n54422), .B(n19126), .X(n19133) );
  nand_x4_sg U61157 ( .A(n54991), .B(n20676), .X(n20636) );
  nand_x1_sg U61158 ( .A(n54990), .B(n20670), .X(n20676) );
  nor_x1_sg U61159 ( .A(n54990), .B(n20670), .X(n20677) );
  nand_x4_sg U61160 ( .A(n52738), .B(n14467), .X(n14427) );
  nand_x1_sg U61161 ( .A(n52737), .B(n14461), .X(n14467) );
  nor_x1_sg U61162 ( .A(n52737), .B(n14461), .X(n14468) );
  nand_x4_sg U61163 ( .A(n16261), .B(n16262), .X(n16207) );
  nand_x1_sg U61164 ( .A(n53309), .B(n16257), .X(n16262) );
  nand_x1_sg U61165 ( .A(n53284), .B(n16256), .X(n16261) );
  nand_x4_sg U61166 ( .A(n20101), .B(n20102), .X(n20050) );
  nand_x1_sg U61167 ( .A(n42429), .B(n20036), .X(n20101) );
  nand_x4_sg U61168 ( .A(n21646), .B(n21647), .X(n21595) );
  nand_x1_sg U61169 ( .A(n42427), .B(n21581), .X(n21646) );
  nand_x4_sg U61170 ( .A(n54138), .B(n18357), .X(n18317) );
  nand_x1_sg U61171 ( .A(n54137), .B(n18351), .X(n18357) );
  nor_x1_sg U61172 ( .A(n54137), .B(n18351), .X(n18358) );
  nand_x4_sg U61173 ( .A(n13118), .B(n13119), .X(n13065) );
  nand_x1_sg U61174 ( .A(n13050), .B(n42454), .X(n13118) );
  nand_x4_sg U61175 ( .A(n15451), .B(n15452), .X(n15398) );
  nand_x1_sg U61176 ( .A(n15383), .B(n42452), .X(n15451) );
  nand_x4_sg U61177 ( .A(n17017), .B(n17018), .X(n16964) );
  nand_x1_sg U61178 ( .A(n16949), .B(n42450), .X(n17017) );
  nand_x1_sg U61179 ( .A(n18490), .B(n43471), .X(n18556) );
  nand_x4_sg U61180 ( .A(n10688), .B(n10689), .X(n10618) );
  nand_x1_sg U61181 ( .A(n51378), .B(n10638), .X(n10689) );
  nand_x4_sg U61182 ( .A(n11469), .B(n11470), .X(n11396) );
  nand_x1_sg U61183 ( .A(n51657), .B(n11417), .X(n11470) );
  nand_x4_sg U61184 ( .A(n13030), .B(n13031), .X(n12957) );
  nand_x1_sg U61185 ( .A(n52213), .B(n12978), .X(n13031) );
  nand_x4_sg U61186 ( .A(n15363), .B(n15364), .X(n15290) );
  nand_x1_sg U61187 ( .A(n53047), .B(n15311), .X(n15364) );
  nand_x4_sg U61188 ( .A(n16929), .B(n16930), .X(n16856) );
  nand_x1_sg U61189 ( .A(n53605), .B(n16877), .X(n16930) );
  nand_x4_sg U61190 ( .A(n13810), .B(n13811), .X(n13737) );
  nand_x1_sg U61191 ( .A(n52490), .B(n13758), .X(n13811) );
  nand_x4_sg U61192 ( .A(n16144), .B(n16145), .X(n16071) );
  nand_x1_sg U61193 ( .A(n53326), .B(n16092), .X(n16145) );
  nand_x4_sg U61194 ( .A(n18479), .B(n54213), .X(n18417) );
  nand_x1_sg U61195 ( .A(n42803), .B(n18468), .X(n18479) );
  nor_x1_sg U61196 ( .A(n18468), .B(n42803), .X(n18480) );
  nand_x4_sg U61197 ( .A(n10775), .B(n10776), .X(n10723) );
  nand_x1_sg U61198 ( .A(n43342), .B(n10709), .X(n10775) );
  nand_x4_sg U61199 ( .A(n12249), .B(n12250), .X(n12176) );
  nand_x1_sg U61200 ( .A(n51938), .B(n12197), .X(n12250) );
  nand_x4_sg U61201 ( .A(n13411), .B(n52395), .X(n8789) );
  nor_x1_sg U61202 ( .A(n13413), .B(n13414), .X(n13412) );
  nand_x4_sg U61203 ( .A(n18596), .B(n18597), .X(n18554) );
  nand_x1_sg U61204 ( .A(n42123), .B(n54279), .X(n18597) );
  nand_x1_sg U61205 ( .A(n40537), .B(n18599), .X(n18596) );
  nand_x4_sg U61206 ( .A(n20142), .B(n54851), .X(n20099) );
  nor_x1_sg U61207 ( .A(n20144), .B(n20145), .X(n20143) );
  nand_x4_sg U61208 ( .A(n21687), .B(n55419), .X(n21644) );
  nor_x1_sg U61209 ( .A(n21689), .B(n21690), .X(n21688) );
  nand_x4_sg U61210 ( .A(n14708), .B(n52881), .X(n14665) );
  nor_x1_sg U61211 ( .A(n14710), .B(n14711), .X(n14709) );
  nand_x4_sg U61212 ( .A(n17829), .B(n54001), .X(n17786) );
  nor_x1_sg U61213 ( .A(n17831), .B(n17832), .X(n17830) );
  nand_x4_sg U61214 ( .A(n19374), .B(n54566), .X(n19331) );
  nor_x1_sg U61215 ( .A(n19376), .B(n19377), .X(n19375) );
  nand_x4_sg U61216 ( .A(n20918), .B(n55134), .X(n20875) );
  nor_x1_sg U61217 ( .A(n20920), .B(n20921), .X(n20919) );
  nand_x4_sg U61218 ( .A(n11398), .B(n51700), .X(n11367) );
  nor_x1_sg U61219 ( .A(n11400), .B(n11401), .X(n11399) );
  nand_x4_sg U61220 ( .A(n12959), .B(n52256), .X(n12928) );
  nor_x1_sg U61221 ( .A(n12961), .B(n12962), .X(n12960) );
  nand_x4_sg U61222 ( .A(n15292), .B(n53090), .X(n15261) );
  nor_x1_sg U61223 ( .A(n15294), .B(n15295), .X(n15293) );
  nand_x4_sg U61224 ( .A(n16858), .B(n53648), .X(n16827) );
  nor_x1_sg U61225 ( .A(n16860), .B(n16861), .X(n16859) );
  nor_x1_sg U61226 ( .A(n52397), .B(n44201), .X(n13525) );
  nand_x4_sg U61227 ( .A(n10866), .B(n10867), .X(n10865) );
  nand_x1_sg U61228 ( .A(n10361), .B(n42094), .X(n10866) );
  nand_x1_sg U61229 ( .A(n42093), .B(n51445), .X(n10867) );
  nand_x4_sg U61230 ( .A(n16321), .B(n16322), .X(n16320) );
  nand_x1_sg U61231 ( .A(n15807), .B(n42088), .X(n16321) );
  nand_x1_sg U61232 ( .A(n42087), .B(n53405), .X(n16322) );
  nand_x4_sg U61233 ( .A(n11646), .B(n11647), .X(n11645) );
  nand_x1_sg U61234 ( .A(n11128), .B(n42092), .X(n11646) );
  nand_x1_sg U61235 ( .A(n42091), .B(n51735), .X(n11647) );
  nand_x4_sg U61236 ( .A(n14758), .B(n14759), .X(n14757) );
  nand_x1_sg U61237 ( .A(n14252), .B(n42090), .X(n14758) );
  nand_x1_sg U61238 ( .A(n42089), .B(n52835), .X(n14759) );
  nand_x4_sg U61239 ( .A(n17879), .B(n17880), .X(n17878) );
  nand_x1_sg U61240 ( .A(n17371), .B(n42086), .X(n17879) );
  nand_x1_sg U61241 ( .A(n42085), .B(n53955), .X(n17880) );
  nand_x4_sg U61242 ( .A(n19424), .B(n19425), .X(n19423) );
  nand_x1_sg U61243 ( .A(n18916), .B(n42084), .X(n19424) );
  nand_x1_sg U61244 ( .A(n42083), .B(n54520), .X(n19425) );
  nand_x4_sg U61245 ( .A(n11596), .B(n11597), .X(n11555) );
  nand_x1_sg U61246 ( .A(n42135), .B(n51767), .X(n11597) );
  nand_x1_sg U61247 ( .A(n40531), .B(n11599), .X(n11596) );
  nand_x4_sg U61248 ( .A(n13157), .B(n13158), .X(n13116) );
  nand_x1_sg U61249 ( .A(n42131), .B(n52323), .X(n13158) );
  nand_x4_sg U61250 ( .A(n13878), .B(n13879), .X(n13848) );
  nand_x1_sg U61251 ( .A(n42105), .B(n52579), .X(n13879) );
  nand_x1_sg U61252 ( .A(n40548), .B(n13881), .X(n13878) );
  nand_x4_sg U61253 ( .A(n13937), .B(n13938), .X(n13896) );
  nand_x1_sg U61254 ( .A(n42129), .B(n52598), .X(n13938) );
  nand_x4_sg U61255 ( .A(n15490), .B(n15491), .X(n15449) );
  nand_x1_sg U61256 ( .A(n42127), .B(n53157), .X(n15491) );
  nand_x4_sg U61257 ( .A(n17056), .B(n17057), .X(n17015) );
  nand_x1_sg U61258 ( .A(n42125), .B(n53715), .X(n17057) );
  nand_x4_sg U61259 ( .A(n18646), .B(n18647), .X(n18645) );
  nand_x1_sg U61260 ( .A(n54239), .B(n42099), .X(n18646) );
  nand_x1_sg U61261 ( .A(n40558), .B(n44329), .X(n18647) );
  nand_x4_sg U61262 ( .A(n20968), .B(n20969), .X(n20967) );
  nand_x1_sg U61263 ( .A(n20460), .B(n42082), .X(n20968) );
  nand_x1_sg U61264 ( .A(n42081), .B(n55088), .X(n20969) );
  nand_x4_sg U61265 ( .A(n20192), .B(n20193), .X(n20191) );
  nand_x1_sg U61266 ( .A(n54804), .B(n42098), .X(n20192) );
  nand_x1_sg U61267 ( .A(n42097), .B(n45417), .X(n20193) );
  nand_x4_sg U61268 ( .A(n21737), .B(n21738), .X(n21736) );
  nand_x1_sg U61269 ( .A(n55372), .B(n42096), .X(n21737) );
  nand_x1_sg U61270 ( .A(n42095), .B(n45415), .X(n21738) );
  nand_x4_sg U61271 ( .A(n12426), .B(n12427), .X(n12425) );
  nand_x1_sg U61272 ( .A(n11911), .B(n42080), .X(n12426) );
  nand_x1_sg U61273 ( .A(n42079), .B(n52013), .X(n12427) );
  nand_x4_sg U61274 ( .A(n13207), .B(n13208), .X(n13206) );
  nand_x1_sg U61275 ( .A(n12689), .B(n42078), .X(n13207) );
  nand_x1_sg U61276 ( .A(n42077), .B(n52290), .X(n13208) );
  nand_x4_sg U61277 ( .A(n13987), .B(n13988), .X(n13986) );
  nand_x1_sg U61278 ( .A(n13473), .B(n42075), .X(n13987) );
  nand_x1_sg U61279 ( .A(n40550), .B(n52565), .X(n13988) );
  nand_x4_sg U61280 ( .A(n15540), .B(n15541), .X(n15539) );
  nand_x1_sg U61281 ( .A(n15022), .B(n42074), .X(n15540) );
  nand_x1_sg U61282 ( .A(n42073), .B(n53124), .X(n15541) );
  nand_x4_sg U61283 ( .A(n17106), .B(n17107), .X(n17105) );
  nand_x1_sg U61284 ( .A(n16588), .B(n42070), .X(n17106) );
  nand_x1_sg U61285 ( .A(n42069), .B(n53682), .X(n17107) );
  nand_x4_sg U61286 ( .A(n10736), .B(n10737), .X(n10668) );
  nand_x1_sg U61287 ( .A(n43100), .B(n51390), .X(n10737) );
  nand_x1_sg U61288 ( .A(n40541), .B(n10739), .X(n10736) );
  nand_x4_sg U61289 ( .A(n11953), .B(n11954), .X(n11852) );
  nand_x1_sg U61290 ( .A(n44327), .B(n51836), .X(n11954) );
  nand_x1_sg U61291 ( .A(n51842), .B(n11956), .X(n11953) );
  nand_x4_sg U61292 ( .A(n15848), .B(n15849), .X(n15747) );
  nand_x1_sg U61293 ( .A(n43141), .B(n53224), .X(n15849) );
  nand_x1_sg U61294 ( .A(n43140), .B(n15851), .X(n15848) );
  nand_x4_sg U61295 ( .A(n16272), .B(n16273), .X(n16226) );
  nand_x1_sg U61296 ( .A(n42120), .B(n53437), .X(n16273) );
  nand_x1_sg U61297 ( .A(n42119), .B(n16275), .X(n16272) );
  nand_x4_sg U61298 ( .A(n11508), .B(n11461), .X(n11506) );
  nand_x4_sg U61299 ( .A(n13069), .B(n13022), .X(n13067) );
  nand_x4_sg U61300 ( .A(n15402), .B(n15355), .X(n15400) );
  nand_x4_sg U61301 ( .A(n16968), .B(n16921), .X(n16966) );
  nand_x4_sg U61302 ( .A(n13414), .B(n13413), .X(n13411) );
  nand_x4_sg U61303 ( .A(n14667), .B(n14668), .X(n14615) );
  nand_x1_sg U61304 ( .A(n43345), .B(n14601), .X(n14667) );
  nand_x4_sg U61305 ( .A(n12296), .B(n12297), .X(n12228) );
  nand_x1_sg U61306 ( .A(n12298), .B(n12299), .X(n12296) );
  nand_x4_sg U61307 ( .A(n13857), .B(n13858), .X(n13789) );
  nand_x1_sg U61308 ( .A(n13859), .B(n13860), .X(n13857) );
  nand_x4_sg U61309 ( .A(n12289), .B(n12225), .X(n12239) );
  nand_x1_sg U61310 ( .A(n51948), .B(n12298), .X(n12289) );
  nand_x4_sg U61311 ( .A(n13850), .B(n13786), .X(n13800) );
  nand_x1_sg U61312 ( .A(n52500), .B(n13859), .X(n13850) );
  nand_x4_sg U61313 ( .A(n20264), .B(n20265), .X(n20263) );
  nand_x1_sg U61314 ( .A(n41895), .B(n20269), .X(n20264) );
  nor_x1_sg U61315 ( .A(n54836), .B(n54791), .X(n20266) );
  nand_x4_sg U61316 ( .A(n21809), .B(n21810), .X(n21808) );
  nand_x1_sg U61317 ( .A(n41889), .B(n21814), .X(n21809) );
  nor_x1_sg U61318 ( .A(n55404), .B(n55359), .X(n21811) );
  nand_x4_sg U61319 ( .A(n16191), .B(n16192), .X(n16123) );
  nand_x1_sg U61320 ( .A(n16193), .B(n16194), .X(n16191) );
  nand_x4_sg U61321 ( .A(n16184), .B(n16120), .X(n16134) );
  nand_x1_sg U61322 ( .A(n53336), .B(n16193), .X(n16184) );
  nand_x4_sg U61323 ( .A(n12337), .B(n12338), .X(n12284) );
  nand_x1_sg U61324 ( .A(n43309), .B(n12270), .X(n12337) );
  nand_x4_sg U61325 ( .A(n18517), .B(n18518), .X(n18450) );
  nand_x1_sg U61326 ( .A(n18519), .B(n18520), .X(n18517) );
  nand_x1_sg U61327 ( .A(n54201), .B(n54179), .X(n18518) );
  nand_x4_sg U61328 ( .A(n11716), .B(n11717), .X(n11715) );
  nand_x1_sg U61329 ( .A(n41917), .B(n11721), .X(n11716) );
  nor_x1_sg U61330 ( .A(n51757), .B(n51707), .X(n11718) );
  nand_x4_sg U61331 ( .A(n52492), .B(n13720), .X(n13709) );
  nand_x1_sg U61332 ( .A(n52485), .B(n52478), .X(n13720) );
  nand_x4_sg U61333 ( .A(n14580), .B(n14581), .X(n14510) );
  nand_x1_sg U61334 ( .A(n52764), .B(n14530), .X(n14581) );
  nand_x4_sg U61335 ( .A(n17701), .B(n17702), .X(n17631) );
  nand_x1_sg U61336 ( .A(n53884), .B(n17651), .X(n17702) );
  nand_x4_sg U61337 ( .A(n19246), .B(n19247), .X(n19176) );
  nand_x1_sg U61338 ( .A(n54449), .B(n19196), .X(n19247) );
  nand_x4_sg U61339 ( .A(n20790), .B(n20791), .X(n20720) );
  nand_x1_sg U61340 ( .A(n55017), .B(n20740), .X(n20791) );
  nand_x4_sg U61341 ( .A(n16123), .B(n16122), .X(n16120) );
  nand_x4_sg U61342 ( .A(n20015), .B(n20016), .X(n19945) );
  nand_x1_sg U61343 ( .A(n54732), .B(n19965), .X(n20016) );
  nand_x4_sg U61344 ( .A(n21560), .B(n21561), .X(n21490) );
  nand_x1_sg U61345 ( .A(n55300), .B(n21510), .X(n21561) );
  nand_x4_sg U61346 ( .A(n17749), .B(n17750), .X(n17681) );
  nand_x1_sg U61347 ( .A(n17751), .B(n43941), .X(n17749) );
  nand_x1_sg U61348 ( .A(n53918), .B(n53899), .X(n17750) );
  nand_x4_sg U61349 ( .A(n19294), .B(n19295), .X(n19226) );
  nand_x1_sg U61350 ( .A(n19296), .B(n43940), .X(n19294) );
  nand_x1_sg U61351 ( .A(n54483), .B(n54464), .X(n19295) );
  nand_x4_sg U61352 ( .A(n20838), .B(n20839), .X(n20770) );
  nand_x1_sg U61353 ( .A(n20840), .B(n43939), .X(n20838) );
  nand_x1_sg U61354 ( .A(n55051), .B(n55032), .X(n20839) );
  nand_x4_sg U61355 ( .A(n13277), .B(n13278), .X(n13276) );
  nand_x1_sg U61356 ( .A(n41915), .B(n13281), .X(n13277) );
  nor_x1_sg U61357 ( .A(n52296), .B(n52263), .X(n13279) );
  nand_x4_sg U61358 ( .A(n14057), .B(n14058), .X(n14056) );
  nand_x1_sg U61359 ( .A(n41914), .B(n14061), .X(n14057) );
  nor_x1_sg U61360 ( .A(n52571), .B(n52539), .X(n14059) );
  nand_x4_sg U61361 ( .A(n15610), .B(n15611), .X(n15609) );
  nand_x1_sg U61362 ( .A(n41910), .B(n15614), .X(n15610) );
  nor_x1_sg U61363 ( .A(n53130), .B(n53097), .X(n15612) );
  nand_x4_sg U61364 ( .A(n17176), .B(n17177), .X(n17175) );
  nand_x1_sg U61365 ( .A(n41909), .B(n17180), .X(n17176) );
  nor_x1_sg U61366 ( .A(n53688), .B(n53655), .X(n17178) );
  nand_x4_sg U61367 ( .A(n13077), .B(n13078), .X(n13009) );
  nand_x1_sg U61368 ( .A(n13079), .B(n13080), .X(n13077) );
  nand_x4_sg U61369 ( .A(n15410), .B(n15411), .X(n15342) );
  nand_x1_sg U61370 ( .A(n15412), .B(n15413), .X(n15410) );
  nand_x4_sg U61371 ( .A(n16976), .B(n16977), .X(n16908) );
  nand_x1_sg U61372 ( .A(n16978), .B(n16979), .X(n16976) );
  nand_x4_sg U61373 ( .A(n13070), .B(n13006), .X(n13020) );
  nand_x1_sg U61374 ( .A(n52223), .B(n13079), .X(n13070) );
  nand_x4_sg U61375 ( .A(n15403), .B(n15339), .X(n15353) );
  nand_x1_sg U61376 ( .A(n53057), .B(n15412), .X(n15403) );
  nand_x4_sg U61377 ( .A(n16969), .B(n16905), .X(n16919) );
  nand_x1_sg U61378 ( .A(n53615), .B(n16978), .X(n16969) );
  nand_x4_sg U61379 ( .A(n20062), .B(n20063), .X(n19995) );
  nand_x1_sg U61380 ( .A(n20064), .B(n20065), .X(n20062) );
  nand_x1_sg U61381 ( .A(n54769), .B(n54746), .X(n20063) );
  nand_x4_sg U61382 ( .A(n21607), .B(n21608), .X(n21540) );
  nand_x1_sg U61383 ( .A(n21609), .B(n21610), .X(n21607) );
  nand_x1_sg U61384 ( .A(n55337), .B(n55314), .X(n21608) );
  nand_x4_sg U61385 ( .A(n11516), .B(n11517), .X(n11448) );
  nand_x1_sg U61386 ( .A(n11518), .B(n11519), .X(n11516) );
  nand_x4_sg U61387 ( .A(n11509), .B(n11445), .X(n11459) );
  nand_x1_sg U61388 ( .A(n51667), .B(n11518), .X(n11509) );
  nand_x4_sg U61389 ( .A(n14628), .B(n14629), .X(n14560) );
  nand_x1_sg U61390 ( .A(n14630), .B(n14631), .X(n14628) );
  nand_x1_sg U61391 ( .A(n52797), .B(n52779), .X(n14629) );
  nand_x4_sg U61392 ( .A(n10668), .B(n10667), .X(n10665) );
  nand_x4_sg U61393 ( .A(n18450), .B(n18449), .X(n18447) );
  nand_x4_sg U61394 ( .A(n19995), .B(n19994), .X(n19992) );
  nand_x4_sg U61395 ( .A(n21540), .B(n21539), .X(n21537) );
  nand_x4_sg U61396 ( .A(n11448), .B(n11447), .X(n11445) );
  nand_x4_sg U61397 ( .A(n13009), .B(n13008), .X(n13006) );
  nand_x4_sg U61398 ( .A(n15342), .B(n15341), .X(n15339) );
  nand_x4_sg U61399 ( .A(n16908), .B(n16907), .X(n16905) );
  nand_x4_sg U61400 ( .A(n14828), .B(n14829), .X(n14827) );
  nand_x1_sg U61401 ( .A(n41913), .B(n14833), .X(n14828) );
  nor_x1_sg U61402 ( .A(n52866), .B(n52808), .X(n14830) );
  nand_x4_sg U61403 ( .A(n18718), .B(n18719), .X(n18717) );
  nand_x1_sg U61404 ( .A(n41901), .B(n18723), .X(n18718) );
  nor_x1_sg U61405 ( .A(n54269), .B(n54224), .X(n18720) );
  nand_x4_sg U61406 ( .A(n12228), .B(n12227), .X(n12225) );
  nand_x4_sg U61407 ( .A(n17418), .B(n17399), .X(n17312) );
  nand_x1_sg U61408 ( .A(n17419), .B(n17420), .X(n17418) );
  nand_x4_sg U61409 ( .A(n18963), .B(n18944), .X(n18857) );
  nand_x1_sg U61410 ( .A(n18964), .B(n18965), .X(n18963) );
  nand_x4_sg U61411 ( .A(n20507), .B(n20488), .X(n20401) );
  nand_x1_sg U61412 ( .A(n20508), .B(n20509), .X(n20507) );
  nand_x4_sg U61413 ( .A(n10816), .B(n10817), .X(n10769) );
  nand_x1_sg U61414 ( .A(n51454), .B(n51488), .X(n10817) );
  nand_x4_sg U61415 ( .A(n11361), .B(n11362), .X(n11332) );
  nand_x4_sg U61416 ( .A(n12141), .B(n12142), .X(n12112) );
  nand_x4_sg U61417 ( .A(n12922), .B(n12923), .X(n12893) );
  nand_x4_sg U61418 ( .A(n13702), .B(n13703), .X(n13673) );
  nand_x4_sg U61419 ( .A(n15255), .B(n15256), .X(n15226) );
  nand_x4_sg U61420 ( .A(n16036), .B(n16037), .X(n16007) );
  nand_x4_sg U61421 ( .A(n16821), .B(n16822), .X(n16792) );
  nand_x4_sg U61422 ( .A(n11368), .B(n11369), .X(n11366) );
  nand_x1_sg U61423 ( .A(n51660), .B(n11363), .X(n11369) );
  nand_x4_sg U61424 ( .A(n12148), .B(n12149), .X(n12146) );
  nand_x1_sg U61425 ( .A(n51941), .B(n12143), .X(n12149) );
  nand_x4_sg U61426 ( .A(n12929), .B(n12930), .X(n12927) );
  nand_x1_sg U61427 ( .A(n52216), .B(n12924), .X(n12930) );
  nand_x4_sg U61428 ( .A(n13709), .B(n13710), .X(n13707) );
  nand_x1_sg U61429 ( .A(n52493), .B(n13704), .X(n13710) );
  nand_x4_sg U61430 ( .A(n15262), .B(n15263), .X(n15260) );
  nand_x1_sg U61431 ( .A(n53050), .B(n15257), .X(n15263) );
  nand_x4_sg U61432 ( .A(n16043), .B(n16044), .X(n16041) );
  nand_x1_sg U61433 ( .A(n53329), .B(n16038), .X(n16044) );
  nand_x4_sg U61434 ( .A(n16828), .B(n16829), .X(n16826) );
  nand_x1_sg U61435 ( .A(n53608), .B(n16823), .X(n16829) );
  nand_x4_sg U61436 ( .A(n11153), .B(n11074), .X(n11080) );
  nand_x4_sg U61437 ( .A(n12714), .B(n12635), .X(n12641) );
  nand_x4_sg U61438 ( .A(n15047), .B(n14968), .X(n14974) );
  nand_x4_sg U61439 ( .A(n16613), .B(n16534), .X(n16540) );
  nand_x4_sg U61440 ( .A(n11223), .B(n11224), .X(n11081) );
  nand_x4_sg U61441 ( .A(n12784), .B(n12785), .X(n12642) );
  nand_x4_sg U61442 ( .A(n13561), .B(n13562), .X(n13426) );
  nand_x4_sg U61443 ( .A(n15895), .B(n15896), .X(n15759) );
  nand_x4_sg U61444 ( .A(n18229), .B(n18230), .X(n18096) );
  nand_x1_sg U61445 ( .A(n54103), .B(n54118), .X(n18230) );
  nand_x4_sg U61446 ( .A(n16683), .B(n16684), .X(n16541) );
  nand_x4_sg U61447 ( .A(n10584), .B(n10585), .X(n10559) );
  nand_x1_sg U61448 ( .A(n51402), .B(n51388), .X(n10585) );
  nand_x4_sg U61449 ( .A(n14476), .B(n14477), .X(n14451) );
  nand_x1_sg U61450 ( .A(n52791), .B(n52776), .X(n14477) );
  nand_x4_sg U61451 ( .A(n17597), .B(n17598), .X(n17571) );
  nand_x1_sg U61452 ( .A(n53911), .B(n53896), .X(n17598) );
  nand_x4_sg U61453 ( .A(n18366), .B(n18367), .X(n18341) );
  nand_x1_sg U61454 ( .A(n54191), .B(n54176), .X(n18367) );
  nand_x4_sg U61455 ( .A(n19142), .B(n19143), .X(n19116) );
  nand_x1_sg U61456 ( .A(n54476), .B(n54461), .X(n19143) );
  nand_x4_sg U61457 ( .A(n19911), .B(n19912), .X(n19886) );
  nand_x1_sg U61458 ( .A(n54758), .B(n54743), .X(n19912) );
  nand_x4_sg U61459 ( .A(n20686), .B(n20687), .X(n20660) );
  nand_x1_sg U61460 ( .A(n55044), .B(n55029), .X(n20687) );
  nand_x4_sg U61461 ( .A(n21456), .B(n21457), .X(n21431) );
  nand_x1_sg U61462 ( .A(n55326), .B(n55311), .X(n21457) );
  nand_x4_sg U61463 ( .A(n12000), .B(n12001), .X(n11864) );
  nand_x4_sg U61464 ( .A(n15117), .B(n15118), .X(n14975) );
  nand_x4_sg U61465 ( .A(n10680), .B(n10681), .X(n10672) );
  nand_x1_sg U61466 ( .A(n51412), .B(n51438), .X(n10681) );
  nand_x4_sg U61467 ( .A(n14572), .B(n14573), .X(n14564) );
  nand_x1_sg U61468 ( .A(n52801), .B(n52827), .X(n14573) );
  nand_x4_sg U61469 ( .A(n17693), .B(n17694), .X(n17685) );
  nand_x1_sg U61470 ( .A(n53922), .B(n53947), .X(n17694) );
  nand_x4_sg U61471 ( .A(n18462), .B(n18463), .X(n18454) );
  nand_x1_sg U61472 ( .A(n54205), .B(n54232), .X(n18463) );
  nand_x4_sg U61473 ( .A(n19238), .B(n19239), .X(n19230) );
  nand_x1_sg U61474 ( .A(n54487), .B(n54512), .X(n19239) );
  nand_x4_sg U61475 ( .A(n20007), .B(n20008), .X(n19999) );
  nand_x1_sg U61476 ( .A(n54773), .B(n54797), .X(n20008) );
  nand_x4_sg U61477 ( .A(n20782), .B(n20783), .X(n20774) );
  nand_x1_sg U61478 ( .A(n55055), .B(n55080), .X(n20783) );
  nand_x4_sg U61479 ( .A(n21552), .B(n21553), .X(n21544) );
  nand_x1_sg U61480 ( .A(n55341), .B(n55365), .X(n21553) );
  nand_x4_sg U61481 ( .A(n20100), .B(n20047), .X(n20098) );
  nand_x4_sg U61482 ( .A(n21645), .B(n21592), .X(n21643) );
  nand_x4_sg U61483 ( .A(n11936), .B(n11857), .X(n11863) );
  nand_x4_sg U61484 ( .A(n15831), .B(n15752), .X(n15758) );
  nor_x1_sg U61485 ( .A(n43850), .B(n52426), .X(n13579) );
  nor_x1_sg U61486 ( .A(n44385), .B(n53822), .X(n17480) );
  nor_x1_sg U61487 ( .A(n44383), .B(n54387), .X(n19025) );
  nor_x1_sg U61488 ( .A(n44381), .B(n54955), .X(n20569) );
  nor_x1_sg U61489 ( .A(n44106), .B(n51314), .X(n10466) );
  nor_x1_sg U61490 ( .A(n43984), .B(n54668), .X(n19793) );
  nor_x1_sg U61491 ( .A(n43982), .B(n55236), .X(n21338) );
  nor_x1_sg U61492 ( .A(n44104), .B(n52703), .X(n14358) );
  nand_x4_sg U61493 ( .A(n10494), .B(n10495), .X(n10470) );
  nand_x1_sg U61494 ( .A(n10496), .B(n10497), .X(n10495) );
  nand_x1_sg U61495 ( .A(n10499), .B(n51343), .X(n10494) );
  nand_x1_sg U61496 ( .A(n51343), .B(n10498), .X(n10497) );
  nand_x4_sg U61497 ( .A(n14385), .B(n14386), .X(n14362) );
  nand_x1_sg U61498 ( .A(n14387), .B(n14388), .X(n14386) );
  nand_x1_sg U61499 ( .A(n14390), .B(n52733), .X(n14385) );
  nand_x1_sg U61500 ( .A(n52733), .B(n14389), .X(n14388) );
  nand_x4_sg U61501 ( .A(n18275), .B(n18276), .X(n18252) );
  nand_x1_sg U61502 ( .A(n18277), .B(n18278), .X(n18276) );
  nand_x1_sg U61503 ( .A(n18281), .B(n18279), .X(n18275) );
  nand_x4_sg U61504 ( .A(n19821), .B(n19822), .X(n19797) );
  nand_x1_sg U61505 ( .A(n19823), .B(n19824), .X(n19822) );
  nand_x1_sg U61506 ( .A(n19826), .B(n54697), .X(n19821) );
  nand_x1_sg U61507 ( .A(n54697), .B(n19825), .X(n19824) );
  nand_x4_sg U61508 ( .A(n21366), .B(n21367), .X(n21342) );
  nand_x1_sg U61509 ( .A(n21368), .B(n21369), .X(n21367) );
  nand_x1_sg U61510 ( .A(n21371), .B(n55265), .X(n21366) );
  nand_x1_sg U61511 ( .A(n55265), .B(n21370), .X(n21369) );
  nand_x4_sg U61512 ( .A(n16089), .B(n16143), .X(n16086) );
  nand_x1_sg U61513 ( .A(n53327), .B(n16144), .X(n16143) );
  nand_x4_sg U61514 ( .A(n10635), .B(n10687), .X(n10632) );
  nand_x1_sg U61515 ( .A(n51379), .B(n10688), .X(n10687) );
  nand_x4_sg U61516 ( .A(n18417), .B(n18469), .X(n18414) );
  nand_x1_sg U61517 ( .A(n54167), .B(n18470), .X(n18469) );
  nand_x4_sg U61518 ( .A(n19962), .B(n20014), .X(n19959) );
  nand_x1_sg U61519 ( .A(n54733), .B(n20015), .X(n20014) );
  nand_x4_sg U61520 ( .A(n21507), .B(n21559), .X(n21504) );
  nand_x1_sg U61521 ( .A(n55301), .B(n21560), .X(n21559) );
  nand_x4_sg U61522 ( .A(n14527), .B(n14579), .X(n14524) );
  nand_x1_sg U61523 ( .A(n52765), .B(n14580), .X(n14579) );
  nand_x4_sg U61524 ( .A(n17648), .B(n17700), .X(n17645) );
  nand_x1_sg U61525 ( .A(n53885), .B(n17701), .X(n17700) );
  nand_x4_sg U61526 ( .A(n19193), .B(n19245), .X(n19190) );
  nand_x1_sg U61527 ( .A(n54450), .B(n19246), .X(n19245) );
  nand_x4_sg U61528 ( .A(n20737), .B(n20789), .X(n20734) );
  nand_x1_sg U61529 ( .A(n55018), .B(n20790), .X(n20789) );
  nand_x4_sg U61530 ( .A(n12194), .B(n12248), .X(n12191) );
  nand_x1_sg U61531 ( .A(n51939), .B(n12249), .X(n12248) );
  nand_x4_sg U61532 ( .A(n53820), .B(n17320), .X(n17317) );
  nand_x4_sg U61533 ( .A(n54385), .B(n18865), .X(n18862) );
  nand_x4_sg U61534 ( .A(n54953), .B(n20409), .X(n20406) );
  nand_x4_sg U61535 ( .A(n10532), .B(n10533), .X(n10525) );
  nor_x1_sg U61536 ( .A(n51340), .B(n10536), .X(n10534) );
  nand_x4_sg U61537 ( .A(n17544), .B(n17545), .X(n17537) );
  nor_x1_sg U61538 ( .A(n53850), .B(n17548), .X(n17546) );
  nand_x4_sg U61539 ( .A(n19089), .B(n19090), .X(n19082) );
  nor_x1_sg U61540 ( .A(n54415), .B(n19093), .X(n19091) );
  nand_x4_sg U61541 ( .A(n20633), .B(n20634), .X(n20626) );
  nor_x1_sg U61542 ( .A(n54983), .B(n20637), .X(n20635) );
  nand_x4_sg U61543 ( .A(n13926), .B(n13927), .X(n13873) );
  nand_x1_sg U61544 ( .A(n52474), .B(n13923), .X(n13927) );
  nand_x1_sg U61545 ( .A(n52450), .B(n13922), .X(n13926) );
  nand_x4_sg U61546 ( .A(n18314), .B(n18315), .X(n18307) );
  nor_x1_sg U61547 ( .A(n54131), .B(n18318), .X(n18316) );
  nand_x4_sg U61548 ( .A(n11759), .B(n11719), .X(n11664) );
  nand_x4_sg U61549 ( .A(n10774), .B(n10720), .X(n10768) );
  nand_x4_sg U61550 ( .A(n14871), .B(n14831), .X(n14776) );
  nand_x4_sg U61551 ( .A(n53961), .B(n17736), .X(n17733) );
  nand_x4_sg U61552 ( .A(n54526), .B(n19281), .X(n19278) );
  nand_x4_sg U61553 ( .A(n55094), .B(n20825), .X(n20822) );
  nand_x4_sg U61554 ( .A(n10386), .B(n10306), .X(n10312) );
  nand_x4_sg U61555 ( .A(n14278), .B(n14198), .X(n14204) );
  nand_x4_sg U61556 ( .A(n18168), .B(n18089), .X(n18095) );
  nand_x4_sg U61557 ( .A(n19713), .B(n19634), .X(n19640) );
  nand_x4_sg U61558 ( .A(n21258), .B(n21179), .X(n21185) );
  nand_x4_sg U61559 ( .A(n18862), .B(n18863), .X(n9212) );
  nand_x4_sg U61560 ( .A(n20406), .B(n20407), .X(n9136) );
  nand_x4_sg U61561 ( .A(n17317), .B(n17318), .X(n9250) );
  nand_x4_sg U61562 ( .A(n52560), .B(n13845), .X(n13842) );
  nand_x4_sg U61563 ( .A(n10726), .B(n10725), .X(n10718) );
  nand_x4_sg U61564 ( .A(n14618), .B(n14617), .X(n14610) );
  nand_x4_sg U61565 ( .A(n17739), .B(n17738), .X(n17731) );
  nand_x4_sg U61566 ( .A(n18508), .B(n18507), .X(n18500) );
  nand_x4_sg U61567 ( .A(n19284), .B(n19283), .X(n19276) );
  nand_x4_sg U61568 ( .A(n20053), .B(n20052), .X(n20045) );
  nand_x4_sg U61569 ( .A(n20828), .B(n20827), .X(n20820) );
  nand_x4_sg U61570 ( .A(n21598), .B(n21597), .X(n21590) );
  nand_x4_sg U61571 ( .A(n11336), .B(n11337), .X(n11334) );
  nand_x4_sg U61572 ( .A(n12897), .B(n12898), .X(n12895) );
  nand_x4_sg U61573 ( .A(n13677), .B(n13678), .X(n13675) );
  nand_x4_sg U61574 ( .A(n15230), .B(n15231), .X(n15228) );
  nand_x4_sg U61575 ( .A(n16796), .B(n16797), .X(n16794) );
  nand_x1_sg U61576 ( .A(n10598), .B(n51385), .X(n10597) );
  nor_x1_sg U61577 ( .A(n10599), .B(n51380), .X(n10598) );
  nand_x1_sg U61578 ( .A(n17611), .B(n53892), .X(n17610) );
  nor_x1_sg U61579 ( .A(n17612), .B(n53886), .X(n17611) );
  nand_x1_sg U61580 ( .A(n19156), .B(n54457), .X(n19155) );
  nor_x1_sg U61581 ( .A(n19157), .B(n54451), .X(n19156) );
  nand_x1_sg U61582 ( .A(n20700), .B(n55025), .X(n20699) );
  nor_x1_sg U61583 ( .A(n20701), .B(n55019), .X(n20700) );
  nand_x4_sg U61584 ( .A(n10535), .B(n10571), .X(n10532) );
  nand_x4_sg U61585 ( .A(n19862), .B(n19898), .X(n19859) );
  nand_x1_sg U61586 ( .A(n54641), .B(n54653), .X(n19899) );
  nand_x4_sg U61587 ( .A(n21407), .B(n21443), .X(n21404) );
  nand_x1_sg U61588 ( .A(n55209), .B(n55221), .X(n21444) );
  nand_x4_sg U61589 ( .A(n17547), .B(n17583), .X(n17544) );
  nand_x4_sg U61590 ( .A(n19092), .B(n19128), .X(n19089) );
  nand_x4_sg U61591 ( .A(n20636), .B(n20672), .X(n20633) );
  nand_x4_sg U61592 ( .A(n14427), .B(n14463), .X(n14424) );
  nand_x1_sg U61593 ( .A(n52677), .B(n52689), .X(n14464) );
  nand_x4_sg U61594 ( .A(n18317), .B(n18353), .X(n18314) );
  nand_x1_sg U61595 ( .A(n18321), .B(n18354), .X(n18353) );
  nand_x4_sg U61596 ( .A(n11507), .B(n11506), .X(n11499) );
  nand_x4_sg U61597 ( .A(n12287), .B(n12286), .X(n12279) );
  nand_x4_sg U61598 ( .A(n13068), .B(n13067), .X(n13060) );
  nand_x4_sg U61599 ( .A(n15401), .B(n15400), .X(n15393) );
  nand_x4_sg U61600 ( .A(n16182), .B(n16181), .X(n16174) );
  nand_x4_sg U61601 ( .A(n16967), .B(n16966), .X(n16959) );
  nand_x4_sg U61602 ( .A(n11591), .B(n51727), .X(n11578) );
  nor_x1_sg U61603 ( .A(n11593), .B(n11594), .X(n11592) );
  nand_x4_sg U61604 ( .A(n12372), .B(n52005), .X(n12359) );
  nor_x1_sg U61605 ( .A(n12374), .B(n12375), .X(n12373) );
  nand_x4_sg U61606 ( .A(n13152), .B(n52283), .X(n13139) );
  nor_x1_sg U61607 ( .A(n13154), .B(n13155), .X(n13153) );
  nand_x4_sg U61608 ( .A(n13932), .B(n52558), .X(n13919) );
  nor_x1_sg U61609 ( .A(n13934), .B(n13935), .X(n13933) );
  nand_x4_sg U61610 ( .A(n15485), .B(n53117), .X(n15472) );
  nor_x1_sg U61611 ( .A(n15487), .B(n15488), .X(n15486) );
  nand_x4_sg U61612 ( .A(n17051), .B(n53675), .X(n17038) );
  nor_x1_sg U61613 ( .A(n17053), .B(n17054), .X(n17052) );
  nand_x4_sg U61614 ( .A(n11405), .B(n11406), .X(n11403) );
  nand_x4_sg U61615 ( .A(n12185), .B(n12186), .X(n12183) );
  nand_x4_sg U61616 ( .A(n12966), .B(n12967), .X(n12964) );
  nand_x4_sg U61617 ( .A(n15299), .B(n15300), .X(n15297) );
  nand_x4_sg U61618 ( .A(n16080), .B(n16081), .X(n16078) );
  nand_x4_sg U61619 ( .A(n16865), .B(n16866), .X(n16863) );
  nand_x4_sg U61620 ( .A(n18591), .B(n54241), .X(n18577) );
  nor_x1_sg U61621 ( .A(n18593), .B(n18594), .X(n18592) );
  nand_x4_sg U61622 ( .A(n19893), .B(n19894), .X(n19888) );
  nand_x4_sg U61623 ( .A(n21438), .B(n21439), .X(n21433) );
  nand_x4_sg U61624 ( .A(n18461), .B(n18460), .X(n18458) );
  nand_x4_sg U61625 ( .A(n13355), .B(n13356), .X(n13318) );
  nand_x1_sg U61626 ( .A(n52323), .B(n40533), .X(n13356) );
  nand_x4_sg U61627 ( .A(n14135), .B(n14136), .X(n14098) );
  nand_x1_sg U61628 ( .A(n52598), .B(n40534), .X(n14136) );
  nand_x4_sg U61629 ( .A(n15688), .B(n15689), .X(n15651) );
  nand_x1_sg U61630 ( .A(n53157), .B(n40535), .X(n15689) );
  nand_x4_sg U61631 ( .A(n17254), .B(n17255), .X(n17217) );
  nand_x1_sg U61632 ( .A(n53715), .B(n40536), .X(n17255) );
  nand_x4_sg U61633 ( .A(n10718), .B(n51469), .X(n10712) );
  nor_x1_sg U61634 ( .A(n10725), .B(n10726), .X(n10724) );
  nand_x4_sg U61635 ( .A(n14610), .B(n52858), .X(n14604) );
  nor_x1_sg U61636 ( .A(n14617), .B(n14618), .X(n14616) );
  nand_x4_sg U61637 ( .A(n17731), .B(n53978), .X(n17725) );
  nor_x1_sg U61638 ( .A(n17738), .B(n17739), .X(n17737) );
  nand_x4_sg U61639 ( .A(n18500), .B(n54262), .X(n18494) );
  nor_x1_sg U61640 ( .A(n18507), .B(n18508), .X(n18506) );
  nand_x4_sg U61641 ( .A(n19276), .B(n54543), .X(n19270) );
  nor_x1_sg U61642 ( .A(n19283), .B(n19284), .X(n19282) );
  nand_x4_sg U61643 ( .A(n20045), .B(n54829), .X(n20039) );
  nor_x1_sg U61644 ( .A(n20052), .B(n20053), .X(n20051) );
  nand_x4_sg U61645 ( .A(n20820), .B(n55111), .X(n20814) );
  nor_x1_sg U61646 ( .A(n20827), .B(n20828), .X(n20826) );
  nand_x4_sg U61647 ( .A(n21590), .B(n55397), .X(n21584) );
  nor_x1_sg U61648 ( .A(n21597), .B(n21598), .X(n21596) );
  nand_x4_sg U61649 ( .A(n13411), .B(n13500), .X(n13418) );
  nand_x4_sg U61650 ( .A(n13805), .B(n13804), .X(n13797) );
  nand_x4_sg U61651 ( .A(n11499), .B(n51749), .X(n11493) );
  nor_x1_sg U61652 ( .A(n11506), .B(n11507), .X(n11505) );
  nand_x4_sg U61653 ( .A(n12279), .B(n52032), .X(n12273) );
  nor_x1_sg U61654 ( .A(n12286), .B(n12287), .X(n12285) );
  nand_x4_sg U61655 ( .A(n13060), .B(n52307), .X(n13054) );
  nor_x1_sg U61656 ( .A(n13067), .B(n13068), .X(n13066) );
  nand_x4_sg U61657 ( .A(n15393), .B(n53141), .X(n15387) );
  nor_x1_sg U61658 ( .A(n15400), .B(n15401), .X(n15399) );
  nand_x4_sg U61659 ( .A(n16174), .B(n53418), .X(n16168) );
  nor_x1_sg U61660 ( .A(n16181), .B(n16182), .X(n16180) );
  nand_x4_sg U61661 ( .A(n16959), .B(n53699), .X(n16953) );
  nor_x1_sg U61662 ( .A(n16966), .B(n16967), .X(n16965) );
  nand_x4_sg U61663 ( .A(n11578), .B(n11583), .X(n11556) );
  nand_x4_sg U61664 ( .A(n13139), .B(n13144), .X(n13117) );
  nand_x4_sg U61665 ( .A(n15472), .B(n15477), .X(n15450) );
  nand_x4_sg U61666 ( .A(n17038), .B(n17043), .X(n17016) );
  nand_x4_sg U61667 ( .A(n14458), .B(n14459), .X(n14453) );
  nand_x4_sg U61668 ( .A(n18577), .B(n18581), .X(n18555) );
  nand_x1_sg U61669 ( .A(n54127), .B(n18583), .X(n18582) );
  nand_x4_sg U61670 ( .A(n18348), .B(n18349), .X(n18343) );
  nand_x4_sg U61671 ( .A(n12244), .B(n12243), .X(n12236) );
  nand_x4_sg U61672 ( .A(n10679), .B(n10678), .X(n10676) );
  nand_x4_sg U61673 ( .A(n20006), .B(n20005), .X(n20003) );
  nand_x4_sg U61674 ( .A(n21551), .B(n21550), .X(n21548) );
  nand_x1_sg U61675 ( .A(n54054), .B(n18076), .X(n18075) );
  nand_x1_sg U61676 ( .A(n54051), .B(n18077), .X(n18074) );
  nand_x4_sg U61677 ( .A(n14571), .B(n14570), .X(n14568) );
  nand_x4_sg U61678 ( .A(n17692), .B(n17691), .X(n17689) );
  nand_x4_sg U61679 ( .A(n19237), .B(n19236), .X(n19234) );
  nand_x4_sg U61680 ( .A(n20781), .B(n20780), .X(n20778) );
  nand_x4_sg U61681 ( .A(n16139), .B(n16138), .X(n16131) );
  nand_x4_sg U61682 ( .A(n18421), .B(n18423), .X(n18377) );
  nand_x1_sg U61683 ( .A(n18424), .B(n18425), .X(n18423) );
  nor_x1_sg U61684 ( .A(n54177), .B(n18426), .X(n18424) );
  nand_x4_sg U61685 ( .A(n10639), .B(n10641), .X(n10595) );
  nand_x1_sg U61686 ( .A(n10642), .B(n10643), .X(n10641) );
  nor_x1_sg U61687 ( .A(n51389), .B(n10644), .X(n10642) );
  nand_x4_sg U61688 ( .A(n19966), .B(n19968), .X(n19922) );
  nand_x1_sg U61689 ( .A(n19969), .B(n19970), .X(n19968) );
  nor_x1_sg U61690 ( .A(n54744), .B(n19971), .X(n19969) );
  nand_x4_sg U61691 ( .A(n21511), .B(n21513), .X(n21467) );
  nand_x1_sg U61692 ( .A(n21514), .B(n21515), .X(n21513) );
  nor_x1_sg U61693 ( .A(n55312), .B(n21516), .X(n21514) );
  nand_x1_sg U61694 ( .A(n20122), .B(n20123), .X(n20121) );
  nor_x1_sg U61695 ( .A(n54777), .B(n20124), .X(n20122) );
  nand_x1_sg U61696 ( .A(n21667), .B(n21668), .X(n21666) );
  nor_x1_sg U61697 ( .A(n55345), .B(n21669), .X(n21667) );
  nand_x1_sg U61698 ( .A(n13543), .B(n13544), .X(n13542) );
  nor_x1_sg U61699 ( .A(n52408), .B(n13545), .X(n13543) );
  nand_x1_sg U61700 ( .A(n16253), .B(n16254), .X(n16252) );
  nor_x1_sg U61701 ( .A(n53379), .B(n16255), .X(n16253) );
  nand_x1_sg U61702 ( .A(n14688), .B(n14689), .X(n14687) );
  nor_x1_sg U61703 ( .A(n52807), .B(n14690), .X(n14688) );
  nand_x4_sg U61704 ( .A(n11152), .B(n11078), .X(n11085) );
  nand_x1_sg U61705 ( .A(n51602), .B(n11225), .X(n11152) );
  nand_x4_sg U61706 ( .A(n13497), .B(n13423), .X(n13430) );
  nand_x1_sg U61707 ( .A(n52434), .B(n13563), .X(n13497) );
  nand_x4_sg U61708 ( .A(n15830), .B(n15756), .X(n15763) );
  nand_x1_sg U61709 ( .A(n53270), .B(n15897), .X(n15830) );
  nand_x4_sg U61710 ( .A(n11935), .B(n11861), .X(n11868) );
  nand_x1_sg U61711 ( .A(n51883), .B(n12002), .X(n11935) );
  nand_x4_sg U61712 ( .A(n12713), .B(n12639), .X(n12646) );
  nand_x1_sg U61713 ( .A(n52160), .B(n12786), .X(n12713) );
  nand_x4_sg U61714 ( .A(n15046), .B(n14972), .X(n14979) );
  nand_x1_sg U61715 ( .A(n52994), .B(n15119), .X(n15046) );
  nand_x4_sg U61716 ( .A(n16612), .B(n16538), .X(n16545) );
  nand_x1_sg U61717 ( .A(n53552), .B(n16685), .X(n16612) );
  nand_x4_sg U61718 ( .A(n12335), .B(n12334), .X(n12328) );
  nand_x4_sg U61719 ( .A(n11460), .B(n11459), .X(n11461) );
  nand_x4_sg U61720 ( .A(n13021), .B(n13020), .X(n13022) );
  nand_x4_sg U61721 ( .A(n15354), .B(n15353), .X(n15355) );
  nand_x4_sg U61722 ( .A(n16920), .B(n16919), .X(n16921) );
  nand_x4_sg U61723 ( .A(n12240), .B(n12239), .X(n12241) );
  nand_x4_sg U61724 ( .A(n16135), .B(n16134), .X(n16136) );
  nand_x4_sg U61725 ( .A(n11368), .B(n11374), .X(n11364) );
  nor_x1_sg U61726 ( .A(n11377), .B(n11378), .X(n11375) );
  nand_x4_sg U61727 ( .A(n12148), .B(n12154), .X(n12144) );
  nor_x1_sg U61728 ( .A(n12157), .B(n12158), .X(n12155) );
  nand_x4_sg U61729 ( .A(n12929), .B(n12935), .X(n12925) );
  nor_x1_sg U61730 ( .A(n12938), .B(n12939), .X(n12936) );
  nand_x4_sg U61731 ( .A(n15262), .B(n15268), .X(n15258) );
  nor_x1_sg U61732 ( .A(n15271), .B(n15272), .X(n15269) );
  nand_x4_sg U61733 ( .A(n16043), .B(n16049), .X(n16039) );
  nor_x1_sg U61734 ( .A(n16052), .B(n16053), .X(n16050) );
  nand_x4_sg U61735 ( .A(n16828), .B(n16834), .X(n16824) );
  nor_x1_sg U61736 ( .A(n16837), .B(n16838), .X(n16835) );
  nand_x4_sg U61737 ( .A(n17733), .B(n17734), .X(n17726) );
  nand_x4_sg U61738 ( .A(n19278), .B(n19279), .X(n19271) );
  nand_x4_sg U61739 ( .A(n20822), .B(n20823), .X(n20815) );
  nand_x4_sg U61740 ( .A(n13842), .B(n13843), .X(n13835) );
  nor_x1_sg U61741 ( .A(n51419), .B(n10798), .X(n10796) );
  nor_x1_sg U61742 ( .A(n44662), .B(n11580), .X(n11577) );
  nor_x1_sg U61743 ( .A(n44661), .B(n13141), .X(n13138) );
  nor_x1_sg U61744 ( .A(n44659), .B(n15474), .X(n15471) );
  nor_x1_sg U61745 ( .A(n44658), .B(n17040), .X(n17037) );
  nor_x1_sg U61746 ( .A(n46587), .B(n26507), .X(\L1_0/n4423 ) );
  nor_x1_sg U61747 ( .A(n18808), .B(n18776), .X(n18806) );
  nand_x1_sg U61748 ( .A(n42885), .B(n46510), .X(n8843) );
  nand_x1_sg U61749 ( .A(n44090), .B(n46419), .X(n9337) );
  nand_x1_sg U61750 ( .A(n42871), .B(n46398), .X(n9301) );
  nand_x1_sg U61751 ( .A(n44084), .B(n46263), .X(n9091) );
  nand_x1_sg U61752 ( .A(n44092), .B(n46465), .X(n9003) );
  nand_x1_sg U61753 ( .A(n41358), .B(n46375), .X(n9263) );
  nand_x1_sg U61754 ( .A(n41356), .B(n46327), .X(n9225) );
  nand_x1_sg U61755 ( .A(n42877), .B(n46442), .X(n8982) );
  nand_x1_sg U61756 ( .A(n41984), .B(n46442), .X(n8984) );
  nand_x1_sg U61757 ( .A(n42875), .B(n46442), .X(n8993) );
  nand_x1_sg U61758 ( .A(n44120), .B(n46442), .X(n8978) );
  nand_x1_sg U61759 ( .A(n44118), .B(n46442), .X(n8964) );
  nand_x1_sg U61760 ( .A(n42891), .B(n46553), .X(n8888) );
  nand_x1_sg U61761 ( .A(n44096), .B(n46531), .X(n8901) );
  nor_x1_sg U61762 ( .A(n11805), .B(n11773), .X(n11803) );
  nand_x4_sg U61763 ( .A(n51377), .B(n46569), .X(n10743) );
  nand_x4_sg U61764 ( .A(n51650), .B(n51543), .X(n11618) );
  nand_x4_sg U61765 ( .A(n51931), .B(n51826), .X(n12399) );
  nand_x4_sg U61766 ( .A(n52206), .B(n52100), .X(n13179) );
  nand_x4_sg U61767 ( .A(n52483), .B(n52378), .X(n13959) );
  nand_x4_sg U61768 ( .A(n53040), .B(n52934), .X(n15512) );
  nand_x4_sg U61769 ( .A(n53214), .B(n53319), .X(n16294) );
  nand_x4_sg U61770 ( .A(n53598), .B(n53492), .X(n17078) );
  nand_x4_sg U61771 ( .A(n46405), .B(n53298), .X(n16256) );
  nand_x4_sg U61772 ( .A(n46517), .B(n46513), .X(n12206) );
  nand_x4_sg U61773 ( .A(n51879), .B(n46513), .X(n12587) );
  nand_x4_sg U61774 ( .A(n46296), .B(n46286), .X(n19972) );
  nand_x4_sg U61775 ( .A(n46251), .B(n46241), .X(n21517) );
  nand_x4_sg U61776 ( .A(n46286), .B(n54660), .X(n20360) );
  nand_x4_sg U61777 ( .A(n46241), .B(n55228), .X(n21905) );
  nor_x1_sg U61778 ( .A(n51396), .B(n10696), .X(n10733) );
  nand_x4_sg U61779 ( .A(n52806), .B(n52648), .X(n14748) );
  nand_x4_sg U61780 ( .A(n53926), .B(n53765), .X(n17869) );
  nand_x4_sg U61781 ( .A(n54491), .B(n54330), .X(n19414) );
  nand_x4_sg U61782 ( .A(n55059), .B(n54898), .X(n20958) );
  nand_x2_sg U61783 ( .A(n16104), .B(n16105), .X(n16103) );
  nand_x1_sg U61784 ( .A(n16107), .B(n16108), .X(n16104) );
  nand_x1_sg U61785 ( .A(n16106), .B(n53298), .X(n16105) );
  nand_x2_sg U61786 ( .A(n14542), .B(n14543), .X(n14541) );
  nand_x1_sg U61787 ( .A(n14545), .B(n14546), .X(n14542) );
  nand_x1_sg U61788 ( .A(n14544), .B(n52742), .X(n14543) );
  nand_x2_sg U61789 ( .A(n17663), .B(n17664), .X(n17662) );
  nand_x1_sg U61790 ( .A(n17666), .B(n17667), .X(n17663) );
  nand_x1_sg U61791 ( .A(n17665), .B(n53862), .X(n17664) );
  nand_x2_sg U61792 ( .A(n19208), .B(n19209), .X(n19207) );
  nand_x1_sg U61793 ( .A(n19211), .B(n19212), .X(n19208) );
  nand_x1_sg U61794 ( .A(n19210), .B(n54427), .X(n19209) );
  nand_x2_sg U61795 ( .A(n20752), .B(n20753), .X(n20751) );
  nand_x1_sg U61796 ( .A(n20755), .B(n20756), .X(n20752) );
  nand_x1_sg U61797 ( .A(n20754), .B(n54995), .X(n20753) );
  nor_x1_sg U61798 ( .A(n13904), .B(n13900), .X(n13902) );
  nor_x1_sg U61799 ( .A(n51893), .B(n12368), .X(n12366) );
  nand_x2_sg U61800 ( .A(n10650), .B(n10651), .X(n10649) );
  nand_x1_sg U61801 ( .A(n10653), .B(n10654), .X(n10650) );
  nand_x2_sg U61802 ( .A(n18432), .B(n18433), .X(n18431) );
  nand_x1_sg U61803 ( .A(n18435), .B(n18436), .X(n18432) );
  nand_x2_sg U61804 ( .A(n19977), .B(n19978), .X(n19976) );
  nand_x1_sg U61805 ( .A(n19980), .B(n19981), .X(n19977) );
  nand_x2_sg U61806 ( .A(n21522), .B(n21523), .X(n21521) );
  nand_x1_sg U61807 ( .A(n21525), .B(n21526), .X(n21522) );
  nand_x2_sg U61808 ( .A(n12209), .B(n12210), .X(n12208) );
  nand_x1_sg U61809 ( .A(n12212), .B(n12213), .X(n12209) );
  nand_x2_sg U61810 ( .A(n13770), .B(n13771), .X(n13769) );
  nand_x1_sg U61811 ( .A(n13773), .B(n13774), .X(n13770) );
  nor_x1_sg U61812 ( .A(n51277), .B(n51288), .X(n10440) );
  nand_x2_sg U61813 ( .A(n11429), .B(n11430), .X(n11428) );
  nand_x1_sg U61814 ( .A(n11432), .B(n11433), .X(n11429) );
  nand_x2_sg U61815 ( .A(n12990), .B(n12991), .X(n12989) );
  nand_x1_sg U61816 ( .A(n12993), .B(n12994), .X(n12990) );
  nand_x2_sg U61817 ( .A(n15323), .B(n15324), .X(n15322) );
  nand_x1_sg U61818 ( .A(n15326), .B(n15327), .X(n15323) );
  nand_x2_sg U61819 ( .A(n16889), .B(n16890), .X(n16888) );
  nand_x1_sg U61820 ( .A(n16892), .B(n16893), .X(n16889) );
  nand_x4_sg U61821 ( .A(n46567), .B(n51377), .X(n10838) );
  nand_x4_sg U61822 ( .A(n52763), .B(n52655), .X(n14730) );
  nand_x4_sg U61823 ( .A(n53883), .B(n46363), .X(n17851) );
  nand_x4_sg U61824 ( .A(n54448), .B(n46316), .X(n19396) );
  nand_x4_sg U61825 ( .A(n55016), .B(n46271), .X(n20940) );
  nand_x4_sg U61826 ( .A(n52806), .B(n52655), .X(n14883) );
  nand_x4_sg U61827 ( .A(n53926), .B(n46363), .X(n18004) );
  nand_x4_sg U61828 ( .A(n54491), .B(n46316), .X(n19549) );
  nand_x4_sg U61829 ( .A(n55059), .B(n46271), .X(n21093) );
  nand_x4_sg U61830 ( .A(n52742), .B(n46450), .X(n14691) );
  nand_x4_sg U61831 ( .A(n53862), .B(n46361), .X(n17812) );
  nand_x4_sg U61832 ( .A(n54427), .B(n46314), .X(n19357) );
  nand_x4_sg U61833 ( .A(n54995), .B(n46269), .X(n20901) );
  nand_x4_sg U61834 ( .A(n14048), .B(n46484), .X(n14148) );
  nand_x4_sg U61835 ( .A(n46567), .B(n46558), .X(n10645) );
  nand_x4_sg U61836 ( .A(n51306), .B(n46558), .X(n11028) );
  nor_x1_sg U61837 ( .A(n10784), .B(n42282), .X(n10783) );
  nor_x1_sg U61838 ( .A(n14743), .B(n41259), .X(n14742) );
  nor_x1_sg U61839 ( .A(n17864), .B(n41257), .X(n17863) );
  nor_x1_sg U61840 ( .A(n19409), .B(n41255), .X(n19408) );
  nor_x1_sg U61841 ( .A(n20953), .B(n41253), .X(n20952) );
  nor_x1_sg U61842 ( .A(n10851), .B(n41239), .X(n10850) );
  nand_x2_sg U61843 ( .A(n46569), .B(n25401), .X(n25400) );
  nand_x1_sg U61844 ( .A(n53266), .B(n53298), .X(n16425) );
  nand_x1_sg U61845 ( .A(n53298), .B(n27412), .X(n27411) );
  nor_x1_sg U61846 ( .A(n46217), .B(n27403), .X(n27412) );
  nand_x4_sg U61847 ( .A(n54776), .B(n54614), .X(n20182) );
  nand_x4_sg U61848 ( .A(n55344), .B(n55182), .X(n21727) );
  nor_x1_sg U61849 ( .A(n17401), .B(n17309), .X(n17311) );
  nor_x1_sg U61850 ( .A(n18946), .B(n18854), .X(n18856) );
  nor_x1_sg U61851 ( .A(n20490), .B(n20398), .X(n20400) );
  nand_x4_sg U61852 ( .A(n54731), .B(n46296), .X(n20164) );
  nand_x4_sg U61853 ( .A(n55299), .B(n46251), .X(n21709) );
  nand_x4_sg U61854 ( .A(n46296), .B(n54776), .X(n20319) );
  nand_x4_sg U61855 ( .A(n46251), .B(n55344), .X(n21864) );
  nand_x1_sg U61856 ( .A(n46285), .B(n46286), .X(n20299) );
  nand_x1_sg U61857 ( .A(n46240), .B(n46241), .X(n21844) );
  nand_x4_sg U61858 ( .A(n46468), .B(n46474), .X(n13767) );
  nand_x4_sg U61859 ( .A(n54751), .B(n54614), .X(n20165) );
  nand_x4_sg U61860 ( .A(n55319), .B(n55182), .X(n21710) );
  nand_x1_sg U61861 ( .A(n51738), .B(n51543), .X(n11708) );
  nand_x1_sg U61862 ( .A(n52848), .B(n52655), .X(n14820) );
  nand_x1_sg U61863 ( .A(n53968), .B(n46363), .X(n17941) );
  nand_x1_sg U61864 ( .A(n54533), .B(n46316), .X(n19486) );
  nand_x1_sg U61865 ( .A(n54818), .B(n46296), .X(n20256) );
  nand_x1_sg U61866 ( .A(n55101), .B(n46271), .X(n21030) );
  nand_x1_sg U61867 ( .A(n55386), .B(n46251), .X(n21801) );
  nand_x4_sg U61868 ( .A(n52249), .B(n46500), .X(n13198) );
  nand_x4_sg U61869 ( .A(n52525), .B(n46478), .X(n13978) );
  nand_x4_sg U61870 ( .A(n53083), .B(n46432), .X(n15531) );
  nand_x4_sg U61871 ( .A(n53641), .B(n46388), .X(n17097) );
  nand_x1_sg U61872 ( .A(n52742), .B(n26853), .X(n26852) );
  nor_x1_sg U61873 ( .A(n46221), .B(n26844), .X(n26853) );
  nand_x1_sg U61874 ( .A(n53862), .B(n27972), .X(n27971) );
  nor_x1_sg U61875 ( .A(n46213), .B(n27963), .X(n27972) );
  nand_x1_sg U61876 ( .A(n54427), .B(n28530), .X(n28529) );
  nor_x1_sg U61877 ( .A(n46209), .B(n28521), .X(n28530) );
  nand_x1_sg U61878 ( .A(n54995), .B(n29089), .X(n29088) );
  nor_x1_sg U61879 ( .A(n46205), .B(n29080), .X(n29089) );
  nor_x1_sg U61880 ( .A(n12542), .B(n52019), .X(n12541) );
  nor_x1_sg U61881 ( .A(n13323), .B(n52295), .X(n13322) );
  nor_x1_sg U61882 ( .A(n14103), .B(n52570), .X(n14102) );
  nor_x1_sg U61883 ( .A(n15656), .B(n53129), .X(n15655) );
  nor_x1_sg U61884 ( .A(n17222), .B(n53687), .X(n17221) );
  nand_x1_sg U61885 ( .A(n12487), .B(n51826), .X(n12488) );
  nand_x1_sg U61886 ( .A(n13268), .B(n52100), .X(n13269) );
  nand_x1_sg U61887 ( .A(n14048), .B(n52378), .X(n14049) );
  nand_x1_sg U61888 ( .A(n15601), .B(n52934), .X(n15602) );
  nand_x1_sg U61889 ( .A(n17167), .B(n53492), .X(n17168) );
  nand_x1_sg U61890 ( .A(n46557), .B(n46558), .X(n10967) );
  nand_x1_sg U61891 ( .A(n51435), .B(n25487), .X(n25486) );
  nor_x1_sg U61892 ( .A(n46231), .B(n25478), .X(n25487) );
  nand_x1_sg U61893 ( .A(n54229), .B(n28280), .X(n28279) );
  nor_x1_sg U61894 ( .A(n46211), .B(n28271), .X(n28280) );
  nor_x1_sg U61895 ( .A(n12915), .B(n46489), .X(n13325) );
  nor_x1_sg U61896 ( .A(n15248), .B(n46421), .X(n15658) );
  nor_x1_sg U61897 ( .A(n16814), .B(n46377), .X(n17224) );
  nor_x1_sg U61898 ( .A(n46367), .B(n53814), .X(n17560) );
  nor_x1_sg U61899 ( .A(n46320), .B(n54379), .X(n19105) );
  nor_x1_sg U61900 ( .A(n46275), .B(n54947), .X(n20649) );
  nand_x4_sg U61901 ( .A(n54184), .B(n46345), .X(n18619) );
  nor_x1_sg U61902 ( .A(n41147), .B(n41215), .X(n10505) );
  nor_x1_sg U61903 ( .A(n41518), .B(n42695), .X(n19832) );
  nor_x1_sg U61904 ( .A(n41514), .B(n42691), .X(n21377) );
  nor_x1_sg U61905 ( .A(n41189), .B(n42701), .X(n14396) );
  nor_x1_sg U61906 ( .A(n41149), .B(n41905), .X(n18287) );
  nand_x1_sg U61907 ( .A(n18333), .B(n18334), .X(n18332) );
  nand_x1_sg U61908 ( .A(n10551), .B(n10552), .X(n10550) );
  nand_x1_sg U61909 ( .A(n14292), .B(n14293), .X(n14291) );
  nor_x1_sg U61910 ( .A(n41598), .B(n19727), .X(n19725) );
  nand_x1_sg U61911 ( .A(n19727), .B(n41598), .X(n19726) );
  nand_x1_sg U61912 ( .A(n21272), .B(n21273), .X(n21271) );
  nor_x1_sg U61913 ( .A(n41602), .B(n11950), .X(n11948) );
  nand_x1_sg U61914 ( .A(n11950), .B(n41602), .X(n11949) );
  nand_x1_sg U61915 ( .A(n10400), .B(n10401), .X(n10399) );
  nor_x1_sg U61916 ( .A(n41596), .B(n15845), .X(n15843) );
  nand_x1_sg U61917 ( .A(n15845), .B(n41596), .X(n15844) );
  nand_x1_sg U61918 ( .A(n19878), .B(n19879), .X(n19877) );
  nand_x1_sg U61919 ( .A(n21423), .B(n21424), .X(n21422) );
  nand_x4_sg U61920 ( .A(n51280), .B(n51334), .X(n10799) );
  nor_x1_sg U61921 ( .A(n19781), .B(n42286), .X(n19780) );
  nor_x1_sg U61922 ( .A(n21326), .B(n42284), .X(n21325) );
  nor_x1_sg U61923 ( .A(n53452), .B(n43172), .X(n16332) );
  nor_x1_sg U61924 ( .A(n52064), .B(n40526), .X(n12438) );
  nor_x1_sg U61925 ( .A(n52341), .B(n40527), .X(n13219) );
  nor_x1_sg U61926 ( .A(n52616), .B(n40528), .X(n13999) );
  nor_x1_sg U61927 ( .A(n53175), .B(n40529), .X(n15552) );
  nor_x1_sg U61928 ( .A(n53733), .B(n40530), .X(n17118) );
  nand_x4_sg U61929 ( .A(n51598), .B(n51543), .X(n11425) );
  nand_x4_sg U61930 ( .A(n52156), .B(n52100), .X(n12986) );
  nand_x4_sg U61931 ( .A(n52990), .B(n52934), .X(n15319) );
  nand_x4_sg U61932 ( .A(n53548), .B(n53492), .X(n16885) );
  nand_x4_sg U61933 ( .A(n53253), .B(n53282), .X(n16452) );
  nor_x1_sg U61934 ( .A(n41584), .B(n10891), .X(n10889) );
  nand_x1_sg U61935 ( .A(n10891), .B(n41584), .X(n10890) );
  nor_x1_sg U61936 ( .A(n41582), .B(n16346), .X(n16344) );
  nand_x1_sg U61937 ( .A(n16346), .B(n41582), .X(n16345) );
  nand_x4_sg U61938 ( .A(n54660), .B(n54647), .X(n20103) );
  nand_x4_sg U61939 ( .A(n55228), .B(n55215), .X(n21648) );
  nand_x4_sg U61940 ( .A(n51839), .B(n51819), .X(n12016) );
  nand_x4_sg U61941 ( .A(n53227), .B(n53207), .X(n15911) );
  nand_x4_sg U61942 ( .A(n54688), .B(n54660), .X(n20326) );
  nand_x4_sg U61943 ( .A(n55256), .B(n55228), .X(n21871) );
  nand_x1_sg U61944 ( .A(n51995), .B(n26043), .X(n26042) );
  nor_x1_sg U61945 ( .A(n46227), .B(n26034), .X(n26043) );
  nand_x1_sg U61946 ( .A(n52271), .B(n26324), .X(n26323) );
  nor_x1_sg U61947 ( .A(n46225), .B(n26315), .X(n26324) );
  nand_x1_sg U61948 ( .A(n52546), .B(n26603), .X(n26602) );
  nor_x1_sg U61949 ( .A(n46223), .B(n26594), .X(n26603) );
  nand_x1_sg U61950 ( .A(n53105), .B(n27160), .X(n27159) );
  nor_x1_sg U61951 ( .A(n46219), .B(n27151), .X(n27160) );
  nand_x1_sg U61952 ( .A(n53663), .B(n27720), .X(n27719) );
  nor_x1_sg U61953 ( .A(n46215), .B(n27711), .X(n27720) );
  nand_x1_sg U61954 ( .A(n54751), .B(n28824), .X(n28823) );
  nor_x1_sg U61955 ( .A(n46207), .B(n28815), .X(n28824) );
  nand_x1_sg U61956 ( .A(n55319), .B(n29385), .X(n29384) );
  nor_x1_sg U61957 ( .A(n46203), .B(n29376), .X(n29385) );
  nor_x1_sg U61958 ( .A(n53446), .B(n53424), .X(n16500) );
  nor_x1_sg U61959 ( .A(n12462), .B(n12601), .X(n12599) );
  nor_x1_sg U61960 ( .A(n52057), .B(n41158), .X(n12600) );
  nor_x1_sg U61961 ( .A(n13243), .B(n13383), .X(n13381) );
  nor_x1_sg U61962 ( .A(n52334), .B(n41157), .X(n13382) );
  nor_x1_sg U61963 ( .A(n14023), .B(n14163), .X(n14161) );
  nor_x1_sg U61964 ( .A(n52609), .B(n41156), .X(n14162) );
  nor_x1_sg U61965 ( .A(n15576), .B(n15716), .X(n15714) );
  nor_x1_sg U61966 ( .A(n53168), .B(n41155), .X(n15715) );
  nor_x1_sg U61967 ( .A(n17142), .B(n17282), .X(n17280) );
  nor_x1_sg U61968 ( .A(n53726), .B(n41154), .X(n17281) );
  nand_x1_sg U61969 ( .A(n13625), .B(n13624), .X(n13626) );
  nand_x1_sg U61970 ( .A(n51717), .B(n25765), .X(n25764) );
  nor_x1_sg U61971 ( .A(n46229), .B(n25756), .X(n25765) );
  nand_x1_sg U61972 ( .A(n53384), .B(n27440), .X(n27439) );
  nor_x1_sg U61973 ( .A(n46217), .B(n27431), .X(n27440) );
  nand_x1_sg U61974 ( .A(n12342), .B(n12339), .X(n12343) );
  nand_x4_sg U61975 ( .A(n54124), .B(n54109), .X(n18656) );
  nand_x4_sg U61976 ( .A(n53266), .B(n53282), .X(n16330) );
  nand_x4_sg U61977 ( .A(n52447), .B(n52430), .X(n13996) );
  nand_x1_sg U61978 ( .A(n10780), .B(n10777), .X(n10781) );
  nand_x1_sg U61979 ( .A(n16237), .B(n16234), .X(n16238) );
  nand_x2_sg U61980 ( .A(n13591), .B(n13585), .X(n13590) );
  nand_x1_sg U61981 ( .A(n20106), .B(n20103), .X(n20107) );
  nand_x1_sg U61982 ( .A(n21651), .B(n21648), .X(n21652) );
  nand_x2_sg U61983 ( .A(n10964), .B(n10965), .X(n10963) );
  nand_x1_sg U61984 ( .A(n51491), .B(n10967), .X(n10964) );
  nand_x1_sg U61985 ( .A(n14672), .B(n14669), .X(n14673) );
  nand_x1_sg U61986 ( .A(n17793), .B(n17790), .X(n17794) );
  nand_x1_sg U61987 ( .A(n19338), .B(n19335), .X(n19339) );
  nand_x1_sg U61988 ( .A(n20882), .B(n20879), .X(n20883) );
  nand_x2_sg U61989 ( .A(n19801), .B(n19799), .X(n19800) );
  nand_x2_sg U61990 ( .A(n21346), .B(n21344), .X(n21345) );
  nand_x2_sg U61991 ( .A(n14366), .B(n14364), .X(n14365) );
  nand_x2_sg U61992 ( .A(n10474), .B(n10472), .X(n10473) );
  nand_x1_sg U61993 ( .A(n12304), .B(n12488), .X(n12484) );
  nand_x1_sg U61994 ( .A(n12486), .B(n12487), .X(n12485) );
  nand_x1_sg U61995 ( .A(n13085), .B(n13269), .X(n13265) );
  nand_x1_sg U61996 ( .A(n13267), .B(n13268), .X(n13266) );
  nand_x1_sg U61997 ( .A(n13865), .B(n14049), .X(n14045) );
  nand_x1_sg U61998 ( .A(n14047), .B(n14048), .X(n14046) );
  nand_x1_sg U61999 ( .A(n15418), .B(n15602), .X(n15598) );
  nand_x1_sg U62000 ( .A(n15600), .B(n15601), .X(n15599) );
  nand_x1_sg U62001 ( .A(n16984), .B(n17168), .X(n17164) );
  nand_x1_sg U62002 ( .A(n17166), .B(n17167), .X(n17165) );
  nand_x1_sg U62003 ( .A(n14841), .B(n14840), .X(n14835) );
  nand_x1_sg U62004 ( .A(n14837), .B(n52806), .X(n14836) );
  nand_x1_sg U62005 ( .A(n18731), .B(n18730), .X(n18725) );
  nand_x1_sg U62006 ( .A(n18727), .B(n54209), .X(n18726) );
  nor_x1_sg U62007 ( .A(n18770), .B(n18805), .X(n18803) );
  nand_x1_sg U62008 ( .A(n18805), .B(n18770), .X(n18804) );
  nand_x4_sg U62009 ( .A(n52447), .B(n46484), .X(n13686) );
  nand_x1_sg U62010 ( .A(n13290), .B(n13289), .X(n13284) );
  nand_x1_sg U62011 ( .A(n13286), .B(n52249), .X(n13285) );
  nand_x1_sg U62012 ( .A(n14070), .B(n14069), .X(n14064) );
  nand_x1_sg U62013 ( .A(n14066), .B(n52525), .X(n14065) );
  nand_x1_sg U62014 ( .A(n15623), .B(n15622), .X(n15617) );
  nand_x1_sg U62015 ( .A(n15619), .B(n53083), .X(n15618) );
  nand_x1_sg U62016 ( .A(n17189), .B(n17188), .X(n17183) );
  nand_x1_sg U62017 ( .A(n17185), .B(n53641), .X(n17184) );
  nand_x2_sg U62018 ( .A(n19936), .B(n19937), .X(n19935) );
  nand_x1_sg U62019 ( .A(n19879), .B(n54712), .X(n19937) );
  nand_x1_sg U62020 ( .A(n54710), .B(n19940), .X(n19936) );
  nand_x2_sg U62021 ( .A(n21481), .B(n21482), .X(n21480) );
  nand_x1_sg U62022 ( .A(n21424), .B(n55280), .X(n21482) );
  nand_x1_sg U62023 ( .A(n55278), .B(n21485), .X(n21481) );
  nand_x2_sg U62024 ( .A(n19809), .B(n19837), .X(n19836) );
  nand_x1_sg U62025 ( .A(n19838), .B(n19805), .X(n19837) );
  nand_x2_sg U62026 ( .A(n21354), .B(n21382), .X(n21381) );
  nand_x1_sg U62027 ( .A(n21383), .B(n21350), .X(n21382) );
  nand_x2_sg U62028 ( .A(n10609), .B(n10610), .X(n10608) );
  nand_x1_sg U62029 ( .A(n51356), .B(n10613), .X(n10609) );
  nand_x1_sg U62030 ( .A(n10552), .B(n51358), .X(n10610) );
  nand_x2_sg U62031 ( .A(n14501), .B(n14502), .X(n14500) );
  nand_x1_sg U62032 ( .A(n52708), .B(n14443), .X(n14502) );
  nand_x1_sg U62033 ( .A(n14506), .B(n14504), .X(n14501) );
  nand_x1_sg U62034 ( .A(n20277), .B(n20276), .X(n20271) );
  nand_x1_sg U62035 ( .A(n21822), .B(n21821), .X(n21816) );
  nand_x2_sg U62036 ( .A(n11705), .B(n11706), .X(n11704) );
  nand_x1_sg U62037 ( .A(n11524), .B(n11708), .X(n11705) );
  nand_x1_sg U62038 ( .A(n11707), .B(n51738), .X(n11706) );
  nand_x2_sg U62039 ( .A(n14817), .B(n14818), .X(n14816) );
  nand_x1_sg U62040 ( .A(n14636), .B(n14820), .X(n14817) );
  nand_x1_sg U62041 ( .A(n14819), .B(n52848), .X(n14818) );
  nand_x2_sg U62042 ( .A(n17938), .B(n17939), .X(n17937) );
  nand_x1_sg U62043 ( .A(n17757), .B(n17941), .X(n17938) );
  nand_x1_sg U62044 ( .A(n17940), .B(n53968), .X(n17939) );
  nand_x2_sg U62045 ( .A(n18707), .B(n18708), .X(n18706) );
  nand_x1_sg U62046 ( .A(n18525), .B(n18710), .X(n18707) );
  nand_x1_sg U62047 ( .A(n18709), .B(n54250), .X(n18708) );
  nand_x2_sg U62048 ( .A(n19483), .B(n19484), .X(n19482) );
  nand_x1_sg U62049 ( .A(n19302), .B(n19486), .X(n19483) );
  nand_x1_sg U62050 ( .A(n19485), .B(n54533), .X(n19484) );
  nand_x2_sg U62051 ( .A(n20253), .B(n20254), .X(n20252) );
  nand_x1_sg U62052 ( .A(n20070), .B(n20256), .X(n20253) );
  nand_x1_sg U62053 ( .A(n20255), .B(n54818), .X(n20254) );
  nand_x2_sg U62054 ( .A(n21027), .B(n21028), .X(n21026) );
  nand_x1_sg U62055 ( .A(n20846), .B(n21030), .X(n21027) );
  nand_x1_sg U62056 ( .A(n21029), .B(n55101), .X(n21028) );
  nand_x2_sg U62057 ( .A(n21798), .B(n21799), .X(n21797) );
  nand_x1_sg U62058 ( .A(n21615), .B(n21801), .X(n21798) );
  nand_x1_sg U62059 ( .A(n21800), .B(n55386), .X(n21799) );
  nand_x1_sg U62060 ( .A(n11729), .B(n11728), .X(n11723) );
  nand_x1_sg U62061 ( .A(n11725), .B(n51693), .X(n11724) );
  nand_x2_sg U62062 ( .A(n17622), .B(n17623), .X(n17621) );
  nand_x1_sg U62063 ( .A(n53835), .B(n17563), .X(n17623) );
  nand_x1_sg U62064 ( .A(n17627), .B(n17625), .X(n17622) );
  nand_x2_sg U62065 ( .A(n19167), .B(n19168), .X(n19166) );
  nand_x1_sg U62066 ( .A(n54400), .B(n19108), .X(n19168) );
  nand_x1_sg U62067 ( .A(n19172), .B(n19170), .X(n19167) );
  nand_x2_sg U62068 ( .A(n20711), .B(n20712), .X(n20710) );
  nand_x1_sg U62069 ( .A(n54968), .B(n20652), .X(n20712) );
  nand_x1_sg U62070 ( .A(n20716), .B(n20714), .X(n20711) );
  nand_x2_sg U62071 ( .A(n11731), .B(n11732), .X(n11730) );
  nand_x1_sg U62072 ( .A(n43049), .B(n11734), .X(n11732) );
  nand_x1_sg U62073 ( .A(n11736), .B(n11735), .X(n11731) );
  nand_x2_sg U62074 ( .A(n12511), .B(n12512), .X(n12510) );
  nand_x1_sg U62075 ( .A(n43047), .B(n12514), .X(n12512) );
  nand_x1_sg U62076 ( .A(n12516), .B(n12515), .X(n12511) );
  nand_x2_sg U62077 ( .A(n13292), .B(n13293), .X(n13291) );
  nand_x1_sg U62078 ( .A(n43045), .B(n13295), .X(n13293) );
  nand_x1_sg U62079 ( .A(n13297), .B(n13296), .X(n13292) );
  nand_x2_sg U62080 ( .A(n14072), .B(n14073), .X(n14071) );
  nand_x1_sg U62081 ( .A(n43043), .B(n14075), .X(n14073) );
  nand_x1_sg U62082 ( .A(n14077), .B(n14076), .X(n14072) );
  nand_x2_sg U62083 ( .A(n15625), .B(n15626), .X(n15624) );
  nand_x1_sg U62084 ( .A(n43041), .B(n15628), .X(n15626) );
  nand_x1_sg U62085 ( .A(n15630), .B(n15629), .X(n15625) );
  nand_x2_sg U62086 ( .A(n17191), .B(n17192), .X(n17190) );
  nand_x1_sg U62087 ( .A(n43037), .B(n17194), .X(n17192) );
  nand_x1_sg U62088 ( .A(n17196), .B(n17195), .X(n17191) );
  nand_x2_sg U62089 ( .A(n18733), .B(n18734), .X(n18732) );
  nand_x1_sg U62090 ( .A(n43943), .B(n18736), .X(n18734) );
  nand_x1_sg U62091 ( .A(n18738), .B(n18737), .X(n18733) );
  nand_x2_sg U62092 ( .A(n20279), .B(n20280), .X(n20278) );
  nand_x1_sg U62093 ( .A(n43847), .B(n20282), .X(n20280) );
  nand_x1_sg U62094 ( .A(n20284), .B(n20283), .X(n20279) );
  nand_x2_sg U62095 ( .A(n21824), .B(n21825), .X(n21823) );
  nand_x1_sg U62096 ( .A(n43845), .B(n21827), .X(n21825) );
  nand_x1_sg U62097 ( .A(n21829), .B(n21828), .X(n21824) );
  nand_x2_sg U62098 ( .A(n18391), .B(n18392), .X(n18390) );
  nand_x1_sg U62099 ( .A(n18334), .B(n54147), .X(n18392) );
  nand_x1_sg U62100 ( .A(n54145), .B(n18395), .X(n18391) );
  nand_x2_sg U62101 ( .A(n16422), .B(n16423), .X(n16421) );
  nand_x1_sg U62102 ( .A(n53440), .B(n16425), .X(n16422) );
  nand_x4_sg U62103 ( .A(n51834), .B(n11994), .X(n12012) );
  nand_x4_sg U62104 ( .A(n13555), .B(n52386), .X(n13573) );
  nand_x4_sg U62105 ( .A(n53222), .B(n15889), .X(n15907) );
  nand_x4_sg U62106 ( .A(n46285), .B(n54660), .X(n20288) );
  nand_x4_sg U62107 ( .A(n46240), .B(n55228), .X(n21833) );
  nand_x4_sg U62108 ( .A(n46557), .B(n51306), .X(n10956) );
  nand_x1_sg U62109 ( .A(n17884), .B(n17885), .X(n17883) );
  nand_x1_sg U62110 ( .A(n19429), .B(n19430), .X(n19428) );
  nand_x1_sg U62111 ( .A(n20973), .B(n20974), .X(n20972) );
  nand_x1_sg U62112 ( .A(n11651), .B(n11652), .X(n11650) );
  nand_x1_sg U62113 ( .A(n13212), .B(n13213), .X(n13211) );
  nand_x1_sg U62114 ( .A(n15545), .B(n15546), .X(n15544) );
  nand_x1_sg U62115 ( .A(n17111), .B(n17112), .X(n17110) );
  nand_x1_sg U62116 ( .A(n16326), .B(n16327), .X(n16325) );
  nand_x1_sg U62117 ( .A(n14763), .B(n14764), .X(n14762) );
  nor_x1_sg U62118 ( .A(n11611), .B(n11612), .X(n11609) );
  nand_x1_sg U62119 ( .A(n11611), .B(n11612), .X(n11610) );
  nor_x1_sg U62120 ( .A(n14723), .B(n14724), .X(n14721) );
  nand_x1_sg U62121 ( .A(n14723), .B(n14724), .X(n14722) );
  nor_x1_sg U62122 ( .A(n16287), .B(n16288), .X(n16285) );
  nand_x1_sg U62123 ( .A(n16287), .B(n16288), .X(n16286) );
  nor_x1_sg U62124 ( .A(n12392), .B(n12393), .X(n12390) );
  nand_x1_sg U62125 ( .A(n12392), .B(n12393), .X(n12391) );
  nor_x1_sg U62126 ( .A(n13172), .B(n13173), .X(n13170) );
  nand_x1_sg U62127 ( .A(n13172), .B(n13173), .X(n13171) );
  nor_x1_sg U62128 ( .A(n13952), .B(n13953), .X(n13950) );
  nand_x1_sg U62129 ( .A(n13952), .B(n13953), .X(n13951) );
  nor_x1_sg U62130 ( .A(n15505), .B(n15506), .X(n15503) );
  nand_x1_sg U62131 ( .A(n15505), .B(n15506), .X(n15504) );
  nor_x1_sg U62132 ( .A(n17071), .B(n17072), .X(n17069) );
  nand_x1_sg U62133 ( .A(n17071), .B(n17072), .X(n17070) );
  nor_x1_sg U62134 ( .A(n18653), .B(n18652), .X(n18650) );
  nand_x1_sg U62135 ( .A(n18652), .B(n18653), .X(n18651) );
  nand_x1_sg U62136 ( .A(n12431), .B(n12432), .X(n12430) );
  nor_x1_sg U62137 ( .A(n12548), .B(n12577), .X(n12575) );
  nand_x1_sg U62138 ( .A(n12577), .B(n12548), .X(n12576) );
  nor_x1_sg U62139 ( .A(n13993), .B(n13992), .X(n13990) );
  nand_x1_sg U62140 ( .A(n13992), .B(n13993), .X(n13991) );
  nand_x1_sg U62141 ( .A(n10871), .B(n10872), .X(n10870) );
  nor_x1_sg U62142 ( .A(n13329), .B(n13359), .X(n13357) );
  nand_x1_sg U62143 ( .A(n13359), .B(n13329), .X(n13358) );
  nor_x1_sg U62144 ( .A(n15662), .B(n15692), .X(n15690) );
  nand_x1_sg U62145 ( .A(n15692), .B(n15662), .X(n15691) );
  nor_x1_sg U62146 ( .A(n17228), .B(n17258), .X(n17256) );
  nand_x1_sg U62147 ( .A(n17258), .B(n17228), .X(n17257) );
  nand_x1_sg U62148 ( .A(n20198), .B(n20199), .X(n20197) );
  nand_x1_sg U62149 ( .A(n21743), .B(n21744), .X(n21742) );
  nor_x1_sg U62150 ( .A(n14109), .B(n14139), .X(n14137) );
  nand_x1_sg U62151 ( .A(n14139), .B(n14109), .X(n14138) );
  nor_x1_sg U62152 ( .A(n11776), .B(n11802), .X(n11800) );
  nand_x1_sg U62153 ( .A(n11802), .B(n11776), .X(n11801) );
  nor_x1_sg U62154 ( .A(n17844), .B(n17845), .X(n17842) );
  nand_x1_sg U62155 ( .A(n17844), .B(n17845), .X(n17843) );
  nor_x1_sg U62156 ( .A(n19389), .B(n19390), .X(n19387) );
  nand_x1_sg U62157 ( .A(n19389), .B(n19390), .X(n19388) );
  nor_x1_sg U62158 ( .A(n20933), .B(n20934), .X(n20931) );
  nand_x1_sg U62159 ( .A(n20933), .B(n20934), .X(n20932) );
  nand_x2_sg U62160 ( .A(n25474), .B(n46235), .X(n25469) );
  nand_x2_sg U62161 ( .A(n25471), .B(n25472), .X(n25470) );
  nand_x1_sg U62162 ( .A(n11784), .B(n11783), .X(n11818) );
  nand_x1_sg U62163 ( .A(n13337), .B(n13336), .X(n13375) );
  nand_x1_sg U62164 ( .A(n15670), .B(n15669), .X(n15708) );
  nand_x1_sg U62165 ( .A(n17236), .B(n17235), .X(n17274) );
  nand_x4_sg U62166 ( .A(n27942), .B(n53814), .X(n27949) );
  nand_x4_sg U62167 ( .A(n28500), .B(n54379), .X(n28507) );
  nand_x4_sg U62168 ( .A(n29059), .B(n54947), .X(n29066) );
  nand_x1_sg U62169 ( .A(n18445), .B(n18446), .X(n18444) );
  nand_x4_sg U62170 ( .A(n54688), .B(n54634), .X(n20125) );
  nand_x4_sg U62171 ( .A(n55256), .B(n55202), .X(n21670) );
  nand_x1_sg U62172 ( .A(n10663), .B(n10664), .X(n10662) );
  nand_x1_sg U62173 ( .A(n16459), .B(n16458), .X(n16493) );
  nand_x1_sg U62174 ( .A(n12556), .B(n12555), .X(n12593) );
  nand_x1_sg U62175 ( .A(n14897), .B(n14896), .X(n14930) );
  nand_x1_sg U62176 ( .A(n18018), .B(n18017), .X(n18051) );
  nand_x1_sg U62177 ( .A(n19563), .B(n19562), .X(n19596) );
  nand_x1_sg U62178 ( .A(n21107), .B(n21106), .X(n21140) );
  nand_x1_sg U62179 ( .A(n19990), .B(n19991), .X(n19989) );
  nand_x1_sg U62180 ( .A(n21535), .B(n21536), .X(n21534) );
  nand_x2_sg U62181 ( .A(n25460), .B(n46235), .X(n25454) );
  nand_x2_sg U62182 ( .A(n25456), .B(n25457), .X(n25455) );
  nand_x2_sg U62183 ( .A(n28253), .B(n46235), .X(n28247) );
  nand_x2_sg U62184 ( .A(n28249), .B(n28250), .X(n28248) );
  nand_x1_sg U62185 ( .A(n13808), .B(n13807), .X(n13820) );
  nand_x2_sg U62186 ( .A(n27952), .B(n46235), .X(n27947) );
  nand_x2_sg U62187 ( .A(n27949), .B(n27950), .X(n27948) );
  nand_x2_sg U62188 ( .A(n28510), .B(n46235), .X(n28505) );
  nand_x2_sg U62189 ( .A(n28507), .B(n28508), .X(n28506) );
  nand_x2_sg U62190 ( .A(n29069), .B(n46235), .X(n29064) );
  nand_x2_sg U62191 ( .A(n29066), .B(n29067), .X(n29065) );
  nand_x2_sg U62192 ( .A(n28811), .B(n46235), .X(n28805) );
  nand_x2_sg U62193 ( .A(n28807), .B(n28808), .X(n28806) );
  nand_x2_sg U62194 ( .A(n29372), .B(n46235), .X(n29366) );
  nand_x2_sg U62195 ( .A(n29368), .B(n29369), .X(n29367) );
  nand_x2_sg U62196 ( .A(n28231), .B(n46235), .X(n28226) );
  nand_x2_sg U62197 ( .A(n28228), .B(n28229), .X(n28227) );
  nand_x2_sg U62198 ( .A(n25717), .B(n46235), .X(n25712) );
  nand_x2_sg U62199 ( .A(n25714), .B(n25715), .X(n25713) );
  nand_x2_sg U62200 ( .A(n26276), .B(n46235), .X(n26271) );
  nand_x2_sg U62201 ( .A(n26273), .B(n26274), .X(n26272) );
  nand_x2_sg U62202 ( .A(n27112), .B(n46235), .X(n27107) );
  nand_x2_sg U62203 ( .A(n27109), .B(n27110), .X(n27108) );
  nand_x2_sg U62204 ( .A(n27672), .B(n46235), .X(n27667) );
  nand_x2_sg U62205 ( .A(n27669), .B(n27670), .X(n27668) );
  nand_x1_sg U62206 ( .A(n11221), .B(n11222), .X(n11220) );
  nand_x1_sg U62207 ( .A(n12782), .B(n12783), .X(n12781) );
  nand_x1_sg U62208 ( .A(n15115), .B(n15116), .X(n15114) );
  nand_x1_sg U62209 ( .A(n16681), .B(n16682), .X(n16680) );
  nor_x1_sg U62210 ( .A(n44421), .B(n41510), .X(n11340) );
  nor_x1_sg U62211 ( .A(n44152), .B(n41506), .X(n12120) );
  nor_x1_sg U62212 ( .A(n42813), .B(n41229), .X(n12901) );
  nor_x1_sg U62213 ( .A(n42809), .B(n41225), .X(n15234) );
  nor_x1_sg U62214 ( .A(n44419), .B(n41498), .X(n16015) );
  nor_x1_sg U62215 ( .A(n42807), .B(n41221), .X(n16800) );
  nand_x2_sg U62216 ( .A(n25442), .B(n51526), .X(n25441) );
  nand_x2_sg U62217 ( .A(n25445), .B(n46235), .X(n25440) );
  nand_x2_sg U62218 ( .A(n25721), .B(n51808), .X(n25720) );
  nand_x2_sg U62219 ( .A(n25724), .B(n46235), .X(n25719) );
  nand_x2_sg U62220 ( .A(n25999), .B(n52084), .X(n25998) );
  nand_x2_sg U62221 ( .A(n26002), .B(n46235), .X(n25997) );
  nand_x2_sg U62222 ( .A(n26280), .B(n52362), .X(n26279) );
  nand_x2_sg U62223 ( .A(n26283), .B(n46235), .X(n26278) );
  nand_x2_sg U62224 ( .A(n27116), .B(n53196), .X(n27115) );
  nand_x2_sg U62225 ( .A(n27119), .B(n46235), .X(n27114) );
  nand_x2_sg U62226 ( .A(n27396), .B(n53476), .X(n27395) );
  nand_x2_sg U62227 ( .A(n27399), .B(n46235), .X(n27394) );
  nand_x2_sg U62228 ( .A(n27676), .B(n53754), .X(n27675) );
  nand_x2_sg U62229 ( .A(n27679), .B(n46235), .X(n27674) );
  nand_x2_sg U62230 ( .A(n28235), .B(n54319), .X(n28234) );
  nand_x2_sg U62231 ( .A(n28238), .B(n46235), .X(n28233) );
  nand_x2_sg U62232 ( .A(n28793), .B(n54887), .X(n28792) );
  nand_x2_sg U62233 ( .A(n28796), .B(n46235), .X(n28791) );
  nand_x2_sg U62234 ( .A(n29354), .B(n55455), .X(n29353) );
  nand_x2_sg U62235 ( .A(n29357), .B(n46235), .X(n29352) );
  nand_x2_sg U62236 ( .A(n26559), .B(n52637), .X(n26558) );
  nand_x2_sg U62237 ( .A(n26562), .B(n46235), .X(n26557) );
  nor_x1_sg U62238 ( .A(n46546), .B(n46533), .X(n11321) );
  nor_x1_sg U62239 ( .A(n46502), .B(n46489), .X(n12882) );
  nor_x1_sg U62240 ( .A(n46434), .B(n46421), .X(n15215) );
  nor_x1_sg U62241 ( .A(n46390), .B(n46377), .X(n16781) );
  nand_x1_sg U62242 ( .A(n46567), .B(n51458), .X(n10924) );
  nand_x4_sg U62243 ( .A(n28221), .B(n54097), .X(n28228) );
  nor_x1_sg U62244 ( .A(n12752), .B(n46502), .X(n12854) );
  nor_x1_sg U62245 ( .A(n15085), .B(n46434), .X(n15187) );
  nor_x1_sg U62246 ( .A(n16651), .B(n46390), .X(n16753) );
  nor_x1_sg U62247 ( .A(n51476), .B(n10856), .X(n10984) );
  nand_x4_sg U62248 ( .A(n52391), .B(n46478), .X(n13577) );
  nand_x1_sg U62249 ( .A(n54184), .B(n28266), .X(n28265) );
  nor_x1_sg U62250 ( .A(n46211), .B(n28257), .X(n28266) );
  nor_x1_sg U62251 ( .A(n46508), .B(n12741), .X(n12827) );
  nor_x1_sg U62252 ( .A(n46440), .B(n15074), .X(n15160) );
  nor_x1_sg U62253 ( .A(n46396), .B(n16640), .X(n16726) );
  nor_x1_sg U62254 ( .A(n17421), .B(n17491), .X(n17489) );
  nor_x1_sg U62255 ( .A(n18966), .B(n19036), .X(n19034) );
  nor_x1_sg U62256 ( .A(n20510), .B(n20580), .X(n20578) );
  nand_x4_sg U62257 ( .A(n52695), .B(n46450), .X(n14538) );
  nand_x4_sg U62258 ( .A(n46443), .B(n52695), .X(n14890) );
  nand_x2_sg U62259 ( .A(n17421), .B(n53761), .X(n17420) );
  nand_x2_sg U62260 ( .A(n18966), .B(n54326), .X(n18965) );
  nand_x2_sg U62261 ( .A(n20510), .B(n54894), .X(n20509) );
  nor_x1_sg U62262 ( .A(n13530), .B(n46480), .X(n13634) );
  nor_x1_sg U62263 ( .A(n10418), .B(n46566), .X(n10514) );
  nor_x1_sg U62264 ( .A(n19745), .B(n46300), .X(n19841) );
  nor_x1_sg U62265 ( .A(n21290), .B(n46255), .X(n21386) );
  nand_x1_sg U62266 ( .A(n54794), .B(n28838), .X(n28837) );
  nor_x1_sg U62267 ( .A(n46207), .B(n28829), .X(n28838) );
  nand_x1_sg U62268 ( .A(n55362), .B(n29399), .X(n29398) );
  nor_x1_sg U62269 ( .A(n46203), .B(n29390), .X(n29399) );
  nor_x1_sg U62270 ( .A(n11969), .B(n46519), .X(n12073) );
  nand_x2_sg U62271 ( .A(n51543), .B(n25687), .X(n25686) );
  nand_x2_sg U62272 ( .A(n52100), .B(n26246), .X(n26245) );
  nand_x2_sg U62273 ( .A(n52934), .B(n27082), .X(n27081) );
  nand_x2_sg U62274 ( .A(n53492), .B(n27642), .X(n27641) );
  nand_x4_sg U62275 ( .A(n25707), .B(n46533), .X(n25714) );
  nand_x4_sg U62276 ( .A(n26266), .B(n46489), .X(n26273) );
  nand_x4_sg U62277 ( .A(n27102), .B(n46421), .X(n27109) );
  nand_x4_sg U62278 ( .A(n27662), .B(n46377), .X(n27669) );
  nand_x2_sg U62279 ( .A(n51537), .B(n25680), .X(n25679) );
  nand_x2_sg U62280 ( .A(n51819), .B(n25958), .X(n25957) );
  nand_x2_sg U62281 ( .A(n53207), .B(n27355), .X(n27354) );
  nand_x2_sg U62282 ( .A(n51826), .B(n25965), .X(n25964) );
  nand_x2_sg U62283 ( .A(n53214), .B(n27362), .X(n27361) );
  nand_x2_sg U62284 ( .A(n53765), .B(n27915), .X(n27914) );
  nand_x2_sg U62285 ( .A(n54330), .B(n28473), .X(n28472) );
  nand_x2_sg U62286 ( .A(n54898), .B(n29032), .X(n29031) );
  nand_x2_sg U62287 ( .A(n52648), .B(n26796), .X(n26795) );
  nand_x4_sg U62288 ( .A(n11217), .B(n51569), .X(n11234) );
  nand_x4_sg U62289 ( .A(n51896), .B(n51879), .X(n12435) );
  nand_x2_sg U62290 ( .A(n14076), .B(n46484), .X(n14168) );
  nand_x4_sg U62291 ( .A(n12778), .B(n52126), .X(n12795) );
  nand_x4_sg U62292 ( .A(n15111), .B(n52960), .X(n15128) );
  nand_x4_sg U62293 ( .A(n16677), .B(n53518), .X(n16694) );
  nand_x2_sg U62294 ( .A(n13392), .B(n13393), .X(n13391) );
  nand_x2_sg U62295 ( .A(n14172), .B(n13393), .X(n14171) );
  nand_x2_sg U62296 ( .A(n21926), .B(n13393), .X(n21925) );
  nand_x4_sg U62297 ( .A(n51911), .B(n51839), .X(n12561) );
  nand_x4_sg U62298 ( .A(n52463), .B(n52391), .X(n14123) );
  nand_x4_sg U62299 ( .A(n52391), .B(n46484), .X(n13538) );
  nand_x4_sg U62300 ( .A(n46517), .B(n51839), .X(n12123) );
  nand_x4_sg U62301 ( .A(n52391), .B(n46474), .X(n13684) );
  nand_x4_sg U62302 ( .A(n46405), .B(n53227), .X(n16018) );
  nor_x1_sg U62303 ( .A(n18525), .B(n46344), .X(n18709) );
  nand_x4_sg U62304 ( .A(n51598), .B(n11595), .X(n11593) );
  nand_x4_sg U62305 ( .A(n51879), .B(n12376), .X(n12374) );
  nand_x4_sg U62306 ( .A(n52156), .B(n13156), .X(n13154) );
  nand_x4_sg U62307 ( .A(n52430), .B(n13936), .X(n13934) );
  nand_x4_sg U62308 ( .A(n52990), .B(n15489), .X(n15487) );
  nand_x4_sg U62309 ( .A(n53266), .B(n16271), .X(n16268) );
  nand_x4_sg U62310 ( .A(n53548), .B(n17055), .X(n17053) );
  nand_x4_sg U62311 ( .A(n51598), .B(n46532), .X(n11655) );
  nand_x4_sg U62312 ( .A(n52156), .B(n46488), .X(n13216) );
  nand_x4_sg U62313 ( .A(n52990), .B(n46420), .X(n15549) );
  nand_x4_sg U62314 ( .A(n53548), .B(n46376), .X(n17115) );
  nand_x4_sg U62315 ( .A(n52430), .B(n46484), .X(n13637) );
  nand_x1_sg U62316 ( .A(n52783), .B(n26867), .X(n26866) );
  nor_x1_sg U62317 ( .A(n46221), .B(n26858), .X(n26867) );
  nand_x4_sg U62318 ( .A(n51630), .B(n46540), .X(n11581) );
  nand_x4_sg U62319 ( .A(n52187), .B(n46496), .X(n13142) );
  nand_x4_sg U62320 ( .A(n53021), .B(n46428), .X(n15475) );
  nand_x4_sg U62321 ( .A(n53579), .B(n46384), .X(n17041) );
  nand_x1_sg U62322 ( .A(n51952), .B(n26029), .X(n26028) );
  nor_x1_sg U62323 ( .A(n46227), .B(n26020), .X(n26029) );
  nand_x1_sg U62324 ( .A(n52227), .B(n26310), .X(n26309) );
  nor_x1_sg U62325 ( .A(n46225), .B(n26301), .X(n26310) );
  nand_x1_sg U62326 ( .A(n52504), .B(n26589), .X(n26588) );
  nor_x1_sg U62327 ( .A(n46223), .B(n26580), .X(n26589) );
  nand_x1_sg U62328 ( .A(n53061), .B(n27146), .X(n27145) );
  nor_x1_sg U62329 ( .A(n46219), .B(n27137), .X(n27146) );
  nand_x1_sg U62330 ( .A(n53619), .B(n27706), .X(n27705) );
  nor_x1_sg U62331 ( .A(n46215), .B(n27697), .X(n27706) );
  nand_x1_sg U62332 ( .A(n53903), .B(n27986), .X(n27985) );
  nor_x1_sg U62333 ( .A(n46213), .B(n27977), .X(n27986) );
  nand_x1_sg U62334 ( .A(n54468), .B(n28544), .X(n28543) );
  nor_x1_sg U62335 ( .A(n46209), .B(n28535), .X(n28544) );
  nand_x1_sg U62336 ( .A(n55036), .B(n29103), .X(n29102) );
  nor_x1_sg U62337 ( .A(n46205), .B(n29094), .X(n29103) );
  nor_x1_sg U62338 ( .A(n46416), .B(n16066), .X(n16065) );
  nor_x1_sg U62339 ( .A(n46528), .B(n12171), .X(n12170) );
  nor_x1_sg U62340 ( .A(n18571), .B(n46340), .X(n18570) );
  nand_x4_sg U62341 ( .A(n46557), .B(n51280), .X(n11006) );
  nand_x1_sg U62342 ( .A(n52824), .B(n26881), .X(n26880) );
  nor_x1_sg U62343 ( .A(n46221), .B(n26872), .X(n26881) );
  nand_x1_sg U62344 ( .A(n53944), .B(n28000), .X(n27999) );
  nor_x1_sg U62345 ( .A(n46213), .B(n27991), .X(n28000) );
  nand_x1_sg U62346 ( .A(n54509), .B(n28558), .X(n28557) );
  nor_x1_sg U62347 ( .A(n46209), .B(n28549), .X(n28558) );
  nand_x1_sg U62348 ( .A(n55077), .B(n29117), .X(n29116) );
  nor_x1_sg U62349 ( .A(n46205), .B(n29108), .X(n29117) );
  nand_x4_sg U62350 ( .A(n46536), .B(n46540), .X(n11267) );
  nor_x1_sg U62351 ( .A(n17477), .B(n46367), .X(n17476) );
  nor_x1_sg U62352 ( .A(n19022), .B(n46320), .X(n19021) );
  nor_x1_sg U62353 ( .A(n20566), .B(n46275), .X(n20565) );
  nor_x1_sg U62354 ( .A(n46373), .B(n17922), .X(n17920) );
  nor_x1_sg U62355 ( .A(n46326), .B(n19467), .X(n19465) );
  nor_x1_sg U62356 ( .A(n46281), .B(n21011), .X(n21009) );
  nand_x2_sg U62357 ( .A(n51839), .B(n25979), .X(n25978) );
  nand_x2_sg U62358 ( .A(n52391), .B(n26539), .X(n26538) );
  nand_x2_sg U62359 ( .A(n52670), .B(n26817), .X(n26816) );
  nand_x2_sg U62360 ( .A(n53227), .B(n27376), .X(n27375) );
  nand_x2_sg U62361 ( .A(n54070), .B(n28215), .X(n28214) );
  nand_x2_sg U62362 ( .A(n54634), .B(n28773), .X(n28772) );
  nand_x2_sg U62363 ( .A(n55202), .B(n29334), .X(n29333) );
  nand_x2_sg U62364 ( .A(n46536), .B(n25702), .X(n25709) );
  nand_x2_sg U62365 ( .A(n52133), .B(n26261), .X(n26268) );
  nand_x2_sg U62366 ( .A(n52406), .B(n26540), .X(n26547) );
  nand_x2_sg U62367 ( .A(n52683), .B(n26818), .X(n26825) );
  nand_x2_sg U62368 ( .A(n52967), .B(n27097), .X(n27104) );
  nand_x2_sg U62369 ( .A(n53525), .B(n27657), .X(n27664) );
  nand_x2_sg U62370 ( .A(n54084), .B(n28216), .X(n28223) );
  nand_x2_sg U62371 ( .A(n54647), .B(n28774), .X(n28781) );
  nand_x2_sg U62372 ( .A(n55215), .B(n29335), .X(n29342) );
  nand_x2_sg U62373 ( .A(n52378), .B(n26525), .X(n26524) );
  nand_x2_sg U62374 ( .A(n52655), .B(n26803), .X(n26802) );
  nor_x1_sg U62375 ( .A(n46552), .B(n11689), .X(n11687) );
  nor_x1_sg U62376 ( .A(n46508), .B(n13249), .X(n13247) );
  nor_x1_sg U62377 ( .A(n46440), .B(n15582), .X(n15580) );
  nor_x1_sg U62378 ( .A(n46396), .B(n17148), .X(n17146) );
  nor_x1_sg U62379 ( .A(n18476), .B(n46341), .X(n18475) );
  nor_x1_sg U62380 ( .A(n11637), .B(n51714), .X(n11769) );
  nor_x1_sg U62381 ( .A(n18637), .B(n54226), .X(n18772) );
  nor_x1_sg U62382 ( .A(n46227), .B(n26006), .X(n26015) );
  nor_x1_sg U62383 ( .A(n46223), .B(n26566), .X(n26575) );
  nand_x2_sg U62384 ( .A(n54614), .B(n28752), .X(n28751) );
  nand_x2_sg U62385 ( .A(n55182), .B(n29313), .X(n29312) );
  nand_x4_sg U62386 ( .A(n51337), .B(n10979), .X(n10937) );
  nand_x1_sg U62387 ( .A(n10984), .B(n10985), .X(n10980) );
  nand_x4_sg U62388 ( .A(n42276), .B(n12540), .X(n12499) );
  nor_x1_sg U62389 ( .A(n16312), .B(n16357), .X(n16443) );
  nor_x1_sg U62390 ( .A(n19980), .B(n46300), .X(n19979) );
  nor_x1_sg U62391 ( .A(n21525), .B(n46255), .X(n21524) );
  nor_x1_sg U62392 ( .A(n46573), .B(n10908), .X(n10906) );
  nor_x1_sg U62393 ( .A(n46416), .B(n16363), .X(n16361) );
  nor_x1_sg U62394 ( .A(n46528), .B(n12468), .X(n12466) );
  nor_x1_sg U62395 ( .A(n12570), .B(n46519), .X(n12569) );
  nor_x1_sg U62396 ( .A(n12212), .B(n46519), .X(n12211) );
  nand_x4_sg U62397 ( .A(n14304), .B(n44473), .X(n14301) );
  nor_x1_sg U62398 ( .A(n10653), .B(n46566), .X(n10652) );
  nor_x1_sg U62399 ( .A(n18435), .B(n46341), .X(n18434) );
  nand_x4_sg U62400 ( .A(n54128), .B(n18765), .X(n18722) );
  nand_x4_sg U62401 ( .A(n53285), .B(n16437), .X(n16395) );
  nand_x1_sg U62402 ( .A(n16443), .B(n16444), .X(n16438) );
  nor_x1_sg U62403 ( .A(n14132), .B(n46480), .X(n14131) );
  nor_x1_sg U62404 ( .A(n13773), .B(n46480), .X(n13772) );
  nor_x1_sg U62405 ( .A(n16107), .B(n46407), .X(n16106) );
  nand_x1_sg U62406 ( .A(n51671), .B(n25751), .X(n25750) );
  nor_x1_sg U62407 ( .A(n46229), .B(n25742), .X(n25751) );
  nand_x1_sg U62408 ( .A(n53340), .B(n27426), .X(n27425) );
  nor_x1_sg U62409 ( .A(n46217), .B(n27417), .X(n27426) );
  nand_x4_sg U62410 ( .A(n54691), .B(n20311), .X(n20268) );
  nand_x4_sg U62411 ( .A(n55259), .B(n21856), .X(n21813) );
  nor_x1_sg U62412 ( .A(n11319), .B(n46546), .X(n11318) );
  nor_x1_sg U62413 ( .A(n12099), .B(n46519), .X(n12098) );
  nor_x1_sg U62414 ( .A(n15994), .B(n46407), .X(n15993) );
  nor_x1_sg U62415 ( .A(n11432), .B(n46546), .X(n11431) );
  nor_x1_sg U62416 ( .A(n13660), .B(n46480), .X(n13659) );
  nand_x4_sg U62417 ( .A(n18192), .B(n45457), .X(n18189) );
  nand_x4_sg U62418 ( .A(n17425), .B(n44209), .X(n17422) );
  nand_x4_sg U62419 ( .A(n18970), .B(n44207), .X(n18967) );
  nand_x4_sg U62420 ( .A(n19739), .B(n44471), .X(n19736) );
  nand_x4_sg U62421 ( .A(n20514), .B(n44205), .X(n20511) );
  nand_x4_sg U62422 ( .A(n21284), .B(n44469), .X(n21281) );
  nor_x1_sg U62423 ( .A(n11161), .B(n46546), .X(n11160) );
  nand_x4_sg U62424 ( .A(n10412), .B(n44475), .X(n10409) );
  nor_x1_sg U62425 ( .A(n13816), .B(n46480), .X(n13815) );
  nor_x1_sg U62426 ( .A(n12880), .B(n46502), .X(n12879) );
  nor_x1_sg U62427 ( .A(n15213), .B(n46434), .X(n15212) );
  nor_x1_sg U62428 ( .A(n16779), .B(n46390), .X(n16778) );
  nor_x1_sg U62429 ( .A(n46306), .B(n20237), .X(n20235) );
  nor_x1_sg U62430 ( .A(n46261), .B(n21782), .X(n21780) );
  nor_x1_sg U62431 ( .A(n13352), .B(n46502), .X(n13351) );
  nor_x1_sg U62432 ( .A(n15685), .B(n46434), .X(n15684) );
  nor_x1_sg U62433 ( .A(n17251), .B(n46390), .X(n17250) );
  nand_x2_sg U62434 ( .A(n46564), .B(n10992), .X(n10991) );
  nor_x1_sg U62435 ( .A(n12993), .B(n46502), .X(n12992) );
  nor_x1_sg U62436 ( .A(n15326), .B(n46434), .X(n15325) );
  nor_x1_sg U62437 ( .A(n16892), .B(n46390), .X(n16891) );
  nor_x1_sg U62438 ( .A(n14354), .B(n46452), .X(n14353) );
  nor_x1_sg U62439 ( .A(n14545), .B(n46452), .X(n14544) );
  nor_x1_sg U62440 ( .A(n12255), .B(n46519), .X(n12254) );
  nor_x1_sg U62441 ( .A(n14586), .B(n46452), .X(n14585) );
  nor_x1_sg U62442 ( .A(n46463), .B(n14801), .X(n14799) );
  nor_x1_sg U62443 ( .A(n18244), .B(n46341), .X(n18243) );
  nand_x2_sg U62444 ( .A(n51280), .B(n25422), .X(n25421) );
  nor_x1_sg U62445 ( .A(n16150), .B(n46407), .X(n16149) );
  nor_x1_sg U62446 ( .A(n17406), .B(n46367), .X(n17405) );
  nor_x1_sg U62447 ( .A(n18951), .B(n46320), .X(n18950) );
  nor_x1_sg U62448 ( .A(n20495), .B(n46275), .X(n20494) );
  nand_x4_sg U62449 ( .A(n52727), .B(n14875), .X(n14832) );
  nor_x1_sg U62450 ( .A(n11171), .B(n46546), .X(n11170) );
  nor_x1_sg U62451 ( .A(n12732), .B(n46502), .X(n12731) );
  nor_x1_sg U62452 ( .A(n15065), .B(n46434), .X(n15064) );
  nor_x1_sg U62453 ( .A(n16631), .B(n46390), .X(n16630) );
  nor_x1_sg U62454 ( .A(n17666), .B(n46367), .X(n17665) );
  nor_x1_sg U62455 ( .A(n19211), .B(n46320), .X(n19210) );
  nor_x1_sg U62456 ( .A(n20755), .B(n46275), .X(n20754) );
  nor_x1_sg U62457 ( .A(n46353), .B(n18691), .X(n18689) );
  nor_x1_sg U62458 ( .A(n18703), .B(n46340), .X(n18702) );
  nor_x1_sg U62459 ( .A(n19722), .B(n46300), .X(n19721) );
  nor_x1_sg U62460 ( .A(n21267), .B(n46255), .X(n21266) );
  nor_x1_sg U62461 ( .A(n10462), .B(n46566), .X(n10461) );
  nor_x1_sg U62462 ( .A(n11945), .B(n46519), .X(n11944) );
  nor_x1_sg U62463 ( .A(n15840), .B(n46407), .X(n15839) );
  nor_x1_sg U62464 ( .A(n18587), .B(n46341), .X(n18586) );
  nand_x4_sg U62465 ( .A(n54109), .B(n18595), .X(n18593) );
  nor_x1_sg U62466 ( .A(n10694), .B(n46566), .X(n10693) );
  nor_x1_sg U62467 ( .A(n20021), .B(n46300), .X(n20020) );
  nor_x1_sg U62468 ( .A(n21566), .B(n46255), .X(n21565) );
  nor_x1_sg U62469 ( .A(n19789), .B(n46300), .X(n19788) );
  nor_x1_sg U62470 ( .A(n21334), .B(n46255), .X(n21333) );
  nor_x1_sg U62471 ( .A(n20133), .B(n46300), .X(n20132) );
  nor_x1_sg U62472 ( .A(n21678), .B(n46255), .X(n21677) );
  nand_x4_sg U62473 ( .A(n51618), .B(n11763), .X(n11720) );
  nand_x1_sg U62474 ( .A(n11766), .B(n41162), .X(n11765) );
  nor_x1_sg U62475 ( .A(n14287), .B(n46452), .X(n14286) );
  nor_x1_sg U62476 ( .A(n43051), .B(n46407), .X(n16410) );
  nor_x1_sg U62477 ( .A(n43847), .B(n46300), .X(n20284) );
  nor_x1_sg U62478 ( .A(n43845), .B(n46255), .X(n21829) );
  nor_x1_sg U62479 ( .A(n43049), .B(n46546), .X(n11736) );
  nor_x1_sg U62480 ( .A(n43045), .B(n46502), .X(n13297) );
  nor_x1_sg U62481 ( .A(n43041), .B(n46434), .X(n15630) );
  nor_x1_sg U62482 ( .A(n43037), .B(n46390), .X(n17196) );
  nor_x1_sg U62483 ( .A(n43043), .B(n46480), .X(n14077) );
  nor_x1_sg U62484 ( .A(n43047), .B(n46519), .X(n12516) );
  nand_x2_sg U62485 ( .A(n52809), .B(n52843), .X(n14917) );
  nand_x2_sg U62486 ( .A(n14886), .B(n14883), .X(n14916) );
  nand_x2_sg U62487 ( .A(n53929), .B(n53963), .X(n18038) );
  nand_x2_sg U62488 ( .A(n18007), .B(n18004), .X(n18037) );
  nand_x2_sg U62489 ( .A(n54494), .B(n54528), .X(n19583) );
  nand_x2_sg U62490 ( .A(n19552), .B(n19549), .X(n19582) );
  nand_x2_sg U62491 ( .A(n55062), .B(n55096), .X(n21127) );
  nand_x2_sg U62492 ( .A(n21096), .B(n21093), .X(n21126) );
  nor_x1_sg U62493 ( .A(n43798), .B(n46566), .X(n10952) );
  nor_x1_sg U62494 ( .A(n43943), .B(n46341), .X(n18738) );
  nand_x2_sg U62495 ( .A(n54778), .B(n54813), .X(n20353) );
  nand_x2_sg U62496 ( .A(n20322), .B(n20319), .X(n20352) );
  nand_x2_sg U62497 ( .A(n55346), .B(n55381), .X(n21898) );
  nand_x2_sg U62498 ( .A(n21867), .B(n21864), .X(n21897) );
  nand_x4_sg U62499 ( .A(n11566), .B(n11565), .X(n11558) );
  nand_x4_sg U62500 ( .A(n16242), .B(n16241), .X(n16233) );
  nand_x4_sg U62501 ( .A(n53847), .B(n17996), .X(n17953) );
  nand_x4_sg U62502 ( .A(n54412), .B(n19541), .X(n19498) );
  nand_x4_sg U62503 ( .A(n54980), .B(n21085), .X(n21042) );
  nand_x4_sg U62504 ( .A(n20111), .B(n20110), .X(n20102) );
  nand_x4_sg U62505 ( .A(n21656), .B(n21655), .X(n21647) );
  nand_x4_sg U62506 ( .A(n42282), .B(n10784), .X(n10776) );
  nand_x4_sg U62507 ( .A(n46536), .B(n11427), .X(n11373) );
  nand_x1_sg U62508 ( .A(n51637), .B(n51560), .X(n11427) );
  nand_x4_sg U62509 ( .A(n52133), .B(n12988), .X(n12934) );
  nand_x1_sg U62510 ( .A(n52193), .B(n52117), .X(n12988) );
  nand_x4_sg U62511 ( .A(n52967), .B(n15321), .X(n15267) );
  nand_x1_sg U62512 ( .A(n53027), .B(n52951), .X(n15321) );
  nand_x4_sg U62513 ( .A(n53525), .B(n16887), .X(n16833) );
  nand_x1_sg U62514 ( .A(n53585), .B(n53509), .X(n16887) );
  nand_x4_sg U62515 ( .A(n44437), .B(n13347), .X(n13338) );
  nand_x4_sg U62516 ( .A(n44435), .B(n14127), .X(n14118) );
  nand_x4_sg U62517 ( .A(n44433), .B(n15680), .X(n15671) );
  nand_x4_sg U62518 ( .A(n44431), .B(n17246), .X(n17237) );
  nand_x4_sg U62519 ( .A(n18595), .B(n18633), .X(n18631) );
  nand_x1_sg U62520 ( .A(n14370), .B(n52678), .X(n14367) );
  nand_x1_sg U62521 ( .A(n19805), .B(n54642), .X(n19802) );
  nand_x1_sg U62522 ( .A(n21350), .B(n55210), .X(n21347) );
  nor_x1_sg U62523 ( .A(n10902), .B(n46555), .X(n10901) );
  nor_x1_sg U62524 ( .A(n18271), .B(n46344), .X(n18270) );
  nand_x4_sg U62525 ( .A(n10747), .B(n44467), .X(n10727) );
  nand_x4_sg U62526 ( .A(n20073), .B(n44465), .X(n20054) );
  nand_x4_sg U62527 ( .A(n21618), .B(n44463), .X(n21599) );
  nand_x4_sg U62528 ( .A(n14639), .B(n44447), .X(n14619) );
  nand_x4_sg U62529 ( .A(n17760), .B(n44445), .X(n17740) );
  nand_x4_sg U62530 ( .A(n18528), .B(n44211), .X(n18509) );
  nand_x4_sg U62531 ( .A(n19305), .B(n44443), .X(n19285) );
  nand_x4_sg U62532 ( .A(n20849), .B(n44441), .X(n20829) );
  nand_x4_sg U62533 ( .A(n53877), .B(n17619), .X(n17576) );
  nand_x1_sg U62534 ( .A(n53876), .B(n17620), .X(n17619) );
  nand_x4_sg U62535 ( .A(n54442), .B(n19164), .X(n19121) );
  nand_x1_sg U62536 ( .A(n54441), .B(n19165), .X(n19164) );
  nand_x4_sg U62537 ( .A(n55010), .B(n20708), .X(n20665) );
  nand_x1_sg U62538 ( .A(n55009), .B(n20709), .X(n20708) );
  nand_x4_sg U62539 ( .A(n51645), .B(n11384), .X(n11360) );
  nand_x1_sg U62540 ( .A(n51644), .B(n11385), .X(n11384) );
  nand_x4_sg U62541 ( .A(n51925), .B(n12164), .X(n12140) );
  nand_x1_sg U62542 ( .A(n51924), .B(n12165), .X(n12164) );
  nand_x4_sg U62543 ( .A(n52201), .B(n12945), .X(n12921) );
  nand_x1_sg U62544 ( .A(n52200), .B(n12946), .X(n12945) );
  nand_x4_sg U62545 ( .A(n53035), .B(n15278), .X(n15254) );
  nand_x1_sg U62546 ( .A(n53034), .B(n15279), .X(n15278) );
  nand_x4_sg U62547 ( .A(n53313), .B(n16059), .X(n16035) );
  nand_x1_sg U62548 ( .A(n53312), .B(n16060), .X(n16059) );
  nand_x4_sg U62549 ( .A(n53593), .B(n16844), .X(n16820) );
  nand_x1_sg U62550 ( .A(n53592), .B(n16845), .X(n16844) );
  nand_x4_sg U62551 ( .A(n51360), .B(n10606), .X(n10564) );
  nand_x1_sg U62552 ( .A(n51359), .B(n10607), .X(n10606) );
  nand_x4_sg U62553 ( .A(n41259), .B(n14743), .X(n14717) );
  nand_x4_sg U62554 ( .A(n41257), .B(n17864), .X(n17838) );
  nand_x4_sg U62555 ( .A(n41255), .B(n19409), .X(n19383) );
  nand_x4_sg U62556 ( .A(n41253), .B(n20953), .X(n20927) );
  nand_x4_sg U62557 ( .A(n41239), .B(n10851), .X(n10825) );
  nand_x4_sg U62558 ( .A(n14350), .B(n14349), .X(n14344) );
  nand_x4_sg U62559 ( .A(n17470), .B(n17469), .X(n17467) );
  nand_x4_sg U62560 ( .A(n19015), .B(n19014), .X(n19012) );
  nand_x4_sg U62561 ( .A(n20559), .B(n20558), .X(n20556) );
  nand_x4_sg U62562 ( .A(n10455), .B(n10454), .X(n10452) );
  nand_x4_sg U62563 ( .A(n42286), .B(n19781), .X(n19779) );
  nand_x4_sg U62564 ( .A(n42284), .B(n21326), .X(n21324) );
  nand_x4_sg U62565 ( .A(n14677), .B(n14676), .X(n14668) );
  nand_x4_sg U62566 ( .A(n12347), .B(n12346), .X(n12338) );
  nand_x4_sg U62567 ( .A(n13127), .B(n13126), .X(n13119) );
  nand_x4_sg U62568 ( .A(n15460), .B(n15459), .X(n15452) );
  nand_x4_sg U62569 ( .A(n17026), .B(n17025), .X(n17018) );
  nand_x4_sg U62570 ( .A(n20141), .B(n20179), .X(n20177) );
  nand_x1_sg U62571 ( .A(n46286), .B(n20139), .X(n20179) );
  nand_x4_sg U62572 ( .A(n21686), .B(n21724), .X(n21722) );
  nand_x1_sg U62573 ( .A(n46241), .B(n21684), .X(n21724) );
  nand_x1_sg U62574 ( .A(n11175), .B(n11195), .X(n11192) );
  nor_x1_sg U62575 ( .A(n11175), .B(n46546), .X(n11194) );
  nand_x1_sg U62576 ( .A(n12736), .B(n12756), .X(n12753) );
  nor_x1_sg U62577 ( .A(n12736), .B(n46502), .X(n12755) );
  nand_x1_sg U62578 ( .A(n15069), .B(n15089), .X(n15086) );
  nor_x1_sg U62579 ( .A(n15069), .B(n46434), .X(n15088) );
  nand_x1_sg U62580 ( .A(n16635), .B(n16655), .X(n16652) );
  nor_x1_sg U62581 ( .A(n16635), .B(n46390), .X(n16654) );
  nand_x4_sg U62582 ( .A(n53400), .B(n16478), .X(n16451) );
  nand_x1_sg U62583 ( .A(n16444), .B(n16479), .X(n16478) );
  nor_x1_sg U62584 ( .A(n16479), .B(n16444), .X(n16480) );
  nand_x4_sg U62585 ( .A(n51339), .B(n10521), .X(n10538) );
  nand_x4_sg U62586 ( .A(n51275), .B(n10295), .X(n9034) );
  nand_x1_sg U62587 ( .A(n43773), .B(n44140), .X(n10295) );
  nand_x1_sg U62588 ( .A(n43755), .B(n43157), .X(n11846) );
  nand_x4_sg U62589 ( .A(n52664), .B(n14187), .X(n8940) );
  nand_x1_sg U62590 ( .A(n43802), .B(n44405), .X(n14187) );
  nand_x1_sg U62591 ( .A(n43771), .B(n43143), .X(n15741) );
  nand_x1_sg U62592 ( .A(n41594), .B(n43149), .X(n19623) );
  nand_x4_sg U62593 ( .A(n55197), .B(n21168), .X(n9119) );
  nand_x1_sg U62594 ( .A(n42815), .B(n44138), .X(n21168) );
  nand_x1_sg U62595 ( .A(n43973), .B(n44403), .X(n18078) );
  nand_x1_sg U62596 ( .A(n43800), .B(n43153), .X(n13408) );
  nand_x4_sg U62597 ( .A(n42192), .B(n11309), .X(n11302) );
  nand_x1_sg U62598 ( .A(n41510), .B(n44421), .X(n11309) );
  nand_x4_sg U62599 ( .A(n42190), .B(n12089), .X(n12082) );
  nand_x1_sg U62600 ( .A(n41506), .B(n44152), .X(n12089) );
  nand_x4_sg U62601 ( .A(n41709), .B(n12870), .X(n12863) );
  nand_x1_sg U62602 ( .A(n41229), .B(n42813), .X(n12870) );
  nand_x4_sg U62603 ( .A(n41705), .B(n15203), .X(n15196) );
  nand_x1_sg U62604 ( .A(n41225), .B(n42809), .X(n15203) );
  nand_x4_sg U62605 ( .A(n42188), .B(n15984), .X(n15977) );
  nand_x1_sg U62606 ( .A(n41498), .B(n44419), .X(n15984) );
  nand_x4_sg U62607 ( .A(n41703), .B(n16769), .X(n16762) );
  nand_x1_sg U62608 ( .A(n41221), .B(n42807), .X(n16769) );
  nand_x4_sg U62609 ( .A(n46452), .B(n46463), .X(n26796) );
  nand_x4_sg U62610 ( .A(n46341), .B(n46353), .X(n28194) );
  nand_x4_sg U62611 ( .A(n46566), .B(n46573), .X(n25401) );
  nand_x4_sg U62612 ( .A(n17462), .B(n44461), .X(n17460) );
  nand_x4_sg U62613 ( .A(n19007), .B(n44459), .X(n19005) );
  nand_x4_sg U62614 ( .A(n20551), .B(n44457), .X(n20549) );
  nor_x1_sg U62615 ( .A(n46229), .B(n25728), .X(n25737) );
  nor_x1_sg U62616 ( .A(n46225), .B(n26287), .X(n26296) );
  nor_x1_sg U62617 ( .A(n46219), .B(n27123), .X(n27132) );
  nor_x1_sg U62618 ( .A(n46215), .B(n27683), .X(n27692) );
  nand_x1_sg U62619 ( .A(n10841), .B(n51381), .X(n10840) );
  nor_x1_sg U62620 ( .A(n16312), .B(n16313), .X(n16311) );
  nor_x1_sg U62621 ( .A(n12417), .B(n12416), .X(n12418) );
  nand_x4_sg U62622 ( .A(n10854), .B(n51447), .X(n10814) );
  nand_x1_sg U62623 ( .A(n10857), .B(n10856), .X(n10854) );
  nor_x1_sg U62624 ( .A(n10856), .B(n10857), .X(n10855) );
  nand_x4_sg U62625 ( .A(n46546), .B(n46552), .X(n25680) );
  nand_x4_sg U62626 ( .A(n46502), .B(n46508), .X(n26239) );
  nand_x4_sg U62627 ( .A(n46434), .B(n46440), .X(n27075) );
  nand_x4_sg U62628 ( .A(n46390), .B(n46396), .X(n27635) );
  nand_x4_sg U62629 ( .A(n46300), .B(n46306), .X(n28752) );
  nand_x4_sg U62630 ( .A(n46255), .B(n46261), .X(n29313) );
  nand_x4_sg U62631 ( .A(n51452), .B(n11019), .X(n10992) );
  nand_x1_sg U62632 ( .A(n10985), .B(n11020), .X(n11019) );
  nor_x1_sg U62633 ( .A(n11020), .B(n10985), .X(n11021) );
  nand_x4_sg U62634 ( .A(n54693), .B(n19848), .X(n19865) );
  nand_x4_sg U62635 ( .A(n55261), .B(n21393), .X(n21410) );
  nor_x1_sg U62636 ( .A(n14748), .B(n14747), .X(n14749) );
  nand_x4_sg U62637 ( .A(n12477), .B(n12478), .X(n12476) );
  nand_x1_sg U62638 ( .A(n12480), .B(n12481), .X(n12477) );
  nand_x1_sg U62639 ( .A(n12479), .B(n51995), .X(n12478) );
  nand_x1_sg U62640 ( .A(n51995), .B(n46517), .X(n12481) );
  nand_x4_sg U62641 ( .A(n13258), .B(n13259), .X(n13257) );
  nand_x1_sg U62642 ( .A(n13261), .B(n13262), .X(n13258) );
  nand_x1_sg U62643 ( .A(n13260), .B(n52271), .X(n13259) );
  nand_x1_sg U62644 ( .A(n52271), .B(n46496), .X(n13262) );
  nand_x4_sg U62645 ( .A(n14038), .B(n14039), .X(n14037) );
  nand_x1_sg U62646 ( .A(n14041), .B(n14042), .X(n14038) );
  nand_x1_sg U62647 ( .A(n14040), .B(n52546), .X(n14039) );
  nand_x1_sg U62648 ( .A(n52546), .B(n46474), .X(n14042) );
  nand_x4_sg U62649 ( .A(n15591), .B(n15592), .X(n15590) );
  nand_x1_sg U62650 ( .A(n15594), .B(n15595), .X(n15591) );
  nand_x1_sg U62651 ( .A(n15593), .B(n53105), .X(n15592) );
  nand_x1_sg U62652 ( .A(n53105), .B(n46428), .X(n15595) );
  nand_x4_sg U62653 ( .A(n17157), .B(n17158), .X(n17156) );
  nand_x1_sg U62654 ( .A(n17160), .B(n17161), .X(n17157) );
  nand_x1_sg U62655 ( .A(n17159), .B(n53663), .X(n17158) );
  nand_x1_sg U62656 ( .A(n53663), .B(n46384), .X(n17161) );
  nand_x4_sg U62657 ( .A(n20223), .B(n20224), .X(n20221) );
  nand_x1_sg U62658 ( .A(n20225), .B(n20226), .X(n20224) );
  nand_x1_sg U62659 ( .A(n20230), .B(n54751), .X(n20223) );
  nor_x1_sg U62660 ( .A(n20227), .B(n20228), .X(n20225) );
  nand_x4_sg U62661 ( .A(n21768), .B(n21769), .X(n21766) );
  nand_x1_sg U62662 ( .A(n21770), .B(n21771), .X(n21769) );
  nand_x1_sg U62663 ( .A(n21775), .B(n55319), .X(n21768) );
  nor_x1_sg U62664 ( .A(n21772), .B(n21773), .X(n21770) );
  nor_x1_sg U62665 ( .A(n17869), .B(n17868), .X(n17870) );
  nor_x1_sg U62666 ( .A(n19414), .B(n19413), .X(n19415) );
  nor_x1_sg U62667 ( .A(n20958), .B(n20957), .X(n20959) );
  nor_x1_sg U62668 ( .A(n20182), .B(n20181), .X(n20183) );
  nor_x1_sg U62669 ( .A(n21727), .B(n21726), .X(n21728) );
  nand_x4_sg U62670 ( .A(n10844), .B(n10845), .X(n10754) );
  nand_x1_sg U62671 ( .A(n51381), .B(n51406), .X(n10845) );
  nand_x1_sg U62672 ( .A(n10841), .B(n10838), .X(n10844) );
  nor_x1_sg U62673 ( .A(n18741), .B(n54160), .X(n18745) );
  nor_x1_sg U62674 ( .A(n53869), .B(n17625), .X(n17626) );
  nor_x1_sg U62675 ( .A(n54434), .B(n19170), .X(n19171) );
  nor_x1_sg U62676 ( .A(n55002), .B(n20714), .X(n20715) );
  nand_x4_sg U62677 ( .A(n46519), .B(n46528), .X(n25958) );
  nand_x4_sg U62678 ( .A(n46407), .B(n46416), .X(n27355) );
  nor_x1_sg U62679 ( .A(n52749), .B(n14504), .X(n14505) );
  nand_x4_sg U62680 ( .A(n18624), .B(n18625), .X(n18535) );
  nand_x4_sg U62681 ( .A(n53849), .B(n17533), .X(n17550) );
  nand_x4_sg U62682 ( .A(n54414), .B(n19078), .X(n19095) );
  nand_x4_sg U62683 ( .A(n54982), .B(n20622), .X(n20639) );
  nand_x4_sg U62684 ( .A(n52729), .B(n14413), .X(n14431) );
  nand_x4_sg U62685 ( .A(n44156), .B(n17451), .X(n17397) );
  nand_x4_sg U62686 ( .A(n44155), .B(n18996), .X(n18942) );
  nand_x4_sg U62687 ( .A(n44154), .B(n20540), .X(n20486) );
  nand_x4_sg U62688 ( .A(n18678), .B(n18679), .X(n18676) );
  nand_x1_sg U62689 ( .A(n18680), .B(n18681), .X(n18679) );
  nand_x1_sg U62690 ( .A(n18684), .B(n54184), .X(n18678) );
  nor_x1_sg U62691 ( .A(n18682), .B(n18683), .X(n18680) );
  nor_x1_sg U62692 ( .A(n11238), .B(n11239), .X(n11237) );
  nand_x1_sg U62693 ( .A(n11522), .B(n51666), .X(n11521) );
  nand_x1_sg U62694 ( .A(n11523), .B(n51684), .X(n11520) );
  nand_x1_sg U62695 ( .A(n16197), .B(n53335), .X(n16196) );
  nand_x1_sg U62696 ( .A(n16198), .B(n53353), .X(n16195) );
  nand_x4_sg U62697 ( .A(n11698), .B(n11699), .X(n11697) );
  nand_x1_sg U62698 ( .A(n11701), .B(n11702), .X(n11698) );
  nand_x1_sg U62699 ( .A(n11700), .B(n51717), .X(n11699) );
  nand_x1_sg U62700 ( .A(n51717), .B(n46540), .X(n11702) );
  nor_x1_sg U62701 ( .A(n13198), .B(n13199), .X(n13197) );
  nor_x1_sg U62702 ( .A(n13978), .B(n13979), .X(n13977) );
  nor_x1_sg U62703 ( .A(n15531), .B(n15532), .X(n15530) );
  nor_x1_sg U62704 ( .A(n17097), .B(n17098), .X(n17096) );
  nor_x1_sg U62705 ( .A(n12799), .B(n12800), .X(n12798) );
  nor_x1_sg U62706 ( .A(n15132), .B(n15133), .X(n15131) );
  nor_x1_sg U62707 ( .A(n16698), .B(n16699), .X(n16697) );
  nand_x1_sg U62708 ( .A(n17755), .B(n53898), .X(n17754) );
  nand_x1_sg U62709 ( .A(n17756), .B(n53916), .X(n17753) );
  nand_x1_sg U62710 ( .A(n19300), .B(n54463), .X(n19299) );
  nand_x1_sg U62711 ( .A(n19301), .B(n54481), .X(n19298) );
  nand_x1_sg U62712 ( .A(n20844), .B(n55031), .X(n20843) );
  nand_x1_sg U62713 ( .A(n20845), .B(n55049), .X(n20842) );
  nand_x4_sg U62714 ( .A(n12719), .B(n12720), .X(n12622) );
  nand_x1_sg U62715 ( .A(n12722), .B(n12723), .X(n12719) );
  nor_x1_sg U62716 ( .A(n12722), .B(n46502), .X(n12721) );
  nand_x4_sg U62717 ( .A(n15052), .B(n15053), .X(n14955) );
  nand_x1_sg U62718 ( .A(n15055), .B(n15056), .X(n15052) );
  nor_x1_sg U62719 ( .A(n15055), .B(n46434), .X(n15054) );
  nand_x4_sg U62720 ( .A(n16618), .B(n16619), .X(n16521) );
  nand_x1_sg U62721 ( .A(n16621), .B(n16622), .X(n16618) );
  nor_x1_sg U62722 ( .A(n16621), .B(n46390), .X(n16620) );
  nand_x1_sg U62723 ( .A(n20068), .B(n54745), .X(n20067) );
  nand_x1_sg U62724 ( .A(n20069), .B(n54767), .X(n20066) );
  nand_x1_sg U62725 ( .A(n21613), .B(n55313), .X(n21612) );
  nand_x1_sg U62726 ( .A(n21614), .B(n55335), .X(n21611) );
  nand_x1_sg U62727 ( .A(n16416), .B(n53316), .X(n16415) );
  nand_x1_sg U62728 ( .A(n16417), .B(n53403), .X(n16414) );
  nand_x4_sg U62729 ( .A(n16379), .B(n16380), .X(n16372) );
  nand_x1_sg U62730 ( .A(n16199), .B(n16382), .X(n16379) );
  nand_x1_sg U62731 ( .A(n16381), .B(n53408), .X(n16380) );
  nand_x1_sg U62732 ( .A(n53408), .B(n53214), .X(n16382) );
  nand_x4_sg U62733 ( .A(n46478), .B(n46484), .X(n13399) );
  nand_x1_sg U62734 ( .A(n11743), .B(n51733), .X(n11740) );
  nand_x1_sg U62735 ( .A(n11742), .B(n51647), .X(n11741) );
  nand_x1_sg U62736 ( .A(n13304), .B(n52288), .X(n13301) );
  nand_x1_sg U62737 ( .A(n13303), .B(n52203), .X(n13302) );
  nand_x1_sg U62738 ( .A(n15637), .B(n53122), .X(n15634) );
  nand_x1_sg U62739 ( .A(n15636), .B(n53037), .X(n15635) );
  nand_x1_sg U62740 ( .A(n17203), .B(n53680), .X(n17200) );
  nand_x1_sg U62741 ( .A(n17202), .B(n53595), .X(n17201) );
  nand_x4_sg U62742 ( .A(n17973), .B(n17974), .X(n17889) );
  nand_x1_sg U62743 ( .A(n17976), .B(n53953), .X(n17973) );
  nand_x1_sg U62744 ( .A(n17975), .B(n53880), .X(n17974) );
  nand_x4_sg U62745 ( .A(n19518), .B(n19519), .X(n19434) );
  nand_x1_sg U62746 ( .A(n19521), .B(n54518), .X(n19518) );
  nand_x1_sg U62747 ( .A(n19520), .B(n54445), .X(n19519) );
  nand_x4_sg U62748 ( .A(n21062), .B(n21063), .X(n20978) );
  nand_x1_sg U62749 ( .A(n21065), .B(n55086), .X(n21062) );
  nand_x1_sg U62750 ( .A(n21064), .B(n55013), .X(n21063) );
  nand_x1_sg U62751 ( .A(n12523), .B(n52011), .X(n12520) );
  nand_x1_sg U62752 ( .A(n12522), .B(n51928), .X(n12521) );
  nand_x1_sg U62753 ( .A(n14084), .B(n52563), .X(n14081) );
  nand_x1_sg U62754 ( .A(n14083), .B(n52480), .X(n14082) );
  nand_x4_sg U62755 ( .A(n14852), .B(n14853), .X(n14768) );
  nand_x1_sg U62756 ( .A(n14855), .B(n52833), .X(n14852) );
  nand_x1_sg U62757 ( .A(n14854), .B(n52760), .X(n14853) );
  nand_x4_sg U62758 ( .A(n11214), .B(n51571), .X(n11211) );
  nand_x1_sg U62759 ( .A(n11217), .B(n11216), .X(n11214) );
  nor_x1_sg U62760 ( .A(n11216), .B(n11217), .X(n11215) );
  nand_x2_sg U62761 ( .A(n51287), .B(n10537), .X(n10574) );
  nand_x2_sg U62762 ( .A(n51299), .B(n10493), .X(n10573) );
  nor_x1_sg U62763 ( .A(n55660), .B(n46585), .X(\L1_0/n4502 ) );
  nor_x1_sg U62764 ( .A(n55720), .B(n46591), .X(\L1_0/n4022 ) );
  nor_x1_sg U62765 ( .A(n46591), .B(n27939), .X(\L1_0/n4003 ) );
  nor_x1_sg U62766 ( .A(n55725), .B(n46591), .X(\L1_0/n4002 ) );
  nor_x1_sg U62767 ( .A(n46591), .B(n27960), .X(\L1_0/n3991 ) );
  nor_x1_sg U62768 ( .A(n55726), .B(n46591), .X(\L1_0/n3990 ) );
  nor_x1_sg U62769 ( .A(n46591), .B(n55584), .X(\L1_0/n3987 ) );
  nor_x1_sg U62770 ( .A(n43914), .B(n46591), .X(\L1_0/n3986 ) );
  nor_x1_sg U62771 ( .A(n46591), .B(n27974), .X(\L1_0/n3983 ) );
  nor_x1_sg U62772 ( .A(n55727), .B(n46591), .X(\L1_0/n3982 ) );
  nor_x1_sg U62773 ( .A(n46591), .B(n55585), .X(\L1_0/n3979 ) );
  nor_x1_sg U62774 ( .A(n43823), .B(n46591), .X(\L1_0/n3978 ) );
  nor_x1_sg U62775 ( .A(n46591), .B(n27988), .X(\L1_0/n3975 ) );
  nor_x1_sg U62776 ( .A(n55728), .B(n46591), .X(\L1_0/n3974 ) );
  nor_x1_sg U62777 ( .A(n46591), .B(n55586), .X(\L1_0/n3971 ) );
  nor_x1_sg U62778 ( .A(n43794), .B(n46591), .X(\L1_0/n3970 ) );
  nor_x1_sg U62779 ( .A(n28459), .B(n28497), .X(\L1_0/n3843 ) );
  nor_x1_sg U62780 ( .A(n55770), .B(n46596), .X(\L1_0/n3622 ) );
  nand_x4_sg U62781 ( .A(n12775), .B(n52128), .X(n12772) );
  nand_x1_sg U62782 ( .A(n12778), .B(n12777), .X(n12775) );
  nor_x1_sg U62783 ( .A(n12777), .B(n12778), .X(n12776) );
  nand_x4_sg U62784 ( .A(n15108), .B(n52962), .X(n15105) );
  nand_x1_sg U62785 ( .A(n15111), .B(n15110), .X(n15108) );
  nor_x1_sg U62786 ( .A(n15110), .B(n15111), .X(n15109) );
  nand_x4_sg U62787 ( .A(n16674), .B(n53520), .X(n16671) );
  nand_x1_sg U62788 ( .A(n16677), .B(n16676), .X(n16674) );
  nor_x1_sg U62789 ( .A(n16676), .B(n16677), .X(n16675) );
  nor_x1_sg U62790 ( .A(n46585), .B(n26263), .X(\L1_0/n4483 ) );
  nor_x1_sg U62791 ( .A(n55665), .B(n46585), .X(\L1_0/n4482 ) );
  nor_x1_sg U62792 ( .A(n46585), .B(n26284), .X(\L1_0/n4471 ) );
  nor_x1_sg U62793 ( .A(n55666), .B(n46585), .X(\L1_0/n4470 ) );
  nor_x1_sg U62794 ( .A(n46585), .B(n55537), .X(\L1_0/n4467 ) );
  nor_x1_sg U62795 ( .A(n44239), .B(n46585), .X(\L1_0/n4466 ) );
  nor_x1_sg U62796 ( .A(n46585), .B(n26298), .X(\L1_0/n4463 ) );
  nor_x1_sg U62797 ( .A(n55667), .B(n46585), .X(\L1_0/n4462 ) );
  nor_x1_sg U62798 ( .A(n46585), .B(n55538), .X(\L1_0/n4459 ) );
  nor_x1_sg U62799 ( .A(n43831), .B(n46585), .X(\L1_0/n4458 ) );
  nor_x1_sg U62800 ( .A(n46585), .B(n26312), .X(\L1_0/n4455 ) );
  nor_x1_sg U62801 ( .A(n55668), .B(n46585), .X(\L1_0/n4454 ) );
  nor_x1_sg U62802 ( .A(n46585), .B(n55539), .X(\L1_0/n4451 ) );
  nor_x1_sg U62803 ( .A(n43928), .B(n46585), .X(\L1_0/n4450 ) );
  nor_x1_sg U62804 ( .A(n46587), .B(n26542), .X(\L1_0/n4403 ) );
  nor_x1_sg U62805 ( .A(n55675), .B(n46587), .X(\L1_0/n4402 ) );
  nor_x1_sg U62806 ( .A(n46587), .B(n55543), .X(\L1_0/n4399 ) );
  nor_x1_sg U62807 ( .A(n44056), .B(n46587), .X(\L1_0/n4398 ) );
  nor_x1_sg U62808 ( .A(n46587), .B(n26563), .X(\L1_0/n4391 ) );
  nor_x1_sg U62809 ( .A(n55676), .B(n46587), .X(\L1_0/n4390 ) );
  nor_x1_sg U62810 ( .A(n46587), .B(n55545), .X(\L1_0/n4387 ) );
  nor_x1_sg U62811 ( .A(n43926), .B(n46587), .X(\L1_0/n4386 ) );
  nor_x1_sg U62812 ( .A(n46587), .B(n26577), .X(\L1_0/n4383 ) );
  nor_x1_sg U62813 ( .A(n55677), .B(n46587), .X(\L1_0/n4382 ) );
  nor_x1_sg U62814 ( .A(n46587), .B(n55546), .X(\L1_0/n4379 ) );
  nor_x1_sg U62815 ( .A(n43924), .B(n46587), .X(\L1_0/n4378 ) );
  nor_x1_sg U62816 ( .A(n46587), .B(n26591), .X(\L1_0/n4375 ) );
  nor_x1_sg U62817 ( .A(n55678), .B(n46587), .X(\L1_0/n4374 ) );
  nor_x1_sg U62818 ( .A(n46587), .B(n55547), .X(\L1_0/n4371 ) );
  nor_x1_sg U62819 ( .A(n44237), .B(n46587), .X(\L1_0/n4370 ) );
  nor_x1_sg U62820 ( .A(n55690), .B(n46589), .X(\L1_0/n4262 ) );
  nor_x1_sg U62821 ( .A(n55745), .B(n28459), .X(\L1_0/n3842 ) );
  nor_x1_sg U62822 ( .A(n28459), .B(n28518), .X(\L1_0/n3831 ) );
  nor_x1_sg U62823 ( .A(n55746), .B(n28459), .X(\L1_0/n3830 ) );
  nor_x1_sg U62824 ( .A(n28459), .B(n55600), .X(\L1_0/n3827 ) );
  nor_x1_sg U62825 ( .A(n43821), .B(n28459), .X(\L1_0/n3826 ) );
  nor_x1_sg U62826 ( .A(n28459), .B(n28532), .X(\L1_0/n3823 ) );
  nor_x1_sg U62827 ( .A(n55747), .B(n28459), .X(\L1_0/n3822 ) );
  nor_x1_sg U62828 ( .A(n28459), .B(n55601), .X(\L1_0/n3819 ) );
  nor_x1_sg U62829 ( .A(n43819), .B(n28459), .X(\L1_0/n3818 ) );
  nor_x1_sg U62830 ( .A(n28459), .B(n28546), .X(\L1_0/n3815 ) );
  nor_x1_sg U62831 ( .A(n55748), .B(n28459), .X(\L1_0/n3814 ) );
  nor_x1_sg U62832 ( .A(n28459), .B(n55602), .X(\L1_0/n3811 ) );
  nor_x1_sg U62833 ( .A(n43906), .B(n28459), .X(\L1_0/n3810 ) );
  nor_x1_sg U62834 ( .A(n28459), .B(n28560), .X(\L1_0/n3807 ) );
  nor_x1_sg U62835 ( .A(n46596), .B(n29337), .X(\L1_0/n3603 ) );
  nor_x1_sg U62836 ( .A(n55775), .B(n46596), .X(\L1_0/n3602 ) );
  nor_x1_sg U62837 ( .A(n46596), .B(n55622), .X(\L1_0/n3599 ) );
  nor_x1_sg U62838 ( .A(n44479), .B(n46596), .X(\L1_0/n3598 ) );
  nor_x1_sg U62839 ( .A(n46596), .B(n29358), .X(\L1_0/n3591 ) );
  nor_x1_sg U62840 ( .A(n55776), .B(n46596), .X(\L1_0/n3590 ) );
  nor_x1_sg U62841 ( .A(n46596), .B(n29373), .X(\L1_0/n3583 ) );
  nor_x1_sg U62842 ( .A(n55777), .B(n46596), .X(\L1_0/n3582 ) );
  nor_x1_sg U62843 ( .A(n46596), .B(n55625), .X(\L1_0/n3579 ) );
  nor_x1_sg U62844 ( .A(n43900), .B(n46596), .X(\L1_0/n3578 ) );
  nor_x1_sg U62845 ( .A(n46596), .B(n29387), .X(\L1_0/n3575 ) );
  nor_x1_sg U62846 ( .A(n55778), .B(n46596), .X(\L1_0/n3574 ) );
  nor_x1_sg U62847 ( .A(n46596), .B(n55626), .X(\L1_0/n3571 ) );
  nor_x1_sg U62848 ( .A(n43815), .B(n46596), .X(\L1_0/n3570 ) );
  nor_x1_sg U62849 ( .A(n55730), .B(n46593), .X(\L1_0/n3942 ) );
  nor_x1_sg U62850 ( .A(n46593), .B(n28189), .X(\L1_0/n3939 ) );
  nor_x1_sg U62851 ( .A(n55731), .B(n46593), .X(\L1_0/n3938 ) );
  nor_x1_sg U62852 ( .A(n46593), .B(n28196), .X(\L1_0/n3935 ) );
  nor_x1_sg U62853 ( .A(n55732), .B(n46593), .X(\L1_0/n3934 ) );
  nor_x1_sg U62854 ( .A(n46593), .B(n28203), .X(\L1_0/n3931 ) );
  nor_x1_sg U62855 ( .A(n55733), .B(n46593), .X(\L1_0/n3930 ) );
  nor_x1_sg U62856 ( .A(n46593), .B(n28210), .X(\L1_0/n3927 ) );
  nor_x1_sg U62857 ( .A(n55734), .B(n46593), .X(\L1_0/n3926 ) );
  nand_x4_sg U62858 ( .A(n10914), .B(n10915), .X(n10912) );
  nand_x1_sg U62859 ( .A(n10917), .B(n10918), .X(n10914) );
  nand_x1_sg U62860 ( .A(n10916), .B(n51435), .X(n10915) );
  nand_x1_sg U62861 ( .A(n51435), .B(n46564), .X(n10918) );
  nor_x1_sg U62862 ( .A(n46573), .B(n9355), .X(\L2_0/n4144 ) );
  nor_x1_sg U62863 ( .A(n9355), .B(n9036), .X(\L2_0/n4136 ) );
  nor_x1_sg U62864 ( .A(n43953), .B(n9355), .X(\L2_0/n4132 ) );
  nor_x1_sg U62865 ( .A(n9355), .B(n9045), .X(\L2_0/n4128 ) );
  nor_x1_sg U62866 ( .A(n46589), .B(n27099), .X(\L1_0/n4243 ) );
  nor_x1_sg U62867 ( .A(n55695), .B(n46589), .X(\L1_0/n4242 ) );
  nor_x1_sg U62868 ( .A(n46589), .B(n27120), .X(\L1_0/n4231 ) );
  nor_x1_sg U62869 ( .A(n55696), .B(n46589), .X(\L1_0/n4230 ) );
  nor_x1_sg U62870 ( .A(n46589), .B(n55561), .X(\L1_0/n4227 ) );
  nor_x1_sg U62871 ( .A(n44233), .B(n46589), .X(\L1_0/n4226 ) );
  nor_x1_sg U62872 ( .A(n46589), .B(n27134), .X(\L1_0/n4223 ) );
  nor_x1_sg U62873 ( .A(n55697), .B(n46589), .X(\L1_0/n4222 ) );
  nor_x1_sg U62874 ( .A(n46589), .B(n55562), .X(\L1_0/n4219 ) );
  nor_x1_sg U62875 ( .A(n43827), .B(n46589), .X(\L1_0/n4218 ) );
  nor_x1_sg U62876 ( .A(n46589), .B(n27148), .X(\L1_0/n4215 ) );
  nor_x1_sg U62877 ( .A(n55698), .B(n46589), .X(\L1_0/n4214 ) );
  nor_x1_sg U62878 ( .A(n46589), .B(n55563), .X(\L1_0/n4211 ) );
  nor_x1_sg U62879 ( .A(n43918), .B(n46589), .X(\L1_0/n4210 ) );
  nor_x1_sg U62880 ( .A(n46593), .B(n28218), .X(\L1_0/n3923 ) );
  nor_x1_sg U62881 ( .A(n55735), .B(n46593), .X(\L1_0/n3922 ) );
  nor_x1_sg U62882 ( .A(n46593), .B(n55590), .X(\L1_0/n3919 ) );
  nor_x1_sg U62883 ( .A(n43912), .B(n46593), .X(\L1_0/n3918 ) );
  nor_x1_sg U62884 ( .A(n46593), .B(n55591), .X(\L1_0/n3915 ) );
  nor_x1_sg U62885 ( .A(n44485), .B(n46593), .X(\L1_0/n3914 ) );
  nor_x1_sg U62886 ( .A(n46593), .B(n28239), .X(\L1_0/n3911 ) );
  nor_x1_sg U62887 ( .A(n55736), .B(n46593), .X(\L1_0/n3910 ) );
  nor_x1_sg U62888 ( .A(n46593), .B(n55592), .X(\L1_0/n3907 ) );
  nor_x1_sg U62889 ( .A(n44483), .B(n46593), .X(\L1_0/n3906 ) );
  nor_x1_sg U62890 ( .A(n46593), .B(n28254), .X(\L1_0/n3903 ) );
  nor_x1_sg U62891 ( .A(n55737), .B(n46593), .X(\L1_0/n3902 ) );
  nor_x1_sg U62892 ( .A(n46593), .B(n55593), .X(\L1_0/n3899 ) );
  nor_x1_sg U62893 ( .A(n43910), .B(n46593), .X(\L1_0/n3898 ) );
  nor_x1_sg U62894 ( .A(n46593), .B(n28268), .X(\L1_0/n3895 ) );
  nor_x1_sg U62895 ( .A(n55738), .B(n46593), .X(\L1_0/n3894 ) );
  nor_x1_sg U62896 ( .A(n46593), .B(n55594), .X(\L1_0/n3891 ) );
  nor_x1_sg U62897 ( .A(n44227), .B(n46593), .X(\L1_0/n3890 ) );
  nand_x4_sg U62898 ( .A(n16373), .B(n16374), .X(n16371) );
  nand_x1_sg U62899 ( .A(n16376), .B(n16377), .X(n16373) );
  nand_x1_sg U62900 ( .A(n16375), .B(n53384), .X(n16374) );
  nand_x1_sg U62901 ( .A(n53384), .B(n46405), .X(n16377) );
  nor_x1_sg U62902 ( .A(n46616), .B(n29056), .X(\L1_0/n3683 ) );
  nor_x1_sg U62903 ( .A(n55765), .B(n46616), .X(\L1_0/n3682 ) );
  nor_x1_sg U62904 ( .A(n46616), .B(n29077), .X(\L1_0/n3671 ) );
  nor_x1_sg U62905 ( .A(n55766), .B(n46616), .X(\L1_0/n3670 ) );
  nor_x1_sg U62906 ( .A(n46616), .B(n55616), .X(\L1_0/n3667 ) );
  nor_x1_sg U62907 ( .A(n43904), .B(n46616), .X(\L1_0/n3666 ) );
  nor_x1_sg U62908 ( .A(n46616), .B(n29091), .X(\L1_0/n3663 ) );
  nor_x1_sg U62909 ( .A(n55767), .B(n46616), .X(\L1_0/n3662 ) );
  nor_x1_sg U62910 ( .A(n46616), .B(n55617), .X(\L1_0/n3659 ) );
  nor_x1_sg U62911 ( .A(n43902), .B(n46616), .X(\L1_0/n3658 ) );
  nor_x1_sg U62912 ( .A(n46616), .B(n29105), .X(\L1_0/n3655 ) );
  nor_x1_sg U62913 ( .A(n46615), .B(n25389), .X(\L1_0/n4743 ) );
  nor_x1_sg U62914 ( .A(n46615), .B(n55630), .X(\L1_0/n4742 ) );
  nor_x1_sg U62915 ( .A(n46615), .B(n25425), .X(\L1_0/n4723 ) );
  nor_x1_sg U62916 ( .A(n46615), .B(n55635), .X(\L1_0/n4722 ) );
  nor_x1_sg U62917 ( .A(n46615), .B(n55513), .X(\L1_0/n4719 ) );
  nor_x1_sg U62918 ( .A(n46615), .B(n44501), .X(\L1_0/n4718 ) );
  nor_x1_sg U62919 ( .A(n46615), .B(n25446), .X(\L1_0/n4711 ) );
  nor_x1_sg U62920 ( .A(n46615), .B(n55636), .X(\L1_0/n4710 ) );
  nor_x1_sg U62921 ( .A(n46615), .B(n25461), .X(\L1_0/n4703 ) );
  nor_x1_sg U62922 ( .A(n46615), .B(n55637), .X(\L1_0/n4702 ) );
  nor_x1_sg U62923 ( .A(n46615), .B(n25475), .X(\L1_0/n4695 ) );
  nor_x1_sg U62924 ( .A(n46615), .B(n55638), .X(\L1_0/n4694 ) );
  nor_x1_sg U62925 ( .A(n46615), .B(n55517), .X(\L1_0/n4691 ) );
  nor_x1_sg U62926 ( .A(n46615), .B(n43835), .X(\L1_0/n4690 ) );
  nor_x1_sg U62927 ( .A(n46615), .B(n25489), .X(\L1_0/n4687 ) );
  nor_x1_sg U62928 ( .A(n46615), .B(n55639), .X(\L1_0/n4686 ) );
  nor_x1_sg U62929 ( .A(n46615), .B(n25496), .X(\L1_0/n4683 ) );
  nor_x1_sg U62930 ( .A(n46615), .B(n55518), .X(\L1_0/n4682 ) );
  nor_x1_sg U62931 ( .A(n46615), .B(n25501), .X(\L1_0/n4679 ) );
  nor_x1_sg U62932 ( .A(n46615), .B(n55519), .X(\L1_0/n4678 ) );
  nor_x1_sg U62933 ( .A(n46612), .B(n25982), .X(\L1_0/n4563 ) );
  nor_x1_sg U62934 ( .A(n55655), .B(n46612), .X(\L1_0/n4562 ) );
  nor_x1_sg U62935 ( .A(n46612), .B(n55528), .X(\L1_0/n4559 ) );
  nor_x1_sg U62936 ( .A(n44497), .B(n46612), .X(\L1_0/n4558 ) );
  nor_x1_sg U62937 ( .A(n46612), .B(n26003), .X(\L1_0/n4551 ) );
  nor_x1_sg U62938 ( .A(n55656), .B(n46612), .X(\L1_0/n4550 ) );
  nor_x1_sg U62939 ( .A(n46612), .B(n55530), .X(\L1_0/n4547 ) );
  nor_x1_sg U62940 ( .A(n43930), .B(n46612), .X(\L1_0/n4546 ) );
  nor_x1_sg U62941 ( .A(n46612), .B(n26017), .X(\L1_0/n4543 ) );
  nor_x1_sg U62942 ( .A(n55657), .B(n46612), .X(\L1_0/n4542 ) );
  nor_x1_sg U62943 ( .A(n46612), .B(n55531), .X(\L1_0/n4539 ) );
  nor_x1_sg U62944 ( .A(n43833), .B(n46612), .X(\L1_0/n4538 ) );
  nor_x1_sg U62945 ( .A(n46612), .B(n26031), .X(\L1_0/n4535 ) );
  nor_x1_sg U62946 ( .A(n46625), .B(n26820), .X(\L1_0/n4323 ) );
  nor_x1_sg U62947 ( .A(n46625), .B(n55685), .X(\L1_0/n4322 ) );
  nor_x1_sg U62948 ( .A(n46625), .B(n55551), .X(\L1_0/n4319 ) );
  nor_x1_sg U62949 ( .A(n46625), .B(n43922), .X(\L1_0/n4318 ) );
  nor_x1_sg U62950 ( .A(n46625), .B(n26841), .X(\L1_0/n4311 ) );
  nor_x1_sg U62951 ( .A(n46625), .B(n55686), .X(\L1_0/n4310 ) );
  nor_x1_sg U62952 ( .A(n46625), .B(n55553), .X(\L1_0/n4307 ) );
  nor_x1_sg U62953 ( .A(n46625), .B(n44054), .X(\L1_0/n4306 ) );
  nor_x1_sg U62954 ( .A(n46625), .B(n26855), .X(\L1_0/n4303 ) );
  nor_x1_sg U62955 ( .A(n46625), .B(n55687), .X(\L1_0/n4302 ) );
  nor_x1_sg U62956 ( .A(n46625), .B(n55554), .X(\L1_0/n4299 ) );
  nor_x1_sg U62957 ( .A(n46625), .B(n43920), .X(\L1_0/n4298 ) );
  nor_x1_sg U62958 ( .A(n46625), .B(n26869), .X(\L1_0/n4295 ) );
  nor_x1_sg U62959 ( .A(n46625), .B(n55688), .X(\L1_0/n4294 ) );
  nor_x1_sg U62960 ( .A(n46611), .B(n25704), .X(\L1_0/n4643 ) );
  nor_x1_sg U62961 ( .A(n46611), .B(n55645), .X(\L1_0/n4642 ) );
  nor_x1_sg U62962 ( .A(n46611), .B(n25725), .X(\L1_0/n4631 ) );
  nor_x1_sg U62963 ( .A(n46611), .B(n55646), .X(\L1_0/n4630 ) );
  nor_x1_sg U62964 ( .A(n46611), .B(n55523), .X(\L1_0/n4627 ) );
  nor_x1_sg U62965 ( .A(n46611), .B(n43932), .X(\L1_0/n4626 ) );
  nor_x1_sg U62966 ( .A(n46611), .B(n25739), .X(\L1_0/n4623 ) );
  nor_x1_sg U62967 ( .A(n46611), .B(n55647), .X(\L1_0/n4622 ) );
  nor_x1_sg U62968 ( .A(n46611), .B(n55524), .X(\L1_0/n4619 ) );
  nor_x1_sg U62969 ( .A(n46611), .B(n44060), .X(\L1_0/n4618 ) );
  nor_x1_sg U62970 ( .A(n46611), .B(n25753), .X(\L1_0/n4615 ) );
  nor_x1_sg U62971 ( .A(n46611), .B(n55648), .X(\L1_0/n4614 ) );
  nor_x1_sg U62972 ( .A(n46623), .B(n27379), .X(\L1_0/n4163 ) );
  nor_x1_sg U62973 ( .A(n46623), .B(n55705), .X(\L1_0/n4162 ) );
  nor_x1_sg U62974 ( .A(n46623), .B(n55567), .X(\L1_0/n4159 ) );
  nor_x1_sg U62975 ( .A(n46623), .B(n44489), .X(\L1_0/n4158 ) );
  nor_x1_sg U62976 ( .A(n46623), .B(n27400), .X(\L1_0/n4151 ) );
  nor_x1_sg U62977 ( .A(n46623), .B(n55706), .X(\L1_0/n4150 ) );
  nor_x1_sg U62978 ( .A(n46623), .B(n55569), .X(\L1_0/n4147 ) );
  nor_x1_sg U62979 ( .A(n46623), .B(n43916), .X(\L1_0/n4146 ) );
  nor_x1_sg U62980 ( .A(n46623), .B(n27414), .X(\L1_0/n4143 ) );
  nor_x1_sg U62981 ( .A(n46623), .B(n55707), .X(\L1_0/n4142 ) );
  nor_x1_sg U62982 ( .A(n46623), .B(n55570), .X(\L1_0/n4139 ) );
  nor_x1_sg U62983 ( .A(n46623), .B(n43825), .X(\L1_0/n4138 ) );
  nor_x1_sg U62984 ( .A(n46623), .B(n27428), .X(\L1_0/n4135 ) );
  nor_x1_sg U62985 ( .A(n46623), .B(n55708), .X(\L1_0/n4134 ) );
  nor_x1_sg U62986 ( .A(n46621), .B(n27659), .X(\L1_0/n4083 ) );
  nor_x1_sg U62987 ( .A(n46621), .B(n55715), .X(\L1_0/n4082 ) );
  nor_x1_sg U62988 ( .A(n46621), .B(n27680), .X(\L1_0/n4071 ) );
  nor_x1_sg U62989 ( .A(n46621), .B(n55716), .X(\L1_0/n4070 ) );
  nor_x1_sg U62990 ( .A(n46621), .B(n55576), .X(\L1_0/n4067 ) );
  nor_x1_sg U62991 ( .A(n46621), .B(n44231), .X(\L1_0/n4066 ) );
  nor_x1_sg U62992 ( .A(n46621), .B(n27694), .X(\L1_0/n4063 ) );
  nor_x1_sg U62993 ( .A(n46621), .B(n55717), .X(\L1_0/n4062 ) );
  nor_x1_sg U62994 ( .A(n46621), .B(n55577), .X(\L1_0/n4059 ) );
  nor_x1_sg U62995 ( .A(n46621), .B(n43796), .X(\L1_0/n4058 ) );
  nor_x1_sg U62996 ( .A(n46621), .B(n27708), .X(\L1_0/n4055 ) );
  nor_x1_sg U62997 ( .A(n46621), .B(n55718), .X(\L1_0/n4054 ) );
  nor_x1_sg U62998 ( .A(n46619), .B(n28776), .X(\L1_0/n3763 ) );
  nor_x1_sg U62999 ( .A(n46619), .B(n55755), .X(\L1_0/n3762 ) );
  nor_x1_sg U63000 ( .A(n46619), .B(n55606), .X(\L1_0/n3759 ) );
  nor_x1_sg U63001 ( .A(n46619), .B(n44481), .X(\L1_0/n3758 ) );
  nor_x1_sg U63002 ( .A(n46619), .B(n28797), .X(\L1_0/n3751 ) );
  nor_x1_sg U63003 ( .A(n46619), .B(n55756), .X(\L1_0/n3750 ) );
  nor_x1_sg U63004 ( .A(n46619), .B(n28812), .X(\L1_0/n3743 ) );
  nor_x1_sg U63005 ( .A(n46619), .B(n55757), .X(\L1_0/n3742 ) );
  nor_x1_sg U63006 ( .A(n46619), .B(n55609), .X(\L1_0/n3739 ) );
  nor_x1_sg U63007 ( .A(n46619), .B(n44221), .X(\L1_0/n3738 ) );
  nor_x1_sg U63008 ( .A(n46619), .B(n28826), .X(\L1_0/n3735 ) );
  nor_x1_sg U63009 ( .A(n46619), .B(n55758), .X(\L1_0/n3734 ) );
  nor_x1_sg U63010 ( .A(n46585), .B(n26334), .X(\L1_0/n4443 ) );
  nor_x1_sg U63011 ( .A(n55540), .B(n46585), .X(\L1_0/n4442 ) );
  nor_x1_sg U63012 ( .A(n46585), .B(n26339), .X(\L1_0/n4439 ) );
  nor_x1_sg U63013 ( .A(n55541), .B(n46585), .X(\L1_0/n4438 ) );
  nor_x1_sg U63014 ( .A(n46587), .B(n26613), .X(\L1_0/n4363 ) );
  nor_x1_sg U63015 ( .A(n55548), .B(n46587), .X(\L1_0/n4362 ) );
  nor_x1_sg U63016 ( .A(n46587), .B(n26618), .X(\L1_0/n4359 ) );
  nor_x1_sg U63017 ( .A(n55549), .B(n46587), .X(\L1_0/n4358 ) );
  nor_x1_sg U63018 ( .A(n46591), .B(n28002), .X(\L1_0/n3967 ) );
  nor_x1_sg U63019 ( .A(n55729), .B(n46591), .X(\L1_0/n3966 ) );
  nor_x1_sg U63020 ( .A(n46591), .B(n28009), .X(\L1_0/n3963 ) );
  nor_x1_sg U63021 ( .A(n55587), .B(n46591), .X(\L1_0/n3962 ) );
  nor_x1_sg U63022 ( .A(n46591), .B(n28014), .X(\L1_0/n3959 ) );
  nor_x1_sg U63023 ( .A(n55588), .B(n46591), .X(\L1_0/n3958 ) );
  nor_x1_sg U63024 ( .A(n55749), .B(n28459), .X(\L1_0/n3806 ) );
  nor_x1_sg U63025 ( .A(n28459), .B(n28567), .X(\L1_0/n3803 ) );
  nor_x1_sg U63026 ( .A(n55603), .B(n28459), .X(\L1_0/n3802 ) );
  nor_x1_sg U63027 ( .A(n28459), .B(n28572), .X(\L1_0/n3799 ) );
  nor_x1_sg U63028 ( .A(n55604), .B(n28459), .X(\L1_0/n3798 ) );
  nor_x1_sg U63029 ( .A(n46596), .B(n29401), .X(\L1_0/n3567 ) );
  nor_x1_sg U63030 ( .A(n55779), .B(n46596), .X(\L1_0/n3566 ) );
  nor_x1_sg U63031 ( .A(n46596), .B(n29408), .X(\L1_0/n3563 ) );
  nor_x1_sg U63032 ( .A(n55627), .B(n46596), .X(\L1_0/n3562 ) );
  nor_x1_sg U63033 ( .A(n46596), .B(n29413), .X(\L1_0/n3559 ) );
  nor_x1_sg U63034 ( .A(n55628), .B(n46596), .X(\L1_0/n3558 ) );
  nor_x1_sg U63035 ( .A(n55768), .B(n46616), .X(\L1_0/n3654 ) );
  nor_x1_sg U63036 ( .A(n46616), .B(n55618), .X(\L1_0/n3651 ) );
  nor_x1_sg U63037 ( .A(n43817), .B(n46616), .X(\L1_0/n3650 ) );
  nor_x1_sg U63038 ( .A(n46616), .B(n29119), .X(\L1_0/n3647 ) );
  nor_x1_sg U63039 ( .A(n55769), .B(n46616), .X(\L1_0/n3646 ) );
  nor_x1_sg U63040 ( .A(n46616), .B(n29126), .X(\L1_0/n3643 ) );
  nor_x1_sg U63041 ( .A(n55619), .B(n46616), .X(\L1_0/n3642 ) );
  nor_x1_sg U63042 ( .A(n46616), .B(n29131), .X(\L1_0/n3639 ) );
  nor_x1_sg U63043 ( .A(n55620), .B(n46616), .X(\L1_0/n3638 ) );
  nor_x1_sg U63044 ( .A(n55658), .B(n46612), .X(\L1_0/n4534 ) );
  nor_x1_sg U63045 ( .A(n46612), .B(n41605), .X(\L1_0/n4531 ) );
  nor_x1_sg U63046 ( .A(n41606), .B(n46612), .X(\L1_0/n4530 ) );
  nor_x1_sg U63047 ( .A(n46612), .B(n26053), .X(\L1_0/n4523 ) );
  nor_x1_sg U63048 ( .A(n55532), .B(n46612), .X(\L1_0/n4522 ) );
  nor_x1_sg U63049 ( .A(n46612), .B(n26058), .X(\L1_0/n4519 ) );
  nor_x1_sg U63050 ( .A(n55533), .B(n46612), .X(\L1_0/n4518 ) );
  nor_x1_sg U63051 ( .A(n46625), .B(n55555), .X(\L1_0/n4291 ) );
  nor_x1_sg U63052 ( .A(n46625), .B(n43829), .X(\L1_0/n4290 ) );
  nor_x1_sg U63053 ( .A(n46625), .B(n26883), .X(\L1_0/n4287 ) );
  nor_x1_sg U63054 ( .A(n46625), .B(n55689), .X(\L1_0/n4286 ) );
  nor_x1_sg U63055 ( .A(n46625), .B(n26890), .X(\L1_0/n4283 ) );
  nor_x1_sg U63056 ( .A(n46625), .B(n55556), .X(\L1_0/n4282 ) );
  nor_x1_sg U63057 ( .A(n46625), .B(n26895), .X(\L1_0/n4279 ) );
  nor_x1_sg U63058 ( .A(n46625), .B(n55557), .X(\L1_0/n4278 ) );
  nor_x1_sg U63059 ( .A(n46611), .B(n41607), .X(\L1_0/n4611 ) );
  nor_x1_sg U63060 ( .A(n46611), .B(n41608), .X(\L1_0/n4610 ) );
  nor_x1_sg U63061 ( .A(n46611), .B(n25767), .X(\L1_0/n4607 ) );
  nor_x1_sg U63062 ( .A(n46611), .B(n55649), .X(\L1_0/n4606 ) );
  nor_x1_sg U63063 ( .A(n46611), .B(n25774), .X(\L1_0/n4603 ) );
  nor_x1_sg U63064 ( .A(n46611), .B(n55525), .X(\L1_0/n4602 ) );
  nor_x1_sg U63065 ( .A(n46611), .B(n25779), .X(\L1_0/n4599 ) );
  nor_x1_sg U63066 ( .A(n46611), .B(n55526), .X(\L1_0/n4598 ) );
  nor_x1_sg U63067 ( .A(n46623), .B(n41603), .X(\L1_0/n4131 ) );
  nor_x1_sg U63068 ( .A(n46623), .B(n41604), .X(\L1_0/n4130 ) );
  nor_x1_sg U63069 ( .A(n46623), .B(n27442), .X(\L1_0/n4127 ) );
  nor_x1_sg U63070 ( .A(n46623), .B(n55709), .X(\L1_0/n4126 ) );
  nor_x1_sg U63071 ( .A(n46623), .B(n27449), .X(\L1_0/n4123 ) );
  nor_x1_sg U63072 ( .A(n46623), .B(n55571), .X(\L1_0/n4122 ) );
  nor_x1_sg U63073 ( .A(n46623), .B(n27454), .X(\L1_0/n4119 ) );
  nor_x1_sg U63074 ( .A(n46623), .B(n55572), .X(\L1_0/n4118 ) );
  nor_x1_sg U63075 ( .A(n46621), .B(n55578), .X(\L1_0/n4051 ) );
  nor_x1_sg U63076 ( .A(n46621), .B(n43769), .X(\L1_0/n4050 ) );
  nor_x1_sg U63077 ( .A(n46621), .B(n27730), .X(\L1_0/n4043 ) );
  nor_x1_sg U63078 ( .A(n46621), .B(n55579), .X(\L1_0/n4042 ) );
  nor_x1_sg U63079 ( .A(n46621), .B(n27735), .X(\L1_0/n4039 ) );
  nor_x1_sg U63080 ( .A(n46621), .B(n55580), .X(\L1_0/n4038 ) );
  nor_x1_sg U63081 ( .A(n46619), .B(n55610), .X(\L1_0/n3731 ) );
  nor_x1_sg U63082 ( .A(n46619), .B(n44044), .X(\L1_0/n3730 ) );
  nor_x1_sg U63083 ( .A(n46619), .B(n28840), .X(\L1_0/n3727 ) );
  nor_x1_sg U63084 ( .A(n46619), .B(n55759), .X(\L1_0/n3726 ) );
  nor_x1_sg U63085 ( .A(n46619), .B(n28847), .X(\L1_0/n3723 ) );
  nor_x1_sg U63086 ( .A(n46619), .B(n55611), .X(\L1_0/n3722 ) );
  nor_x1_sg U63087 ( .A(n46619), .B(n28852), .X(\L1_0/n3719 ) );
  nor_x1_sg U63088 ( .A(n46619), .B(n55612), .X(\L1_0/n3718 ) );
  nand_x4_sg U63089 ( .A(n11046), .B(n11047), .X(n10879) );
  nand_x1_sg U63090 ( .A(n11048), .B(n51498), .X(n11047) );
  nand_x1_sg U63091 ( .A(n10899), .B(n51476), .X(n11046) );
  nor_x1_sg U63092 ( .A(n11973), .B(n46519), .X(n11972) );
  nand_x2_sg U63093 ( .A(n15867), .B(n46405), .X(n15866) );
  nand_x2_sg U63094 ( .A(n15868), .B(n15869), .X(n15865) );
  nor_x1_sg U63095 ( .A(n15868), .B(n46407), .X(n15867) );
  nor_x1_sg U63096 ( .A(n46589), .B(n27162), .X(\L1_0/n4207 ) );
  nor_x1_sg U63097 ( .A(n55699), .B(n46589), .X(\L1_0/n4206 ) );
  nor_x1_sg U63098 ( .A(n46589), .B(n27170), .X(\L1_0/n4203 ) );
  nor_x1_sg U63099 ( .A(n55564), .B(n46589), .X(\L1_0/n4202 ) );
  nor_x1_sg U63100 ( .A(n46589), .B(n27175), .X(\L1_0/n4199 ) );
  nor_x1_sg U63101 ( .A(n55565), .B(n46589), .X(\L1_0/n4198 ) );
  nand_x4_sg U63102 ( .A(n10730), .B(n10731), .X(n10667) );
  nand_x1_sg U63103 ( .A(n10664), .B(n51398), .X(n10730) );
  nand_x1_sg U63104 ( .A(n10732), .B(n10696), .X(n10731) );
  nand_x4_sg U63105 ( .A(n18512), .B(n18513), .X(n18449) );
  nand_x1_sg U63106 ( .A(n18446), .B(n54187), .X(n18512) );
  nand_x1_sg U63107 ( .A(n54185), .B(n18478), .X(n18513) );
  nand_x4_sg U63108 ( .A(n20057), .B(n20058), .X(n19994) );
  nand_x1_sg U63109 ( .A(n19991), .B(n54754), .X(n20057) );
  nand_x1_sg U63110 ( .A(n54752), .B(n20023), .X(n20058) );
  nand_x4_sg U63111 ( .A(n21602), .B(n21603), .X(n21539) );
  nand_x1_sg U63112 ( .A(n21536), .B(n55322), .X(n21602) );
  nand_x1_sg U63113 ( .A(n55320), .B(n21568), .X(n21603) );
  nor_x1_sg U63114 ( .A(n29020), .B(n46616), .X(\L1_0/n3706 ) );
  nor_x1_sg U63115 ( .A(n46616), .B(n29021), .X(\L1_0/n3703 ) );
  nor_x1_sg U63116 ( .A(n55760), .B(n46616), .X(\L1_0/n3702 ) );
  nor_x1_sg U63117 ( .A(n25946), .B(n46612), .X(\L1_0/n4586 ) );
  nor_x1_sg U63118 ( .A(n46612), .B(n25947), .X(\L1_0/n4583 ) );
  nor_x1_sg U63119 ( .A(n55650), .B(n46612), .X(\L1_0/n4582 ) );
  nor_x1_sg U63120 ( .A(n46611), .B(n25668), .X(\L1_0/n4666 ) );
  nor_x1_sg U63121 ( .A(n46611), .B(n25669), .X(\L1_0/n4663 ) );
  nor_x1_sg U63122 ( .A(n46611), .B(n55640), .X(\L1_0/n4662 ) );
  nor_x1_sg U63123 ( .A(n46625), .B(n26784), .X(\L1_0/n4346 ) );
  nor_x1_sg U63124 ( .A(n46625), .B(n26785), .X(\L1_0/n4343 ) );
  nor_x1_sg U63125 ( .A(n46625), .B(n55680), .X(\L1_0/n4342 ) );
  nor_x1_sg U63126 ( .A(n46623), .B(n27343), .X(\L1_0/n4186 ) );
  nor_x1_sg U63127 ( .A(n46623), .B(n27344), .X(\L1_0/n4183 ) );
  nor_x1_sg U63128 ( .A(n46623), .B(n55700), .X(\L1_0/n4182 ) );
  nor_x1_sg U63129 ( .A(n46621), .B(n27623), .X(\L1_0/n4106 ) );
  nor_x1_sg U63130 ( .A(n46621), .B(n27624), .X(\L1_0/n4103 ) );
  nor_x1_sg U63131 ( .A(n46621), .B(n55710), .X(\L1_0/n4102 ) );
  nor_x1_sg U63132 ( .A(n46619), .B(n28740), .X(\L1_0/n3786 ) );
  nor_x1_sg U63133 ( .A(n46619), .B(n28741), .X(\L1_0/n3783 ) );
  nor_x1_sg U63134 ( .A(n46619), .B(n55750), .X(\L1_0/n3782 ) );
  nor_x1_sg U63135 ( .A(n13534), .B(n46480), .X(n13533) );
  nand_x4_sg U63136 ( .A(n16185), .B(n16186), .X(n16122) );
  nand_x1_sg U63137 ( .A(n16117), .B(n16119), .X(n16185) );
  nand_x1_sg U63138 ( .A(n16187), .B(n16152), .X(n16186) );
  nand_x4_sg U63139 ( .A(n46367), .B(n46373), .X(n27915) );
  nand_x4_sg U63140 ( .A(n46320), .B(n46326), .X(n28473) );
  nand_x4_sg U63141 ( .A(n46275), .B(n46281), .X(n29032) );
  nand_x4_sg U63142 ( .A(n51478), .B(n10976), .X(n10936) );
  nand_x4_sg U63143 ( .A(n53427), .B(n16434), .X(n16394) );
  nand_x4_sg U63144 ( .A(n53987), .B(n17993), .X(n17952) );
  nand_x4_sg U63145 ( .A(n54552), .B(n19538), .X(n19497) );
  nand_x4_sg U63146 ( .A(n55120), .B(n21082), .X(n21041) );
  nand_x4_sg U63147 ( .A(n14788), .B(n14789), .X(n14786) );
  nand_x1_sg U63148 ( .A(n14790), .B(n14791), .X(n14789) );
  nand_x1_sg U63149 ( .A(n14794), .B(n52783), .X(n14788) );
  nor_x1_sg U63150 ( .A(n14792), .B(n14793), .X(n14790) );
  nand_x4_sg U63151 ( .A(n20246), .B(n20247), .X(n20245) );
  nand_x1_sg U63152 ( .A(n20249), .B(n20250), .X(n20246) );
  nand_x1_sg U63153 ( .A(n20248), .B(n54794), .X(n20247) );
  nand_x1_sg U63154 ( .A(n54794), .B(n46294), .X(n20250) );
  nand_x4_sg U63155 ( .A(n21791), .B(n21792), .X(n21790) );
  nand_x1_sg U63156 ( .A(n21794), .B(n21795), .X(n21791) );
  nand_x1_sg U63157 ( .A(n21793), .B(n55362), .X(n21792) );
  nand_x1_sg U63158 ( .A(n55362), .B(n46249), .X(n21795) );
  nand_x4_sg U63159 ( .A(n11510), .B(n11511), .X(n11447) );
  nand_x1_sg U63160 ( .A(n11442), .B(n11444), .X(n11510) );
  nand_x1_sg U63161 ( .A(n11512), .B(n11477), .X(n11511) );
  nand_x4_sg U63162 ( .A(n13071), .B(n13072), .X(n13008) );
  nand_x1_sg U63163 ( .A(n13003), .B(n13005), .X(n13071) );
  nand_x1_sg U63164 ( .A(n13073), .B(n13038), .X(n13072) );
  nand_x4_sg U63165 ( .A(n15404), .B(n15405), .X(n15341) );
  nand_x1_sg U63166 ( .A(n15336), .B(n15338), .X(n15404) );
  nand_x1_sg U63167 ( .A(n15406), .B(n15371), .X(n15405) );
  nand_x4_sg U63168 ( .A(n16970), .B(n16971), .X(n16907) );
  nand_x1_sg U63169 ( .A(n16902), .B(n16904), .X(n16970) );
  nand_x1_sg U63170 ( .A(n16972), .B(n16937), .X(n16971) );
  nor_x1_sg U63171 ( .A(n14559), .B(n14560), .X(n14558) );
  nor_x1_sg U63172 ( .A(n17680), .B(n17681), .X(n17679) );
  nor_x1_sg U63173 ( .A(n19225), .B(n19226), .X(n19224) );
  nor_x1_sg U63174 ( .A(n20769), .B(n20770), .X(n20768) );
  nor_x1_sg U63175 ( .A(n13788), .B(n13789), .X(n13787) );
  nand_x4_sg U63176 ( .A(n12290), .B(n12291), .X(n12227) );
  nand_x1_sg U63177 ( .A(n12222), .B(n12224), .X(n12290) );
  nand_x1_sg U63178 ( .A(n12292), .B(n12257), .X(n12291) );
  nand_x4_sg U63179 ( .A(n10483), .B(n10484), .X(n10472) );
  nor_x1_sg U63180 ( .A(n10485), .B(n46566), .X(n10484) );
  nor_x1_sg U63181 ( .A(n10493), .B(n51300), .X(n10483) );
  nand_x2_sg U63182 ( .A(n52697), .B(n14537), .X(n14550) );
  nand_x2_sg U63183 ( .A(n52709), .B(n14538), .X(n14551) );
  nand_x2_sg U63184 ( .A(n53824), .B(n17658), .X(n17671) );
  nand_x2_sg U63185 ( .A(n53836), .B(n17659), .X(n17672) );
  nand_x2_sg U63186 ( .A(n54389), .B(n19203), .X(n19216) );
  nand_x2_sg U63187 ( .A(n54401), .B(n19204), .X(n19217) );
  nand_x2_sg U63188 ( .A(n54957), .B(n20747), .X(n20760) );
  nand_x2_sg U63189 ( .A(n54969), .B(n20748), .X(n20761) );
  nand_x4_sg U63190 ( .A(n14404), .B(n14405), .X(n14372) );
  nand_x1_sg U63191 ( .A(n14310), .B(n14407), .X(n14404) );
  nor_x1_sg U63192 ( .A(n14310), .B(n46452), .X(n14406) );
  nand_x4_sg U63193 ( .A(n13237), .B(n13238), .X(n13235) );
  nand_x1_sg U63194 ( .A(n13239), .B(n52313), .X(n13238) );
  nand_x1_sg U63195 ( .A(n13241), .B(n52227), .X(n13237) );
  nor_x1_sg U63196 ( .A(n13240), .B(n52334), .X(n13239) );
  nand_x4_sg U63197 ( .A(n14017), .B(n14018), .X(n14015) );
  nand_x1_sg U63198 ( .A(n14019), .B(n52588), .X(n14018) );
  nand_x1_sg U63199 ( .A(n14021), .B(n52504), .X(n14017) );
  nor_x1_sg U63200 ( .A(n14020), .B(n52609), .X(n14019) );
  nand_x4_sg U63201 ( .A(n15570), .B(n15571), .X(n15568) );
  nand_x1_sg U63202 ( .A(n15572), .B(n53147), .X(n15571) );
  nand_x1_sg U63203 ( .A(n15574), .B(n53061), .X(n15570) );
  nor_x1_sg U63204 ( .A(n15573), .B(n53168), .X(n15572) );
  nand_x4_sg U63205 ( .A(n17136), .B(n17137), .X(n17134) );
  nand_x1_sg U63206 ( .A(n17138), .B(n53705), .X(n17137) );
  nand_x1_sg U63207 ( .A(n17140), .B(n53619), .X(n17136) );
  nor_x1_sg U63208 ( .A(n17139), .B(n53726), .X(n17138) );
  nand_x4_sg U63209 ( .A(n19810), .B(n19811), .X(n19799) );
  nor_x1_sg U63210 ( .A(n19812), .B(n46300), .X(n19811) );
  nor_x1_sg U63211 ( .A(n19820), .B(n54654), .X(n19810) );
  nand_x4_sg U63212 ( .A(n21355), .B(n21356), .X(n21344) );
  nor_x1_sg U63213 ( .A(n21357), .B(n46255), .X(n21356) );
  nor_x1_sg U63214 ( .A(n21365), .B(n55222), .X(n21355) );
  nand_x4_sg U63215 ( .A(n15966), .B(n15967), .X(n15928) );
  nand_x1_sg U63216 ( .A(n15864), .B(n15969), .X(n15966) );
  nor_x1_sg U63217 ( .A(n15864), .B(n46407), .X(n15968) );
  nand_x4_sg U63218 ( .A(n13911), .B(n13912), .X(n13823) );
  nand_x1_sg U63219 ( .A(n13914), .B(n13915), .X(n13911) );
  nor_x1_sg U63220 ( .A(n52863), .B(n14921), .X(n14919) );
  nor_x1_sg U63221 ( .A(n53983), .B(n18042), .X(n18040) );
  nor_x1_sg U63222 ( .A(n54548), .B(n19587), .X(n19585) );
  nor_x1_sg U63223 ( .A(n55116), .B(n21131), .X(n21129) );
  nor_x1_sg U63224 ( .A(n11415), .B(n11416), .X(n11413) );
  nor_x1_sg U63225 ( .A(n12976), .B(n12977), .X(n12974) );
  nor_x1_sg U63226 ( .A(n15309), .B(n15310), .X(n15307) );
  nor_x1_sg U63227 ( .A(n16875), .B(n16876), .X(n16873) );
  nand_x2_sg U63228 ( .A(n54106), .B(n18427), .X(n18440) );
  nand_x2_sg U63229 ( .A(n54110), .B(n18428), .X(n18441) );
  nand_x2_sg U63230 ( .A(n46517), .B(n25972), .X(n25971) );
  nand_x4_sg U63231 ( .A(n16271), .B(n16309), .X(n16307) );
  nand_x4_sg U63232 ( .A(n16204), .B(n53377), .X(n16202) );
  nand_x1_sg U63233 ( .A(n16206), .B(n53310), .X(n16204) );
  nor_x1_sg U63234 ( .A(n53310), .B(n16206), .X(n16205) );
  nand_x1_sg U63235 ( .A(n14635), .B(n52795), .X(n14632) );
  nand_x1_sg U63236 ( .A(n14634), .B(n52778), .X(n14633) );
  nand_x1_sg U63237 ( .A(n51339), .B(n10951), .X(n11040) );
  nand_x4_sg U63238 ( .A(n16497), .B(n16498), .X(n16419) );
  nand_x1_sg U63239 ( .A(n53452), .B(n43172), .X(n16497) );
  nand_x1_sg U63240 ( .A(n16409), .B(n53287), .X(n16498) );
  nand_x4_sg U63241 ( .A(n12376), .B(n12414), .X(n12412) );
  nand_x1_sg U63242 ( .A(n18523), .B(n54178), .X(n18522) );
  nand_x1_sg U63243 ( .A(n18524), .B(n54199), .X(n18521) );
  nand_x1_sg U63244 ( .A(n12303), .B(n51964), .X(n12300) );
  nand_x1_sg U63245 ( .A(n12302), .B(n51947), .X(n12301) );
  nand_x1_sg U63246 ( .A(n13083), .B(n52222), .X(n13082) );
  nand_x1_sg U63247 ( .A(n13084), .B(n52239), .X(n13081) );
  nand_x1_sg U63248 ( .A(n13863), .B(n52499), .X(n13862) );
  nand_x1_sg U63249 ( .A(n13864), .B(n52516), .X(n13861) );
  nand_x1_sg U63250 ( .A(n15416), .B(n53056), .X(n15415) );
  nand_x1_sg U63251 ( .A(n15417), .B(n53073), .X(n15414) );
  nand_x1_sg U63252 ( .A(n16982), .B(n53614), .X(n16981) );
  nand_x1_sg U63253 ( .A(n16983), .B(n53631), .X(n16980) );
  nor_x1_sg U63254 ( .A(n17888), .B(n17889), .X(n17887) );
  nor_x1_sg U63255 ( .A(n19433), .B(n19434), .X(n19432) );
  nor_x1_sg U63256 ( .A(n20977), .B(n20978), .X(n20976) );
  nand_x4_sg U63257 ( .A(n10829), .B(n10830), .X(n10757) );
  nand_x1_sg U63258 ( .A(n51393), .B(n10831), .X(n10830) );
  nand_x1_sg U63259 ( .A(n10832), .B(n51413), .X(n10829) );
  nand_x4_sg U63260 ( .A(n14810), .B(n14811), .X(n14809) );
  nand_x1_sg U63261 ( .A(n14813), .B(n14814), .X(n14810) );
  nand_x1_sg U63262 ( .A(n14812), .B(n52824), .X(n14811) );
  nand_x1_sg U63263 ( .A(n52824), .B(n46450), .X(n14814) );
  nand_x4_sg U63264 ( .A(n17931), .B(n17932), .X(n17930) );
  nand_x1_sg U63265 ( .A(n17934), .B(n17935), .X(n17931) );
  nand_x1_sg U63266 ( .A(n17933), .B(n53944), .X(n17932) );
  nand_x1_sg U63267 ( .A(n53944), .B(n46361), .X(n17935) );
  nand_x4_sg U63268 ( .A(n19476), .B(n19477), .X(n19475) );
  nand_x1_sg U63269 ( .A(n19479), .B(n19480), .X(n19476) );
  nand_x1_sg U63270 ( .A(n19478), .B(n54509), .X(n19477) );
  nand_x1_sg U63271 ( .A(n54509), .B(n46314), .X(n19480) );
  nand_x4_sg U63272 ( .A(n21020), .B(n21021), .X(n21019) );
  nand_x1_sg U63273 ( .A(n21023), .B(n21024), .X(n21020) );
  nand_x1_sg U63274 ( .A(n21022), .B(n55077), .X(n21021) );
  nand_x1_sg U63275 ( .A(n55077), .B(n46269), .X(n21024) );
  nor_x1_sg U63276 ( .A(n14767), .B(n14768), .X(n14766) );
  nor_x1_sg U63277 ( .A(n44668), .B(n20358), .X(n20355) );
  nor_x1_sg U63278 ( .A(n44667), .B(n21903), .X(n21900) );
  nand_x4_sg U63279 ( .A(n18355), .B(n18356), .X(n18304) );
  nand_x1_sg U63280 ( .A(n54077), .B(n18320), .X(n18356) );
  nand_x1_sg U63281 ( .A(n54091), .B(n18319), .X(n18355) );
  nand_x4_sg U63282 ( .A(n10516), .B(n51324), .X(n10481) );
  nand_x1_sg U63283 ( .A(n10511), .B(n51300), .X(n10516) );
  nor_x1_sg U63284 ( .A(n51300), .B(n10511), .X(n10517) );
  nand_x4_sg U63285 ( .A(n19843), .B(n54678), .X(n19808) );
  nand_x1_sg U63286 ( .A(n19838), .B(n54654), .X(n19843) );
  nor_x1_sg U63287 ( .A(n54654), .B(n19838), .X(n19844) );
  nand_x4_sg U63288 ( .A(n21388), .B(n55246), .X(n21353) );
  nand_x1_sg U63289 ( .A(n21383), .B(n55222), .X(n21388) );
  nor_x1_sg U63290 ( .A(n55222), .B(n21383), .X(n21389) );
  nand_x4_sg U63291 ( .A(n11595), .B(n11633), .X(n11631) );
  nand_x4_sg U63292 ( .A(n53343), .B(n16188), .X(n16119) );
  nand_x1_sg U63293 ( .A(n16152), .B(n53342), .X(n16188) );
  nor_x1_sg U63294 ( .A(n53342), .B(n16152), .X(n16189) );
  nor_x1_sg U63295 ( .A(n46573), .B(n24473), .X(\L1_0/n4747 ) );
  nand_x4_sg U63296 ( .A(n53780), .B(n17409), .X(n17308) );
  nand_x1_sg U63297 ( .A(n17401), .B(n17410), .X(n17409) );
  nor_x1_sg U63298 ( .A(n17410), .B(n17401), .X(n17411) );
  nand_x4_sg U63299 ( .A(n54345), .B(n18954), .X(n18853) );
  nand_x1_sg U63300 ( .A(n18946), .B(n18955), .X(n18954) );
  nor_x1_sg U63301 ( .A(n18955), .B(n18946), .X(n18956) );
  nand_x4_sg U63302 ( .A(n54913), .B(n20498), .X(n20397) );
  nand_x1_sg U63303 ( .A(n20490), .B(n20499), .X(n20498) );
  nor_x1_sg U63304 ( .A(n20499), .B(n20490), .X(n20500) );
  nand_x4_sg U63305 ( .A(n11660), .B(n11822), .X(n11747) );
  nand_x1_sg U63306 ( .A(n11735), .B(n51620), .X(n11822) );
  nand_x4_sg U63307 ( .A(n12597), .B(n12598), .X(n12527) );
  nand_x1_sg U63308 ( .A(n52064), .B(n40526), .X(n12597) );
  nand_x1_sg U63309 ( .A(n12515), .B(n51902), .X(n12598) );
  nand_x4_sg U63310 ( .A(n13379), .B(n13380), .X(n13308) );
  nand_x1_sg U63311 ( .A(n52341), .B(n40527), .X(n13379) );
  nand_x1_sg U63312 ( .A(n13296), .B(n52179), .X(n13380) );
  nand_x4_sg U63313 ( .A(n14159), .B(n14160), .X(n14088) );
  nand_x1_sg U63314 ( .A(n52616), .B(n40528), .X(n14159) );
  nand_x1_sg U63315 ( .A(n14076), .B(n52454), .X(n14160) );
  nand_x4_sg U63316 ( .A(n14770), .B(n14934), .X(n14859) );
  nand_x1_sg U63317 ( .A(n14847), .B(n52729), .X(n14934) );
  nand_x4_sg U63318 ( .A(n15712), .B(n15713), .X(n15641) );
  nand_x1_sg U63319 ( .A(n53175), .B(n40529), .X(n15712) );
  nand_x1_sg U63320 ( .A(n15629), .B(n53013), .X(n15713) );
  nand_x4_sg U63321 ( .A(n17278), .B(n17279), .X(n17207) );
  nand_x1_sg U63322 ( .A(n53733), .B(n40530), .X(n17278) );
  nand_x1_sg U63323 ( .A(n17195), .B(n53571), .X(n17279) );
  nand_x4_sg U63324 ( .A(n17891), .B(n18055), .X(n17980) );
  nand_x1_sg U63325 ( .A(n17968), .B(n53849), .X(n18055) );
  nand_x4_sg U63326 ( .A(n18660), .B(n18827), .X(n18749) );
  nand_x1_sg U63327 ( .A(n18737), .B(n54130), .X(n18827) );
  nand_x4_sg U63328 ( .A(n19436), .B(n19600), .X(n19525) );
  nand_x1_sg U63329 ( .A(n19513), .B(n54414), .X(n19600) );
  nand_x4_sg U63330 ( .A(n20205), .B(n20372), .X(n20295) );
  nand_x1_sg U63331 ( .A(n20283), .B(n54693), .X(n20372) );
  nand_x4_sg U63332 ( .A(n20980), .B(n21144), .X(n21069) );
  nand_x1_sg U63333 ( .A(n21057), .B(n54982), .X(n21144) );
  nand_x4_sg U63334 ( .A(n21750), .B(n21917), .X(n21840) );
  nand_x1_sg U63335 ( .A(n21828), .B(n55261), .X(n21917) );
  nand_x4_sg U63336 ( .A(n52465), .B(n13653), .X(n13644) );
  nand_x1_sg U63337 ( .A(n44074), .B(n13655), .X(n13653) );
  nand_x4_sg U63338 ( .A(n42370), .B(n18322), .X(n18308) );
  nand_x1_sg U63339 ( .A(n43223), .B(n41794), .X(n18322) );
  nand_x4_sg U63340 ( .A(n10532), .B(n10568), .X(n10567) );
  nand_x1_sg U63341 ( .A(n10569), .B(n10570), .X(n10568) );
  nand_x4_sg U63342 ( .A(n43248), .B(n14432), .X(n14418) );
  nand_x1_sg U63343 ( .A(n42365), .B(n41802), .X(n14432) );
  nor_x1_sg U63344 ( .A(n46281), .B(n46278), .X(\L2_0/n3104 ) );
  nor_x1_sg U63345 ( .A(n46278), .B(n9163), .X(\L2_0/n3088 ) );
  nor_x1_sg U63346 ( .A(n46552), .B(n46549), .X(\L2_0/n4064 ) );
  nor_x1_sg U63347 ( .A(n46549), .B(n8897), .X(\L2_0/n4048 ) );
  nor_x1_sg U63348 ( .A(n46508), .B(n46505), .X(\L2_0/n3904 ) );
  nor_x1_sg U63349 ( .A(n46505), .B(n8846), .X(\L2_0/n3888 ) );
  nor_x1_sg U63350 ( .A(n46463), .B(n46460), .X(\L2_0/n3744 ) );
  nor_x1_sg U63351 ( .A(n46460), .B(n9011), .X(\L2_0/n3728 ) );
  nor_x1_sg U63352 ( .A(n46416), .B(n46415), .X(\L2_0/n3584 ) );
  nor_x1_sg U63353 ( .A(n46415), .B(n9326), .X(\L2_0/n3568 ) );
  nor_x1_sg U63354 ( .A(n46373), .B(n46370), .X(\L2_0/n3424 ) );
  nor_x1_sg U63355 ( .A(n46370), .B(n9277), .X(\L2_0/n3408 ) );
  nor_x1_sg U63356 ( .A(n46326), .B(n46323), .X(\L2_0/n3264 ) );
  nor_x1_sg U63357 ( .A(n46323), .B(n9239), .X(\L2_0/n3248 ) );
  nor_x1_sg U63358 ( .A(n46528), .B(n46527), .X(\L2_0/n3984 ) );
  nor_x1_sg U63359 ( .A(n46527), .B(n8931), .X(\L2_0/n3968 ) );
  nor_x1_sg U63360 ( .A(n46306), .B(n46303), .X(\L2_0/n3184 ) );
  nor_x1_sg U63361 ( .A(n46303), .B(n9181), .X(\L2_0/n3168 ) );
  nor_x1_sg U63362 ( .A(n46303), .B(n9177), .X(\L2_0/n3156 ) );
  nor_x1_sg U63363 ( .A(n41970), .B(n46303), .X(\L2_0/n3144 ) );
  nor_x1_sg U63364 ( .A(n46303), .B(n9187), .X(\L2_0/n3132 ) );
  nor_x1_sg U63365 ( .A(n44391), .B(n46303), .X(\L2_0/n3120 ) );
  nor_x1_sg U63366 ( .A(n46303), .B(n9179), .X(\L2_0/n3108 ) );
  nor_x1_sg U63367 ( .A(n46440), .B(n46437), .X(\L2_0/n3664 ) );
  nor_x1_sg U63368 ( .A(n46437), .B(n8988), .X(\L2_0/n3648 ) );
  nor_x1_sg U63369 ( .A(n46353), .B(n46350), .X(\L2_0/n3344 ) );
  nor_x1_sg U63370 ( .A(n46350), .B(n9071), .X(\L2_0/n3328 ) );
  nor_x1_sg U63371 ( .A(n46350), .B(n9085), .X(\L2_0/n3316 ) );
  nor_x1_sg U63372 ( .A(n44108), .B(n46350), .X(\L2_0/n3304 ) );
  nor_x1_sg U63373 ( .A(n46350), .B(n9073), .X(\L2_0/n3292 ) );
  nor_x1_sg U63374 ( .A(n44395), .B(n46350), .X(\L2_0/n3280 ) );
  nor_x1_sg U63375 ( .A(n46350), .B(n9087), .X(\L2_0/n3268 ) );
  nor_x1_sg U63376 ( .A(n46483), .B(n8805), .X(\L2_0/n3808 ) );
  nor_x1_sg U63377 ( .A(n46396), .B(n46393), .X(\L2_0/n3504 ) );
  nor_x1_sg U63378 ( .A(n46393), .B(n9313), .X(\L2_0/n3488 ) );
  nor_x1_sg U63379 ( .A(n46261), .B(n46258), .X(\L2_0/n3024 ) );
  nor_x1_sg U63380 ( .A(n46258), .B(n9101), .X(\L2_0/n3008 ) );
  nand_x4_sg U63381 ( .A(n42368), .B(n10539), .X(n10526) );
  nand_x1_sg U63382 ( .A(n43221), .B(n41788), .X(n10539) );
  nand_x4_sg U63383 ( .A(n43234), .B(n19866), .X(n19853) );
  nand_x1_sg U63384 ( .A(n42357), .B(n41792), .X(n19866) );
  nand_x4_sg U63385 ( .A(n43232), .B(n21411), .X(n21398) );
  nand_x1_sg U63386 ( .A(n42355), .B(n41790), .X(n21411) );
  nand_x4_sg U63387 ( .A(n51913), .B(n12092), .X(n12083) );
  nand_x1_sg U63388 ( .A(n12093), .B(n12094), .X(n12092) );
  nand_x4_sg U63389 ( .A(n53300), .B(n15987), .X(n15978) );
  nand_x1_sg U63390 ( .A(n15988), .B(n15989), .X(n15987) );
  nand_x2_sg U63391 ( .A(n46296), .B(n28759), .X(n28758) );
  nand_x2_sg U63392 ( .A(n46251), .B(n29320), .X(n29319) );
  nand_x4_sg U63393 ( .A(n53781), .B(n17306), .X(n9242) );
  nand_x1_sg U63394 ( .A(n17307), .B(n17308), .X(n17306) );
  nand_x4_sg U63395 ( .A(n54346), .B(n18851), .X(n9204) );
  nand_x1_sg U63396 ( .A(n18852), .B(n18853), .X(n18851) );
  nand_x4_sg U63397 ( .A(n54914), .B(n20395), .X(n9128) );
  nand_x1_sg U63398 ( .A(n20396), .B(n20397), .X(n20395) );
  nand_x4_sg U63399 ( .A(n51674), .B(n11513), .X(n11444) );
  nand_x1_sg U63400 ( .A(n11477), .B(n51673), .X(n11513) );
  nor_x1_sg U63401 ( .A(n51673), .B(n11477), .X(n11514) );
  nand_x4_sg U63402 ( .A(n52230), .B(n13074), .X(n13005) );
  nand_x1_sg U63403 ( .A(n13038), .B(n52229), .X(n13074) );
  nor_x1_sg U63404 ( .A(n52229), .B(n13038), .X(n13075) );
  nand_x4_sg U63405 ( .A(n53064), .B(n15407), .X(n15338) );
  nand_x1_sg U63406 ( .A(n15371), .B(n53063), .X(n15407) );
  nor_x1_sg U63407 ( .A(n53063), .B(n15371), .X(n15408) );
  nand_x4_sg U63408 ( .A(n53622), .B(n16973), .X(n16904) );
  nand_x1_sg U63409 ( .A(n16937), .B(n53621), .X(n16973) );
  nor_x1_sg U63410 ( .A(n53621), .B(n16937), .X(n16974) );
  nand_x4_sg U63411 ( .A(n51955), .B(n12293), .X(n12224) );
  nand_x1_sg U63412 ( .A(n12257), .B(n51954), .X(n12293) );
  nor_x1_sg U63413 ( .A(n51954), .B(n12257), .X(n12294) );
  nand_x4_sg U63414 ( .A(n25397), .B(n25398), .X(n25396) );
  nor_x1_sg U63415 ( .A(n51263), .B(n25399), .X(n25398) );
  nor_x1_sg U63416 ( .A(n25402), .B(n46236), .X(n25397) );
  nand_x4_sg U63417 ( .A(n11676), .B(n11677), .X(n11674) );
  nand_x1_sg U63418 ( .A(n11678), .B(n11679), .X(n11677) );
  nand_x1_sg U63419 ( .A(n11682), .B(n51671), .X(n11676) );
  nor_x1_sg U63420 ( .A(n11680), .B(n11681), .X(n11678) );
  nand_x4_sg U63421 ( .A(n52537), .B(n13828), .X(n13805) );
  nand_x1_sg U63422 ( .A(n41846), .B(n13830), .X(n13828) );
  nor_x1_sg U63423 ( .A(n13830), .B(n41846), .X(n13831) );
  nand_x4_sg U63424 ( .A(n52507), .B(n13854), .X(n13785) );
  nand_x1_sg U63425 ( .A(n13818), .B(n52506), .X(n13854) );
  nor_x1_sg U63426 ( .A(n52506), .B(n13818), .X(n13855) );
  nand_x4_sg U63427 ( .A(n52786), .B(n14625), .X(n14556) );
  nand_x1_sg U63428 ( .A(n14588), .B(n52785), .X(n14625) );
  nor_x1_sg U63429 ( .A(n52785), .B(n14588), .X(n14626) );
  nand_x4_sg U63430 ( .A(n53906), .B(n17746), .X(n17677) );
  nand_x1_sg U63431 ( .A(n17709), .B(n53905), .X(n17746) );
  nor_x1_sg U63432 ( .A(n53905), .B(n17709), .X(n17747) );
  nand_x4_sg U63433 ( .A(n54471), .B(n19291), .X(n19222) );
  nand_x1_sg U63434 ( .A(n19254), .B(n54470), .X(n19291) );
  nor_x1_sg U63435 ( .A(n54470), .B(n19254), .X(n19292) );
  nand_x4_sg U63436 ( .A(n55039), .B(n20835), .X(n20766) );
  nand_x1_sg U63437 ( .A(n20798), .B(n55038), .X(n20835) );
  nor_x1_sg U63438 ( .A(n55038), .B(n20798), .X(n20836) );
  nand_x4_sg U63439 ( .A(n13332), .B(n13333), .X(n13321) );
  nand_x1_sg U63440 ( .A(n13336), .B(n52220), .X(n13332) );
  nand_x1_sg U63441 ( .A(n13334), .B(n13335), .X(n13333) );
  nand_x4_sg U63442 ( .A(n15665), .B(n15666), .X(n15654) );
  nand_x1_sg U63443 ( .A(n15669), .B(n53054), .X(n15665) );
  nand_x1_sg U63444 ( .A(n15667), .B(n15668), .X(n15666) );
  nand_x4_sg U63445 ( .A(n17231), .B(n17232), .X(n17220) );
  nand_x1_sg U63446 ( .A(n17235), .B(n53612), .X(n17231) );
  nand_x1_sg U63447 ( .A(n17233), .B(n17234), .X(n17232) );
  nand_x4_sg U63448 ( .A(n25404), .B(n25405), .X(n25403) );
  nor_x1_sg U63449 ( .A(n51270), .B(n25406), .X(n25405) );
  nor_x1_sg U63450 ( .A(n25409), .B(n46236), .X(n25404) );
  nand_x4_sg U63451 ( .A(n25411), .B(n25412), .X(n25410) );
  nor_x1_sg U63452 ( .A(n51278), .B(n25413), .X(n25412) );
  nor_x1_sg U63453 ( .A(n25416), .B(n46236), .X(n25411) );
  nand_x4_sg U63454 ( .A(n25418), .B(n25419), .X(n25417) );
  nor_x1_sg U63455 ( .A(n51290), .B(n25420), .X(n25419) );
  nor_x1_sg U63456 ( .A(n25424), .B(n46236), .X(n25418) );
  nand_x4_sg U63457 ( .A(n25676), .B(n25677), .X(n25675) );
  nor_x1_sg U63458 ( .A(n51539), .B(n25678), .X(n25677) );
  nor_x1_sg U63459 ( .A(n25681), .B(n46236), .X(n25676) );
  nand_x4_sg U63460 ( .A(n25683), .B(n25684), .X(n25682) );
  nor_x1_sg U63461 ( .A(n51548), .B(n25685), .X(n25684) );
  nor_x1_sg U63462 ( .A(n25688), .B(n46236), .X(n25683) );
  nand_x4_sg U63463 ( .A(n25690), .B(n25691), .X(n25689) );
  nor_x1_sg U63464 ( .A(n51556), .B(n25692), .X(n25691) );
  nor_x1_sg U63465 ( .A(n25695), .B(n46236), .X(n25690) );
  nand_x4_sg U63466 ( .A(n25697), .B(n25698), .X(n25696) );
  nor_x1_sg U63467 ( .A(n51561), .B(n25699), .X(n25698) );
  nor_x1_sg U63468 ( .A(n25703), .B(n46236), .X(n25697) );
  nand_x4_sg U63469 ( .A(n25954), .B(n25955), .X(n25953) );
  nor_x1_sg U63470 ( .A(n51822), .B(n25956), .X(n25955) );
  nor_x1_sg U63471 ( .A(n25959), .B(n46236), .X(n25954) );
  nand_x4_sg U63472 ( .A(n25961), .B(n25962), .X(n25960) );
  nor_x1_sg U63473 ( .A(n51830), .B(n25963), .X(n25962) );
  nor_x1_sg U63474 ( .A(n25966), .B(n46236), .X(n25961) );
  nand_x4_sg U63475 ( .A(n25968), .B(n25969), .X(n25967) );
  nor_x1_sg U63476 ( .A(n51837), .B(n25970), .X(n25969) );
  nor_x1_sg U63477 ( .A(n25973), .B(n46236), .X(n25968) );
  nand_x4_sg U63478 ( .A(n25975), .B(n25976), .X(n25974) );
  nor_x1_sg U63479 ( .A(n51851), .B(n25977), .X(n25976) );
  nor_x1_sg U63480 ( .A(n25981), .B(n46236), .X(n25975) );
  nand_x4_sg U63481 ( .A(n26046), .B(n26047), .X(n26045) );
  nor_x1_sg U63482 ( .A(n42485), .B(n26049), .X(n26047) );
  nor_x1_sg U63483 ( .A(n26052), .B(n46236), .X(n26046) );
  nand_x4_sg U63484 ( .A(n26235), .B(n26236), .X(n26234) );
  nor_x1_sg U63485 ( .A(n52096), .B(n26237), .X(n26236) );
  nor_x1_sg U63486 ( .A(n26240), .B(n46236), .X(n26235) );
  nand_x4_sg U63487 ( .A(n26242), .B(n26243), .X(n26241) );
  nor_x1_sg U63488 ( .A(n52105), .B(n26244), .X(n26243) );
  nor_x1_sg U63489 ( .A(n26247), .B(n46236), .X(n26242) );
  nand_x4_sg U63490 ( .A(n26249), .B(n26250), .X(n26248) );
  nor_x1_sg U63491 ( .A(n52113), .B(n26251), .X(n26250) );
  nor_x1_sg U63492 ( .A(n26254), .B(n46236), .X(n26249) );
  nand_x4_sg U63493 ( .A(n26256), .B(n26257), .X(n26255) );
  nor_x1_sg U63494 ( .A(n52118), .B(n26258), .X(n26257) );
  nor_x1_sg U63495 ( .A(n26262), .B(n46236), .X(n26256) );
  nand_x4_sg U63496 ( .A(n26327), .B(n26328), .X(n26326) );
  nor_x1_sg U63497 ( .A(n42483), .B(n26330), .X(n26328) );
  nor_x1_sg U63498 ( .A(n26333), .B(n46236), .X(n26327) );
  nand_x4_sg U63499 ( .A(n26508), .B(n26509), .X(n26507) );
  nor_x1_sg U63500 ( .A(n52367), .B(n26510), .X(n26509) );
  nor_x1_sg U63501 ( .A(n26511), .B(n46236), .X(n26508) );
  nand_x4_sg U63502 ( .A(n26514), .B(n26515), .X(n26513) );
  nor_x1_sg U63503 ( .A(n52374), .B(n26516), .X(n26515) );
  nor_x1_sg U63504 ( .A(n26519), .B(n46236), .X(n26514) );
  nand_x4_sg U63505 ( .A(n26521), .B(n26522), .X(n26520) );
  nor_x1_sg U63506 ( .A(n52382), .B(n26523), .X(n26522) );
  nor_x1_sg U63507 ( .A(n26526), .B(n46236), .X(n26521) );
  nand_x4_sg U63508 ( .A(n26528), .B(n26529), .X(n26527) );
  nor_x1_sg U63509 ( .A(n52389), .B(n26530), .X(n26529) );
  nor_x1_sg U63510 ( .A(n26533), .B(n46236), .X(n26528) );
  nand_x4_sg U63511 ( .A(n26535), .B(n26536), .X(n26534) );
  nor_x1_sg U63512 ( .A(n52403), .B(n26537), .X(n26536) );
  nor_x1_sg U63513 ( .A(n26541), .B(n46236), .X(n26535) );
  nand_x4_sg U63514 ( .A(n26606), .B(n26607), .X(n26605) );
  nor_x1_sg U63515 ( .A(n42481), .B(n26609), .X(n26607) );
  nor_x1_sg U63516 ( .A(n26612), .B(n46236), .X(n26606) );
  nand_x4_sg U63517 ( .A(n26792), .B(n26793), .X(n26791) );
  nor_x1_sg U63518 ( .A(n52651), .B(n26794), .X(n26793) );
  nor_x1_sg U63519 ( .A(n26797), .B(n46236), .X(n26792) );
  nand_x4_sg U63520 ( .A(n26799), .B(n26800), .X(n26798) );
  nor_x1_sg U63521 ( .A(n52659), .B(n26801), .X(n26800) );
  nor_x1_sg U63522 ( .A(n26804), .B(n46236), .X(n26799) );
  nand_x4_sg U63523 ( .A(n26806), .B(n26807), .X(n26805) );
  nor_x1_sg U63524 ( .A(n52667), .B(n26808), .X(n26807) );
  nor_x1_sg U63525 ( .A(n26811), .B(n46236), .X(n26806) );
  nand_x4_sg U63526 ( .A(n26813), .B(n26814), .X(n26812) );
  nor_x1_sg U63527 ( .A(n52680), .B(n26815), .X(n26814) );
  nor_x1_sg U63528 ( .A(n26819), .B(n46236), .X(n26813) );
  nand_x4_sg U63529 ( .A(n27071), .B(n27072), .X(n27070) );
  nor_x1_sg U63530 ( .A(n52930), .B(n27073), .X(n27072) );
  nor_x1_sg U63531 ( .A(n27076), .B(n46236), .X(n27071) );
  nand_x4_sg U63532 ( .A(n27078), .B(n27079), .X(n27077) );
  nor_x1_sg U63533 ( .A(n52939), .B(n27080), .X(n27079) );
  nor_x1_sg U63534 ( .A(n27083), .B(n46236), .X(n27078) );
  nand_x4_sg U63535 ( .A(n27085), .B(n27086), .X(n27084) );
  nor_x1_sg U63536 ( .A(n52947), .B(n27087), .X(n27086) );
  nor_x1_sg U63537 ( .A(n27090), .B(n46236), .X(n27085) );
  nand_x4_sg U63538 ( .A(n27092), .B(n27093), .X(n27091) );
  nor_x1_sg U63539 ( .A(n52952), .B(n27094), .X(n27093) );
  nor_x1_sg U63540 ( .A(n27098), .B(n46236), .X(n27092) );
  nand_x4_sg U63541 ( .A(n27163), .B(n27164), .X(n27162) );
  nor_x1_sg U63542 ( .A(n42479), .B(n27166), .X(n27164) );
  nor_x1_sg U63543 ( .A(n27169), .B(n46236), .X(n27163) );
  nand_x4_sg U63544 ( .A(n27351), .B(n27352), .X(n27350) );
  nor_x1_sg U63545 ( .A(n53210), .B(n27353), .X(n27352) );
  nor_x1_sg U63546 ( .A(n27356), .B(n46236), .X(n27351) );
  nand_x4_sg U63547 ( .A(n27358), .B(n27359), .X(n27357) );
  nor_x1_sg U63548 ( .A(n53218), .B(n27360), .X(n27359) );
  nor_x1_sg U63549 ( .A(n27363), .B(n46236), .X(n27358) );
  nand_x4_sg U63550 ( .A(n27365), .B(n27366), .X(n27364) );
  nor_x1_sg U63551 ( .A(n53225), .B(n27367), .X(n27366) );
  nor_x1_sg U63552 ( .A(n27370), .B(n46236), .X(n27365) );
  nand_x4_sg U63553 ( .A(n27372), .B(n27373), .X(n27371) );
  nor_x1_sg U63554 ( .A(n53237), .B(n27374), .X(n27373) );
  nor_x1_sg U63555 ( .A(n27378), .B(n46236), .X(n27372) );
  nand_x4_sg U63556 ( .A(n27631), .B(n27632), .X(n27630) );
  nor_x1_sg U63557 ( .A(n53488), .B(n27633), .X(n27632) );
  nor_x1_sg U63558 ( .A(n27636), .B(n46236), .X(n27631) );
  nand_x4_sg U63559 ( .A(n27638), .B(n27639), .X(n27637) );
  nor_x1_sg U63560 ( .A(n53497), .B(n27640), .X(n27639) );
  nor_x1_sg U63561 ( .A(n27643), .B(n46236), .X(n27638) );
  nand_x4_sg U63562 ( .A(n27645), .B(n27646), .X(n27644) );
  nor_x1_sg U63563 ( .A(n53505), .B(n27647), .X(n27646) );
  nor_x1_sg U63564 ( .A(n27650), .B(n46236), .X(n27645) );
  nand_x4_sg U63565 ( .A(n27652), .B(n27653), .X(n27651) );
  nor_x1_sg U63566 ( .A(n53510), .B(n27654), .X(n27653) );
  nor_x1_sg U63567 ( .A(n27658), .B(n46236), .X(n27652) );
  nand_x4_sg U63568 ( .A(n27723), .B(n27724), .X(n27722) );
  nor_x1_sg U63569 ( .A(n42475), .B(n27726), .X(n27724) );
  nor_x1_sg U63570 ( .A(n27729), .B(n46236), .X(n27723) );
  nand_x4_sg U63571 ( .A(n27911), .B(n27912), .X(n27910) );
  nor_x1_sg U63572 ( .A(n53768), .B(n27913), .X(n27912) );
  nor_x1_sg U63573 ( .A(n27916), .B(n46236), .X(n27911) );
  nand_x4_sg U63574 ( .A(n27918), .B(n27919), .X(n27917) );
  nor_x1_sg U63575 ( .A(n53775), .B(n27920), .X(n27919) );
  nor_x1_sg U63576 ( .A(n27923), .B(n46236), .X(n27918) );
  nand_x4_sg U63577 ( .A(n27925), .B(n27926), .X(n27924) );
  nor_x1_sg U63578 ( .A(n53784), .B(n27927), .X(n27926) );
  nor_x1_sg U63579 ( .A(n27930), .B(n46236), .X(n27925) );
  nand_x4_sg U63580 ( .A(n27932), .B(n27933), .X(n27931) );
  nor_x1_sg U63581 ( .A(n53789), .B(n27934), .X(n27933) );
  nor_x1_sg U63582 ( .A(n27938), .B(n46236), .X(n27932) );
  nand_x4_sg U63583 ( .A(n28190), .B(n28191), .X(n28189) );
  nor_x1_sg U63584 ( .A(n54052), .B(n28192), .X(n28191) );
  nor_x1_sg U63585 ( .A(n28195), .B(n46236), .X(n28190) );
  nand_x4_sg U63586 ( .A(n28197), .B(n28198), .X(n28196) );
  nor_x1_sg U63587 ( .A(n54056), .B(n28199), .X(n28198) );
  nor_x1_sg U63588 ( .A(n28202), .B(n46236), .X(n28197) );
  nand_x4_sg U63589 ( .A(n28204), .B(n28205), .X(n28203) );
  nor_x1_sg U63590 ( .A(n54066), .B(n28206), .X(n28205) );
  nor_x1_sg U63591 ( .A(n28209), .B(n46236), .X(n28204) );
  nand_x4_sg U63592 ( .A(n28211), .B(n28212), .X(n28210) );
  nor_x1_sg U63593 ( .A(n54080), .B(n28213), .X(n28212) );
  nor_x1_sg U63594 ( .A(n28217), .B(n46236), .X(n28211) );
  nand_x4_sg U63595 ( .A(n28469), .B(n28470), .X(n28468) );
  nor_x1_sg U63596 ( .A(n54333), .B(n28471), .X(n28470) );
  nor_x1_sg U63597 ( .A(n28474), .B(n46236), .X(n28469) );
  nand_x4_sg U63598 ( .A(n28476), .B(n28477), .X(n28475) );
  nor_x1_sg U63599 ( .A(n54340), .B(n28478), .X(n28477) );
  nor_x1_sg U63600 ( .A(n28481), .B(n46236), .X(n28476) );
  nand_x4_sg U63601 ( .A(n28483), .B(n28484), .X(n28482) );
  nor_x1_sg U63602 ( .A(n54349), .B(n28485), .X(n28484) );
  nor_x1_sg U63603 ( .A(n28488), .B(n46236), .X(n28483) );
  nand_x4_sg U63604 ( .A(n28490), .B(n28491), .X(n28489) );
  nor_x1_sg U63605 ( .A(n54354), .B(n28492), .X(n28491) );
  nor_x1_sg U63606 ( .A(n28496), .B(n46236), .X(n28490) );
  nand_x4_sg U63607 ( .A(n28748), .B(n28749), .X(n28747) );
  nor_x1_sg U63608 ( .A(n54617), .B(n28750), .X(n28749) );
  nor_x1_sg U63609 ( .A(n28753), .B(n46236), .X(n28748) );
  nand_x4_sg U63610 ( .A(n28755), .B(n28756), .X(n28754) );
  nor_x1_sg U63611 ( .A(n54624), .B(n28757), .X(n28756) );
  nor_x1_sg U63612 ( .A(n28760), .B(n46236), .X(n28755) );
  nand_x4_sg U63613 ( .A(n28762), .B(n28763), .X(n28761) );
  nor_x1_sg U63614 ( .A(n54632), .B(n28764), .X(n28763) );
  nor_x1_sg U63615 ( .A(n28767), .B(n46236), .X(n28762) );
  nand_x4_sg U63616 ( .A(n28769), .B(n28770), .X(n28768) );
  nor_x1_sg U63617 ( .A(n54644), .B(n28771), .X(n28770) );
  nor_x1_sg U63618 ( .A(n28775), .B(n46236), .X(n28769) );
  nand_x4_sg U63619 ( .A(n29028), .B(n29029), .X(n29027) );
  nor_x1_sg U63620 ( .A(n54901), .B(n29030), .X(n29029) );
  nor_x1_sg U63621 ( .A(n29033), .B(n46236), .X(n29028) );
  nand_x4_sg U63622 ( .A(n29035), .B(n29036), .X(n29034) );
  nor_x1_sg U63623 ( .A(n54908), .B(n29037), .X(n29036) );
  nor_x1_sg U63624 ( .A(n29040), .B(n46236), .X(n29035) );
  nand_x4_sg U63625 ( .A(n29042), .B(n29043), .X(n29041) );
  nor_x1_sg U63626 ( .A(n54917), .B(n29044), .X(n29043) );
  nor_x1_sg U63627 ( .A(n29047), .B(n46236), .X(n29042) );
  nand_x4_sg U63628 ( .A(n29049), .B(n29050), .X(n29048) );
  nor_x1_sg U63629 ( .A(n54922), .B(n29051), .X(n29050) );
  nor_x1_sg U63630 ( .A(n29055), .B(n46236), .X(n29049) );
  nand_x4_sg U63631 ( .A(n29309), .B(n29310), .X(n29308) );
  nor_x1_sg U63632 ( .A(n55185), .B(n29311), .X(n29310) );
  nor_x1_sg U63633 ( .A(n29314), .B(n46236), .X(n29309) );
  nand_x4_sg U63634 ( .A(n29316), .B(n29317), .X(n29315) );
  nor_x1_sg U63635 ( .A(n55192), .B(n29318), .X(n29317) );
  nor_x1_sg U63636 ( .A(n29321), .B(n46236), .X(n29316) );
  nand_x4_sg U63637 ( .A(n29323), .B(n29324), .X(n29322) );
  nor_x1_sg U63638 ( .A(n55200), .B(n29325), .X(n29324) );
  nor_x1_sg U63639 ( .A(n29328), .B(n46236), .X(n29323) );
  nand_x2_sg U63640 ( .A(n46361), .B(n27929), .X(n27928) );
  nand_x2_sg U63641 ( .A(n46314), .B(n28487), .X(n28486) );
  nand_x2_sg U63642 ( .A(n46269), .B(n29046), .X(n29045) );
  nand_x2_sg U63643 ( .A(n46567), .B(n25408), .X(n25407) );
  nand_x2_sg U63644 ( .A(n46450), .B(n26810), .X(n26809) );
  nor_x1_sg U63645 ( .A(n44096), .B(n46527), .X(\L2_0/n3972 ) );
  nor_x1_sg U63646 ( .A(n44090), .B(n46415), .X(\L2_0/n3572 ) );
  nor_x1_sg U63647 ( .A(n44092), .B(n46460), .X(\L2_0/n3732 ) );
  nor_x1_sg U63648 ( .A(n41358), .B(n46370), .X(\L2_0/n3412 ) );
  nor_x1_sg U63649 ( .A(n41356), .B(n46323), .X(\L2_0/n3252 ) );
  nor_x1_sg U63650 ( .A(n41352), .B(n46278), .X(\L2_0/n3092 ) );
  nor_x1_sg U63651 ( .A(n42891), .B(n46549), .X(\L2_0/n4052 ) );
  nor_x1_sg U63652 ( .A(n42885), .B(n46505), .X(\L2_0/n3892 ) );
  nor_x1_sg U63653 ( .A(n42877), .B(n46437), .X(\L2_0/n3652 ) );
  nor_x1_sg U63654 ( .A(n42871), .B(n46393), .X(\L2_0/n3492 ) );
  nor_x1_sg U63655 ( .A(n44086), .B(n46303), .X(\L2_0/n3172 ) );
  nor_x1_sg U63656 ( .A(n44084), .B(n46258), .X(\L2_0/n3012 ) );
  nor_x1_sg U63657 ( .A(n42865), .B(n46350), .X(\L2_0/n3288 ) );
  nor_x1_sg U63658 ( .A(n42861), .B(n46303), .X(\L2_0/n3128 ) );
  nor_x1_sg U63659 ( .A(n44088), .B(n46350), .X(\L2_0/n3332 ) );
  nand_x4_sg U63660 ( .A(n52431), .B(n13636), .X(n13588) );
  nand_x1_sg U63661 ( .A(n13630), .B(n13637), .X(n13636) );
  nor_x1_sg U63662 ( .A(n13637), .B(n13630), .X(n13638) );
  nand_x2_sg U63663 ( .A(n46540), .B(n25694), .X(n25693) );
  nand_x2_sg U63664 ( .A(n46496), .B(n26253), .X(n26252) );
  nand_x2_sg U63665 ( .A(n46428), .B(n27089), .X(n27088) );
  nand_x2_sg U63666 ( .A(n46384), .B(n27649), .X(n27648) );
  nand_x2_sg U63667 ( .A(n46294), .B(n28766), .X(n28765) );
  nand_x2_sg U63668 ( .A(n46249), .B(n29327), .X(n29326) );
  nand_x4_sg U63669 ( .A(n18565), .B(n18566), .X(n18563) );
  nand_x1_sg U63670 ( .A(n18573), .B(n18571), .X(n18565) );
  nor_x1_sg U63671 ( .A(n42603), .B(n46344), .X(n18567) );
  nand_x4_sg U63672 ( .A(n10809), .B(n10810), .X(n10750) );
  nand_x1_sg U63673 ( .A(n51336), .B(n51355), .X(n10809) );
  nand_x1_sg U63674 ( .A(n10803), .B(n10799), .X(n10810) );
  nand_x4_sg U63675 ( .A(n20135), .B(n20136), .X(n20076) );
  nand_x1_sg U63676 ( .A(n54690), .B(n54709), .X(n20135) );
  nand_x1_sg U63677 ( .A(n20129), .B(n20125), .X(n20136) );
  nand_x4_sg U63678 ( .A(n21680), .B(n21681), .X(n21621) );
  nand_x1_sg U63679 ( .A(n55258), .B(n55277), .X(n21680) );
  nand_x1_sg U63680 ( .A(n21674), .B(n21670), .X(n21681) );
  nand_x4_sg U63681 ( .A(n17544), .B(n17580), .X(n17579) );
  nand_x1_sg U63682 ( .A(n17581), .B(n17582), .X(n17580) );
  nand_x4_sg U63683 ( .A(n19089), .B(n19125), .X(n19124) );
  nand_x1_sg U63684 ( .A(n19126), .B(n19127), .X(n19125) );
  nand_x4_sg U63685 ( .A(n20633), .B(n20669), .X(n20668) );
  nand_x1_sg U63686 ( .A(n20670), .B(n20671), .X(n20669) );
  nand_x4_sg U63687 ( .A(n17497), .B(n17498), .X(n17486) );
  nor_x1_sg U63688 ( .A(n17499), .B(n46367), .X(n17498) );
  nor_x1_sg U63689 ( .A(n17505), .B(n17492), .X(n17497) );
  nand_x4_sg U63690 ( .A(n19042), .B(n19043), .X(n19031) );
  nor_x1_sg U63691 ( .A(n19044), .B(n46320), .X(n19043) );
  nor_x1_sg U63692 ( .A(n19050), .B(n19037), .X(n19042) );
  nand_x4_sg U63693 ( .A(n20586), .B(n20587), .X(n20575) );
  nor_x1_sg U63694 ( .A(n20588), .B(n46275), .X(n20587) );
  nor_x1_sg U63695 ( .A(n20594), .B(n20581), .X(n20586) );
  nand_x4_sg U63696 ( .A(n11823), .B(n11824), .X(n11659) );
  nand_x1_sg U63697 ( .A(n51755), .B(n51777), .X(n11823) );
  nand_x1_sg U63698 ( .A(n11679), .B(n11681), .X(n11824) );
  nand_x4_sg U63699 ( .A(n14935), .B(n14936), .X(n14772) );
  nand_x1_sg U63700 ( .A(n52864), .B(n52887), .X(n14936) );
  nand_x1_sg U63701 ( .A(n14791), .B(n14793), .X(n14935) );
  nand_x4_sg U63702 ( .A(n18056), .B(n18057), .X(n17893) );
  nand_x1_sg U63703 ( .A(n53984), .B(n54007), .X(n18057) );
  nand_x1_sg U63704 ( .A(n17912), .B(n17914), .X(n18056) );
  nand_x4_sg U63705 ( .A(n18828), .B(n18829), .X(n18662) );
  nand_x1_sg U63706 ( .A(n54267), .B(n54289), .X(n18829) );
  nand_x1_sg U63707 ( .A(n18681), .B(n18683), .X(n18828) );
  nand_x4_sg U63708 ( .A(n19601), .B(n19602), .X(n19438) );
  nand_x1_sg U63709 ( .A(n54549), .B(n54572), .X(n19602) );
  nand_x1_sg U63710 ( .A(n19457), .B(n19459), .X(n19601) );
  nand_x4_sg U63711 ( .A(n20373), .B(n20374), .X(n20207) );
  nand_x1_sg U63712 ( .A(n54834), .B(n54857), .X(n20374) );
  nand_x1_sg U63713 ( .A(n20226), .B(n20228), .X(n20373) );
  nand_x4_sg U63714 ( .A(n21145), .B(n21146), .X(n20982) );
  nand_x1_sg U63715 ( .A(n55117), .B(n55140), .X(n21146) );
  nand_x1_sg U63716 ( .A(n21001), .B(n21003), .X(n21145) );
  nand_x4_sg U63717 ( .A(n21918), .B(n21919), .X(n21752) );
  nand_x1_sg U63718 ( .A(n55402), .B(n55425), .X(n21919) );
  nand_x1_sg U63719 ( .A(n21771), .B(n21773), .X(n21918) );
  nand_x4_sg U63720 ( .A(n13752), .B(n13806), .X(n13804) );
  nand_x1_sg U63721 ( .A(n52528), .B(n13807), .X(n13806) );
  nand_x4_sg U63722 ( .A(n17437), .B(n53779), .X(n17425) );
  nand_x1_sg U63723 ( .A(n17440), .B(n17439), .X(n17437) );
  nor_x1_sg U63724 ( .A(n17439), .B(n17440), .X(n17438) );
  nand_x4_sg U63725 ( .A(n18982), .B(n54344), .X(n18970) );
  nand_x1_sg U63726 ( .A(n18985), .B(n18984), .X(n18982) );
  nor_x1_sg U63727 ( .A(n18984), .B(n18985), .X(n18983) );
  nand_x4_sg U63728 ( .A(n20526), .B(n54912), .X(n20514) );
  nand_x1_sg U63729 ( .A(n20529), .B(n20528), .X(n20526) );
  nor_x1_sg U63730 ( .A(n20528), .B(n20529), .X(n20527) );
  nand_x4_sg U63731 ( .A(n18414), .B(n18466), .X(n18460) );
  nand_x1_sg U63732 ( .A(n42802), .B(n18468), .X(n18466) );
  nand_x4_sg U63733 ( .A(n11322), .B(n51631), .X(n11314) );
  nor_x1_sg U63734 ( .A(n11324), .B(n11325), .X(n11323) );
  nand_x4_sg U63735 ( .A(n12191), .B(n12245), .X(n12243) );
  nand_x1_sg U63736 ( .A(n43311), .B(n12247), .X(n12245) );
  nand_x4_sg U63737 ( .A(n54065), .B(n18203), .X(n18192) );
  nand_x1_sg U63738 ( .A(n18204), .B(n18205), .X(n18203) );
  nor_x1_sg U63739 ( .A(n18205), .B(n18204), .X(n18206) );
  nand_x4_sg U63740 ( .A(n12528), .B(n12529), .X(n12526) );
  nand_x1_sg U63741 ( .A(n41588), .B(n12531), .X(n12528) );
  nand_x4_sg U63742 ( .A(n14089), .B(n14090), .X(n14087) );
  nand_x1_sg U63743 ( .A(n42769), .B(n14092), .X(n14089) );
  nand_x4_sg U63744 ( .A(n10422), .B(n51273), .X(n10412) );
  nand_x1_sg U63745 ( .A(n10425), .B(n10424), .X(n10422) );
  nor_x1_sg U63746 ( .A(n10424), .B(n10425), .X(n10423) );
  nand_x4_sg U63747 ( .A(n19904), .B(n19905), .X(n19897) );
  nand_x1_sg U63748 ( .A(n19907), .B(n54700), .X(n19904) );
  nand_x1_sg U63749 ( .A(n19906), .B(n54655), .X(n19905) );
  nand_x4_sg U63750 ( .A(n21449), .B(n21450), .X(n21442) );
  nand_x1_sg U63751 ( .A(n21452), .B(n55268), .X(n21449) );
  nand_x1_sg U63752 ( .A(n21451), .B(n55223), .X(n21450) );
  nand_x4_sg U63753 ( .A(n12883), .B(n52188), .X(n12875) );
  nor_x1_sg U63754 ( .A(n12885), .B(n12886), .X(n12884) );
  nand_x4_sg U63755 ( .A(n13663), .B(n52464), .X(n13655) );
  nor_x1_sg U63756 ( .A(n13665), .B(n13666), .X(n13664) );
  nand_x4_sg U63757 ( .A(n15216), .B(n53022), .X(n15208) );
  nor_x1_sg U63758 ( .A(n15218), .B(n15219), .X(n15217) );
  nand_x4_sg U63759 ( .A(n16782), .B(n53580), .X(n16774) );
  nor_x1_sg U63760 ( .A(n16784), .B(n16785), .X(n16783) );
  nand_x4_sg U63761 ( .A(n19749), .B(n54627), .X(n19739) );
  nand_x1_sg U63762 ( .A(n19752), .B(n19751), .X(n19749) );
  nor_x1_sg U63763 ( .A(n19751), .B(n19752), .X(n19750) );
  nand_x4_sg U63764 ( .A(n21294), .B(n55195), .X(n21284) );
  nand_x1_sg U63765 ( .A(n21297), .B(n21296), .X(n21294) );
  nor_x1_sg U63766 ( .A(n21296), .B(n21297), .X(n21295) );
  nand_x4_sg U63767 ( .A(n14469), .B(n14470), .X(n14462) );
  nand_x1_sg U63768 ( .A(n14472), .B(n52736), .X(n14469) );
  nand_x1_sg U63769 ( .A(n14471), .B(n52691), .X(n14470) );
  nand_x4_sg U63770 ( .A(n18359), .B(n18360), .X(n18352) );
  nand_x1_sg U63771 ( .A(n18362), .B(n54136), .X(n18359) );
  nand_x1_sg U63772 ( .A(n18361), .B(n54093), .X(n18360) );
  nand_x4_sg U63773 ( .A(n13338), .B(n52297), .X(n13203) );
  nor_x1_sg U63774 ( .A(n13347), .B(n44437), .X(n13346) );
  nand_x4_sg U63775 ( .A(n14118), .B(n52572), .X(n13983) );
  nor_x1_sg U63776 ( .A(n14127), .B(n44435), .X(n14126) );
  nand_x4_sg U63777 ( .A(n15671), .B(n53131), .X(n15536) );
  nor_x1_sg U63778 ( .A(n15680), .B(n44433), .X(n15679) );
  nand_x4_sg U63779 ( .A(n17237), .B(n53689), .X(n17102) );
  nor_x1_sg U63780 ( .A(n17246), .B(n44431), .X(n17245) );
  nand_x4_sg U63781 ( .A(n54156), .B(n18363), .X(n18348) );
  nand_x1_sg U63782 ( .A(n54155), .B(n18364), .X(n18363) );
  nor_x1_sg U63783 ( .A(n18364), .B(n54155), .X(n18365) );
  nand_x4_sg U63784 ( .A(n54721), .B(n19908), .X(n19893) );
  nand_x1_sg U63785 ( .A(n54720), .B(n19909), .X(n19908) );
  nor_x1_sg U63786 ( .A(n19909), .B(n54720), .X(n19910) );
  nand_x4_sg U63787 ( .A(n55289), .B(n21453), .X(n21438) );
  nand_x1_sg U63788 ( .A(n55288), .B(n21454), .X(n21453) );
  nor_x1_sg U63789 ( .A(n21454), .B(n55288), .X(n21455) );
  nand_x4_sg U63790 ( .A(n51553), .B(n11165), .X(n11065) );
  nand_x1_sg U63791 ( .A(n51547), .B(n11166), .X(n11165) );
  nor_x1_sg U63792 ( .A(n11166), .B(n51547), .X(n11167) );
  nand_x4_sg U63793 ( .A(n52110), .B(n12726), .X(n12626) );
  nand_x1_sg U63794 ( .A(n52104), .B(n12727), .X(n12726) );
  nor_x1_sg U63795 ( .A(n12727), .B(n52104), .X(n12728) );
  nand_x4_sg U63796 ( .A(n52944), .B(n15059), .X(n14959) );
  nand_x1_sg U63797 ( .A(n52938), .B(n15060), .X(n15059) );
  nor_x1_sg U63798 ( .A(n15060), .B(n52938), .X(n15061) );
  nand_x4_sg U63799 ( .A(n53502), .B(n16625), .X(n16525) );
  nand_x1_sg U63800 ( .A(n53496), .B(n16626), .X(n16625) );
  nor_x1_sg U63801 ( .A(n16626), .B(n53496), .X(n16627) );
  nand_x4_sg U63802 ( .A(n11748), .B(n11749), .X(n11746) );
  nand_x1_sg U63803 ( .A(n51770), .B(n11751), .X(n11748) );
  nand_x4_sg U63804 ( .A(n13309), .B(n13310), .X(n13307) );
  nand_x1_sg U63805 ( .A(n42771), .B(n13312), .X(n13309) );
  nand_x4_sg U63806 ( .A(n15642), .B(n15643), .X(n15640) );
  nand_x1_sg U63807 ( .A(n42767), .B(n15645), .X(n15642) );
  nand_x4_sg U63808 ( .A(n17208), .B(n17209), .X(n17206) );
  nand_x1_sg U63809 ( .A(n42763), .B(n17211), .X(n17208) );
  nand_x4_sg U63810 ( .A(n14301), .B(n52672), .X(n14298) );
  nor_x1_sg U63811 ( .A(n44473), .B(n14304), .X(n14302) );
  nand_x4_sg U63812 ( .A(n51638), .B(n11355), .X(n11336) );
  nand_x1_sg U63813 ( .A(n51637), .B(n11356), .X(n11355) );
  nor_x1_sg U63814 ( .A(n11356), .B(n51637), .X(n11357) );
  nand_x4_sg U63815 ( .A(n52194), .B(n12916), .X(n12897) );
  nand_x1_sg U63816 ( .A(n52193), .B(n12917), .X(n12916) );
  nor_x1_sg U63817 ( .A(n12917), .B(n52193), .X(n12918) );
  nand_x4_sg U63818 ( .A(n53028), .B(n15249), .X(n15230) );
  nand_x1_sg U63819 ( .A(n53027), .B(n15250), .X(n15249) );
  nor_x1_sg U63820 ( .A(n15250), .B(n53027), .X(n15251) );
  nand_x4_sg U63821 ( .A(n53586), .B(n16815), .X(n16796) );
  nand_x1_sg U63822 ( .A(n53585), .B(n16816), .X(n16815) );
  nor_x1_sg U63823 ( .A(n16816), .B(n53585), .X(n16817) );
  nand_x4_sg U63824 ( .A(n12036), .B(n12037), .X(n12024) );
  nor_x1_sg U63825 ( .A(n12046), .B(n12016), .X(n12036) );
  nor_x1_sg U63826 ( .A(n12038), .B(n46519), .X(n12037) );
  nand_x4_sg U63827 ( .A(n15931), .B(n15932), .X(n15919) );
  nor_x1_sg U63828 ( .A(n15941), .B(n15911), .X(n15931) );
  nor_x1_sg U63829 ( .A(n15933), .B(n46407), .X(n15932) );
  nand_x4_sg U63830 ( .A(n10632), .B(n10684), .X(n10678) );
  nand_x1_sg U63831 ( .A(n43315), .B(n10686), .X(n10684) );
  nand_x4_sg U63832 ( .A(n19959), .B(n20011), .X(n20005) );
  nand_x1_sg U63833 ( .A(n43323), .B(n20013), .X(n20011) );
  nand_x4_sg U63834 ( .A(n21504), .B(n21556), .X(n21550) );
  nand_x1_sg U63835 ( .A(n43319), .B(n21558), .X(n21556) );
  nand_x4_sg U63836 ( .A(n17822), .B(n17823), .X(n17763) );
  nand_x1_sg U63837 ( .A(n53867), .B(n17813), .X(n17823) );
  nand_x1_sg U63838 ( .A(n53846), .B(n17812), .X(n17822) );
  nand_x4_sg U63839 ( .A(n19367), .B(n19368), .X(n19308) );
  nand_x1_sg U63840 ( .A(n54432), .B(n19358), .X(n19368) );
  nand_x1_sg U63841 ( .A(n54411), .B(n19357), .X(n19367) );
  nand_x4_sg U63842 ( .A(n20911), .B(n20912), .X(n20852) );
  nand_x1_sg U63843 ( .A(n55000), .B(n20902), .X(n20912) );
  nand_x1_sg U63844 ( .A(n54979), .B(n20901), .X(n20911) );
  nand_x4_sg U63845 ( .A(n18189), .B(n54072), .X(n18187) );
  nor_x1_sg U63846 ( .A(n45457), .B(n18192), .X(n18190) );
  nand_x4_sg U63847 ( .A(n19736), .B(n54636), .X(n19733) );
  nor_x1_sg U63848 ( .A(n44471), .B(n19739), .X(n19737) );
  nand_x4_sg U63849 ( .A(n21281), .B(n55204), .X(n21278) );
  nor_x1_sg U63850 ( .A(n44469), .B(n21284), .X(n21282) );
  nand_x4_sg U63851 ( .A(n10409), .B(n51282), .X(n10406) );
  nor_x1_sg U63852 ( .A(n44475), .B(n10412), .X(n10410) );
  nand_x4_sg U63853 ( .A(n14524), .B(n14576), .X(n14570) );
  nand_x1_sg U63854 ( .A(n43339), .B(n14578), .X(n14576) );
  nand_x2_sg U63855 ( .A(n46405), .B(n27369), .X(n27368) );
  nand_x4_sg U63856 ( .A(n52471), .B(n13696), .X(n13677) );
  nand_x1_sg U63857 ( .A(n52470), .B(n13697), .X(n13696) );
  nor_x1_sg U63858 ( .A(n13697), .B(n52470), .X(n13698) );
  nand_x4_sg U63859 ( .A(n17645), .B(n17697), .X(n17691) );
  nand_x1_sg U63860 ( .A(n43335), .B(n17699), .X(n17697) );
  nand_x4_sg U63861 ( .A(n19190), .B(n19242), .X(n19236) );
  nand_x1_sg U63862 ( .A(n43331), .B(n19244), .X(n19242) );
  nand_x4_sg U63863 ( .A(n20734), .B(n20786), .X(n20780) );
  nand_x1_sg U63864 ( .A(n43327), .B(n20788), .X(n20786) );
  nand_x4_sg U63865 ( .A(n17719), .B(n17720), .X(n17692) );
  nand_x1_sg U63866 ( .A(n53932), .B(n42435), .X(n17720) );
  nand_x4_sg U63867 ( .A(n19264), .B(n19265), .X(n19237) );
  nand_x1_sg U63868 ( .A(n54497), .B(n42433), .X(n19265) );
  nand_x4_sg U63869 ( .A(n20808), .B(n20809), .X(n20781) );
  nand_x1_sg U63870 ( .A(n55065), .B(n42431), .X(n20809) );
  nand_x4_sg U63871 ( .A(n16086), .B(n16140), .X(n16138) );
  nand_x1_sg U63872 ( .A(n43305), .B(n16142), .X(n16140) );
  nor_x1_sg U63873 ( .A(n18260), .B(n18223), .X(n18259) );
  nor_x1_sg U63874 ( .A(n46278), .B(n9155), .X(\L2_0/n3096 ) );
  nor_x1_sg U63875 ( .A(n46549), .B(n8893), .X(\L2_0/n4056 ) );
  nor_x1_sg U63876 ( .A(n46505), .B(n8853), .X(\L2_0/n3896 ) );
  nor_x1_sg U63877 ( .A(n46460), .B(n9007), .X(\L2_0/n3736 ) );
  nor_x1_sg U63878 ( .A(n46415), .B(n9343), .X(\L2_0/n3576 ) );
  nor_x1_sg U63879 ( .A(n46370), .B(n9269), .X(\L2_0/n3416 ) );
  nor_x1_sg U63880 ( .A(n46323), .B(n9231), .X(\L2_0/n3256 ) );
  nor_x1_sg U63881 ( .A(n46527), .B(n8919), .X(\L2_0/n3976 ) );
  nor_x1_sg U63882 ( .A(n46303), .B(n9191), .X(\L2_0/n3176 ) );
  nor_x1_sg U63883 ( .A(n46303), .B(n41354), .X(\L2_0/n3164 ) );
  nor_x1_sg U63884 ( .A(n46303), .B(n9195), .X(\L2_0/n3160 ) );
  nor_x1_sg U63885 ( .A(n46303), .B(n9173), .X(\L2_0/n3152 ) );
  nor_x1_sg U63886 ( .A(n46303), .B(n9193), .X(\L2_0/n3148 ) );
  nor_x1_sg U63887 ( .A(n46303), .B(n9183), .X(\L2_0/n3140 ) );
  nor_x1_sg U63888 ( .A(n46303), .B(n9201), .X(\L2_0/n3136 ) );
  nor_x1_sg U63889 ( .A(n46303), .B(n9199), .X(\L2_0/n3124 ) );
  nor_x1_sg U63890 ( .A(n46303), .B(n9171), .X(\L2_0/n3116 ) );
  nor_x1_sg U63891 ( .A(n46303), .B(n9166), .X(\L2_0/n3112 ) );
  nor_x1_sg U63892 ( .A(n46437), .B(n8996), .X(\L2_0/n3656 ) );
  nor_x1_sg U63893 ( .A(n46350), .B(n9077), .X(\L2_0/n3336 ) );
  nor_x1_sg U63894 ( .A(n46350), .B(n42629), .X(\L2_0/n3324 ) );
  nor_x1_sg U63895 ( .A(n46350), .B(n9063), .X(\L2_0/n3320 ) );
  nor_x1_sg U63896 ( .A(n46350), .B(n9069), .X(\L2_0/n3312 ) );
  nor_x1_sg U63897 ( .A(n46350), .B(n9061), .X(\L2_0/n3308 ) );
  nor_x1_sg U63898 ( .A(n46350), .B(n9075), .X(\L2_0/n3300 ) );
  nor_x1_sg U63899 ( .A(n46350), .B(n9067), .X(\L2_0/n3296 ) );
  nor_x1_sg U63900 ( .A(n46350), .B(n9065), .X(\L2_0/n3284 ) );
  nor_x1_sg U63901 ( .A(n46350), .B(n9081), .X(\L2_0/n3276 ) );
  nor_x1_sg U63902 ( .A(n46350), .B(n9054), .X(\L2_0/n3272 ) );
  nor_x1_sg U63903 ( .A(n46483), .B(n8809), .X(\L2_0/n3816 ) );
  nor_x1_sg U63904 ( .A(n46393), .B(n9307), .X(\L2_0/n3496 ) );
  nor_x1_sg U63905 ( .A(n46258), .B(n9103), .X(\L2_0/n3016 ) );
  nand_x4_sg U63906 ( .A(n51766), .B(n11813), .X(n11798) );
  nand_x1_sg U63907 ( .A(n51744), .B(n51609), .X(n11814) );
  nand_x4_sg U63908 ( .A(n52322), .B(n13370), .X(n13355) );
  nand_x1_sg U63909 ( .A(n52301), .B(n52167), .X(n13371) );
  nand_x4_sg U63910 ( .A(n53156), .B(n15703), .X(n15688) );
  nand_x1_sg U63911 ( .A(n53135), .B(n53001), .X(n15704) );
  nand_x4_sg U63912 ( .A(n53714), .B(n17269), .X(n17254) );
  nand_x1_sg U63913 ( .A(n53693), .B(n53559), .X(n17270) );
  nand_x4_sg U63914 ( .A(n52597), .B(n14150), .X(n14135) );
  nand_x1_sg U63915 ( .A(n52576), .B(n52441), .X(n14151) );
  nand_x4_sg U63916 ( .A(n53436), .B(n16488), .X(n16473) );
  nand_x1_sg U63917 ( .A(n53413), .B(n53277), .X(n16489) );
  nand_x4_sg U63918 ( .A(n52875), .B(n14925), .X(n14911) );
  nand_x4_sg U63919 ( .A(n53995), .B(n18046), .X(n18032) );
  nand_x4_sg U63920 ( .A(n54560), .B(n19591), .X(n19577) );
  nand_x4_sg U63921 ( .A(n55128), .B(n21135), .X(n21121) );
  nand_x4_sg U63922 ( .A(n51698), .B(n11468), .X(n11411) );
  nand_x1_sg U63923 ( .A(n51658), .B(n11469), .X(n11468) );
  nand_x4_sg U63924 ( .A(n52254), .B(n13029), .X(n12972) );
  nand_x1_sg U63925 ( .A(n52214), .B(n13030), .X(n13029) );
  nand_x4_sg U63926 ( .A(n53088), .B(n15362), .X(n15305) );
  nand_x1_sg U63927 ( .A(n53048), .B(n15363), .X(n15362) );
  nand_x4_sg U63928 ( .A(n53646), .B(n16928), .X(n16871) );
  nand_x1_sg U63929 ( .A(n53606), .B(n16929), .X(n16928) );
  nand_x4_sg U63930 ( .A(n13597), .B(n13598), .X(n13585) );
  nor_x1_sg U63931 ( .A(n13577), .B(n13607), .X(n13597) );
  nor_x1_sg U63932 ( .A(n13599), .B(n46480), .X(n13598) );
  nand_x4_sg U63933 ( .A(n54810), .B(n20127), .X(n20100) );
  nand_x1_sg U63934 ( .A(n54690), .B(n20129), .X(n20128) );
  nand_x4_sg U63935 ( .A(n55378), .B(n21672), .X(n21645) );
  nand_x1_sg U63936 ( .A(n55258), .B(n21674), .X(n21673) );
  nand_x4_sg U63937 ( .A(n51591), .B(n11209), .X(n11153) );
  nand_x4_sg U63938 ( .A(n52149), .B(n12770), .X(n12714) );
  nand_x4_sg U63939 ( .A(n52983), .B(n15103), .X(n15047) );
  nand_x4_sg U63940 ( .A(n53541), .B(n16669), .X(n16613) );
  nand_x4_sg U63941 ( .A(n54259), .B(n18620), .X(n18607) );
  nand_x1_sg U63942 ( .A(n54195), .B(n54169), .X(n18621) );
  nand_x4_sg U63943 ( .A(n53975), .B(n17853), .X(n17840) );
  nand_x1_sg U63944 ( .A(n53904), .B(n53887), .X(n17854) );
  nand_x4_sg U63945 ( .A(n54540), .B(n19398), .X(n19385) );
  nand_x1_sg U63946 ( .A(n54469), .B(n54452), .X(n19399) );
  nand_x4_sg U63947 ( .A(n55108), .B(n20942), .X(n20929) );
  nand_x1_sg U63948 ( .A(n55037), .B(n55020), .X(n20943) );
  nand_x4_sg U63949 ( .A(n53415), .B(n16296), .X(n16283) );
  nand_x1_sg U63950 ( .A(n53341), .B(n53330), .X(n16297) );
  nand_x4_sg U63951 ( .A(n54826), .B(n20166), .X(n20153) );
  nand_x1_sg U63952 ( .A(n54762), .B(n54735), .X(n20167) );
  nand_x4_sg U63953 ( .A(n55394), .B(n21711), .X(n21698) );
  nand_x1_sg U63954 ( .A(n55330), .B(n55303), .X(n21712) );
  nand_x4_sg U63955 ( .A(n52028), .B(n12401), .X(n12388) );
  nand_x1_sg U63956 ( .A(n51953), .B(n51942), .X(n12402) );
  nand_x4_sg U63957 ( .A(n53258), .B(n15883), .X(n15831) );
  nand_x4_sg U63958 ( .A(n51871), .B(n11988), .X(n11936) );
  nand_x4_sg U63959 ( .A(n52855), .B(n14732), .X(n14719) );
  nand_x1_sg U63960 ( .A(n52784), .B(n52767), .X(n14733) );
  nand_x4_sg U63961 ( .A(n54170), .B(n18822), .X(n18787) );
  nand_x1_sg U63962 ( .A(n18785), .B(n18823), .X(n18822) );
  nor_x1_sg U63963 ( .A(n18823), .B(n18785), .X(n18824) );
  nand_x4_sg U63964 ( .A(n54736), .B(n20367), .X(n20333) );
  nand_x1_sg U63965 ( .A(n20331), .B(n20368), .X(n20367) );
  nor_x1_sg U63966 ( .A(n20368), .B(n20331), .X(n20369) );
  nand_x4_sg U63967 ( .A(n55304), .B(n21912), .X(n21878) );
  nand_x1_sg U63968 ( .A(n21876), .B(n21913), .X(n21912) );
  nor_x1_sg U63969 ( .A(n21913), .B(n21876), .X(n21914) );
  nand_x4_sg U63970 ( .A(n51746), .B(n11620), .X(n11607) );
  nand_x1_sg U63971 ( .A(n51672), .B(n51661), .X(n11621) );
  nand_x4_sg U63972 ( .A(n52303), .B(n13181), .X(n13168) );
  nand_x1_sg U63973 ( .A(n52228), .B(n52217), .X(n13182) );
  nand_x4_sg U63974 ( .A(n53137), .B(n15514), .X(n15501) );
  nand_x1_sg U63975 ( .A(n53062), .B(n53051), .X(n15515) );
  nand_x4_sg U63976 ( .A(n53695), .B(n17080), .X(n17067) );
  nand_x1_sg U63977 ( .A(n53620), .B(n53609), .X(n17081) );
  nand_x4_sg U63978 ( .A(n52744), .B(n14473), .X(n14458) );
  nand_x1_sg U63979 ( .A(n52743), .B(n14474), .X(n14473) );
  nor_x1_sg U63980 ( .A(n14474), .B(n52743), .X(n14475) );
  nand_x2_sg U63981 ( .A(n46363), .B(n27922), .X(n27921) );
  nand_x2_sg U63982 ( .A(n46316), .B(n28480), .X(n28479) );
  nand_x2_sg U63983 ( .A(n46271), .B(n29039), .X(n29038) );
  nand_x4_sg U63984 ( .A(n12034), .B(n12033), .X(n12035) );
  nor_x1_sg U63985 ( .A(n10989), .B(n10990), .X(n10986) );
  nand_x1_sg U63986 ( .A(n10988), .B(n10985), .X(n10987) );
  nand_x4_sg U63987 ( .A(n53848), .B(n17860), .X(n18045) );
  nand_x4_sg U63988 ( .A(n54413), .B(n19405), .X(n19590) );
  nand_x4_sg U63989 ( .A(n54981), .B(n20949), .X(n21134) );
  nand_x4_sg U63990 ( .A(n52014), .B(n12566), .X(n12557) );
  nand_x4_sg U63991 ( .A(n53286), .B(n16303), .X(n16487) );
  nand_x1_sg U63992 ( .A(n43953), .B(n8050), .X(n9048) );
  nand_x1_sg U63993 ( .A(n44401), .B(n8050), .X(n9042) );
  nand_x1_sg U63994 ( .A(n11062), .B(n11061), .X(n11059) );
  nor_x1_sg U63995 ( .A(n11061), .B(n11062), .X(n11060) );
  nand_x4_sg U63996 ( .A(n11779), .B(n11780), .X(n11760) );
  nand_x1_sg U63997 ( .A(n11783), .B(n51664), .X(n11779) );
  nand_x1_sg U63998 ( .A(n11781), .B(n11782), .X(n11780) );
  nand_x4_sg U63999 ( .A(n18298), .B(n54115), .X(n18263) );
  nand_x1_sg U64000 ( .A(n18300), .B(n18260), .X(n18298) );
  nor_x1_sg U64001 ( .A(n18260), .B(n18300), .X(n18299) );
  nor_x1_sg U64002 ( .A(n46231), .B(n25464), .X(n25473) );
  nor_x1_sg U64003 ( .A(n44209), .B(n17425), .X(n17423) );
  nor_x1_sg U64004 ( .A(n44207), .B(n18970), .X(n18968) );
  nor_x1_sg U64005 ( .A(n44205), .B(n20514), .X(n20512) );
  nand_x2_sg U64006 ( .A(n46564), .B(n25415), .X(n25414) );
  nand_x1_sg U64007 ( .A(n12623), .B(n12622), .X(n12620) );
  nor_x1_sg U64008 ( .A(n12622), .B(n12623), .X(n12621) );
  nand_x1_sg U64009 ( .A(n14956), .B(n14955), .X(n14953) );
  nor_x1_sg U64010 ( .A(n14955), .B(n14956), .X(n14954) );
  nand_x1_sg U64011 ( .A(n16522), .B(n16521), .X(n16519) );
  nor_x1_sg U64012 ( .A(n16521), .B(n16522), .X(n16520) );
  nand_x4_sg U64013 ( .A(n11669), .B(n51800), .X(n11667) );
  nand_x1_sg U64014 ( .A(n11672), .B(n44341), .X(n11669) );
  nor_x1_sg U64015 ( .A(n44341), .B(n11672), .X(n11670) );
  nand_x4_sg U64016 ( .A(n12449), .B(n52076), .X(n12447) );
  nand_x1_sg U64017 ( .A(n12452), .B(n44339), .X(n12449) );
  nor_x1_sg U64018 ( .A(n44339), .B(n12452), .X(n12450) );
  nand_x4_sg U64019 ( .A(n13230), .B(n52354), .X(n13228) );
  nand_x1_sg U64020 ( .A(n13233), .B(n43971), .X(n13230) );
  nor_x1_sg U64021 ( .A(n43971), .B(n13233), .X(n13231) );
  nand_x4_sg U64022 ( .A(n14010), .B(n52629), .X(n14008) );
  nand_x1_sg U64023 ( .A(n14013), .B(n43969), .X(n14010) );
  nor_x1_sg U64024 ( .A(n43969), .B(n14013), .X(n14011) );
  nand_x4_sg U64025 ( .A(n14781), .B(n52910), .X(n14779) );
  nand_x1_sg U64026 ( .A(n14784), .B(n44337), .X(n14781) );
  nor_x1_sg U64027 ( .A(n44337), .B(n14784), .X(n14782) );
  nand_x4_sg U64028 ( .A(n15563), .B(n53188), .X(n15561) );
  nand_x1_sg U64029 ( .A(n15566), .B(n43967), .X(n15563) );
  nor_x1_sg U64030 ( .A(n43967), .B(n15566), .X(n15564) );
  nand_x4_sg U64031 ( .A(n17129), .B(n53746), .X(n17127) );
  nand_x1_sg U64032 ( .A(n17132), .B(n43965), .X(n17129) );
  nor_x1_sg U64033 ( .A(n43965), .B(n17132), .X(n17130) );
  nand_x4_sg U64034 ( .A(n17902), .B(n54030), .X(n17900) );
  nand_x1_sg U64035 ( .A(n17905), .B(n43963), .X(n17902) );
  nor_x1_sg U64036 ( .A(n43963), .B(n17905), .X(n17903) );
  nand_x4_sg U64037 ( .A(n18671), .B(n54311), .X(n18669) );
  nand_x1_sg U64038 ( .A(n18674), .B(n44335), .X(n18671) );
  nor_x1_sg U64039 ( .A(n44335), .B(n18674), .X(n18672) );
  nand_x4_sg U64040 ( .A(n19447), .B(n54595), .X(n19445) );
  nand_x1_sg U64041 ( .A(n19450), .B(n43961), .X(n19447) );
  nor_x1_sg U64042 ( .A(n43961), .B(n19450), .X(n19448) );
  nand_x4_sg U64043 ( .A(n20216), .B(n54879), .X(n20214) );
  nand_x1_sg U64044 ( .A(n20219), .B(n43959), .X(n20216) );
  nor_x1_sg U64045 ( .A(n43959), .B(n20219), .X(n20217) );
  nand_x4_sg U64046 ( .A(n20991), .B(n55163), .X(n20989) );
  nand_x1_sg U64047 ( .A(n20994), .B(n43957), .X(n20991) );
  nor_x1_sg U64048 ( .A(n43957), .B(n20994), .X(n20992) );
  nand_x4_sg U64049 ( .A(n21761), .B(n55447), .X(n21759) );
  nand_x1_sg U64050 ( .A(n21764), .B(n43955), .X(n21761) );
  nor_x1_sg U64051 ( .A(n43955), .B(n21764), .X(n21762) );
  nand_x4_sg U64052 ( .A(n14909), .B(n14910), .X(n14907) );
  nand_x1_sg U64053 ( .A(n52727), .B(n14891), .X(n14910) );
  nand_x4_sg U64054 ( .A(n16471), .B(n16472), .X(n16470) );
  nand_x1_sg U64055 ( .A(n53285), .B(n16453), .X(n16472) );
  nand_x4_sg U64056 ( .A(n18030), .B(n18031), .X(n18028) );
  nand_x1_sg U64057 ( .A(n53847), .B(n18012), .X(n18031) );
  nand_x4_sg U64058 ( .A(n19575), .B(n19576), .X(n19573) );
  nand_x1_sg U64059 ( .A(n54412), .B(n19557), .X(n19576) );
  nand_x4_sg U64060 ( .A(n20345), .B(n20346), .X(n20343) );
  nand_x1_sg U64061 ( .A(n54691), .B(n20327), .X(n20346) );
  nand_x4_sg U64062 ( .A(n21119), .B(n21120), .X(n21117) );
  nand_x1_sg U64063 ( .A(n54980), .B(n21101), .X(n21120) );
  nand_x4_sg U64064 ( .A(n21890), .B(n21891), .X(n21888) );
  nand_x1_sg U64065 ( .A(n55259), .B(n21872), .X(n21891) );
  nand_x4_sg U64066 ( .A(n18264), .B(n18292), .X(n18285) );
  nor_x1_sg U64067 ( .A(n46353), .B(n18260), .X(n18293) );
  nand_x4_sg U64068 ( .A(n14892), .B(n14893), .X(n14872) );
  nand_x1_sg U64069 ( .A(n14896), .B(n52770), .X(n14892) );
  nand_x1_sg U64070 ( .A(n14894), .B(n14895), .X(n14893) );
  nand_x4_sg U64071 ( .A(n11587), .B(n11588), .X(n11531) );
  nand_x1_sg U64072 ( .A(n11590), .B(n51708), .X(n11587) );
  nand_x1_sg U64073 ( .A(n11589), .B(n51612), .X(n11588) );
  nand_x4_sg U64074 ( .A(n13148), .B(n13149), .X(n13092) );
  nand_x1_sg U64075 ( .A(n13151), .B(n52264), .X(n13148) );
  nand_x1_sg U64076 ( .A(n13150), .B(n52170), .X(n13149) );
  nand_x4_sg U64077 ( .A(n13928), .B(n13929), .X(n13872) );
  nand_x1_sg U64078 ( .A(n13931), .B(n52540), .X(n13928) );
  nand_x1_sg U64079 ( .A(n13930), .B(n52444), .X(n13929) );
  nand_x4_sg U64080 ( .A(n15481), .B(n15482), .X(n15425) );
  nand_x1_sg U64081 ( .A(n15484), .B(n53098), .X(n15481) );
  nand_x1_sg U64082 ( .A(n15483), .B(n53004), .X(n15482) );
  nand_x4_sg U64083 ( .A(n17047), .B(n17048), .X(n16991) );
  nand_x1_sg U64084 ( .A(n17050), .B(n53656), .X(n17047) );
  nand_x1_sg U64085 ( .A(n17049), .B(n53562), .X(n17048) );
  nand_x4_sg U64086 ( .A(n18697), .B(n54274), .X(n18674) );
  nand_x1_sg U64087 ( .A(n54251), .B(n18699), .X(n18697) );
  nor_x1_sg U64088 ( .A(n18699), .B(n54251), .X(n18698) );
  nand_x4_sg U64089 ( .A(n14825), .B(n52892), .X(n14823) );
  nand_x1_sg U64090 ( .A(n52891), .B(n14827), .X(n14825) );
  nor_x1_sg U64091 ( .A(n14827), .B(n52891), .X(n14826) );
  nand_x4_sg U64092 ( .A(n17946), .B(n54012), .X(n17944) );
  nand_x1_sg U64093 ( .A(n54011), .B(n17948), .X(n17946) );
  nor_x1_sg U64094 ( .A(n17948), .B(n54011), .X(n17947) );
  nand_x4_sg U64095 ( .A(n19491), .B(n54577), .X(n19489) );
  nand_x1_sg U64096 ( .A(n54576), .B(n19493), .X(n19491) );
  nor_x1_sg U64097 ( .A(n19493), .B(n54576), .X(n19492) );
  nand_x4_sg U64098 ( .A(n21035), .B(n55145), .X(n21033) );
  nand_x1_sg U64099 ( .A(n55144), .B(n21037), .X(n21035) );
  nor_x1_sg U64100 ( .A(n21037), .B(n55144), .X(n21036) );
  nor_x1_sg U64101 ( .A(n18777), .B(n18778), .X(n18773) );
  nand_x1_sg U64102 ( .A(n18775), .B(n18776), .X(n18774) );
  nor_x1_sg U64103 ( .A(n16448), .B(n16449), .X(n16445) );
  nand_x1_sg U64104 ( .A(n16447), .B(n16444), .X(n16446) );
  nand_x4_sg U64105 ( .A(n54277), .B(n18820), .X(n18811) );
  nand_x1_sg U64106 ( .A(n54171), .B(n18786), .X(n18820) );
  nor_x1_sg U64107 ( .A(n54171), .B(n18786), .X(n18821) );
  nand_x4_sg U64108 ( .A(n54844), .B(n20365), .X(n20356) );
  nand_x1_sg U64109 ( .A(n54737), .B(n20332), .X(n20365) );
  nor_x1_sg U64110 ( .A(n54737), .B(n20332), .X(n20366) );
  nand_x4_sg U64111 ( .A(n55412), .B(n21910), .X(n21901) );
  nand_x1_sg U64112 ( .A(n55305), .B(n21877), .X(n21910) );
  nor_x1_sg U64113 ( .A(n55305), .B(n21877), .X(n21911) );
  nor_x1_sg U64114 ( .A(n20323), .B(n20324), .X(n20320) );
  nand_x1_sg U64115 ( .A(n20322), .B(n54778), .X(n20321) );
  nor_x1_sg U64116 ( .A(n21868), .B(n21869), .X(n21865) );
  nand_x1_sg U64117 ( .A(n21867), .B(n55346), .X(n21866) );
  nand_x4_sg U64118 ( .A(n17412), .B(n17413), .X(n17410) );
  nand_x1_sg U64119 ( .A(n17415), .B(n17416), .X(n17412) );
  nor_x1_sg U64120 ( .A(n17415), .B(n46367), .X(n17414) );
  nand_x4_sg U64121 ( .A(n18957), .B(n18958), .X(n18955) );
  nand_x1_sg U64122 ( .A(n18960), .B(n18961), .X(n18957) );
  nor_x1_sg U64123 ( .A(n18960), .B(n46320), .X(n18959) );
  nand_x4_sg U64124 ( .A(n20501), .B(n20502), .X(n20499) );
  nand_x1_sg U64125 ( .A(n20504), .B(n20505), .X(n20501) );
  nor_x1_sg U64126 ( .A(n20504), .B(n46275), .X(n20503) );
  nand_x4_sg U64127 ( .A(n29330), .B(n29331), .X(n29329) );
  nor_x1_sg U64128 ( .A(n55212), .B(n29332), .X(n29331) );
  nor_x1_sg U64129 ( .A(n29336), .B(n46236), .X(n29330) );
  nand_x4_sg U64130 ( .A(n52509), .B(n13782), .X(n13763) );
  nand_x1_sg U64131 ( .A(n52508), .B(n13783), .X(n13782) );
  nor_x1_sg U64132 ( .A(n52508), .B(n13783), .X(n13784) );
  nand_x4_sg U64133 ( .A(n14642), .B(n14641), .X(n14693) );
  nand_x4_sg U64134 ( .A(n17763), .B(n17762), .X(n17814) );
  nand_x4_sg U64135 ( .A(n18531), .B(n18530), .X(n18580) );
  nand_x4_sg U64136 ( .A(n19308), .B(n19307), .X(n19359) );
  nand_x4_sg U64137 ( .A(n20852), .B(n20851), .X(n20903) );
  nand_x1_sg U64138 ( .A(n42435), .B(n17722), .X(n17788) );
  nand_x1_sg U64139 ( .A(n42433), .B(n19267), .X(n19333) );
  nand_x1_sg U64140 ( .A(n42431), .B(n20811), .X(n20877) );
  nand_x4_sg U64141 ( .A(n51486), .B(n11033), .X(n11024) );
  nand_x1_sg U64142 ( .A(n51383), .B(n10999), .X(n11033) );
  nor_x1_sg U64143 ( .A(n51383), .B(n10999), .X(n11034) );
  nand_x4_sg U64144 ( .A(n51957), .B(n12221), .X(n12202) );
  nand_x1_sg U64145 ( .A(n51956), .B(n12222), .X(n12221) );
  nor_x1_sg U64146 ( .A(n51956), .B(n12222), .X(n12223) );
  nand_x4_sg U64147 ( .A(n14314), .B(n14315), .X(n14304) );
  nand_x1_sg U64148 ( .A(n14317), .B(n14316), .X(n14314) );
  nand_x1_sg U64149 ( .A(n52662), .B(n52658), .X(n14315) );
  nand_x4_sg U64150 ( .A(n53345), .B(n16116), .X(n16097) );
  nand_x1_sg U64151 ( .A(n53344), .B(n16117), .X(n16116) );
  nor_x1_sg U64152 ( .A(n53344), .B(n16117), .X(n16118) );
  nand_x4_sg U64153 ( .A(n51676), .B(n11441), .X(n11422) );
  nand_x1_sg U64154 ( .A(n51675), .B(n11442), .X(n11441) );
  nor_x1_sg U64155 ( .A(n51675), .B(n11442), .X(n11443) );
  nand_x4_sg U64156 ( .A(n52232), .B(n13002), .X(n12983) );
  nand_x1_sg U64157 ( .A(n52231), .B(n13003), .X(n13002) );
  nor_x1_sg U64158 ( .A(n52231), .B(n13003), .X(n13004) );
  nand_x4_sg U64159 ( .A(n53066), .B(n15335), .X(n15316) );
  nand_x1_sg U64160 ( .A(n53065), .B(n15336), .X(n15335) );
  nor_x1_sg U64161 ( .A(n53065), .B(n15336), .X(n15337) );
  nand_x4_sg U64162 ( .A(n53624), .B(n16901), .X(n16882) );
  nand_x1_sg U64163 ( .A(n53623), .B(n16902), .X(n16901) );
  nor_x1_sg U64164 ( .A(n53623), .B(n16902), .X(n16903) );
  nand_x1_sg U64165 ( .A(n14886), .B(n52809), .X(n14885) );
  nor_x1_sg U64166 ( .A(n14887), .B(n14888), .X(n14884) );
  nand_x1_sg U64167 ( .A(n13830), .B(n41845), .X(n13898) );
  nand_x4_sg U64168 ( .A(n18470), .B(n18471), .X(n18400) );
  nand_x1_sg U64169 ( .A(n54166), .B(n18420), .X(n18471) );
  nand_x4_sg U64170 ( .A(n12258), .B(n12259), .X(n12194) );
  nand_x1_sg U64171 ( .A(n43310), .B(n12247), .X(n12258) );
  nand_x1_sg U64172 ( .A(n51927), .B(n43311), .X(n12259) );
  nand_x4_sg U64173 ( .A(n52728), .B(n14739), .X(n14924) );
  nand_x1_sg U64174 ( .A(n42006), .B(n8050), .X(n9025) );
  nand_x1_sg U64175 ( .A(n42893), .B(n46577), .X(n9021) );
  nand_x4_sg U64176 ( .A(n42624), .B(n17313), .X(n17320) );
  nand_x4_sg U64177 ( .A(n18169), .B(n18085), .X(n18092) );
  nand_x4_sg U64178 ( .A(n42622), .B(n18858), .X(n18865) );
  nand_x4_sg U64179 ( .A(n42620), .B(n20402), .X(n20409) );
  nor_x1_sg U64180 ( .A(n11774), .B(n11775), .X(n11770) );
  nand_x1_sg U64181 ( .A(n11772), .B(n11773), .X(n11771) );
  nand_x4_sg U64182 ( .A(n14279), .B(n14194), .X(n14201) );
  nand_x4_sg U64183 ( .A(n11937), .B(n11853), .X(n11860) );
  nand_x4_sg U64184 ( .A(n15832), .B(n15748), .X(n15755) );
  nand_x4_sg U64185 ( .A(n42617), .B(n11070), .X(n11077) );
  nand_x4_sg U64186 ( .A(n42615), .B(n12631), .X(n12638) );
  nand_x4_sg U64187 ( .A(n42613), .B(n14964), .X(n14971) );
  nand_x4_sg U64188 ( .A(n42611), .B(n16530), .X(n16537) );
  nand_x4_sg U64189 ( .A(n42605), .B(n10302), .X(n10309) );
  nand_x4_sg U64190 ( .A(n42609), .B(n19630), .X(n19637) );
  nand_x4_sg U64191 ( .A(n42607), .B(n21175), .X(n21182) );
  nand_x4_sg U64192 ( .A(n11537), .B(n11538), .X(n11507) );
  nand_x1_sg U64193 ( .A(n42111), .B(n51747), .X(n11538) );
  nand_x1_sg U64194 ( .A(n40543), .B(n11540), .X(n11537) );
  nand_x4_sg U64195 ( .A(n14647), .B(n14648), .X(n14618) );
  nand_x1_sg U64196 ( .A(n42121), .B(n52856), .X(n14648) );
  nand_x1_sg U64197 ( .A(n40551), .B(n14650), .X(n14647) );
  nand_x4_sg U64198 ( .A(n16212), .B(n16213), .X(n16182) );
  nand_x1_sg U64199 ( .A(n42071), .B(n53416), .X(n16213) );
  nand_x1_sg U64200 ( .A(n40554), .B(n16215), .X(n16212) );
  nand_x4_sg U64201 ( .A(n12317), .B(n12318), .X(n12287) );
  nand_x1_sg U64202 ( .A(n42109), .B(n52029), .X(n12318) );
  nand_x1_sg U64203 ( .A(n40544), .B(n12320), .X(n12317) );
  nand_x4_sg U64204 ( .A(n12377), .B(n12378), .X(n12335) );
  nand_x1_sg U64205 ( .A(n42133), .B(n52047), .X(n12378) );
  nand_x1_sg U64206 ( .A(n40532), .B(n12380), .X(n12377) );
  nand_x4_sg U64207 ( .A(n13098), .B(n13099), .X(n13068) );
  nand_x1_sg U64208 ( .A(n42107), .B(n52304), .X(n13099) );
  nand_x1_sg U64209 ( .A(n40546), .B(n13101), .X(n13098) );
  nand_x4_sg U64210 ( .A(n15431), .B(n15432), .X(n15401) );
  nand_x1_sg U64211 ( .A(n42103), .B(n53138), .X(n15432) );
  nand_x1_sg U64212 ( .A(n40552), .B(n15434), .X(n15431) );
  nand_x4_sg U64213 ( .A(n16997), .B(n16998), .X(n16967) );
  nand_x1_sg U64214 ( .A(n42101), .B(n53696), .X(n16998) );
  nand_x1_sg U64215 ( .A(n40555), .B(n17000), .X(n16997) );
  nand_x4_sg U64216 ( .A(n17768), .B(n17769), .X(n17739) );
  nand_x1_sg U64217 ( .A(n42117), .B(n53976), .X(n17769) );
  nand_x1_sg U64218 ( .A(n40557), .B(n17771), .X(n17768) );
  nand_x4_sg U64219 ( .A(n19313), .B(n19314), .X(n19284) );
  nand_x1_sg U64220 ( .A(n42115), .B(n54541), .X(n19314) );
  nand_x1_sg U64221 ( .A(n40559), .B(n19316), .X(n19313) );
  nand_x4_sg U64222 ( .A(n20857), .B(n20858), .X(n20828) );
  nand_x1_sg U64223 ( .A(n42113), .B(n55109), .X(n20858) );
  nand_x1_sg U64224 ( .A(n40560), .B(n20860), .X(n20857) );
  nand_x4_sg U64225 ( .A(n13514), .B(n13515), .X(n13414) );
  nand_x1_sg U64226 ( .A(n44325), .B(n52388), .X(n13515) );
  nand_x1_sg U64227 ( .A(n52394), .B(n13517), .X(n13514) );
  nand_x4_sg U64228 ( .A(n14619), .B(n52826), .X(n14575) );
  nor_x1_sg U64229 ( .A(n44447), .B(n14639), .X(n14637) );
  nand_x4_sg U64230 ( .A(n17740), .B(n53946), .X(n17696) );
  nor_x1_sg U64231 ( .A(n44445), .B(n17760), .X(n17758) );
  nand_x4_sg U64232 ( .A(n18509), .B(n54231), .X(n18465) );
  nor_x1_sg U64233 ( .A(n44211), .B(n18528), .X(n18526) );
  nand_x4_sg U64234 ( .A(n19285), .B(n54511), .X(n19241) );
  nor_x1_sg U64235 ( .A(n44443), .B(n19305), .X(n19303) );
  nand_x4_sg U64236 ( .A(n20829), .B(n55079), .X(n20785) );
  nor_x1_sg U64237 ( .A(n44441), .B(n20849), .X(n20847) );
  nand_x4_sg U64238 ( .A(n20054), .B(n54796), .X(n20010) );
  nor_x1_sg U64239 ( .A(n44465), .B(n20073), .X(n20071) );
  nand_x4_sg U64240 ( .A(n21599), .B(n55364), .X(n21555) );
  nor_x1_sg U64241 ( .A(n44463), .B(n21618), .X(n21616) );
  nand_x4_sg U64242 ( .A(n10727), .B(n51437), .X(n10683) );
  nor_x1_sg U64243 ( .A(n44467), .B(n10747), .X(n10745) );
  nand_x4_sg U64244 ( .A(n11525), .B(n11526), .X(n11460) );
  nand_x1_sg U64245 ( .A(n51711), .B(n45413), .X(n11526) );
  nand_x1_sg U64246 ( .A(n51719), .B(n44150), .X(n11525) );
  nand_x4_sg U64247 ( .A(n13086), .B(n13087), .X(n13021) );
  nand_x1_sg U64248 ( .A(n52267), .B(n45411), .X(n13087) );
  nand_x1_sg U64249 ( .A(n52273), .B(n44148), .X(n13086) );
  nand_x4_sg U64250 ( .A(n15419), .B(n15420), .X(n15354) );
  nand_x1_sg U64251 ( .A(n53101), .B(n45407), .X(n15420) );
  nand_x1_sg U64252 ( .A(n53107), .B(n44144), .X(n15419) );
  nand_x4_sg U64253 ( .A(n16985), .B(n16986), .X(n16920) );
  nand_x1_sg U64254 ( .A(n53659), .B(n45405), .X(n16986) );
  nand_x1_sg U64255 ( .A(n53665), .B(n44142), .X(n16985) );
  nor_x1_sg U64256 ( .A(n18008), .B(n18009), .X(n18005) );
  nand_x1_sg U64257 ( .A(n18007), .B(n53929), .X(n18006) );
  nor_x1_sg U64258 ( .A(n19553), .B(n19554), .X(n19550) );
  nand_x1_sg U64259 ( .A(n19552), .B(n54494), .X(n19551) );
  nor_x1_sg U64260 ( .A(n21097), .B(n21098), .X(n21094) );
  nand_x1_sg U64261 ( .A(n21096), .B(n55062), .X(n21095) );
  nand_x4_sg U64262 ( .A(n12496), .B(n12497), .X(n12495) );
  nand_x1_sg U64263 ( .A(n41916), .B(n12500), .X(n12496) );
  nor_x1_sg U64264 ( .A(n52020), .B(n51992), .X(n12498) );
  nand_x4_sg U64265 ( .A(n20076), .B(n20075), .X(n20126) );
  nand_x4_sg U64266 ( .A(n21621), .B(n21620), .X(n21671) );
  nand_x2_sg U64267 ( .A(n46474), .B(n26532), .X(n26531) );
  nor_x1_sg U64268 ( .A(n43139), .B(n18228), .X(n18226) );
  nand_x4_sg U64269 ( .A(n10697), .B(n10698), .X(n10635) );
  nand_x1_sg U64270 ( .A(n43314), .B(n10686), .X(n10697) );
  nand_x1_sg U64271 ( .A(n51371), .B(n43315), .X(n10698) );
  nand_x4_sg U64272 ( .A(n20024), .B(n20025), .X(n19962) );
  nand_x1_sg U64273 ( .A(n43322), .B(n20013), .X(n20024) );
  nand_x1_sg U64274 ( .A(n54725), .B(n43323), .X(n20025) );
  nand_x4_sg U64275 ( .A(n21569), .B(n21570), .X(n21507) );
  nand_x1_sg U64276 ( .A(n43318), .B(n21558), .X(n21569) );
  nand_x1_sg U64277 ( .A(n55293), .B(n43319), .X(n21570) );
  nand_x4_sg U64278 ( .A(n17949), .B(n17950), .X(n17948) );
  nand_x1_sg U64279 ( .A(n41908), .B(n17954), .X(n17949) );
  nor_x1_sg U64280 ( .A(n53986), .B(n53928), .X(n17951) );
  nand_x4_sg U64281 ( .A(n19494), .B(n19495), .X(n19493) );
  nand_x1_sg U64282 ( .A(n41900), .B(n19499), .X(n19494) );
  nor_x1_sg U64283 ( .A(n54551), .B(n54493), .X(n19496) );
  nand_x4_sg U64284 ( .A(n21038), .B(n21039), .X(n21037) );
  nand_x1_sg U64285 ( .A(n41894), .B(n21043), .X(n21038) );
  nor_x1_sg U64286 ( .A(n55119), .B(n55061), .X(n21040) );
  nor_x1_sg U64287 ( .A(n42853), .B(n10447), .X(n10445) );
  nor_x1_sg U64288 ( .A(n42855), .B(n14339), .X(n14337) );
  nor_x1_sg U64289 ( .A(n43135), .B(n19774), .X(n19772) );
  nor_x1_sg U64290 ( .A(n43131), .B(n21319), .X(n21317) );
  nand_x4_sg U64291 ( .A(n13789), .B(n13788), .X(n13786) );
  nand_x4_sg U64292 ( .A(n14560), .B(n14559), .X(n14557) );
  nand_x4_sg U64293 ( .A(n17681), .B(n17680), .X(n17678) );
  nand_x4_sg U64294 ( .A(n19226), .B(n19225), .X(n19223) );
  nand_x4_sg U64295 ( .A(n20770), .B(n20769), .X(n20767) );
  nand_x4_sg U64296 ( .A(n12557), .B(n12564), .X(n12422) );
  nand_x1_sg U64297 ( .A(n52021), .B(n12565), .X(n12564) );
  nand_x4_sg U64298 ( .A(n13588), .B(n13587), .X(n13589) );
  nand_x4_sg U64299 ( .A(n53805), .B(n45420), .X(n17313) );
  nand_x4_sg U64300 ( .A(n54370), .B(n45419), .X(n18858) );
  nand_x4_sg U64301 ( .A(n54938), .B(n45418), .X(n20402) );
  nand_x4_sg U64302 ( .A(n14589), .B(n14590), .X(n14527) );
  nand_x1_sg U64303 ( .A(n43338), .B(n14578), .X(n14589) );
  nand_x1_sg U64304 ( .A(n52759), .B(n43339), .X(n14590) );
  nand_x4_sg U64305 ( .A(n51578), .B(n11073), .X(n11070) );
  nand_x4_sg U64306 ( .A(n52136), .B(n12634), .X(n12631) );
  nand_x4_sg U64307 ( .A(n52970), .B(n14967), .X(n14964) );
  nand_x4_sg U64308 ( .A(n53528), .B(n16533), .X(n16530) );
  nand_x4_sg U64309 ( .A(n10755), .B(n10756), .X(n10726) );
  nand_x1_sg U64310 ( .A(n51414), .B(n51467), .X(n10756) );
  nand_x4_sg U64311 ( .A(n18536), .B(n18537), .X(n18508) );
  nand_x1_sg U64312 ( .A(n54198), .B(n54260), .X(n18537) );
  nand_x4_sg U64313 ( .A(n20081), .B(n20082), .X(n20053) );
  nand_x1_sg U64314 ( .A(n54765), .B(n54827), .X(n20082) );
  nand_x4_sg U64315 ( .A(n21626), .B(n21627), .X(n21598) );
  nand_x1_sg U64316 ( .A(n55333), .B(n55395), .X(n21627) );
  nand_x4_sg U64317 ( .A(n17313), .B(n17314), .X(n9273) );
  nand_x4_sg U64318 ( .A(n18858), .B(n18859), .X(n9235) );
  nand_x4_sg U64319 ( .A(n20402), .B(n20403), .X(n9159) );
  nand_x4_sg U64320 ( .A(n11070), .B(n11071), .X(n8886) );
  nand_x4_sg U64321 ( .A(n12631), .B(n12632), .X(n8857) );
  nand_x4_sg U64322 ( .A(n14964), .B(n14965), .X(n8990) );
  nand_x4_sg U64323 ( .A(n16530), .B(n16531), .X(n9311) );
  nor_x1_sg U64324 ( .A(n43994), .B(n51874), .X(n12018) );
  nand_x4_sg U64325 ( .A(n17710), .B(n17711), .X(n17648) );
  nand_x1_sg U64326 ( .A(n43334), .B(n17699), .X(n17710) );
  nand_x1_sg U64327 ( .A(n53879), .B(n43335), .X(n17711) );
  nand_x4_sg U64328 ( .A(n19255), .B(n19256), .X(n19193) );
  nand_x1_sg U64329 ( .A(n43330), .B(n19244), .X(n19255) );
  nand_x1_sg U64330 ( .A(n54444), .B(n43331), .X(n19256) );
  nand_x4_sg U64331 ( .A(n20799), .B(n20800), .X(n20737) );
  nand_x1_sg U64332 ( .A(n43326), .B(n20788), .X(n20799) );
  nand_x1_sg U64333 ( .A(n55012), .B(n43327), .X(n20800) );
  nor_x1_sg U64334 ( .A(n43992), .B(n52152), .X(n12803) );
  nor_x1_sg U64335 ( .A(n43990), .B(n52986), .X(n15136) );
  nor_x1_sg U64336 ( .A(n43986), .B(n53544), .X(n16702) );
  nand_x4_sg U64337 ( .A(n16153), .B(n16154), .X(n16089) );
  nand_x1_sg U64338 ( .A(n43304), .B(n16142), .X(n16153) );
  nand_x1_sg U64339 ( .A(n53315), .B(n43305), .X(n16154) );
  nor_x1_sg U64340 ( .A(n43996), .B(n51594), .X(n11242) );
  nor_x1_sg U64341 ( .A(n43988), .B(n53261), .X(n15913) );
  nor_x1_sg U64342 ( .A(n44477), .B(n54104), .X(n18248) );
  nand_x4_sg U64343 ( .A(n11268), .B(n11269), .X(n11246) );
  nand_x1_sg U64344 ( .A(n44076), .B(n11271), .X(n11269) );
  nand_x1_sg U64345 ( .A(n11273), .B(n51622), .X(n11268) );
  nand_x4_sg U64346 ( .A(n12829), .B(n12830), .X(n12807) );
  nand_x1_sg U64347 ( .A(n44283), .B(n12832), .X(n12830) );
  nand_x1_sg U64348 ( .A(n12834), .B(n52181), .X(n12829) );
  nand_x4_sg U64349 ( .A(n15162), .B(n15163), .X(n15140) );
  nand_x1_sg U64350 ( .A(n44281), .B(n15165), .X(n15163) );
  nand_x1_sg U64351 ( .A(n15167), .B(n53015), .X(n15162) );
  nand_x4_sg U64352 ( .A(n16728), .B(n16729), .X(n16706) );
  nand_x1_sg U64353 ( .A(n44279), .B(n16731), .X(n16729) );
  nand_x1_sg U64354 ( .A(n16733), .B(n53573), .X(n16728) );
  nand_x4_sg U64355 ( .A(n12047), .B(n12048), .X(n12022) );
  nand_x1_sg U64356 ( .A(n45529), .B(n12050), .X(n12048) );
  nand_x1_sg U64357 ( .A(n12052), .B(n51904), .X(n12047) );
  nand_x4_sg U64358 ( .A(n13608), .B(n13609), .X(n13583) );
  nand_x1_sg U64359 ( .A(n41734), .B(n13611), .X(n13609) );
  nand_x1_sg U64360 ( .A(n13613), .B(n52457), .X(n13608) );
  nand_x1_sg U64361 ( .A(n52457), .B(n13612), .X(n13611) );
  nand_x4_sg U64362 ( .A(n15942), .B(n15943), .X(n15917) );
  nand_x1_sg U64363 ( .A(n44695), .B(n15945), .X(n15943) );
  nand_x1_sg U64364 ( .A(n15947), .B(n53289), .X(n15942) );
  nand_x4_sg U64365 ( .A(n51619), .B(n11627), .X(n11812) );
  nand_x4_sg U64366 ( .A(n52178), .B(n13188), .X(n13369) );
  nand_x4_sg U64367 ( .A(n53012), .B(n15521), .X(n15702) );
  nand_x4_sg U64368 ( .A(n53570), .B(n17087), .X(n17268) );
  nand_x4_sg U64369 ( .A(n17506), .B(n17507), .X(n17484) );
  nand_x1_sg U64370 ( .A(n17508), .B(n17509), .X(n17507) );
  nand_x1_sg U64371 ( .A(n17511), .B(n53853), .X(n17506) );
  nand_x1_sg U64372 ( .A(n53853), .B(n17510), .X(n17509) );
  nand_x4_sg U64373 ( .A(n19051), .B(n19052), .X(n19029) );
  nand_x1_sg U64374 ( .A(n19053), .B(n19054), .X(n19052) );
  nand_x1_sg U64375 ( .A(n19056), .B(n54418), .X(n19051) );
  nand_x1_sg U64376 ( .A(n54418), .B(n19055), .X(n19054) );
  nand_x4_sg U64377 ( .A(n20595), .B(n20596), .X(n20573) );
  nand_x1_sg U64378 ( .A(n20597), .B(n20598), .X(n20596) );
  nand_x1_sg U64379 ( .A(n20600), .B(n54986), .X(n20595) );
  nand_x1_sg U64380 ( .A(n54986), .B(n20599), .X(n20598) );
  nand_x4_sg U64381 ( .A(n16206), .B(n16207), .X(n16258) );
  nor_x1_sg U64382 ( .A(n46231), .B(n25449), .X(n25458) );
  nor_x1_sg U64383 ( .A(n46211), .B(n28242), .X(n28251) );
  nand_x4_sg U64384 ( .A(n51296), .B(n10305), .X(n10302) );
  nand_x4_sg U64385 ( .A(n51857), .B(n11856), .X(n11853) );
  nand_x4_sg U64386 ( .A(n52686), .B(n14197), .X(n14194) );
  nand_x4_sg U64387 ( .A(n53243), .B(n15751), .X(n15748) );
  nand_x4_sg U64388 ( .A(n54087), .B(n18088), .X(n18085) );
  nand_x4_sg U64389 ( .A(n54650), .B(n19633), .X(n19630) );
  nand_x4_sg U64390 ( .A(n55218), .B(n21178), .X(n21175) );
  nand_x4_sg U64391 ( .A(n54101), .B(n18217), .X(n18168) );
  nand_x4_sg U64392 ( .A(n51311), .B(n10436), .X(n10386) );
  nand_x4_sg U64393 ( .A(n52700), .B(n14328), .X(n14278) );
  nand_x4_sg U64394 ( .A(n54665), .B(n19763), .X(n19713) );
  nand_x4_sg U64395 ( .A(n55233), .B(n21308), .X(n21258) );
  nand_x4_sg U64396 ( .A(n10811), .B(n51448), .X(n10797) );
  nand_x1_sg U64397 ( .A(n10814), .B(n10813), .X(n10811) );
  nor_x1_sg U64398 ( .A(n10813), .B(n10814), .X(n10812) );
  nand_x4_sg U64399 ( .A(n10975), .B(n10936), .X(n10884) );
  nand_x4_sg U64400 ( .A(n18761), .B(n18721), .X(n18666) );
  nand_x4_sg U64401 ( .A(n20307), .B(n20267), .X(n20211) );
  nand_x4_sg U64402 ( .A(n21852), .B(n21812), .X(n21756) );
  nand_x4_sg U64403 ( .A(n16433), .B(n16394), .X(n16339) );
  nand_x4_sg U64404 ( .A(n17992), .B(n17952), .X(n17897) );
  nand_x4_sg U64405 ( .A(n19537), .B(n19497), .X(n19442) );
  nand_x4_sg U64406 ( .A(n21081), .B(n21041), .X(n20986) );
  nand_x4_sg U64407 ( .A(n51592), .B(n11077), .X(n11074) );
  nand_x4_sg U64408 ( .A(n52150), .B(n12638), .X(n12635) );
  nand_x4_sg U64409 ( .A(n52984), .B(n14971), .X(n14968) );
  nand_x4_sg U64410 ( .A(n53542), .B(n16537), .X(n16534) );
  nand_x4_sg U64411 ( .A(n51872), .B(n11860), .X(n11857) );
  nand_x4_sg U64412 ( .A(n53259), .B(n15755), .X(n15752) );
  nand_x4_sg U64413 ( .A(n11282), .B(n11283), .X(n11281) );
  nand_x1_sg U64414 ( .A(n51606), .B(n11284), .X(n11283) );
  nand_x1_sg U64415 ( .A(n51587), .B(n11285), .X(n11282) );
  nand_x4_sg U64416 ( .A(n12843), .B(n12844), .X(n12842) );
  nand_x1_sg U64417 ( .A(n52164), .B(n12845), .X(n12844) );
  nand_x1_sg U64418 ( .A(n52145), .B(n12846), .X(n12843) );
  nand_x4_sg U64419 ( .A(n15176), .B(n15177), .X(n15175) );
  nand_x1_sg U64420 ( .A(n52998), .B(n15178), .X(n15177) );
  nand_x1_sg U64421 ( .A(n52979), .B(n15179), .X(n15176) );
  nand_x4_sg U64422 ( .A(n16742), .B(n16743), .X(n16741) );
  nand_x1_sg U64423 ( .A(n53556), .B(n16744), .X(n16743) );
  nand_x1_sg U64424 ( .A(n53537), .B(n16745), .X(n16742) );
  nand_x4_sg U64425 ( .A(n10306), .B(n10307), .X(n9047) );
  nand_x4_sg U64426 ( .A(n11074), .B(n11075), .X(n8870) );
  nand_x4_sg U64427 ( .A(n11857), .B(n11858), .X(n8923) );
  nand_x4_sg U64428 ( .A(n12635), .B(n12636), .X(n8832) );
  nand_x4_sg U64429 ( .A(n14198), .B(n14199), .X(n8938) );
  nand_x4_sg U64430 ( .A(n18089), .B(n18090), .X(n9069) );
  nand_x4_sg U64431 ( .A(n14968), .B(n14969), .X(n8971) );
  nand_x4_sg U64432 ( .A(n15752), .B(n15753), .X(n9347) );
  nand_x4_sg U64433 ( .A(n16534), .B(n16535), .X(n9288) );
  nand_x4_sg U64434 ( .A(n19634), .B(n19635), .X(n9173) );
  nand_x4_sg U64435 ( .A(n21179), .B(n21180), .X(n9107) );
  nand_x4_sg U64436 ( .A(n10302), .B(n10303), .X(n9030) );
  nand_x4_sg U64437 ( .A(n11853), .B(n11854), .X(n8933) );
  nand_x4_sg U64438 ( .A(n14194), .B(n14195), .X(n8960) );
  nand_x4_sg U64439 ( .A(n15748), .B(n15749), .X(n9322) );
  nand_x4_sg U64440 ( .A(n18085), .B(n18086), .X(n9085) );
  nand_x4_sg U64441 ( .A(n19630), .B(n19631), .X(n9177) );
  nand_x4_sg U64442 ( .A(n21175), .B(n21176), .X(n9123) );
  nand_x4_sg U64443 ( .A(n51312), .B(n10309), .X(n10306) );
  nand_x4_sg U64444 ( .A(n52701), .B(n14201), .X(n14198) );
  nand_x4_sg U64445 ( .A(n54102), .B(n18092), .X(n18089) );
  nand_x4_sg U64446 ( .A(n54666), .B(n19637), .X(n19634) );
  nand_x4_sg U64447 ( .A(n55234), .B(n21182), .X(n21179) );
  nand_x4_sg U64448 ( .A(n12062), .B(n12063), .X(n12060) );
  nand_x1_sg U64449 ( .A(n51887), .B(n12064), .X(n12063) );
  nand_x1_sg U64450 ( .A(n51875), .B(n12065), .X(n12062) );
  nand_x4_sg U64451 ( .A(n15957), .B(n15958), .X(n15955) );
  nand_x1_sg U64452 ( .A(n53274), .B(n15959), .X(n15958) );
  nand_x1_sg U64453 ( .A(n53262), .B(n15960), .X(n15957) );
  nor_x1_sg U64454 ( .A(n46207), .B(n28800), .X(n28809) );
  nor_x1_sg U64455 ( .A(n46203), .B(n29361), .X(n29370) );
  nand_x4_sg U64456 ( .A(n12116), .B(n12117), .X(n12114) );
  nand_x4_sg U64457 ( .A(n16011), .B(n16012), .X(n16009) );
  nand_x4_sg U64458 ( .A(n12288), .B(n12241), .X(n12286) );
  nand_x4_sg U64459 ( .A(n16183), .B(n16136), .X(n16181) );
  nor_x1_sg U64460 ( .A(n53804), .B(n17447), .X(n17445) );
  nor_x1_sg U64461 ( .A(n54369), .B(n18992), .X(n18990) );
  nor_x1_sg U64462 ( .A(n54937), .B(n20536), .X(n20534) );
  nand_x4_sg U64463 ( .A(n17495), .B(n17494), .X(n17496) );
  nand_x4_sg U64464 ( .A(n19040), .B(n19039), .X(n19041) );
  nand_x4_sg U64465 ( .A(n20584), .B(n20583), .X(n20585) );
  nand_x4_sg U64466 ( .A(n14535), .B(n14548), .X(n14531) );
  nand_x1_sg U64467 ( .A(n52697), .B(n52709), .X(n14549) );
  nand_x4_sg U64468 ( .A(n17656), .B(n17669), .X(n17652) );
  nand_x1_sg U64469 ( .A(n53824), .B(n53836), .X(n17670) );
  nand_x4_sg U64470 ( .A(n19201), .B(n19214), .X(n19197) );
  nand_x1_sg U64471 ( .A(n54389), .B(n54401), .X(n19215) );
  nand_x4_sg U64472 ( .A(n20745), .B(n20758), .X(n20741) );
  nand_x1_sg U64473 ( .A(n54957), .B(n54969), .X(n20759) );
  nand_x4_sg U64474 ( .A(n10933), .B(n10934), .X(n10931) );
  nand_x1_sg U64475 ( .A(n41925), .B(n10938), .X(n10933) );
  nor_x1_sg U64476 ( .A(n51477), .B(n51432), .X(n10935) );
  nand_x4_sg U64477 ( .A(n16391), .B(n16392), .X(n16389) );
  nand_x1_sg U64478 ( .A(n41924), .B(n16396), .X(n16391) );
  nor_x1_sg U64479 ( .A(n53426), .B(n53381), .X(n16393) );
  nand_x4_sg U64480 ( .A(n10481), .B(n10480), .X(n10482) );
  nand_x4_sg U64481 ( .A(n19808), .B(n19807), .X(n19809) );
  nand_x4_sg U64482 ( .A(n21353), .B(n21352), .X(n21354) );
  nand_x4_sg U64483 ( .A(n18811), .B(n18816), .X(n18801) );
  nand_x4_sg U64484 ( .A(n20356), .B(n20361), .X(n20347) );
  nand_x4_sg U64485 ( .A(n21901), .B(n21906), .X(n21892) );
  nand_x4_sg U64486 ( .A(n13763), .B(n13776), .X(n13759) );
  nand_x1_sg U64487 ( .A(n52419), .B(n52440), .X(n13777) );
  nand_x4_sg U64488 ( .A(n11024), .B(n11029), .X(n11014) );
  nand_x4_sg U64489 ( .A(n10750), .B(n10749), .X(n10800) );
  nand_x4_sg U64490 ( .A(n11585), .B(n11586), .X(n11532) );
  nand_x1_sg U64491 ( .A(n51617), .B(n11581), .X(n11585) );
  nand_x1_sg U64492 ( .A(n51641), .B(n11582), .X(n11586) );
  nand_x4_sg U64493 ( .A(n13146), .B(n13147), .X(n13093) );
  nand_x1_sg U64494 ( .A(n52175), .B(n13142), .X(n13146) );
  nand_x1_sg U64495 ( .A(n52197), .B(n13143), .X(n13147) );
  nand_x4_sg U64496 ( .A(n15479), .B(n15480), .X(n15426) );
  nand_x1_sg U64497 ( .A(n53009), .B(n15475), .X(n15479) );
  nand_x1_sg U64498 ( .A(n53031), .B(n15476), .X(n15480) );
  nand_x4_sg U64499 ( .A(n17045), .B(n17046), .X(n16992) );
  nand_x1_sg U64500 ( .A(n53567), .B(n17041), .X(n17045) );
  nand_x1_sg U64501 ( .A(n53589), .B(n17042), .X(n17046) );
  nand_x4_sg U64502 ( .A(n14373), .B(n14372), .X(n14374) );
  nand_x4_sg U64503 ( .A(n18263), .B(n18262), .X(n18264) );
  nand_x4_sg U64504 ( .A(n15929), .B(n15928), .X(n15930) );
  nand_x4_sg U64505 ( .A(n18174), .B(n18175), .X(n18077) );
  nand_x1_sg U64506 ( .A(n18177), .B(n18178), .X(n18174) );
  nor_x1_sg U64507 ( .A(n18177), .B(n46341), .X(n18176) );
  nand_x4_sg U64508 ( .A(n11007), .B(n11008), .X(n10832) );
  nand_x1_sg U64509 ( .A(n11009), .B(n11006), .X(n11007) );
  nand_x1_sg U64510 ( .A(n51373), .B(n51392), .X(n11008) );
  nor_x1_sg U64511 ( .A(n28461), .B(n28459), .X(\L1_0/n3866 ) );
  nor_x1_sg U64512 ( .A(n28459), .B(n28462), .X(\L1_0/n3863 ) );
  nor_x1_sg U64513 ( .A(n55740), .B(n28459), .X(\L1_0/n3862 ) );
  nand_x4_sg U64514 ( .A(n12305), .B(n12306), .X(n12240) );
  nand_x4_sg U64515 ( .A(n10797), .B(n10801), .X(n10774) );
  nand_x1_sg U64516 ( .A(n51336), .B(n10803), .X(n10802) );
  nand_x4_sg U64517 ( .A(n16200), .B(n16201), .X(n16135) );
  nand_x4_sg U64518 ( .A(n10566), .B(n10567), .X(n10561) );
  nor_x1_sg U64519 ( .A(n26227), .B(n46585), .X(\L1_0/n4506 ) );
  nor_x1_sg U64520 ( .A(n27063), .B(n46589), .X(\L1_0/n4266 ) );
  nor_x1_sg U64521 ( .A(n27903), .B(n46591), .X(\L1_0/n4026 ) );
  nor_x1_sg U64522 ( .A(n28182), .B(n46593), .X(\L1_0/n3946 ) );
  nor_x1_sg U64523 ( .A(n29301), .B(n46596), .X(\L1_0/n3626 ) );
  nand_x4_sg U64524 ( .A(n13025), .B(n13024), .X(n13017) );
  nand_x4_sg U64525 ( .A(n15358), .B(n15357), .X(n15350) );
  nand_x4_sg U64526 ( .A(n16924), .B(n16923), .X(n16916) );
  nand_x4_sg U64527 ( .A(n11464), .B(n11463), .X(n11456) );
  nand_x4_sg U64528 ( .A(n17578), .B(n17579), .X(n17573) );
  nand_x4_sg U64529 ( .A(n19123), .B(n19124), .X(n19118) );
  nand_x4_sg U64530 ( .A(n20667), .B(n20668), .X(n20662) );
  nand_x1_sg U64531 ( .A(n51267), .B(n10293), .X(n10292) );
  nand_x1_sg U64532 ( .A(n51262), .B(n10294), .X(n10291) );
  nand_x1_sg U64533 ( .A(n53772), .B(n17304), .X(n17303) );
  nand_x1_sg U64534 ( .A(n53767), .B(n17305), .X(n17302) );
  nand_x1_sg U64535 ( .A(n54337), .B(n18849), .X(n18848) );
  nand_x1_sg U64536 ( .A(n54332), .B(n18850), .X(n18847) );
  nand_x1_sg U64537 ( .A(n54905), .B(n20393), .X(n20392) );
  nand_x1_sg U64538 ( .A(n54900), .B(n20394), .X(n20391) );
  nand_x1_sg U64539 ( .A(n51828), .B(n11844), .X(n11843) );
  nand_x1_sg U64540 ( .A(n51821), .B(n11845), .X(n11842) );
  nand_x1_sg U64541 ( .A(n53216), .B(n15739), .X(n15738) );
  nand_x1_sg U64542 ( .A(n53209), .B(n15740), .X(n15737) );
  nand_x1_sg U64543 ( .A(n52656), .B(n14185), .X(n14184) );
  nand_x1_sg U64544 ( .A(n52650), .B(n14186), .X(n14183) );
  nand_x1_sg U64545 ( .A(n54621), .B(n19621), .X(n19620) );
  nand_x1_sg U64546 ( .A(n54616), .B(n19622), .X(n19619) );
  nand_x1_sg U64547 ( .A(n55189), .B(n21166), .X(n21165) );
  nand_x1_sg U64548 ( .A(n55184), .B(n21167), .X(n21164) );
  nand_x1_sg U64549 ( .A(n52380), .B(n13406), .X(n13405) );
  nand_x1_sg U64550 ( .A(n52373), .B(n13407), .X(n13404) );
  nand_x4_sg U64551 ( .A(n11798), .B(n11806), .X(n11599) );
  nand_x1_sg U64552 ( .A(n11807), .B(n11808), .X(n11806) );
  nor_x1_sg U64553 ( .A(n51754), .B(n11809), .X(n11807) );
  nand_x4_sg U64554 ( .A(n13355), .B(n13363), .X(n13160) );
  nand_x1_sg U64555 ( .A(n13364), .B(n13365), .X(n13363) );
  nor_x1_sg U64556 ( .A(n52312), .B(n13366), .X(n13364) );
  nand_x4_sg U64557 ( .A(n15688), .B(n15696), .X(n15493) );
  nand_x1_sg U64558 ( .A(n15697), .B(n15698), .X(n15696) );
  nor_x1_sg U64559 ( .A(n53146), .B(n15699), .X(n15697) );
  nand_x4_sg U64560 ( .A(n17254), .B(n17262), .X(n17059) );
  nand_x1_sg U64561 ( .A(n17263), .B(n17264), .X(n17262) );
  nor_x1_sg U64562 ( .A(n53704), .B(n17265), .X(n17263) );
  nand_x4_sg U64563 ( .A(n14135), .B(n14143), .X(n13940) );
  nand_x1_sg U64564 ( .A(n14144), .B(n14145), .X(n14143) );
  nor_x1_sg U64565 ( .A(n52587), .B(n14146), .X(n14144) );
  nand_x4_sg U64566 ( .A(n16473), .B(n16481), .X(n16275) );
  nand_x1_sg U64567 ( .A(n16482), .B(n16483), .X(n16481) );
  nor_x1_sg U64568 ( .A(n53423), .B(n16484), .X(n16482) );
  nand_x4_sg U64569 ( .A(n13948), .B(n13954), .X(n13881) );
  nand_x1_sg U64570 ( .A(n13955), .B(n13956), .X(n13954) );
  nor_x1_sg U64571 ( .A(n43979), .B(n13958), .X(n13955) );
  nand_x1_sg U64572 ( .A(n17809), .B(n17810), .X(n17808) );
  nor_x1_sg U64573 ( .A(n53927), .B(n17811), .X(n17809) );
  nand_x1_sg U64574 ( .A(n19354), .B(n19355), .X(n19353) );
  nor_x1_sg U64575 ( .A(n54492), .B(n19356), .X(n19354) );
  nand_x1_sg U64576 ( .A(n20898), .B(n20899), .X(n20897) );
  nor_x1_sg U64577 ( .A(n55060), .B(n20900), .X(n20898) );
  nand_x4_sg U64578 ( .A(n13709), .B(n13715), .X(n13705) );
  nor_x1_sg U64579 ( .A(n13718), .B(n13719), .X(n13716) );
  nand_x4_sg U64580 ( .A(n14531), .B(n14533), .X(n14487) );
  nor_x1_sg U64581 ( .A(n52777), .B(n14536), .X(n14534) );
  nand_x4_sg U64582 ( .A(n17652), .B(n17654), .X(n17608) );
  nor_x1_sg U64583 ( .A(n53897), .B(n17657), .X(n17655) );
  nand_x4_sg U64584 ( .A(n19197), .B(n19199), .X(n19153) );
  nor_x1_sg U64585 ( .A(n54462), .B(n19202), .X(n19200) );
  nand_x4_sg U64586 ( .A(n20741), .B(n20743), .X(n20697) );
  nor_x1_sg U64587 ( .A(n55030), .B(n20746), .X(n20744) );
  nand_x4_sg U64588 ( .A(n18801), .B(n18809), .X(n18599) );
  nor_x1_sg U64589 ( .A(n44663), .B(n18813), .X(n18810) );
  nand_x4_sg U64590 ( .A(n13759), .B(n13761), .X(n13713) );
  nor_x1_sg U64591 ( .A(n13764), .B(n13765), .X(n13762) );
  nand_x4_sg U64592 ( .A(n11014), .B(n11022), .X(n10819) );
  nor_x1_sg U64593 ( .A(n44664), .B(n11026), .X(n11023) );
  nor_x1_sg U64594 ( .A(n46585), .B(n26228), .X(\L1_0/n4503 ) );
  nor_x1_sg U64595 ( .A(n46587), .B(n26505), .X(\L1_0/n4427 ) );
  nand_x2_sg U64596 ( .A(n46235), .B(n46484), .X(n26505) );
  nor_x1_sg U64597 ( .A(n46591), .B(n27904), .X(\L1_0/n4023 ) );
  nor_x1_sg U64598 ( .A(n46596), .B(n29302), .X(\L1_0/n3623 ) );
  nor_x1_sg U64599 ( .A(n46589), .B(n27064), .X(\L1_0/n4263 ) );
  nor_x1_sg U64600 ( .A(n46593), .B(n28183), .X(\L1_0/n3943 ) );
  inv_x2_sg U64601 ( .A(n46672), .X(n46665) );
  inv_x2_sg U64602 ( .A(n46672), .X(n46664) );
  inv_x2_sg U64603 ( .A(n46672), .X(n46663) );
  inv_x2_sg U64604 ( .A(n46672), .X(n46670) );
  inv_x2_sg U64605 ( .A(n46672), .X(n46669) );
  inv_x2_sg U64606 ( .A(n46672), .X(n46668) );
  inv_x2_sg U64607 ( .A(n46672), .X(n46667) );
  inv_x2_sg U64608 ( .A(n46672), .X(n46666) );
  nand_x1_sg U64609 ( .A(n41352), .B(n46283), .X(n9149) );
  nand_x1_sg U64610 ( .A(n41968), .B(n46283), .X(n9156) );
  nand_x1_sg U64611 ( .A(n42859), .B(n46283), .X(n9152) );
  nand_x1_sg U64612 ( .A(n44389), .B(n46283), .X(n9129) );
  nor_x1_sg U64613 ( .A(n42313), .B(n46514), .X(n12264) );
  nor_x1_sg U64614 ( .A(n13124), .B(n13120), .X(n13122) );
  nor_x1_sg U64615 ( .A(n15457), .B(n15453), .X(n15455) );
  nor_x1_sg U64616 ( .A(n17023), .B(n17019), .X(n17021) );
  nor_x1_sg U64617 ( .A(n11563), .B(n11559), .X(n11561) );
  nand_x4_sg U64618 ( .A(n52848), .B(n46458), .X(n14891) );
  nand_x4_sg U64619 ( .A(n53408), .B(n15728), .X(n16453) );
  nand_x4_sg U64620 ( .A(n53968), .B(n46368), .X(n18012) );
  nand_x4_sg U64621 ( .A(n54533), .B(n46321), .X(n19557) );
  nand_x4_sg U64622 ( .A(n54818), .B(n46301), .X(n20327) );
  nand_x4_sg U64623 ( .A(n55101), .B(n46276), .X(n21101) );
  nand_x4_sg U64624 ( .A(n55386), .B(n46256), .X(n21872) );
  nand_x4_sg U64625 ( .A(n51738), .B(n46547), .X(n11778) );
  nand_x4_sg U64626 ( .A(n54250), .B(n46348), .X(n18781) );
  nor_x1_sg U64627 ( .A(n42323), .B(n46561), .X(n10703) );
  nor_x1_sg U64628 ( .A(n42327), .B(n46289), .X(n20030) );
  nor_x1_sg U64629 ( .A(n42325), .B(n46244), .X(n21575) );
  nor_x1_sg U64630 ( .A(n42335), .B(n46445), .X(n14595) );
  nor_x1_sg U64631 ( .A(n42333), .B(n53814), .X(n17716) );
  nor_x1_sg U64632 ( .A(n42331), .B(n54379), .X(n19261) );
  nor_x1_sg U64633 ( .A(n42329), .B(n54947), .X(n20805) );
  nor_x1_sg U64634 ( .A(n42311), .B(n46402), .X(n16159) );
  nand_x1_sg U64635 ( .A(n53298), .B(n15728), .X(n16108) );
  nor_x1_sg U64636 ( .A(n18327), .B(n46335), .X(n18638) );
  nand_x1_sg U64637 ( .A(n46572), .B(n46569), .X(n10396) );
  nand_x4_sg U64638 ( .A(n54165), .B(n46343), .X(n18618) );
  nand_x1_sg U64639 ( .A(n54250), .B(n46343), .X(n18710) );
  nand_x1_sg U64640 ( .A(n52742), .B(n46458), .X(n14546) );
  nand_x1_sg U64641 ( .A(n53862), .B(n46368), .X(n17667) );
  nand_x1_sg U64642 ( .A(n54427), .B(n46321), .X(n19212) );
  nand_x1_sg U64643 ( .A(n54995), .B(n46276), .X(n20756) );
  nand_x2_sg U64644 ( .A(n12611), .B(n52271), .X(n13354) );
  nand_x2_sg U64645 ( .A(n13395), .B(n52546), .X(n14134) );
  nand_x2_sg U64646 ( .A(n14944), .B(n53105), .X(n15687) );
  nand_x2_sg U64647 ( .A(n16510), .B(n53663), .X(n17253) );
  nor_x1_sg U64648 ( .A(n12134), .B(n46514), .X(n12544) );
  nor_x1_sg U64649 ( .A(n13695), .B(n46469), .X(n14105) );
  nor_x1_sg U64650 ( .A(n46566), .B(n46561), .X(n10548) );
  nor_x1_sg U64651 ( .A(n46300), .B(n46289), .X(n19875) );
  nor_x1_sg U64652 ( .A(n46255), .B(n46244), .X(n21420) );
  nor_x1_sg U64653 ( .A(n11345), .B(n11300), .X(n11341) );
  nor_x1_sg U64654 ( .A(n12125), .B(n12080), .X(n12121) );
  nor_x1_sg U64655 ( .A(n12906), .B(n12861), .X(n12902) );
  nor_x1_sg U64656 ( .A(n15239), .B(n15194), .X(n15235) );
  nor_x1_sg U64657 ( .A(n16020), .B(n15975), .X(n16016) );
  nor_x1_sg U64658 ( .A(n16805), .B(n16760), .X(n16801) );
  nor_x1_sg U64659 ( .A(n41600), .B(n13512), .X(n13510) );
  nand_x1_sg U64660 ( .A(n13512), .B(n41600), .X(n13511) );
  nand_x1_sg U64661 ( .A(n11382), .B(n11381), .X(n11383) );
  nand_x1_sg U64662 ( .A(n12162), .B(n12161), .X(n12163) );
  nand_x1_sg U64663 ( .A(n12943), .B(n12942), .X(n12944) );
  nand_x1_sg U64664 ( .A(n15276), .B(n15275), .X(n15277) );
  nand_x1_sg U64665 ( .A(n16057), .B(n16056), .X(n16058) );
  nand_x1_sg U64666 ( .A(n16842), .B(n16841), .X(n16843) );
  nand_x2_sg U64667 ( .A(n10876), .B(n51334), .X(n10957) );
  nand_x2_sg U64668 ( .A(n18657), .B(n54109), .X(n18743) );
  nand_x2_sg U64669 ( .A(n20202), .B(n46286), .X(n20289) );
  nand_x2_sg U64670 ( .A(n21747), .B(n46241), .X(n21834) );
  nand_x2_sg U64671 ( .A(n12436), .B(n51879), .X(n12519) );
  nand_x2_sg U64672 ( .A(n13997), .B(n52430), .X(n14080) );
  nand_x2_sg U64673 ( .A(n16331), .B(n53282), .X(n16413) );
  nand_x2_sg U64674 ( .A(n11656), .B(n46532), .X(n11739) );
  nand_x2_sg U64675 ( .A(n13217), .B(n46488), .X(n13300) );
  nand_x2_sg U64676 ( .A(n15550), .B(n46420), .X(n15633) );
  nand_x2_sg U64677 ( .A(n17116), .B(n46376), .X(n17199) );
  nand_x2_sg U64678 ( .A(n10521), .B(n10522), .X(n10523) );
  nand_x1_sg U64679 ( .A(n52627), .B(n14015), .X(n14016) );
  nand_x1_sg U64680 ( .A(n52908), .B(n14786), .X(n14787) );
  nand_x1_sg U64681 ( .A(n54309), .B(n18676), .X(n18677) );
  nand_x1_sg U64682 ( .A(n54877), .B(n20221), .X(n20222) );
  nand_x1_sg U64683 ( .A(n55445), .B(n21766), .X(n21767) );
  nand_x1_sg U64684 ( .A(n52074), .B(n12454), .X(n12455) );
  nand_x1_sg U64685 ( .A(n51798), .B(n11674), .X(n11675) );
  nand_x1_sg U64686 ( .A(n52352), .B(n13235), .X(n13236) );
  nand_x1_sg U64687 ( .A(n53186), .B(n15568), .X(n15569) );
  nand_x1_sg U64688 ( .A(n53744), .B(n17134), .X(n17135) );
  nand_x1_sg U64689 ( .A(n54028), .B(n17907), .X(n17908) );
  nand_x1_sg U64690 ( .A(n54593), .B(n19452), .X(n19453) );
  nand_x1_sg U64691 ( .A(n55161), .B(n20996), .X(n20997) );
  nand_x2_sg U64692 ( .A(n19848), .B(n19849), .X(n19850) );
  nand_x2_sg U64693 ( .A(n21393), .B(n21394), .X(n21395) );
  nand_x2_sg U64694 ( .A(n14413), .B(n14414), .X(n14415) );
  nand_x2_sg U64695 ( .A(n46608), .B(n46576), .X(n24471) );
  nand_x2_sg U64696 ( .A(n46484), .B(n13876), .X(n13963) );
  nor_x1_sg U64697 ( .A(n18561), .B(n18558), .X(n18559) );
  nand_x2_sg U64698 ( .A(n12026), .B(n12024), .X(n12025) );
  nand_x2_sg U64699 ( .A(n15921), .B(n15919), .X(n15920) );
  nand_x4_sg U64700 ( .A(n26315), .B(n13184), .X(n26322) );
  nand_x4_sg U64701 ( .A(n26594), .B(n13964), .X(n26601) );
  nand_x4_sg U64702 ( .A(n27151), .B(n15517), .X(n27158) );
  nand_x4_sg U64703 ( .A(n27711), .B(n17083), .X(n27718) );
  nand_x1_sg U64704 ( .A(n17962), .B(n17961), .X(n17956) );
  nand_x1_sg U64705 ( .A(n17958), .B(n53926), .X(n17957) );
  nand_x1_sg U64706 ( .A(n19507), .B(n19506), .X(n19501) );
  nand_x1_sg U64707 ( .A(n19503), .B(n54491), .X(n19502) );
  nand_x1_sg U64708 ( .A(n21051), .B(n21050), .X(n21045) );
  nand_x1_sg U64709 ( .A(n21047), .B(n55059), .X(n21046) );
  nand_x4_sg U64710 ( .A(n51293), .B(n10648), .X(n10596) );
  nand_x1_sg U64711 ( .A(n51366), .B(n10464), .X(n10648) );
  nand_x4_sg U64712 ( .A(n53802), .B(n17661), .X(n17609) );
  nand_x1_sg U64713 ( .A(n53863), .B(n53788), .X(n17661) );
  nand_x4_sg U64714 ( .A(n54367), .B(n19206), .X(n19154) );
  nand_x1_sg U64715 ( .A(n54428), .B(n54353), .X(n19206) );
  nand_x4_sg U64716 ( .A(n54935), .B(n20750), .X(n20698) );
  nand_x1_sg U64717 ( .A(n54996), .B(n54921), .X(n20750) );
  nand_x4_sg U64718 ( .A(n25478), .B(n10843), .X(n25485) );
  nand_x2_sg U64719 ( .A(n10482), .B(n10510), .X(n10509) );
  nand_x1_sg U64720 ( .A(n10511), .B(n10478), .X(n10510) );
  nand_x1_sg U64721 ( .A(n10946), .B(n10945), .X(n10940) );
  nand_x1_sg U64722 ( .A(n12173), .B(n12171), .X(n12167) );
  nor_x1_sg U64723 ( .A(n46528), .B(n12174), .X(n12173) );
  nand_x1_sg U64724 ( .A(n16068), .B(n16066), .X(n16062) );
  nor_x1_sg U64725 ( .A(n46416), .B(n16069), .X(n16068) );
  nand_x1_sg U64726 ( .A(n11393), .B(n11391), .X(n11387) );
  nor_x1_sg U64727 ( .A(n46552), .B(n11394), .X(n11393) );
  nand_x2_sg U64728 ( .A(n12819), .B(n12848), .X(n12847) );
  nand_x1_sg U64729 ( .A(n12849), .B(n12850), .X(n12848) );
  nor_x1_sg U64730 ( .A(n46508), .B(n46491), .X(n12849) );
  nand_x2_sg U64731 ( .A(n15152), .B(n15181), .X(n15180) );
  nand_x1_sg U64732 ( .A(n15182), .B(n15183), .X(n15181) );
  nor_x1_sg U64733 ( .A(n46440), .B(n46423), .X(n15182) );
  nand_x2_sg U64734 ( .A(n16718), .B(n16747), .X(n16746) );
  nand_x1_sg U64735 ( .A(n16748), .B(n16749), .X(n16747) );
  nor_x1_sg U64736 ( .A(n46396), .B(n46379), .X(n16748) );
  nand_x1_sg U64737 ( .A(n12954), .B(n12952), .X(n12948) );
  nor_x1_sg U64738 ( .A(n46508), .B(n12955), .X(n12954) );
  nand_x1_sg U64739 ( .A(n15287), .B(n15285), .X(n15281) );
  nor_x1_sg U64740 ( .A(n46440), .B(n15288), .X(n15287) );
  nand_x1_sg U64741 ( .A(n16853), .B(n16851), .X(n16847) );
  nor_x1_sg U64742 ( .A(n46396), .B(n16854), .X(n16853) );
  nand_x2_sg U64743 ( .A(n11258), .B(n11287), .X(n11286) );
  nand_x1_sg U64744 ( .A(n11288), .B(n11289), .X(n11287) );
  nor_x1_sg U64745 ( .A(n46552), .B(n46535), .X(n11288) );
  nand_x1_sg U64746 ( .A(n12509), .B(n12508), .X(n12503) );
  nand_x2_sg U64747 ( .A(n18256), .B(n18254), .X(n18255) );
  nand_x2_sg U64748 ( .A(n14843), .B(n14844), .X(n14842) );
  nand_x1_sg U64749 ( .A(n43805), .B(n14846), .X(n14844) );
  nand_x1_sg U64750 ( .A(n14848), .B(n14847), .X(n14843) );
  nand_x2_sg U64751 ( .A(n17964), .B(n17965), .X(n17963) );
  nand_x1_sg U64752 ( .A(n43035), .B(n17967), .X(n17965) );
  nand_x1_sg U64753 ( .A(n17969), .B(n17968), .X(n17964) );
  nand_x2_sg U64754 ( .A(n19509), .B(n19510), .X(n19508) );
  nand_x1_sg U64755 ( .A(n43033), .B(n19512), .X(n19510) );
  nand_x1_sg U64756 ( .A(n19514), .B(n19513), .X(n19509) );
  nand_x2_sg U64757 ( .A(n21053), .B(n21054), .X(n21052) );
  nand_x1_sg U64758 ( .A(n43031), .B(n21056), .X(n21054) );
  nand_x1_sg U64759 ( .A(n21058), .B(n21057), .X(n21053) );
  nand_x2_sg U64760 ( .A(n14374), .B(n14402), .X(n14401) );
  nand_x1_sg U64761 ( .A(n14403), .B(n14370), .X(n14402) );
  nand_x2_sg U64762 ( .A(n12035), .B(n12067), .X(n12066) );
  nand_x1_sg U64763 ( .A(n12068), .B(n12069), .X(n12067) );
  nor_x1_sg U64764 ( .A(n46528), .B(n46512), .X(n12068) );
  nand_x2_sg U64765 ( .A(n15930), .B(n15962), .X(n15961) );
  nand_x1_sg U64766 ( .A(n15963), .B(n15964), .X(n15962) );
  nor_x1_sg U64767 ( .A(n46416), .B(n46400), .X(n15963) );
  nand_x1_sg U64768 ( .A(n16404), .B(n16403), .X(n16398) );
  nand_x4_sg U64769 ( .A(n25756), .B(n11623), .X(n25763) );
  nor_x1_sg U64770 ( .A(n17673), .B(n53788), .X(n18015) );
  nor_x1_sg U64771 ( .A(n19218), .B(n54353), .X(n19560) );
  nor_x1_sg U64772 ( .A(n20762), .B(n54921), .X(n21104) );
  nand_x4_sg U64773 ( .A(n53827), .B(n53765), .X(n17564) );
  nand_x4_sg U64774 ( .A(n54392), .B(n54330), .X(n19109) );
  nand_x4_sg U64775 ( .A(n54960), .B(n54898), .X(n20653) );
  nand_x2_sg U64776 ( .A(n27413), .B(n46235), .X(n27408) );
  nand_x2_sg U64777 ( .A(n27410), .B(n27411), .X(n27409) );
  nand_x4_sg U64778 ( .A(n52707), .B(n52648), .X(n14444) );
  nand_x2_sg U64779 ( .A(n26854), .B(n46235), .X(n26849) );
  nand_x2_sg U64780 ( .A(n26851), .B(n26852), .X(n26850) );
  nand_x2_sg U64781 ( .A(n27973), .B(n46235), .X(n27968) );
  nand_x2_sg U64782 ( .A(n27970), .B(n27971), .X(n27969) );
  nand_x2_sg U64783 ( .A(n28531), .B(n46235), .X(n28526) );
  nand_x2_sg U64784 ( .A(n28528), .B(n28529), .X(n28527) );
  nand_x2_sg U64785 ( .A(n29090), .B(n46235), .X(n29085) );
  nand_x2_sg U64786 ( .A(n29087), .B(n29088), .X(n29086) );
  nand_x2_sg U64787 ( .A(n25488), .B(n46235), .X(n25483) );
  nand_x2_sg U64788 ( .A(n25485), .B(n25486), .X(n25484) );
  nand_x2_sg U64789 ( .A(n28281), .B(n46235), .X(n28276) );
  nand_x2_sg U64790 ( .A(n28278), .B(n28279), .X(n28277) );
  nand_x2_sg U64791 ( .A(n25752), .B(n46235), .X(n25747) );
  nand_x2_sg U64792 ( .A(n25749), .B(n25750), .X(n25748) );
  nand_x2_sg U64793 ( .A(n26030), .B(n46235), .X(n26025) );
  nand_x2_sg U64794 ( .A(n26027), .B(n26028), .X(n26026) );
  nand_x2_sg U64795 ( .A(n26311), .B(n46235), .X(n26306) );
  nand_x2_sg U64796 ( .A(n26308), .B(n26309), .X(n26307) );
  nand_x2_sg U64797 ( .A(n26590), .B(n46235), .X(n26585) );
  nand_x2_sg U64798 ( .A(n26587), .B(n26588), .X(n26586) );
  nand_x2_sg U64799 ( .A(n27147), .B(n46235), .X(n27142) );
  nand_x2_sg U64800 ( .A(n27144), .B(n27145), .X(n27143) );
  nand_x2_sg U64801 ( .A(n27427), .B(n46235), .X(n27422) );
  nand_x2_sg U64802 ( .A(n27424), .B(n27425), .X(n27423) );
  nand_x2_sg U64803 ( .A(n27707), .B(n46235), .X(n27702) );
  nand_x2_sg U64804 ( .A(n27704), .B(n27705), .X(n27703) );
  nand_x2_sg U64805 ( .A(n26868), .B(n46235), .X(n26863) );
  nand_x2_sg U64806 ( .A(n26865), .B(n26866), .X(n26864) );
  nand_x2_sg U64807 ( .A(n27987), .B(n46235), .X(n27982) );
  nand_x2_sg U64808 ( .A(n27984), .B(n27985), .X(n27983) );
  nand_x2_sg U64809 ( .A(n28545), .B(n46235), .X(n28540) );
  nand_x2_sg U64810 ( .A(n28542), .B(n28543), .X(n28541) );
  nand_x2_sg U64811 ( .A(n29104), .B(n46235), .X(n29099) );
  nand_x2_sg U64812 ( .A(n29101), .B(n29102), .X(n29100) );
  nand_x4_sg U64813 ( .A(n25428), .B(n46561), .X(n25435) );
  nand_x2_sg U64814 ( .A(n28267), .B(n46235), .X(n28262) );
  nand_x2_sg U64815 ( .A(n28264), .B(n28265), .X(n28263) );
  nand_x2_sg U64816 ( .A(n28825), .B(n46235), .X(n28820) );
  nand_x2_sg U64817 ( .A(n28822), .B(n28823), .X(n28821) );
  nand_x2_sg U64818 ( .A(n29386), .B(n46235), .X(n29381) );
  nand_x2_sg U64819 ( .A(n29383), .B(n29384), .X(n29382) );
  nand_x2_sg U64820 ( .A(n26882), .B(n46235), .X(n26877) );
  nand_x2_sg U64821 ( .A(n26879), .B(n26880), .X(n26878) );
  nand_x2_sg U64822 ( .A(n28001), .B(n46235), .X(n27996) );
  nand_x2_sg U64823 ( .A(n27998), .B(n27999), .X(n27997) );
  nand_x2_sg U64824 ( .A(n28559), .B(n46235), .X(n28554) );
  nand_x2_sg U64825 ( .A(n28556), .B(n28557), .X(n28555) );
  nand_x2_sg U64826 ( .A(n29118), .B(n46235), .X(n29113) );
  nand_x2_sg U64827 ( .A(n29115), .B(n29116), .X(n29114) );
  nand_x2_sg U64828 ( .A(n28839), .B(n46235), .X(n28834) );
  nand_x2_sg U64829 ( .A(n28836), .B(n28837), .X(n28835) );
  nand_x2_sg U64830 ( .A(n29400), .B(n46235), .X(n29395) );
  nand_x2_sg U64831 ( .A(n29397), .B(n29398), .X(n29396) );
  nand_x2_sg U64832 ( .A(n26044), .B(n46235), .X(n26039) );
  nand_x2_sg U64833 ( .A(n26041), .B(n26042), .X(n26040) );
  nand_x2_sg U64834 ( .A(n26325), .B(n46235), .X(n26320) );
  nand_x2_sg U64835 ( .A(n26322), .B(n26323), .X(n26321) );
  nand_x2_sg U64836 ( .A(n26604), .B(n46235), .X(n26599) );
  nand_x2_sg U64837 ( .A(n26601), .B(n26602), .X(n26600) );
  nand_x2_sg U64838 ( .A(n27161), .B(n46235), .X(n27156) );
  nand_x2_sg U64839 ( .A(n27158), .B(n27159), .X(n27157) );
  nand_x2_sg U64840 ( .A(n27721), .B(n46235), .X(n27716) );
  nand_x2_sg U64841 ( .A(n27718), .B(n27719), .X(n27717) );
  nand_x1_sg U64842 ( .A(n14117), .B(n14116), .X(n14155) );
  nand_x2_sg U64843 ( .A(n25766), .B(n46235), .X(n25761) );
  nand_x2_sg U64844 ( .A(n25763), .B(n25764), .X(n25762) );
  nand_x2_sg U64845 ( .A(n27441), .B(n46235), .X(n27436) );
  nand_x2_sg U64846 ( .A(n27438), .B(n27439), .X(n27437) );
  nand_x1_sg U64847 ( .A(n11467), .B(n11466), .X(n11479) );
  nand_x1_sg U64848 ( .A(n13028), .B(n13027), .X(n13040) );
  nand_x1_sg U64849 ( .A(n15361), .B(n15360), .X(n15373) );
  nand_x1_sg U64850 ( .A(n16927), .B(n16926), .X(n16939) );
  nand_x2_sg U64851 ( .A(n26576), .B(n46235), .X(n26571) );
  nand_x2_sg U64852 ( .A(n26573), .B(n26574), .X(n26572) );
  nand_x2_sg U64853 ( .A(n25438), .B(n46235), .X(n25433) );
  nand_x2_sg U64854 ( .A(n25435), .B(n25436), .X(n25434) );
  nand_x2_sg U64855 ( .A(n26016), .B(n46235), .X(n26011) );
  nand_x2_sg U64856 ( .A(n26013), .B(n26014), .X(n26012) );
  nand_x2_sg U64857 ( .A(n25995), .B(n46235), .X(n25990) );
  nand_x2_sg U64858 ( .A(n25992), .B(n25993), .X(n25991) );
  nand_x2_sg U64859 ( .A(n27392), .B(n46235), .X(n27387) );
  nand_x2_sg U64860 ( .A(n27389), .B(n27390), .X(n27388) );
  nand_x2_sg U64861 ( .A(n26833), .B(n46235), .X(n26828) );
  nand_x2_sg U64862 ( .A(n26830), .B(n26831), .X(n26829) );
  nand_x2_sg U64863 ( .A(n28789), .B(n46235), .X(n28784) );
  nand_x2_sg U64864 ( .A(n28786), .B(n28787), .X(n28785) );
  nand_x2_sg U64865 ( .A(n29350), .B(n46235), .X(n29345) );
  nand_x2_sg U64866 ( .A(n29347), .B(n29348), .X(n29346) );
  nand_x2_sg U64867 ( .A(n25738), .B(n46235), .X(n25733) );
  nand_x2_sg U64868 ( .A(n25735), .B(n25736), .X(n25734) );
  nand_x2_sg U64869 ( .A(n26297), .B(n46235), .X(n26292) );
  nand_x2_sg U64870 ( .A(n26294), .B(n26295), .X(n26293) );
  nand_x2_sg U64871 ( .A(n27133), .B(n46235), .X(n27128) );
  nand_x2_sg U64872 ( .A(n27130), .B(n27131), .X(n27129) );
  nand_x2_sg U64873 ( .A(n27693), .B(n46235), .X(n27688) );
  nand_x2_sg U64874 ( .A(n27690), .B(n27691), .X(n27689) );
  nand_x2_sg U64875 ( .A(n26555), .B(n46235), .X(n26550) );
  nand_x2_sg U64876 ( .A(n26552), .B(n26553), .X(n26551) );
  nand_x4_sg U64877 ( .A(n53827), .B(n46358), .X(n18044) );
  nand_x4_sg U64878 ( .A(n54392), .B(n46311), .X(n19589) );
  nand_x4_sg U64879 ( .A(n54960), .B(n46266), .X(n21133) );
  nand_x1_sg U64880 ( .A(n13096), .B(n13095), .X(n13097) );
  nand_x1_sg U64881 ( .A(n15429), .B(n15428), .X(n15430) );
  nand_x1_sg U64882 ( .A(n16995), .B(n16994), .X(n16996) );
  nand_x1_sg U64883 ( .A(n11535), .B(n11534), .X(n11536) );
  nand_x4_sg U64884 ( .A(n25985), .B(n46514), .X(n25992) );
  nand_x4_sg U64885 ( .A(n27382), .B(n46402), .X(n27389) );
  nand_x4_sg U64886 ( .A(n26034), .B(n12404), .X(n26041) );
  nand_x4_sg U64887 ( .A(n27431), .B(n16299), .X(n27438) );
  nand_x4_sg U64888 ( .A(n26823), .B(n46445), .X(n26830) );
  nand_x4_sg U64889 ( .A(n28779), .B(n46289), .X(n28786) );
  nand_x4_sg U64890 ( .A(n29340), .B(n46244), .X(n29347) );
  nor_x1_sg U64891 ( .A(n11180), .B(n11253), .X(n11251) );
  nand_x2_sg U64892 ( .A(n46536), .B(n46547), .X(n11254) );
  nor_x1_sg U64893 ( .A(n12741), .B(n12814), .X(n12812) );
  nand_x2_sg U64894 ( .A(n52133), .B(n46503), .X(n12815) );
  nor_x1_sg U64895 ( .A(n15074), .B(n15147), .X(n15145) );
  nand_x2_sg U64896 ( .A(n52967), .B(n46435), .X(n15148) );
  nor_x1_sg U64897 ( .A(n16640), .B(n16713), .X(n16711) );
  nand_x2_sg U64898 ( .A(n53525), .B(n46391), .X(n16714) );
  nand_x4_sg U64899 ( .A(n52707), .B(n52695), .X(n14923) );
  nand_x4_sg U64900 ( .A(n26545), .B(n46469), .X(n26552) );
  nor_x1_sg U64901 ( .A(n46519), .B(n46514), .X(n12101) );
  nor_x1_sg U64902 ( .A(n46407), .B(n46402), .X(n15996) );
  nand_x4_sg U64903 ( .A(n46230), .B(n25786), .X(n25795) );
  nand_x4_sg U64904 ( .A(n46222), .B(n26902), .X(n26911) );
  nand_x4_sg U64905 ( .A(n46218), .B(n27461), .X(n27470) );
  nand_x4_sg U64906 ( .A(n46214), .B(n28021), .X(n28030) );
  nand_x4_sg U64907 ( .A(n46212), .B(n28301), .X(n28310) );
  nand_x4_sg U64908 ( .A(n46210), .B(n28579), .X(n28588) );
  nand_x4_sg U64909 ( .A(n46208), .B(n28859), .X(n28868) );
  nand_x4_sg U64910 ( .A(n46206), .B(n29138), .X(n29147) );
  nand_x4_sg U64911 ( .A(n46204), .B(n29420), .X(n29429) );
  nand_x4_sg U64912 ( .A(n53827), .B(n17828), .X(n17825) );
  nand_x4_sg U64913 ( .A(n54392), .B(n19373), .X(n19370) );
  nand_x4_sg U64914 ( .A(n54960), .B(n20917), .X(n20914) );
  nand_x4_sg U64915 ( .A(n53827), .B(n46356), .X(n17888) );
  nand_x4_sg U64916 ( .A(n54392), .B(n46309), .X(n19433) );
  nand_x4_sg U64917 ( .A(n54960), .B(n46264), .X(n20977) );
  nand_x4_sg U64918 ( .A(n46228), .B(n26065), .X(n26074) );
  nand_x4_sg U64919 ( .A(n46226), .B(n26346), .X(n26355) );
  nand_x4_sg U64920 ( .A(n46224), .B(n26625), .X(n26634) );
  nand_x4_sg U64921 ( .A(n46220), .B(n27182), .X(n27191) );
  nand_x4_sg U64922 ( .A(n46216), .B(n27742), .X(n27751) );
  nand_x2_sg U64923 ( .A(n13393), .B(n16508), .X(n16507) );
  nand_x1_sg U64924 ( .A(n46576), .B(n46583), .X(n16508) );
  nand_x2_sg U64925 ( .A(n13393), .B(n17291), .X(n17290) );
  nand_x1_sg U64926 ( .A(n55465), .B(n46576), .X(n17291) );
  nand_x2_sg U64927 ( .A(n46405), .B(n16451), .X(n16450) );
  nand_x2_sg U64928 ( .A(n46450), .B(n14880), .X(n14889) );
  nand_x4_sg U64929 ( .A(n51854), .B(n12207), .X(n12153) );
  nand_x1_sg U64930 ( .A(n51918), .B(n12061), .X(n12207) );
  nand_x4_sg U64931 ( .A(n53240), .B(n16102), .X(n16048) );
  nand_x1_sg U64932 ( .A(n53305), .B(n15956), .X(n16102) );
  nand_x4_sg U64933 ( .A(n46230), .B(n51756), .X(n25778) );
  nand_x4_sg U64934 ( .A(n46222), .B(n52865), .X(n26894) );
  nand_x4_sg U64935 ( .A(n46218), .B(n53425), .X(n27453) );
  nand_x4_sg U64936 ( .A(n46214), .B(n53985), .X(n28013) );
  nand_x4_sg U64937 ( .A(n46212), .B(n54268), .X(n28293) );
  nand_x4_sg U64938 ( .A(n46210), .B(n54550), .X(n28571) );
  nand_x4_sg U64939 ( .A(n46208), .B(n54835), .X(n28851) );
  nand_x4_sg U64940 ( .A(n46206), .B(n55118), .X(n29130) );
  nand_x4_sg U64941 ( .A(n46204), .B(n55403), .X(n29412) );
  nand_x4_sg U64942 ( .A(n46232), .B(n51474), .X(n25500) );
  nor_x1_sg U64943 ( .A(n53353), .B(n16442), .X(n16440) );
  nor_x1_sg U64944 ( .A(n51684), .B(n11768), .X(n11766) );
  nor_x1_sg U64945 ( .A(n53916), .B(n18002), .X(n17999) );
  nor_x1_sg U64946 ( .A(n54481), .B(n19547), .X(n19544) );
  nor_x1_sg U64947 ( .A(n55049), .B(n21091), .X(n21088) );
  nor_x1_sg U64948 ( .A(n17757), .B(n46364), .X(n17940) );
  nor_x1_sg U64949 ( .A(n19302), .B(n46317), .X(n19485) );
  nor_x1_sg U64950 ( .A(n20846), .B(n46272), .X(n21029) );
  nor_x1_sg U64951 ( .A(n54767), .B(n20317), .X(n20314) );
  nor_x1_sg U64952 ( .A(n55335), .B(n21862), .X(n21859) );
  nand_x4_sg U64953 ( .A(n52683), .B(n14540), .X(n14488) );
  nand_x1_sg U64954 ( .A(n52743), .B(n14356), .X(n14540) );
  nand_x4_sg U64955 ( .A(n54647), .B(n19975), .X(n19923) );
  nand_x1_sg U64956 ( .A(n54720), .B(n19791), .X(n19975) );
  nand_x4_sg U64957 ( .A(n55215), .B(n21520), .X(n21468) );
  nand_x1_sg U64958 ( .A(n55288), .B(n21336), .X(n21520) );
  nand_x4_sg U64959 ( .A(n54084), .B(n18430), .X(n18378) );
  nand_x1_sg U64960 ( .A(n54155), .B(n18246), .X(n18430) );
  nor_x1_sg U64961 ( .A(n17885), .B(n46362), .X(n17958) );
  nor_x1_sg U64962 ( .A(n19430), .B(n46315), .X(n19503) );
  nor_x1_sg U64963 ( .A(n20974), .B(n46270), .X(n21047) );
  nor_x1_sg U64964 ( .A(n16327), .B(n16239), .X(n16400) );
  nor_x1_sg U64965 ( .A(n11652), .B(n46541), .X(n11725) );
  nor_x1_sg U64966 ( .A(n13213), .B(n46497), .X(n13286) );
  nor_x1_sg U64967 ( .A(n14764), .B(n46451), .X(n14837) );
  nor_x1_sg U64968 ( .A(n15546), .B(n46429), .X(n15619) );
  nor_x1_sg U64969 ( .A(n17112), .B(n46385), .X(n17185) );
  nor_x1_sg U64970 ( .A(n12548), .B(n46518), .X(n12547) );
  nor_x1_sg U64971 ( .A(n12432), .B(n12344), .X(n12505) );
  nor_x1_sg U64972 ( .A(n13993), .B(n46475), .X(n14066) );
  nor_x1_sg U64973 ( .A(n20199), .B(n20108), .X(n20273) );
  nor_x1_sg U64974 ( .A(n21744), .B(n21653), .X(n21818) );
  nor_x1_sg U64975 ( .A(n13329), .B(n46497), .X(n13328) );
  nor_x1_sg U64976 ( .A(n15662), .B(n46429), .X(n15661) );
  nor_x1_sg U64977 ( .A(n17228), .B(n46385), .X(n17227) );
  nor_x1_sg U64978 ( .A(n10872), .B(n10782), .X(n10942) );
  nor_x1_sg U64979 ( .A(n14109), .B(n46475), .X(n14108) );
  nor_x1_sg U64980 ( .A(n20070), .B(n46297), .X(n20255) );
  nor_x1_sg U64981 ( .A(n21615), .B(n46252), .X(n21800) );
  nor_x1_sg U64982 ( .A(n13865), .B(n46477), .X(n14047) );
  nand_x4_sg U64983 ( .A(n46228), .B(n52039), .X(n26057) );
  nand_x4_sg U64984 ( .A(n46226), .B(n52315), .X(n26338) );
  nand_x4_sg U64985 ( .A(n46224), .B(n52590), .X(n26617) );
  nand_x4_sg U64986 ( .A(n46220), .B(n53149), .X(n27174) );
  nand_x4_sg U64987 ( .A(n46216), .B(n53707), .X(n27734) );
  nor_x1_sg U64988 ( .A(n13085), .B(n46499), .X(n13267) );
  nor_x1_sg U64989 ( .A(n15418), .B(n46431), .X(n15600) );
  nor_x1_sg U64990 ( .A(n16984), .B(n46387), .X(n17166) );
  nor_x1_sg U64991 ( .A(n11524), .B(n46543), .X(n11707) );
  nor_x1_sg U64992 ( .A(n12304), .B(n46521), .X(n12486) );
  nor_x1_sg U64993 ( .A(n14636), .B(n46454), .X(n14819) );
  nor_x1_sg U64994 ( .A(n16199), .B(n46409), .X(n16381) );
  nor_x1_sg U64995 ( .A(n53295), .B(n16069), .X(n16245) );
  nor_x1_sg U64996 ( .A(n53440), .B(n16069), .X(n16424) );
  nor_x1_sg U64997 ( .A(n13914), .B(n46475), .X(n13913) );
  nand_x4_sg U64998 ( .A(n18265), .B(n43514), .X(n18254) );
  nor_x1_sg U64999 ( .A(n18266), .B(n46335), .X(n18265) );
  nand_x4_sg U65000 ( .A(n12131), .B(n51890), .X(n12130) );
  nor_x1_sg U65001 ( .A(n46519), .B(n46523), .X(n12131) );
  nand_x4_sg U65002 ( .A(n12912), .B(n52167), .X(n12911) );
  nor_x1_sg U65003 ( .A(n46502), .B(n46501), .X(n12912) );
  nand_x4_sg U65004 ( .A(n15245), .B(n53001), .X(n15244) );
  nor_x1_sg U65005 ( .A(n46434), .B(n46433), .X(n15245) );
  nand_x4_sg U65006 ( .A(n16811), .B(n53559), .X(n16810) );
  nor_x1_sg U65007 ( .A(n46390), .B(n46389), .X(n16811) );
  nand_x4_sg U65008 ( .A(n12039), .B(n12040), .X(n12008) );
  nand_x1_sg U65009 ( .A(n12044), .B(n46513), .X(n12039) );
  nor_x1_sg U65010 ( .A(n12042), .B(n46518), .X(n12041) );
  nand_x2_sg U65011 ( .A(n12572), .B(n12416), .X(n12565) );
  nor_x1_sg U65012 ( .A(n46519), .B(n12404), .X(n12572) );
  nand_x1_sg U65013 ( .A(n11735), .B(n46547), .X(n11734) );
  nand_x1_sg U65014 ( .A(n12515), .B(n46525), .X(n12514) );
  nand_x1_sg U65015 ( .A(n13296), .B(n46503), .X(n13295) );
  nand_x1_sg U65016 ( .A(n14076), .B(n46481), .X(n14075) );
  nand_x1_sg U65017 ( .A(n14847), .B(n46458), .X(n14846) );
  nand_x1_sg U65018 ( .A(n15629), .B(n46435), .X(n15628) );
  nand_x1_sg U65019 ( .A(n17195), .B(n46391), .X(n17194) );
  nand_x1_sg U65020 ( .A(n17968), .B(n46368), .X(n17967) );
  nand_x1_sg U65021 ( .A(n18737), .B(n46348), .X(n18736) );
  nand_x1_sg U65022 ( .A(n19513), .B(n46321), .X(n19512) );
  nand_x1_sg U65023 ( .A(n20283), .B(n46301), .X(n20282) );
  nand_x1_sg U65024 ( .A(n21057), .B(n46276), .X(n21056) );
  nand_x1_sg U65025 ( .A(n21828), .B(n46256), .X(n21827) );
  nand_x4_sg U65026 ( .A(n18836), .B(n13393), .X(n18063) );
  nand_x4_sg U65027 ( .A(n13692), .B(n52441), .X(n13691) );
  nor_x1_sg U65028 ( .A(n46480), .B(n46479), .X(n13692) );
  nand_x2_sg U65029 ( .A(n46539), .B(n25701), .X(n25700) );
  nand_x2_sg U65030 ( .A(n46495), .B(n26260), .X(n26259) );
  nand_x2_sg U65031 ( .A(n46427), .B(n27096), .X(n27095) );
  nand_x2_sg U65032 ( .A(n46383), .B(n27656), .X(n27655) );
  nand_x2_sg U65033 ( .A(n44004), .B(n27936), .X(n27935) );
  nand_x2_sg U65034 ( .A(n44002), .B(n28494), .X(n28493) );
  nand_x2_sg U65035 ( .A(n44000), .B(n29053), .X(n29052) );
  nand_x4_sg U65036 ( .A(n54109), .B(n46333), .X(n18815) );
  nand_x2_sg U65037 ( .A(n51854), .B(n25980), .X(n25987) );
  nand_x2_sg U65038 ( .A(n53240), .B(n27377), .X(n27384) );
  nand_x2_sg U65039 ( .A(n53802), .B(n27937), .X(n27944) );
  nand_x2_sg U65040 ( .A(n54367), .B(n28495), .X(n28502) );
  nand_x2_sg U65041 ( .A(n54935), .B(n29054), .X(n29061) );
  nand_x2_sg U65042 ( .A(n46208), .B(n28793), .X(n28802) );
  nand_x2_sg U65043 ( .A(n46204), .B(n29354), .X(n29363) );
  nand_x2_sg U65044 ( .A(n46232), .B(n25471), .X(n25480) );
  nand_x2_sg U65045 ( .A(n46228), .B(n26027), .X(n26036) );
  nand_x2_sg U65046 ( .A(n46218), .B(n27424), .X(n27433) );
  nand_x2_sg U65047 ( .A(n46228), .B(n25999), .X(n26008) );
  nand_x2_sg U65048 ( .A(n46361), .B(n18001), .X(n18010) );
  nor_x1_sg U65049 ( .A(n46340), .B(n18770), .X(n18779) );
  nand_x2_sg U65050 ( .A(n46314), .B(n19546), .X(n19555) );
  nand_x2_sg U65051 ( .A(n46269), .B(n21090), .X(n21099) );
  nand_x4_sg U65052 ( .A(n11351), .B(n51609), .X(n11350) );
  nor_x1_sg U65053 ( .A(n46546), .B(n46545), .X(n11351) );
  nand_x4_sg U65054 ( .A(n16026), .B(n53277), .X(n16025) );
  nor_x1_sg U65055 ( .A(n46407), .B(n46411), .X(n16026) );
  nor_x1_sg U65056 ( .A(n51408), .B(n46565), .X(n10982) );
  nand_x4_sg U65057 ( .A(n52707), .B(n14707), .X(n14704) );
  nand_x4_sg U65058 ( .A(n52707), .B(n46443), .X(n14767) );
  nand_x2_sg U65059 ( .A(n17504), .B(n46358), .X(n17500) );
  nor_x1_sg U65060 ( .A(n46373), .B(n17421), .X(n17504) );
  nand_x2_sg U65061 ( .A(n19049), .B(n46311), .X(n19045) );
  nor_x1_sg U65062 ( .A(n46326), .B(n18966), .X(n19049) );
  nand_x2_sg U65063 ( .A(n20593), .B(n46266), .X(n20589) );
  nor_x1_sg U65064 ( .A(n46281), .B(n20510), .X(n20593) );
  nand_x2_sg U65065 ( .A(n46232), .B(n25442), .X(n25451) );
  nand_x2_sg U65066 ( .A(n46212), .B(n28235), .X(n28244) );
  nand_x2_sg U65067 ( .A(n43807), .B(n28249), .X(n28259) );
  nand_x2_sg U65068 ( .A(n43852), .B(n28807), .X(n28817) );
  nand_x2_sg U65069 ( .A(n44160), .B(n29368), .X(n29378) );
  nand_x2_sg U65070 ( .A(n46224), .B(n26559), .X(n26568) );
  nand_x2_sg U65071 ( .A(n46218), .B(n27396), .X(n27405) );
  nor_x1_sg U65072 ( .A(n10807), .B(n46566), .X(n10806) );
  nor_x1_sg U65073 ( .A(n17820), .B(n46367), .X(n17819) );
  nor_x1_sg U65074 ( .A(n19365), .B(n46320), .X(n19364) );
  nor_x1_sg U65075 ( .A(n20909), .B(n46275), .X(n20908) );
  nor_x1_sg U65076 ( .A(n51770), .B(n11394), .X(n11750) );
  nor_x1_sg U65077 ( .A(n42771), .B(n12955), .X(n13311) );
  nor_x1_sg U65078 ( .A(n42767), .B(n15288), .X(n15644) );
  nor_x1_sg U65079 ( .A(n42763), .B(n16854), .X(n17210) );
  nor_x1_sg U65080 ( .A(n14699), .B(n46452), .X(n14698) );
  nand_x4_sg U65081 ( .A(n46539), .B(n51630), .X(n11791) );
  nand_x4_sg U65082 ( .A(n46495), .B(n52187), .X(n13343) );
  nand_x4_sg U65083 ( .A(n46427), .B(n53021), .X(n15676) );
  nand_x4_sg U65084 ( .A(n46383), .B(n53579), .X(n17242) );
  nand_x2_sg U65085 ( .A(n51293), .B(n25423), .X(n25430) );
  nand_x4_sg U65086 ( .A(n12071), .B(n12072), .X(n12033) );
  nand_x1_sg U65087 ( .A(n11969), .B(n12074), .X(n12071) );
  nand_x1_sg U65088 ( .A(n12073), .B(n46513), .X(n12072) );
  nand_x1_sg U65089 ( .A(n46513), .B(n46525), .X(n12074) );
  nor_x1_sg U65090 ( .A(n16376), .B(n46406), .X(n16375) );
  nor_x1_sg U65091 ( .A(n11701), .B(n46541), .X(n11700) );
  nor_x1_sg U65092 ( .A(n12480), .B(n46518), .X(n12479) );
  nand_x4_sg U65093 ( .A(n10287), .B(n10288), .X(n9045) );
  nand_x1_sg U65094 ( .A(n46569), .B(n51268), .X(n10288) );
  nor_x1_sg U65095 ( .A(n19982), .B(n46295), .X(n20120) );
  nor_x1_sg U65096 ( .A(n21527), .B(n46250), .X(n21665) );
  nand_x2_sg U65097 ( .A(n46232), .B(n25456), .X(n25466) );
  nand_x2_sg U65098 ( .A(n44166), .B(n25735), .X(n25744) );
  nand_x2_sg U65099 ( .A(n46230), .B(n25749), .X(n25758) );
  nand_x2_sg U65100 ( .A(n44168), .B(n26013), .X(n26022) );
  nand_x2_sg U65101 ( .A(n43792), .B(n26294), .X(n26303) );
  nand_x2_sg U65102 ( .A(n43809), .B(n26573), .X(n26582) );
  nand_x2_sg U65103 ( .A(n43786), .B(n26851), .X(n26860) );
  nand_x2_sg U65104 ( .A(n43790), .B(n27130), .X(n27139) );
  nand_x2_sg U65105 ( .A(n44164), .B(n27410), .X(n27419) );
  nand_x2_sg U65106 ( .A(n43854), .B(n27690), .X(n27699) );
  nand_x2_sg U65107 ( .A(n43767), .B(n27970), .X(n27979) );
  nand_x2_sg U65108 ( .A(n44162), .B(n28528), .X(n28537) );
  nand_x2_sg U65109 ( .A(n46208), .B(n28822), .X(n28831) );
  nand_x2_sg U65110 ( .A(n43788), .B(n29087), .X(n29096) );
  nand_x2_sg U65111 ( .A(n46204), .B(n29383), .X(n29392) );
  nor_x1_sg U65112 ( .A(n14813), .B(n46451), .X(n14812) );
  nand_x4_sg U65113 ( .A(n13600), .B(n13601), .X(n13569) );
  nand_x1_sg U65114 ( .A(n13605), .B(n46468), .X(n13600) );
  nor_x1_sg U65115 ( .A(n13603), .B(n46477), .X(n13602) );
  nor_x1_sg U65116 ( .A(n13261), .B(n46497), .X(n13260) );
  nor_x1_sg U65117 ( .A(n14041), .B(n46475), .X(n14040) );
  nor_x1_sg U65118 ( .A(n15594), .B(n46429), .X(n15593) );
  nor_x1_sg U65119 ( .A(n17160), .B(n46385), .X(n17159) );
  nor_x1_sg U65120 ( .A(n43177), .B(n46406), .X(n16441) );
  nor_x1_sg U65121 ( .A(n52879), .B(n14507), .X(n14862) );
  nor_x1_sg U65122 ( .A(n53999), .B(n17628), .X(n17983) );
  nor_x1_sg U65123 ( .A(n54564), .B(n19173), .X(n19528) );
  nor_x1_sg U65124 ( .A(n55132), .B(n20717), .X(n21072) );
  nand_x2_sg U65125 ( .A(n46294), .B(n20316), .X(n20325) );
  nand_x2_sg U65126 ( .A(n46249), .B(n21861), .X(n21870) );
  nor_x1_sg U65127 ( .A(n17934), .B(n46362), .X(n17933) );
  nor_x1_sg U65128 ( .A(n19479), .B(n46315), .X(n19478) );
  nor_x1_sg U65129 ( .A(n21023), .B(n46270), .X(n21022) );
  nor_x1_sg U65130 ( .A(n10917), .B(n46565), .X(n10916) );
  nor_x1_sg U65131 ( .A(n20249), .B(n46295), .X(n20248) );
  nor_x1_sg U65132 ( .A(n21794), .B(n46250), .X(n21793) );
  nor_x1_sg U65133 ( .A(n52449), .B(n46477), .X(n13910) );
  nor_x1_sg U65134 ( .A(n53845), .B(n46364), .X(n17801) );
  nor_x1_sg U65135 ( .A(n54410), .B(n46317), .X(n19346) );
  nor_x1_sg U65136 ( .A(n54978), .B(n46272), .X(n20890) );
  nor_x1_sg U65137 ( .A(n46291), .B(n20108), .X(n20184) );
  nor_x1_sg U65138 ( .A(n46246), .B(n21653), .X(n21729) );
  nor_x1_sg U65139 ( .A(n52725), .B(n46454), .X(n14680) );
  nor_x1_sg U65140 ( .A(n51908), .B(n46521), .X(n12350) );
  nor_x1_sg U65141 ( .A(n43805), .B(n46452), .X(n14848) );
  nor_x1_sg U65142 ( .A(n43035), .B(n46367), .X(n17969) );
  nor_x1_sg U65143 ( .A(n43033), .B(n46320), .X(n19514) );
  nor_x1_sg U65144 ( .A(n43031), .B(n46275), .X(n21058) );
  nor_x1_sg U65145 ( .A(n51453), .B(n10923), .X(n10983) );
  nor_x1_sg U65146 ( .A(n46565), .B(n10655), .X(n10794) );
  nand_x2_sg U65147 ( .A(n46230), .B(n25721), .X(n25730) );
  nand_x2_sg U65148 ( .A(n46226), .B(n26308), .X(n26317) );
  nand_x2_sg U65149 ( .A(n46224), .B(n26587), .X(n26596) );
  nand_x2_sg U65150 ( .A(n46222), .B(n26837), .X(n26846) );
  nand_x2_sg U65151 ( .A(n46222), .B(n26865), .X(n26874) );
  nand_x2_sg U65152 ( .A(n46220), .B(n27144), .X(n27153) );
  nand_x2_sg U65153 ( .A(n46216), .B(n27704), .X(n27713) );
  nand_x2_sg U65154 ( .A(n46214), .B(n27956), .X(n27965) );
  nand_x2_sg U65155 ( .A(n46214), .B(n27984), .X(n27993) );
  nand_x2_sg U65156 ( .A(n46212), .B(n28264), .X(n28273) );
  nand_x2_sg U65157 ( .A(n46210), .B(n28514), .X(n28523) );
  nand_x2_sg U65158 ( .A(n46210), .B(n28542), .X(n28551) );
  nand_x2_sg U65159 ( .A(n46206), .B(n29073), .X(n29082) );
  nand_x2_sg U65160 ( .A(n46206), .B(n29101), .X(n29110) );
  nand_x4_sg U65161 ( .A(n52406), .B(n13768), .X(n13714) );
  nand_x1_sg U65162 ( .A(n52470), .B(n13622), .X(n13768) );
  nand_x2_sg U65163 ( .A(n46226), .B(n26280), .X(n26289) );
  nand_x2_sg U65164 ( .A(n46220), .B(n27116), .X(n27125) );
  nand_x2_sg U65165 ( .A(n46216), .B(n27676), .X(n27685) );
  nor_x1_sg U65166 ( .A(n41588), .B(n46512), .X(n12530) );
  nor_x1_sg U65167 ( .A(n42769), .B(n46467), .X(n14091) );
  nor_x1_sg U65168 ( .A(n51491), .B(n46559), .X(n10966) );
  nand_x4_sg U65169 ( .A(n12252), .B(n12253), .X(n12251) );
  nand_x1_sg U65170 ( .A(n12255), .B(n12256), .X(n12252) );
  nand_x1_sg U65171 ( .A(n12254), .B(n51931), .X(n12253) );
  nand_x1_sg U65172 ( .A(n51931), .B(n46525), .X(n12256) );
  nand_x4_sg U65173 ( .A(n16147), .B(n16148), .X(n16146) );
  nand_x1_sg U65174 ( .A(n16150), .B(n16151), .X(n16147) );
  nand_x1_sg U65175 ( .A(n16149), .B(n53319), .X(n16148) );
  nand_x1_sg U65176 ( .A(n53319), .B(n46413), .X(n16151) );
  nand_x4_sg U65177 ( .A(n11472), .B(n11473), .X(n11471) );
  nand_x1_sg U65178 ( .A(n11475), .B(n11476), .X(n11472) );
  nand_x1_sg U65179 ( .A(n11474), .B(n51650), .X(n11473) );
  nand_x1_sg U65180 ( .A(n51650), .B(n46547), .X(n11476) );
  nand_x4_sg U65181 ( .A(n13033), .B(n13034), .X(n13032) );
  nand_x1_sg U65182 ( .A(n13036), .B(n13037), .X(n13033) );
  nand_x1_sg U65183 ( .A(n13035), .B(n52206), .X(n13034) );
  nand_x1_sg U65184 ( .A(n52206), .B(n46503), .X(n13037) );
  nand_x4_sg U65185 ( .A(n13813), .B(n13814), .X(n13812) );
  nand_x1_sg U65186 ( .A(n13816), .B(n13817), .X(n13813) );
  nand_x1_sg U65187 ( .A(n13815), .B(n52483), .X(n13814) );
  nand_x1_sg U65188 ( .A(n52483), .B(n46481), .X(n13817) );
  nand_x4_sg U65189 ( .A(n15366), .B(n15367), .X(n15365) );
  nand_x1_sg U65190 ( .A(n15369), .B(n15370), .X(n15366) );
  nand_x1_sg U65191 ( .A(n15368), .B(n53040), .X(n15367) );
  nand_x1_sg U65192 ( .A(n53040), .B(n46435), .X(n15370) );
  nand_x4_sg U65193 ( .A(n16932), .B(n16933), .X(n16931) );
  nand_x1_sg U65194 ( .A(n16935), .B(n16936), .X(n16932) );
  nand_x1_sg U65195 ( .A(n16934), .B(n53598), .X(n16933) );
  nand_x1_sg U65196 ( .A(n53598), .B(n46391), .X(n16936) );
  nand_x4_sg U65197 ( .A(n14678), .B(n14679), .X(n14676) );
  nand_x1_sg U65198 ( .A(n14686), .B(n14684), .X(n14678) );
  nand_x1_sg U65199 ( .A(n14680), .B(n52742), .X(n14679) );
  nor_x1_sg U65200 ( .A(n46451), .B(n14547), .X(n14686) );
  nand_x4_sg U65201 ( .A(n17799), .B(n17800), .X(n17797) );
  nand_x1_sg U65202 ( .A(n17807), .B(n17805), .X(n17799) );
  nand_x1_sg U65203 ( .A(n17801), .B(n53862), .X(n17800) );
  nor_x1_sg U65204 ( .A(n46362), .B(n17668), .X(n17807) );
  nand_x4_sg U65205 ( .A(n19344), .B(n19345), .X(n19342) );
  nand_x1_sg U65206 ( .A(n19352), .B(n19350), .X(n19344) );
  nand_x1_sg U65207 ( .A(n19346), .B(n54427), .X(n19345) );
  nor_x1_sg U65208 ( .A(n46315), .B(n19213), .X(n19352) );
  nand_x4_sg U65209 ( .A(n20888), .B(n20889), .X(n20886) );
  nand_x1_sg U65210 ( .A(n20896), .B(n20894), .X(n20888) );
  nand_x1_sg U65211 ( .A(n20890), .B(n54995), .X(n20889) );
  nor_x1_sg U65212 ( .A(n46270), .B(n20757), .X(n20896) );
  nor_x1_sg U65213 ( .A(n46306), .B(n19819), .X(n19818) );
  nor_x1_sg U65214 ( .A(n46261), .B(n21364), .X(n21363) );
  nand_x1_sg U65215 ( .A(n10478), .B(n51288), .X(n10475) );
  nand_x1_sg U65216 ( .A(n46598), .B(n50321), .X(n10029) );
  nand_x1_sg U65217 ( .A(n49326), .B(n46598), .X(n25283) );
  nand_x1_sg U65218 ( .A(n46607), .B(n50658), .X(n9685) );
  nand_x1_sg U65219 ( .A(n46598), .B(n50508), .X(n9836) );
  nand_x1_sg U65220 ( .A(n46598), .B(n50461), .X(n9884) );
  nand_x1_sg U65221 ( .A(n46598), .B(n50415), .X(n9932) );
  nand_x1_sg U65222 ( .A(n46598), .B(n50185), .X(n10175) );
  nand_x1_sg U65223 ( .A(n46607), .B(n50374), .X(n9972) );
  nand_x1_sg U65224 ( .A(n46607), .B(n50281), .X(n10069) );
  nand_x1_sg U65225 ( .A(n46607), .B(n50235), .X(n10118) );
  nand_x1_sg U65226 ( .A(n49799), .B(n46607), .X(n24793) );
  nand_x1_sg U65227 ( .A(n49649), .B(n46598), .X(n24944) );
  nand_x1_sg U65228 ( .A(n49602), .B(n46598), .X(n24992) );
  nand_x1_sg U65229 ( .A(n49556), .B(n46598), .X(n25040) );
  nand_x1_sg U65230 ( .A(n49462), .B(n46598), .X(n25137) );
  nand_x1_sg U65231 ( .A(n49515), .B(n46607), .X(n25080) );
  nand_x1_sg U65232 ( .A(n49422), .B(n46607), .X(n25177) );
  nand_x1_sg U65233 ( .A(n49376), .B(n46607), .X(n25226) );
  nand_x1_sg U65234 ( .A(n50319), .B(n46608), .X(n10028) );
  nand_x1_sg U65235 ( .A(n49460), .B(n46608), .X(n25136) );
  nand_x4_sg U65236 ( .A(n44195), .B(n18197), .X(n18169) );
  nand_x4_sg U65237 ( .A(n44199), .B(n14309), .X(n14279) );
  nand_x4_sg U65238 ( .A(n52478), .B(n13725), .X(n13701) );
  nand_x1_sg U65239 ( .A(n52477), .B(n13726), .X(n13725) );
  nand_x4_sg U65240 ( .A(n13349), .B(n13350), .X(n13347) );
  nand_x1_sg U65241 ( .A(n13352), .B(n13353), .X(n13349) );
  nand_x1_sg U65242 ( .A(n13351), .B(n13268), .X(n13350) );
  nand_x1_sg U65243 ( .A(n13268), .B(n46503), .X(n13353) );
  nand_x4_sg U65244 ( .A(n14129), .B(n14130), .X(n14127) );
  nand_x1_sg U65245 ( .A(n14132), .B(n14133), .X(n14129) );
  nand_x1_sg U65246 ( .A(n14131), .B(n14048), .X(n14130) );
  nand_x1_sg U65247 ( .A(n14048), .B(n46481), .X(n14133) );
  nand_x4_sg U65248 ( .A(n15682), .B(n15683), .X(n15680) );
  nand_x1_sg U65249 ( .A(n15685), .B(n15686), .X(n15682) );
  nand_x1_sg U65250 ( .A(n15684), .B(n15601), .X(n15683) );
  nand_x1_sg U65251 ( .A(n15601), .B(n46435), .X(n15686) );
  nand_x4_sg U65252 ( .A(n17248), .B(n17249), .X(n17246) );
  nand_x1_sg U65253 ( .A(n17251), .B(n17252), .X(n17248) );
  nand_x1_sg U65254 ( .A(n17250), .B(n17167), .X(n17249) );
  nand_x1_sg U65255 ( .A(n17167), .B(n46391), .X(n17252) );
  nand_x4_sg U65256 ( .A(n44203), .B(n11968), .X(n11937) );
  nand_x4_sg U65257 ( .A(n44197), .B(n15863), .X(n15832) );
  nor_x1_sg U65258 ( .A(n16113), .B(n46404), .X(n16456) );
  nor_x1_sg U65259 ( .A(n46516), .B(n12218), .X(n12553) );
  nor_x1_sg U65260 ( .A(n46473), .B(n13779), .X(n14114) );
  nand_x1_sg U65261 ( .A(n50413), .B(n46608), .X(n9931) );
  nand_x1_sg U65262 ( .A(n49554), .B(n46608), .X(n25039) );
  nand_x1_sg U65263 ( .A(n50183), .B(n46608), .X(n10174) );
  nand_x1_sg U65264 ( .A(n49324), .B(n46608), .X(n25282) );
  nand_x4_sg U65265 ( .A(n46525), .B(n11834), .X(n8919) );
  nand_x4_sg U65266 ( .A(n46458), .B(n14175), .X(n9007) );
  nand_x4_sg U65267 ( .A(n46368), .B(n17294), .X(n9269) );
  nand_x4_sg U65268 ( .A(n46348), .B(n18066), .X(n9077) );
  nand_x4_sg U65269 ( .A(n46321), .B(n18839), .X(n9231) );
  nand_x4_sg U65270 ( .A(n46276), .B(n20383), .X(n9155) );
  nand_x4_sg U65271 ( .A(n10486), .B(n10487), .X(n10458) );
  nor_x1_sg U65272 ( .A(n10489), .B(n46565), .X(n10488) );
  nand_x4_sg U65273 ( .A(n19813), .B(n19814), .X(n19785) );
  nor_x1_sg U65274 ( .A(n19816), .B(n46295), .X(n19815) );
  nand_x4_sg U65275 ( .A(n21358), .B(n21359), .X(n21330) );
  nor_x1_sg U65276 ( .A(n21361), .B(n46250), .X(n21360) );
  nand_x4_sg U65277 ( .A(n14750), .B(n52711), .X(n14707) );
  nor_x1_sg U65278 ( .A(n46447), .B(n14674), .X(n14750) );
  nor_x1_sg U65279 ( .A(n46463), .B(n14384), .X(n14383) );
  nor_x1_sg U65280 ( .A(n46416), .B(n15940), .X(n15939) );
  nand_x4_sg U65281 ( .A(n46413), .B(n15729), .X(n9343) );
  nand_x4_sg U65282 ( .A(n46301), .B(n19611), .X(n9191) );
  nand_x4_sg U65283 ( .A(n46256), .B(n21156), .X(n9103) );
  nand_x4_sg U65284 ( .A(n14696), .B(n14697), .X(n14641) );
  nand_x1_sg U65285 ( .A(n14699), .B(n14700), .X(n14696) );
  nand_x1_sg U65286 ( .A(n14698), .B(n52806), .X(n14697) );
  nand_x1_sg U65287 ( .A(n52806), .B(n46458), .X(n14700) );
  nand_x4_sg U65288 ( .A(n17817), .B(n17818), .X(n17762) );
  nand_x1_sg U65289 ( .A(n17820), .B(n17821), .X(n17817) );
  nand_x1_sg U65290 ( .A(n17819), .B(n53926), .X(n17818) );
  nand_x1_sg U65291 ( .A(n53926), .B(n46368), .X(n17821) );
  nand_x4_sg U65292 ( .A(n18584), .B(n18585), .X(n18530) );
  nand_x1_sg U65293 ( .A(n18587), .B(n18588), .X(n18584) );
  nand_x1_sg U65294 ( .A(n18586), .B(n54209), .X(n18585) );
  nand_x1_sg U65295 ( .A(n54209), .B(n46348), .X(n18588) );
  nand_x4_sg U65296 ( .A(n19362), .B(n19363), .X(n19307) );
  nand_x1_sg U65297 ( .A(n19365), .B(n19366), .X(n19362) );
  nand_x1_sg U65298 ( .A(n19364), .B(n54491), .X(n19363) );
  nand_x1_sg U65299 ( .A(n54491), .B(n46321), .X(n19366) );
  nand_x4_sg U65300 ( .A(n20906), .B(n20907), .X(n20851) );
  nand_x1_sg U65301 ( .A(n20909), .B(n20910), .X(n20906) );
  nand_x1_sg U65302 ( .A(n20908), .B(n55059), .X(n20907) );
  nand_x1_sg U65303 ( .A(n55059), .B(n46276), .X(n20910) );
  nand_x4_sg U65304 ( .A(n10815), .B(n10853), .X(n10851) );
  nand_x1_sg U65305 ( .A(n46558), .B(n10814), .X(n10853) );
  nand_x4_sg U65306 ( .A(n10691), .B(n10692), .X(n10690) );
  nand_x1_sg U65307 ( .A(n10694), .B(n10695), .X(n10691) );
  nand_x1_sg U65308 ( .A(n10693), .B(n51377), .X(n10692) );
  nand_x1_sg U65309 ( .A(n51377), .B(n46572), .X(n10695) );
  nand_x4_sg U65310 ( .A(n14583), .B(n14584), .X(n14582) );
  nand_x1_sg U65311 ( .A(n14586), .B(n14587), .X(n14583) );
  nand_x1_sg U65312 ( .A(n14585), .B(n52763), .X(n14584) );
  nand_x1_sg U65313 ( .A(n52763), .B(n46458), .X(n14587) );
  nand_x4_sg U65314 ( .A(n17704), .B(n17705), .X(n17703) );
  nand_x1_sg U65315 ( .A(n17707), .B(n17708), .X(n17704) );
  nand_x1_sg U65316 ( .A(n17706), .B(n53883), .X(n17705) );
  nand_x1_sg U65317 ( .A(n53883), .B(n46368), .X(n17708) );
  nand_x4_sg U65318 ( .A(n19249), .B(n19250), .X(n19248) );
  nand_x1_sg U65319 ( .A(n19252), .B(n19253), .X(n19249) );
  nand_x1_sg U65320 ( .A(n19251), .B(n54448), .X(n19250) );
  nand_x1_sg U65321 ( .A(n54448), .B(n46321), .X(n19253) );
  nand_x4_sg U65322 ( .A(n20793), .B(n20794), .X(n20792) );
  nand_x1_sg U65323 ( .A(n20796), .B(n20797), .X(n20793) );
  nand_x1_sg U65324 ( .A(n20795), .B(n55016), .X(n20794) );
  nand_x1_sg U65325 ( .A(n55016), .B(n46276), .X(n20797) );
  nor_x1_sg U65326 ( .A(n52334), .B(n13243), .X(n13242) );
  nor_x1_sg U65327 ( .A(n52609), .B(n14023), .X(n14022) );
  nor_x1_sg U65328 ( .A(n53168), .B(n15576), .X(n15575) );
  nor_x1_sg U65329 ( .A(n53726), .B(n17142), .X(n17141) );
  nand_x1_sg U65330 ( .A(n46607), .B(n50149), .X(n10210) );
  nand_x1_sg U65331 ( .A(n49290), .B(n46607), .X(n25318) );
  nand_x4_sg U65332 ( .A(n13632), .B(n13633), .X(n13587) );
  nand_x1_sg U65333 ( .A(n13530), .B(n13635), .X(n13632) );
  nand_x1_sg U65334 ( .A(n13634), .B(n46468), .X(n13633) );
  nand_x1_sg U65335 ( .A(n46468), .B(n46481), .X(n13635) );
  nand_x4_sg U65336 ( .A(n20130), .B(n20131), .X(n20075) );
  nand_x1_sg U65337 ( .A(n20133), .B(n20134), .X(n20130) );
  nand_x1_sg U65338 ( .A(n20132), .B(n54776), .X(n20131) );
  nand_x1_sg U65339 ( .A(n54776), .B(n46301), .X(n20134) );
  nand_x4_sg U65340 ( .A(n21675), .B(n21676), .X(n21620) );
  nand_x1_sg U65341 ( .A(n21678), .B(n21679), .X(n21675) );
  nand_x1_sg U65342 ( .A(n21677), .B(n55344), .X(n21676) );
  nand_x1_sg U65343 ( .A(n55344), .B(n46256), .X(n21679) );
  nor_x1_sg U65344 ( .A(n46541), .B(n11434), .X(n11575) );
  nor_x1_sg U65345 ( .A(n46497), .B(n12995), .X(n13136) );
  nor_x1_sg U65346 ( .A(n46429), .B(n15328), .X(n15469) );
  nor_x1_sg U65347 ( .A(n46385), .B(n16894), .X(n17035) );
  nand_x4_sg U65348 ( .A(n12567), .B(n12568), .X(n12566) );
  nand_x1_sg U65349 ( .A(n12570), .B(n12571), .X(n12567) );
  nand_x1_sg U65350 ( .A(n12569), .B(n12487), .X(n12568) );
  nand_x1_sg U65351 ( .A(n12487), .B(n46525), .X(n12571) );
  nor_x1_sg U65352 ( .A(n53375), .B(n16265), .X(n16264) );
  nand_x4_sg U65353 ( .A(n46329), .B(n46343), .X(n18484) );
  nand_x4_sg U65354 ( .A(n46576), .B(n46672), .X(n25394) );
  nand_x4_sg U65355 ( .A(n18473), .B(n18474), .X(n18472) );
  nand_x1_sg U65356 ( .A(n18476), .B(n18477), .X(n18473) );
  nand_x1_sg U65357 ( .A(n18475), .B(n54165), .X(n18474) );
  nand_x1_sg U65358 ( .A(n54165), .B(n46348), .X(n18477) );
  nand_x4_sg U65359 ( .A(n20018), .B(n20019), .X(n20017) );
  nand_x1_sg U65360 ( .A(n20021), .B(n20022), .X(n20018) );
  nand_x1_sg U65361 ( .A(n20020), .B(n54731), .X(n20019) );
  nand_x1_sg U65362 ( .A(n54731), .B(n46301), .X(n20022) );
  nand_x4_sg U65363 ( .A(n21563), .B(n21564), .X(n21562) );
  nand_x1_sg U65364 ( .A(n21566), .B(n21567), .X(n21563) );
  nand_x1_sg U65365 ( .A(n21565), .B(n55299), .X(n21564) );
  nand_x1_sg U65366 ( .A(n55299), .B(n46256), .X(n21567) );
  nand_x4_sg U65367 ( .A(n14378), .B(n14379), .X(n14347) );
  nor_x1_sg U65368 ( .A(n14381), .B(n46454), .X(n14380) );
  nand_x4_sg U65369 ( .A(n46576), .B(n27899), .X(n27622) );
  nand_x4_sg U65370 ( .A(n25740), .B(n25741), .X(n25739) );
  nor_x1_sg U65371 ( .A(n25745), .B(n46236), .X(n25740) );
  nor_x1_sg U65372 ( .A(n25742), .B(n25743), .X(n25741) );
  nand_x4_sg U65373 ( .A(n26018), .B(n26019), .X(n26017) );
  nor_x1_sg U65374 ( .A(n26023), .B(n46236), .X(n26018) );
  nor_x1_sg U65375 ( .A(n26020), .B(n26021), .X(n26019) );
  nand_x4_sg U65376 ( .A(n26299), .B(n26300), .X(n26298) );
  nor_x1_sg U65377 ( .A(n26304), .B(n46236), .X(n26299) );
  nor_x1_sg U65378 ( .A(n26301), .B(n26302), .X(n26300) );
  nand_x4_sg U65379 ( .A(n26578), .B(n26579), .X(n26577) );
  nor_x1_sg U65380 ( .A(n26583), .B(n46236), .X(n26578) );
  nor_x1_sg U65381 ( .A(n26580), .B(n26581), .X(n26579) );
  nand_x4_sg U65382 ( .A(n27135), .B(n27136), .X(n27134) );
  nor_x1_sg U65383 ( .A(n27140), .B(n46236), .X(n27135) );
  nor_x1_sg U65384 ( .A(n27137), .B(n27138), .X(n27136) );
  nand_x4_sg U65385 ( .A(n27415), .B(n27416), .X(n27414) );
  nor_x1_sg U65386 ( .A(n27420), .B(n46236), .X(n27415) );
  nor_x1_sg U65387 ( .A(n27417), .B(n27418), .X(n27416) );
  nand_x4_sg U65388 ( .A(n27695), .B(n27696), .X(n27694) );
  nor_x1_sg U65389 ( .A(n27700), .B(n46236), .X(n27695) );
  nor_x1_sg U65390 ( .A(n27697), .B(n27698), .X(n27696) );
  nand_x4_sg U65391 ( .A(n46572), .B(n10283), .X(n9036) );
  nand_x4_sg U65392 ( .A(n46547), .B(n11051), .X(n8893) );
  nand_x4_sg U65393 ( .A(n46503), .B(n12612), .X(n8853) );
  nand_x4_sg U65394 ( .A(n46435), .B(n14945), .X(n8996) );
  nand_x4_sg U65395 ( .A(n46391), .B(n16511), .X(n9307) );
  nand_x4_sg U65396 ( .A(n46481), .B(n13396), .X(n8809) );
  nand_x2_sg U65397 ( .A(n46204), .B(n29397), .X(n29406) );
  nand_x4_sg U65398 ( .A(n18700), .B(n18701), .X(n18699) );
  nand_x1_sg U65399 ( .A(n18703), .B(n18704), .X(n18700) );
  nand_x1_sg U65400 ( .A(n18702), .B(n54229), .X(n18701) );
  nand_x1_sg U65401 ( .A(n54229), .B(n46339), .X(n18704) );
  nand_x4_sg U65402 ( .A(n25462), .B(n25463), .X(n25461) );
  nor_x1_sg U65403 ( .A(n25467), .B(n46236), .X(n25462) );
  nor_x1_sg U65404 ( .A(n25464), .B(n25465), .X(n25463) );
  nand_x4_sg U65405 ( .A(n26856), .B(n26857), .X(n26855) );
  nor_x1_sg U65406 ( .A(n26861), .B(n46236), .X(n26856) );
  nor_x1_sg U65407 ( .A(n26858), .B(n26859), .X(n26857) );
  nand_x4_sg U65408 ( .A(n27975), .B(n27976), .X(n27974) );
  nor_x1_sg U65409 ( .A(n27980), .B(n46236), .X(n27975) );
  nor_x1_sg U65410 ( .A(n27977), .B(n27978), .X(n27976) );
  nand_x4_sg U65411 ( .A(n28533), .B(n28534), .X(n28532) );
  nor_x1_sg U65412 ( .A(n28538), .B(n46236), .X(n28533) );
  nor_x1_sg U65413 ( .A(n28535), .B(n28536), .X(n28534) );
  nand_x4_sg U65414 ( .A(n29092), .B(n29093), .X(n29091) );
  nor_x1_sg U65415 ( .A(n29097), .B(n46236), .X(n29092) );
  nor_x1_sg U65416 ( .A(n29094), .B(n29095), .X(n29093) );
  nand_x4_sg U65417 ( .A(n26870), .B(n26871), .X(n26869) );
  nor_x1_sg U65418 ( .A(n26875), .B(n46236), .X(n26870) );
  nor_x1_sg U65419 ( .A(n26872), .B(n26873), .X(n26871) );
  nand_x4_sg U65420 ( .A(n27989), .B(n27990), .X(n27988) );
  nor_x1_sg U65421 ( .A(n27994), .B(n46236), .X(n27989) );
  nor_x1_sg U65422 ( .A(n27991), .B(n27992), .X(n27990) );
  nand_x4_sg U65423 ( .A(n28269), .B(n28270), .X(n28268) );
  nor_x1_sg U65424 ( .A(n28274), .B(n46236), .X(n28269) );
  nor_x1_sg U65425 ( .A(n28271), .B(n28272), .X(n28270) );
  nand_x4_sg U65426 ( .A(n28547), .B(n28548), .X(n28546) );
  nor_x1_sg U65427 ( .A(n28552), .B(n46236), .X(n28547) );
  nor_x1_sg U65428 ( .A(n28549), .B(n28550), .X(n28548) );
  nand_x4_sg U65429 ( .A(n29106), .B(n29107), .X(n29105) );
  nor_x1_sg U65430 ( .A(n29111), .B(n46236), .X(n29106) );
  nor_x1_sg U65431 ( .A(n29108), .B(n29109), .X(n29107) );
  nand_x4_sg U65432 ( .A(n46539), .B(n46540), .X(n11343) );
  nand_x4_sg U65433 ( .A(n46495), .B(n46496), .X(n12904) );
  nand_x4_sg U65434 ( .A(n46427), .B(n46428), .X(n15237) );
  nand_x4_sg U65435 ( .A(n46383), .B(n46384), .X(n16803) );
  nand_x4_sg U65436 ( .A(n17525), .B(n17526), .X(n17494) );
  nand_x1_sg U65437 ( .A(n17431), .B(n17528), .X(n17525) );
  nor_x1_sg U65438 ( .A(n17431), .B(n46367), .X(n17527) );
  nand_x4_sg U65439 ( .A(n19070), .B(n19071), .X(n19039) );
  nand_x1_sg U65440 ( .A(n18976), .B(n19073), .X(n19070) );
  nor_x1_sg U65441 ( .A(n18976), .B(n46320), .X(n19072) );
  nand_x4_sg U65442 ( .A(n20614), .B(n20615), .X(n20583) );
  nand_x1_sg U65443 ( .A(n20520), .B(n20617), .X(n20614) );
  nor_x1_sg U65444 ( .A(n20520), .B(n46275), .X(n20616) );
  nor_x1_sg U65445 ( .A(n46591), .B(n55583), .X(\L1_0/n3995 ) );
  nor_x1_sg U65446 ( .A(n44229), .B(n46591), .X(\L1_0/n3994 ) );
  nand_x4_sg U65447 ( .A(n28255), .B(n28256), .X(n28254) );
  nor_x1_sg U65448 ( .A(n28260), .B(n46236), .X(n28255) );
  nor_x1_sg U65449 ( .A(n28257), .B(n28258), .X(n28256) );
  nand_x4_sg U65450 ( .A(n28813), .B(n28814), .X(n28812) );
  nor_x1_sg U65451 ( .A(n28818), .B(n46236), .X(n28813) );
  nor_x1_sg U65452 ( .A(n28815), .B(n28816), .X(n28814) );
  nand_x4_sg U65453 ( .A(n29374), .B(n29375), .X(n29373) );
  nor_x1_sg U65454 ( .A(n29379), .B(n46236), .X(n29374) );
  nor_x1_sg U65455 ( .A(n29376), .B(n29377), .X(n29375) );
  nand_x4_sg U65456 ( .A(n28827), .B(n28828), .X(n28826) );
  nor_x1_sg U65457 ( .A(n28832), .B(n46236), .X(n28827) );
  nor_x1_sg U65458 ( .A(n28829), .B(n28830), .X(n28828) );
  nand_x4_sg U65459 ( .A(n29388), .B(n29389), .X(n29387) );
  nor_x1_sg U65460 ( .A(n29393), .B(n46236), .X(n29388) );
  nor_x1_sg U65461 ( .A(n29390), .B(n29391), .X(n29389) );
  nor_x1_sg U65462 ( .A(n28459), .B(n55599), .X(\L1_0/n3835 ) );
  nor_x1_sg U65463 ( .A(n43908), .B(n28459), .X(\L1_0/n3834 ) );
  nand_x4_sg U65464 ( .A(n10459), .B(n10460), .X(n10454) );
  nand_x1_sg U65465 ( .A(n10462), .B(n10463), .X(n10459) );
  nand_x4_sg U65466 ( .A(n17474), .B(n17475), .X(n17469) );
  nand_x1_sg U65467 ( .A(n17477), .B(n17478), .X(n17474) );
  nand_x4_sg U65468 ( .A(n19019), .B(n19020), .X(n19014) );
  nand_x1_sg U65469 ( .A(n19022), .B(n19023), .X(n19019) );
  nand_x4_sg U65470 ( .A(n20563), .B(n20564), .X(n20558) );
  nand_x1_sg U65471 ( .A(n20566), .B(n20567), .X(n20563) );
  nand_x4_sg U65472 ( .A(n10896), .B(n10897), .X(n10895) );
  nand_x1_sg U65473 ( .A(n10898), .B(n10899), .X(n10897) );
  nor_x1_sg U65474 ( .A(n10900), .B(n51476), .X(n10898) );
  nand_x4_sg U65475 ( .A(n11168), .B(n11169), .X(n11166) );
  nand_x1_sg U65476 ( .A(n11171), .B(n11172), .X(n11168) );
  nand_x4_sg U65477 ( .A(n12729), .B(n12730), .X(n12727) );
  nand_x1_sg U65478 ( .A(n12732), .B(n12733), .X(n12729) );
  nand_x4_sg U65479 ( .A(n15062), .B(n15063), .X(n15060) );
  nand_x1_sg U65480 ( .A(n15065), .B(n15066), .X(n15062) );
  nand_x4_sg U65481 ( .A(n16628), .B(n16629), .X(n16626) );
  nand_x1_sg U65482 ( .A(n16631), .B(n16632), .X(n16628) );
  nor_x1_sg U65483 ( .A(n9802), .B(n9355), .X(\L2_0/n4184 ) );
  nor_x1_sg U65484 ( .A(n9850), .B(n9355), .X(\L2_0/n4180 ) );
  nor_x1_sg U65485 ( .A(n9898), .B(n9355), .X(\L2_0/n4176 ) );
  nor_x1_sg U65486 ( .A(n9946), .B(n9355), .X(\L2_0/n4172 ) );
  nor_x1_sg U65487 ( .A(n9995), .B(n9355), .X(\L2_0/n4168 ) );
  nor_x1_sg U65488 ( .A(n10043), .B(n9355), .X(\L2_0/n4164 ) );
  nor_x1_sg U65489 ( .A(n10092), .B(n9355), .X(\L2_0/n4160 ) );
  nor_x1_sg U65490 ( .A(n10141), .B(n9355), .X(\L2_0/n4156 ) );
  nor_x1_sg U65491 ( .A(n10188), .B(n9355), .X(\L2_0/n4152 ) );
  nand_x4_sg U65492 ( .A(n11055), .B(n11056), .X(n8897) );
  nand_x4_sg U65493 ( .A(n11838), .B(n11839), .X(n8931) );
  nand_x4_sg U65494 ( .A(n15733), .B(n15734), .X(n9326) );
  nand_x4_sg U65495 ( .A(n17298), .B(n17299), .X(n9277) );
  nand_x4_sg U65496 ( .A(n18843), .B(n18844), .X(n9239) );
  nand_x4_sg U65497 ( .A(n20387), .B(n20388), .X(n9163) );
  nand_x4_sg U65498 ( .A(n16243), .B(n16244), .X(n16241) );
  nand_x1_sg U65499 ( .A(n16251), .B(n16249), .X(n16243) );
  nor_x1_sg U65500 ( .A(n46406), .B(n16109), .X(n16251) );
  nor_x1_sg U65501 ( .A(n46616), .B(n55615), .X(\L1_0/n3675 ) );
  nor_x1_sg U65502 ( .A(n44219), .B(n46616), .X(\L1_0/n3674 ) );
  nor_x1_sg U65503 ( .A(n46615), .B(n25510), .X(\L1_0/n4675 ) );
  nand_x4_sg U65504 ( .A(n15934), .B(n15935), .X(n15903) );
  nor_x1_sg U65505 ( .A(n15937), .B(n46409), .X(n15936) );
  nor_x1_sg U65506 ( .A(n46625), .B(n55552), .X(\L1_0/n4315 ) );
  nor_x1_sg U65507 ( .A(n46625), .B(n44235), .X(\L1_0/n4314 ) );
  nand_x4_sg U65508 ( .A(n14179), .B(n14180), .X(n9011) );
  nand_x4_sg U65509 ( .A(n46329), .B(n46333), .X(n18742) );
  nand_x4_sg U65510 ( .A(n26313), .B(n26314), .X(n26312) );
  nor_x1_sg U65511 ( .A(n26318), .B(n46236), .X(n26313) );
  nor_x1_sg U65512 ( .A(n26315), .B(n26316), .X(n26314) );
  nand_x4_sg U65513 ( .A(n26592), .B(n26593), .X(n26591) );
  nor_x1_sg U65514 ( .A(n26597), .B(n46236), .X(n26592) );
  nor_x1_sg U65515 ( .A(n26594), .B(n26595), .X(n26593) );
  nand_x4_sg U65516 ( .A(n27149), .B(n27150), .X(n27148) );
  nor_x1_sg U65517 ( .A(n27154), .B(n46236), .X(n27149) );
  nor_x1_sg U65518 ( .A(n27151), .B(n27152), .X(n27150) );
  nand_x4_sg U65519 ( .A(n27709), .B(n27710), .X(n27708) );
  nor_x1_sg U65520 ( .A(n27714), .B(n46236), .X(n27709) );
  nor_x1_sg U65521 ( .A(n27711), .B(n27712), .X(n27710) );
  nor_x1_sg U65522 ( .A(n46585), .B(n26348), .X(\L1_0/n4435 ) );
  nor_x1_sg U65523 ( .A(n55542), .B(n46585), .X(\L1_0/n4434 ) );
  nor_x1_sg U65524 ( .A(n46587), .B(n26627), .X(\L1_0/n4355 ) );
  nor_x1_sg U65525 ( .A(n55550), .B(n46587), .X(\L1_0/n4354 ) );
  nor_x1_sg U65526 ( .A(n46591), .B(n28023), .X(\L1_0/n3955 ) );
  nor_x1_sg U65527 ( .A(n55589), .B(n46591), .X(\L1_0/n3954 ) );
  nor_x1_sg U65528 ( .A(n28459), .B(n28581), .X(\L1_0/n3795 ) );
  nor_x1_sg U65529 ( .A(n55605), .B(n28459), .X(\L1_0/n3794 ) );
  nor_x1_sg U65530 ( .A(n46596), .B(n29422), .X(\L1_0/n3555 ) );
  nor_x1_sg U65531 ( .A(n55629), .B(n46596), .X(\L1_0/n3554 ) );
  nor_x1_sg U65532 ( .A(n46625), .B(n26904), .X(\L1_0/n4275 ) );
  nor_x1_sg U65533 ( .A(n46611), .B(n25788), .X(\L1_0/n4595 ) );
  nor_x1_sg U65534 ( .A(n46623), .B(n27463), .X(\L1_0/n4115 ) );
  nor_x1_sg U65535 ( .A(n46621), .B(n27744), .X(\L1_0/n4035 ) );
  nor_x1_sg U65536 ( .A(n46619), .B(n28861), .X(\L1_0/n3715 ) );
  nand_x4_sg U65537 ( .A(n10512), .B(n10513), .X(n10480) );
  nand_x1_sg U65538 ( .A(n10418), .B(n10515), .X(n10512) );
  nand_x4_sg U65539 ( .A(n19839), .B(n19840), .X(n19807) );
  nand_x1_sg U65540 ( .A(n19745), .B(n19842), .X(n19839) );
  nand_x4_sg U65541 ( .A(n21384), .B(n21385), .X(n21352) );
  nand_x1_sg U65542 ( .A(n21290), .B(n21387), .X(n21384) );
  nand_x4_sg U65543 ( .A(n10804), .B(n10805), .X(n10749) );
  nand_x1_sg U65544 ( .A(n10807), .B(n10808), .X(n10804) );
  nand_x1_sg U65545 ( .A(n10806), .B(n51418), .X(n10805) );
  nand_x1_sg U65546 ( .A(n51418), .B(n46572), .X(n10808) );
  nor_x1_sg U65547 ( .A(n9354), .B(n9355), .X(\L2_0/n4220 ) );
  nor_x1_sg U65548 ( .A(n9416), .B(n9355), .X(\L2_0/n4216 ) );
  nor_x1_sg U65549 ( .A(n9465), .B(n9355), .X(\L2_0/n4212 ) );
  nor_x1_sg U65550 ( .A(n9514), .B(n9355), .X(\L2_0/n4208 ) );
  nor_x1_sg U65551 ( .A(n9563), .B(n9355), .X(\L2_0/n4204 ) );
  nor_x1_sg U65552 ( .A(n9611), .B(n9355), .X(\L2_0/n4200 ) );
  nor_x1_sg U65553 ( .A(n9659), .B(n9355), .X(\L2_0/n4196 ) );
  nor_x1_sg U65554 ( .A(n9706), .B(n9355), .X(\L2_0/n4192 ) );
  nor_x1_sg U65555 ( .A(n9754), .B(n9355), .X(\L2_0/n4188 ) );
  nand_x4_sg U65556 ( .A(n25426), .B(n25427), .X(n25425) );
  nor_x1_sg U65557 ( .A(n25431), .B(n46236), .X(n25426) );
  nor_x1_sg U65558 ( .A(n25428), .B(n25429), .X(n25427) );
  nand_x4_sg U65559 ( .A(n27940), .B(n27941), .X(n27939) );
  nor_x1_sg U65560 ( .A(n27945), .B(n46236), .X(n27940) );
  nor_x1_sg U65561 ( .A(n27942), .B(n27943), .X(n27941) );
  nand_x4_sg U65562 ( .A(n28498), .B(n28499), .X(n28497) );
  nor_x1_sg U65563 ( .A(n28503), .B(n46236), .X(n28498) );
  nor_x1_sg U65564 ( .A(n28500), .B(n28501), .X(n28499) );
  nand_x4_sg U65565 ( .A(n29057), .B(n29058), .X(n29056) );
  nor_x1_sg U65566 ( .A(n29062), .B(n46236), .X(n29057) );
  nor_x1_sg U65567 ( .A(n29059), .B(n29060), .X(n29058) );
  nor_x1_sg U65568 ( .A(n46589), .B(n27184), .X(\L1_0/n4195 ) );
  nor_x1_sg U65569 ( .A(n55566), .B(n46589), .X(\L1_0/n4194 ) );
  nor_x1_sg U65570 ( .A(n46593), .B(n28282), .X(\L1_0/n3887 ) );
  nor_x1_sg U65571 ( .A(n55739), .B(n46593), .X(\L1_0/n3886 ) );
  nor_x1_sg U65572 ( .A(n46593), .B(n28289), .X(\L1_0/n3883 ) );
  nor_x1_sg U65573 ( .A(n55595), .B(n46593), .X(\L1_0/n3882 ) );
  nor_x1_sg U65574 ( .A(n46593), .B(n28294), .X(\L1_0/n3879 ) );
  nor_x1_sg U65575 ( .A(n55596), .B(n46593), .X(\L1_0/n3878 ) );
  nor_x1_sg U65576 ( .A(n46593), .B(n28303), .X(\L1_0/n3875 ) );
  nor_x1_sg U65577 ( .A(n55597), .B(n46593), .X(\L1_0/n3874 ) );
  nand_x4_sg U65578 ( .A(n25447), .B(n25448), .X(n25446) );
  nor_x1_sg U65579 ( .A(n25452), .B(n46236), .X(n25447) );
  nor_x1_sg U65580 ( .A(n25449), .B(n25450), .X(n25448) );
  nand_x4_sg U65581 ( .A(n28240), .B(n28241), .X(n28239) );
  nor_x1_sg U65582 ( .A(n28245), .B(n46236), .X(n28240) );
  nor_x1_sg U65583 ( .A(n28242), .B(n28243), .X(n28241) );
  nand_x4_sg U65584 ( .A(n26564), .B(n26565), .X(n26563) );
  nor_x1_sg U65585 ( .A(n26569), .B(n46236), .X(n26564) );
  nor_x1_sg U65586 ( .A(n26566), .B(n26567), .X(n26565) );
  nand_x4_sg U65587 ( .A(n27401), .B(n27402), .X(n27400) );
  nor_x1_sg U65588 ( .A(n27406), .B(n46236), .X(n27401) );
  nor_x1_sg U65589 ( .A(n27403), .B(n27404), .X(n27402) );
  nand_x4_sg U65590 ( .A(n25476), .B(n25477), .X(n25475) );
  nor_x1_sg U65591 ( .A(n25481), .B(n46236), .X(n25476) );
  nor_x1_sg U65592 ( .A(n25478), .B(n25479), .X(n25477) );
  nand_x4_sg U65593 ( .A(n25754), .B(n25755), .X(n25753) );
  nor_x1_sg U65594 ( .A(n25759), .B(n46236), .X(n25754) );
  nor_x1_sg U65595 ( .A(n25756), .B(n25757), .X(n25755) );
  nand_x4_sg U65596 ( .A(n25983), .B(n25984), .X(n25982) );
  nor_x1_sg U65597 ( .A(n25988), .B(n46236), .X(n25983) );
  nor_x1_sg U65598 ( .A(n25985), .B(n25986), .X(n25984) );
  nand_x4_sg U65599 ( .A(n27380), .B(n27381), .X(n27379) );
  nor_x1_sg U65600 ( .A(n27385), .B(n46236), .X(n27380) );
  nor_x1_sg U65601 ( .A(n27382), .B(n27383), .X(n27381) );
  inv_x4_sg U65602 ( .A(n44169), .X(n46618) );
  nand_x4_sg U65603 ( .A(n28798), .B(n28799), .X(n28797) );
  nor_x1_sg U65604 ( .A(n28803), .B(n46236), .X(n28798) );
  nor_x1_sg U65605 ( .A(n28800), .B(n28801), .X(n28799) );
  nand_x4_sg U65606 ( .A(n29359), .B(n29360), .X(n29358) );
  nor_x1_sg U65607 ( .A(n29364), .B(n46236), .X(n29359) );
  nor_x1_sg U65608 ( .A(n29361), .B(n29362), .X(n29360) );
  nand_x4_sg U65609 ( .A(n13851), .B(n13852), .X(n13788) );
  nand_x1_sg U65610 ( .A(n13783), .B(n13785), .X(n13851) );
  nand_x1_sg U65611 ( .A(n13853), .B(n13818), .X(n13852) );
  nand_x4_sg U65612 ( .A(n14622), .B(n14623), .X(n14559) );
  nand_x1_sg U65613 ( .A(n14554), .B(n14556), .X(n14622) );
  nand_x1_sg U65614 ( .A(n14624), .B(n14588), .X(n14623) );
  nand_x4_sg U65615 ( .A(n17743), .B(n17744), .X(n17680) );
  nand_x1_sg U65616 ( .A(n17675), .B(n17677), .X(n17743) );
  nand_x1_sg U65617 ( .A(n17745), .B(n17709), .X(n17744) );
  nand_x4_sg U65618 ( .A(n19288), .B(n19289), .X(n19225) );
  nand_x1_sg U65619 ( .A(n19220), .B(n19222), .X(n19288) );
  nand_x1_sg U65620 ( .A(n19290), .B(n19254), .X(n19289) );
  nand_x4_sg U65621 ( .A(n20832), .B(n20833), .X(n20769) );
  nand_x1_sg U65622 ( .A(n20764), .B(n20766), .X(n20832) );
  nand_x1_sg U65623 ( .A(n20834), .B(n20798), .X(n20833) );
  nand_x4_sg U65624 ( .A(n26004), .B(n26005), .X(n26003) );
  nor_x1_sg U65625 ( .A(n26009), .B(n46236), .X(n26004) );
  nor_x1_sg U65626 ( .A(n26006), .B(n26007), .X(n26005) );
  inv_x4_sg U65627 ( .A(n29627), .X(n46610) );
  nand_x4_sg U65628 ( .A(n18568), .B(n18569), .X(n18483) );
  nand_x1_sg U65629 ( .A(n18571), .B(n18572), .X(n18568) );
  nand_x4_sg U65630 ( .A(n12545), .B(n12546), .X(n12542) );
  nand_x1_sg U65631 ( .A(n12549), .B(n12550), .X(n12545) );
  nand_x1_sg U65632 ( .A(n12547), .B(n51952), .X(n12546) );
  nor_x1_sg U65633 ( .A(n46523), .B(n12404), .X(n12549) );
  nand_x4_sg U65634 ( .A(n13326), .B(n13327), .X(n13323) );
  nand_x1_sg U65635 ( .A(n13330), .B(n13331), .X(n13326) );
  nand_x1_sg U65636 ( .A(n13328), .B(n52227), .X(n13327) );
  nor_x1_sg U65637 ( .A(n46501), .B(n13184), .X(n13330) );
  nand_x4_sg U65638 ( .A(n14106), .B(n14107), .X(n14103) );
  nand_x1_sg U65639 ( .A(n14110), .B(n14111), .X(n14106) );
  nand_x1_sg U65640 ( .A(n14108), .B(n52504), .X(n14107) );
  nor_x1_sg U65641 ( .A(n46479), .B(n13964), .X(n14110) );
  nand_x4_sg U65642 ( .A(n15659), .B(n15660), .X(n15656) );
  nand_x1_sg U65643 ( .A(n15663), .B(n15664), .X(n15659) );
  nand_x1_sg U65644 ( .A(n15661), .B(n53061), .X(n15660) );
  nor_x1_sg U65645 ( .A(n46433), .B(n15517), .X(n15663) );
  nand_x4_sg U65646 ( .A(n17225), .B(n17226), .X(n17222) );
  nand_x1_sg U65647 ( .A(n17229), .B(n17230), .X(n17225) );
  nand_x1_sg U65648 ( .A(n17227), .B(n53619), .X(n17226) );
  nor_x1_sg U65649 ( .A(n46389), .B(n17083), .X(n17229) );
  nand_x4_sg U65650 ( .A(n12456), .B(n12457), .X(n12454) );
  nand_x1_sg U65651 ( .A(n12458), .B(n52037), .X(n12457) );
  nand_x1_sg U65652 ( .A(n12460), .B(n51952), .X(n12456) );
  nor_x1_sg U65653 ( .A(n12459), .B(n52057), .X(n12458) );
  nand_x4_sg U65654 ( .A(n17909), .B(n17910), .X(n17907) );
  nand_x1_sg U65655 ( .A(n17911), .B(n17912), .X(n17910) );
  nand_x1_sg U65656 ( .A(n17915), .B(n53903), .X(n17909) );
  nor_x1_sg U65657 ( .A(n17913), .B(n17914), .X(n17911) );
  nand_x4_sg U65658 ( .A(n19454), .B(n19455), .X(n19452) );
  nand_x1_sg U65659 ( .A(n19456), .B(n19457), .X(n19455) );
  nand_x1_sg U65660 ( .A(n19460), .B(n54468), .X(n19454) );
  nor_x1_sg U65661 ( .A(n19458), .B(n19459), .X(n19456) );
  nand_x4_sg U65662 ( .A(n20998), .B(n20999), .X(n20996) );
  nand_x1_sg U65663 ( .A(n21000), .B(n21001), .X(n20999) );
  nand_x1_sg U65664 ( .A(n21004), .B(n55036), .X(n20998) );
  nor_x1_sg U65665 ( .A(n21002), .B(n21003), .X(n21000) );
  nand_x4_sg U65666 ( .A(n26821), .B(n26822), .X(n26820) );
  nor_x1_sg U65667 ( .A(n26826), .B(n46236), .X(n26821) );
  nor_x1_sg U65668 ( .A(n26823), .B(n26824), .X(n26822) );
  nand_x4_sg U65669 ( .A(n28219), .B(n28220), .X(n28218) );
  nor_x1_sg U65670 ( .A(n28224), .B(n46236), .X(n28219) );
  nor_x1_sg U65671 ( .A(n28221), .B(n28222), .X(n28220) );
  nand_x4_sg U65672 ( .A(n28777), .B(n28778), .X(n28776) );
  nor_x1_sg U65673 ( .A(n28782), .B(n46236), .X(n28777) );
  nor_x1_sg U65674 ( .A(n28779), .B(n28780), .X(n28778) );
  nand_x4_sg U65675 ( .A(n29338), .B(n29339), .X(n29337) );
  nor_x1_sg U65676 ( .A(n29343), .B(n46236), .X(n29338) );
  nor_x1_sg U65677 ( .A(n29340), .B(n29341), .X(n29339) );
  nand_x4_sg U65678 ( .A(n18294), .B(n18295), .X(n18262) );
  nand_x1_sg U65679 ( .A(n18198), .B(n18297), .X(n18294) );
  nor_x1_sg U65680 ( .A(n18198), .B(n46341), .X(n18296) );
  nand_x4_sg U65681 ( .A(n14375), .B(n14376), .X(n14364) );
  nor_x1_sg U65682 ( .A(n14377), .B(n46449), .X(n14376) );
  nor_x1_sg U65683 ( .A(n14316), .B(n52690), .X(n14375) );
  nand_x4_sg U65684 ( .A(n16502), .B(n16503), .X(n16335) );
  nand_x1_sg U65685 ( .A(n16109), .B(n16504), .X(n16502) );
  nand_x4_sg U65686 ( .A(n14166), .B(n14167), .X(n14001) );
  nor_x1_sg U65687 ( .A(n46559), .B(n25444), .X(n25443) );
  nand_x2_sg U65688 ( .A(n46232), .B(n25435), .X(n25444) );
  nor_x1_sg U65689 ( .A(n29577), .B(n46233), .X(\L1_0/n3507 ) );
  nor_x1_sg U65690 ( .A(n24472), .B(n46233), .X(\L1_0/n4823 ) );
  nor_x1_sg U65691 ( .A(n24622), .B(n46233), .X(\L1_0/n4811 ) );
  nor_x1_sg U65692 ( .A(n24767), .B(n46233), .X(\L1_0/n4799 ) );
  nor_x1_sg U65693 ( .A(n24910), .B(n46233), .X(\L1_0/n4787 ) );
  nor_x1_sg U65694 ( .A(n25054), .B(n46233), .X(\L1_0/n4775 ) );
  nor_x1_sg U65695 ( .A(n25200), .B(n46233), .X(\L1_0/n4763 ) );
  nor_x1_sg U65696 ( .A(n12315), .B(n12316), .X(n12314) );
  nor_x1_sg U65697 ( .A(n16210), .B(n16211), .X(n16209) );
  nand_x4_sg U65698 ( .A(n26032), .B(n26033), .X(n26031) );
  nor_x1_sg U65699 ( .A(n26037), .B(n46236), .X(n26032) );
  nor_x1_sg U65700 ( .A(n26034), .B(n26035), .X(n26033) );
  nand_x4_sg U65701 ( .A(n27429), .B(n27430), .X(n27428) );
  nor_x1_sg U65702 ( .A(n27434), .B(n46236), .X(n27429) );
  nor_x1_sg U65703 ( .A(n27431), .B(n27432), .X(n27430) );
  nand_x4_sg U65704 ( .A(n25705), .B(n25706), .X(n25704) );
  nor_x1_sg U65705 ( .A(n25710), .B(n46236), .X(n25705) );
  nor_x1_sg U65706 ( .A(n25707), .B(n25708), .X(n25706) );
  nand_x4_sg U65707 ( .A(n26264), .B(n26265), .X(n26263) );
  nor_x1_sg U65708 ( .A(n26269), .B(n46236), .X(n26264) );
  nor_x1_sg U65709 ( .A(n26266), .B(n26267), .X(n26265) );
  nand_x4_sg U65710 ( .A(n26543), .B(n26544), .X(n26542) );
  nor_x1_sg U65711 ( .A(n26548), .B(n46236), .X(n26543) );
  nor_x1_sg U65712 ( .A(n26545), .B(n26546), .X(n26544) );
  nand_x4_sg U65713 ( .A(n27100), .B(n27101), .X(n27099) );
  nor_x1_sg U65714 ( .A(n27105), .B(n46236), .X(n27100) );
  nor_x1_sg U65715 ( .A(n27102), .B(n27103), .X(n27101) );
  nand_x4_sg U65716 ( .A(n27660), .B(n27661), .X(n27659) );
  nor_x1_sg U65717 ( .A(n27665), .B(n46236), .X(n27660) );
  nor_x1_sg U65718 ( .A(n27662), .B(n27663), .X(n27661) );
  nor_x1_sg U65719 ( .A(n46512), .B(n26001), .X(n26000) );
  nand_x2_sg U65720 ( .A(n46228), .B(n25992), .X(n26001) );
  nor_x1_sg U65721 ( .A(n46467), .B(n26561), .X(n26560) );
  nand_x2_sg U65722 ( .A(n46224), .B(n26552), .X(n26561) );
  nor_x1_sg U65723 ( .A(n46400), .B(n27398), .X(n27397) );
  nand_x2_sg U65724 ( .A(n46218), .B(n27389), .X(n27398) );
  nor_x1_sg U65725 ( .A(n46287), .B(n28795), .X(n28794) );
  nand_x2_sg U65726 ( .A(n46208), .B(n28786), .X(n28795) );
  nor_x1_sg U65727 ( .A(n46242), .B(n29356), .X(n29355) );
  nand_x2_sg U65728 ( .A(n46204), .B(n29347), .X(n29356) );
  nor_x1_sg U65729 ( .A(n46535), .B(n25723), .X(n25722) );
  nand_x2_sg U65730 ( .A(n46230), .B(n25714), .X(n25723) );
  nor_x1_sg U65731 ( .A(n46491), .B(n26282), .X(n26281) );
  nand_x2_sg U65732 ( .A(n46226), .B(n26273), .X(n26282) );
  nor_x1_sg U65733 ( .A(n46423), .B(n27118), .X(n27117) );
  nand_x2_sg U65734 ( .A(n46220), .B(n27109), .X(n27118) );
  nor_x1_sg U65735 ( .A(n46379), .B(n27678), .X(n27677) );
  nand_x2_sg U65736 ( .A(n46216), .B(n27669), .X(n27678) );
  nor_x1_sg U65737 ( .A(n46331), .B(n28237), .X(n28236) );
  nand_x2_sg U65738 ( .A(n46212), .B(n28228), .X(n28237) );
  nand_x4_sg U65739 ( .A(n25768), .B(n25769), .X(n25767) );
  nor_x1_sg U65740 ( .A(n42487), .B(n25771), .X(n25769) );
  nor_x1_sg U65741 ( .A(n25773), .B(n46236), .X(n25768) );
  nand_x4_sg U65742 ( .A(n26884), .B(n26885), .X(n26883) );
  nor_x1_sg U65743 ( .A(n26886), .B(n26887), .X(n26885) );
  nor_x1_sg U65744 ( .A(n26889), .B(n46236), .X(n26884) );
  nand_x4_sg U65745 ( .A(n27443), .B(n27444), .X(n27442) );
  nor_x1_sg U65746 ( .A(n42477), .B(n27446), .X(n27444) );
  nor_x1_sg U65747 ( .A(n27448), .B(n46236), .X(n27443) );
  nand_x4_sg U65748 ( .A(n28003), .B(n28004), .X(n28002) );
  nor_x1_sg U65749 ( .A(n28005), .B(n28006), .X(n28004) );
  nor_x1_sg U65750 ( .A(n28008), .B(n46236), .X(n28003) );
  nand_x4_sg U65751 ( .A(n28283), .B(n28284), .X(n28282) );
  nor_x1_sg U65752 ( .A(n28285), .B(n28286), .X(n28284) );
  nor_x1_sg U65753 ( .A(n28288), .B(n46236), .X(n28283) );
  nand_x4_sg U65754 ( .A(n28561), .B(n28562), .X(n28560) );
  nor_x1_sg U65755 ( .A(n28563), .B(n28564), .X(n28562) );
  nor_x1_sg U65756 ( .A(n28566), .B(n46236), .X(n28561) );
  nand_x4_sg U65757 ( .A(n28841), .B(n28842), .X(n28840) );
  nor_x1_sg U65758 ( .A(n28843), .B(n28844), .X(n28842) );
  nor_x1_sg U65759 ( .A(n28846), .B(n46236), .X(n28841) );
  nand_x4_sg U65760 ( .A(n29120), .B(n29121), .X(n29119) );
  nor_x1_sg U65761 ( .A(n29122), .B(n29123), .X(n29121) );
  nor_x1_sg U65762 ( .A(n29125), .B(n46236), .X(n29120) );
  nand_x4_sg U65763 ( .A(n29402), .B(n29403), .X(n29401) );
  nor_x1_sg U65764 ( .A(n29407), .B(n46236), .X(n29402) );
  nor_x1_sg U65765 ( .A(n29404), .B(n29405), .X(n29403) );
  nand_x4_sg U65766 ( .A(n25726), .B(n25727), .X(n25725) );
  nor_x1_sg U65767 ( .A(n25731), .B(n46236), .X(n25726) );
  nor_x1_sg U65768 ( .A(n25728), .B(n25729), .X(n25727) );
  nand_x4_sg U65769 ( .A(n26842), .B(n26843), .X(n26841) );
  nor_x1_sg U65770 ( .A(n26847), .B(n46236), .X(n26842) );
  nor_x1_sg U65771 ( .A(n26844), .B(n26845), .X(n26843) );
  nand_x4_sg U65772 ( .A(n27961), .B(n27962), .X(n27960) );
  nor_x1_sg U65773 ( .A(n27966), .B(n46236), .X(n27961) );
  nor_x1_sg U65774 ( .A(n27963), .B(n27964), .X(n27962) );
  nand_x4_sg U65775 ( .A(n28519), .B(n28520), .X(n28518) );
  nor_x1_sg U65776 ( .A(n28524), .B(n46236), .X(n28519) );
  nor_x1_sg U65777 ( .A(n28521), .B(n28522), .X(n28520) );
  nand_x4_sg U65778 ( .A(n29078), .B(n29079), .X(n29077) );
  nor_x1_sg U65779 ( .A(n29083), .B(n46236), .X(n29078) );
  nor_x1_sg U65780 ( .A(n29080), .B(n29081), .X(n29079) );
  nand_x4_sg U65781 ( .A(n26285), .B(n26286), .X(n26284) );
  nor_x1_sg U65782 ( .A(n26290), .B(n46236), .X(n26285) );
  nor_x1_sg U65783 ( .A(n26287), .B(n26288), .X(n26286) );
  nand_x4_sg U65784 ( .A(n27121), .B(n27122), .X(n27120) );
  nor_x1_sg U65785 ( .A(n27126), .B(n46236), .X(n27121) );
  nor_x1_sg U65786 ( .A(n27123), .B(n27124), .X(n27122) );
  nand_x4_sg U65787 ( .A(n27681), .B(n27682), .X(n27680) );
  nor_x1_sg U65788 ( .A(n27686), .B(n46236), .X(n27681) );
  nor_x1_sg U65789 ( .A(n27683), .B(n27684), .X(n27682) );
  nand_x4_sg U65790 ( .A(n18268), .B(n18269), .X(n18240) );
  nor_x1_sg U65791 ( .A(n46353), .B(n18274), .X(n18272) );
  nand_x4_sg U65792 ( .A(n11942), .B(n11943), .X(n11845) );
  nand_x1_sg U65793 ( .A(n11945), .B(n11946), .X(n11942) );
  nand_x4_sg U65794 ( .A(n15837), .B(n15838), .X(n15740) );
  nand_x1_sg U65795 ( .A(n15840), .B(n15841), .X(n15837) );
  nand_x4_sg U65796 ( .A(n17403), .B(n17404), .X(n17305) );
  nand_x1_sg U65797 ( .A(n17406), .B(n17407), .X(n17403) );
  nand_x4_sg U65798 ( .A(n18948), .B(n18949), .X(n18850) );
  nand_x1_sg U65799 ( .A(n18951), .B(n18952), .X(n18948) );
  nand_x4_sg U65800 ( .A(n20492), .B(n20493), .X(n20394) );
  nand_x1_sg U65801 ( .A(n20495), .B(n20496), .X(n20492) );
  nand_x4_sg U65802 ( .A(n14284), .B(n14285), .X(n14186) );
  nand_x1_sg U65803 ( .A(n14287), .B(n14288), .X(n14284) );
  nand_x4_sg U65804 ( .A(n25497), .B(n46235), .X(n25496) );
  nor_x1_sg U65805 ( .A(n25498), .B(n25499), .X(n25497) );
  nand_x4_sg U65806 ( .A(n25502), .B(n46235), .X(n25501) );
  nor_x1_sg U65807 ( .A(n25503), .B(n25504), .X(n25502) );
  nand_x4_sg U65808 ( .A(n25775), .B(n46235), .X(n25774) );
  nor_x1_sg U65809 ( .A(n25776), .B(n25777), .X(n25775) );
  nand_x4_sg U65810 ( .A(n25780), .B(n46235), .X(n25779) );
  nor_x1_sg U65811 ( .A(n25781), .B(n25782), .X(n25780) );
  nand_x4_sg U65812 ( .A(n26054), .B(n46235), .X(n26053) );
  nor_x1_sg U65813 ( .A(n26055), .B(n26056), .X(n26054) );
  nand_x4_sg U65814 ( .A(n26059), .B(n46235), .X(n26058) );
  nor_x1_sg U65815 ( .A(n26060), .B(n26061), .X(n26059) );
  nand_x4_sg U65816 ( .A(n26335), .B(n46235), .X(n26334) );
  nor_x1_sg U65817 ( .A(n26336), .B(n26337), .X(n26335) );
  nand_x4_sg U65818 ( .A(n26340), .B(n46235), .X(n26339) );
  nor_x1_sg U65819 ( .A(n26341), .B(n26342), .X(n26340) );
  nand_x4_sg U65820 ( .A(n26891), .B(n46235), .X(n26890) );
  nor_x1_sg U65821 ( .A(n26892), .B(n26893), .X(n26891) );
  nand_x4_sg U65822 ( .A(n27171), .B(n46235), .X(n27170) );
  nor_x1_sg U65823 ( .A(n27172), .B(n27173), .X(n27171) );
  nand_x4_sg U65824 ( .A(n27176), .B(n46235), .X(n27175) );
  nor_x1_sg U65825 ( .A(n27177), .B(n27178), .X(n27176) );
  nand_x4_sg U65826 ( .A(n27450), .B(n46235), .X(n27449) );
  nor_x1_sg U65827 ( .A(n27451), .B(n27452), .X(n27450) );
  nand_x4_sg U65828 ( .A(n27455), .B(n46235), .X(n27454) );
  nor_x1_sg U65829 ( .A(n27456), .B(n27457), .X(n27455) );
  nand_x4_sg U65830 ( .A(n27731), .B(n46235), .X(n27730) );
  nor_x1_sg U65831 ( .A(n27732), .B(n27733), .X(n27731) );
  nand_x4_sg U65832 ( .A(n27736), .B(n46235), .X(n27735) );
  nor_x1_sg U65833 ( .A(n27737), .B(n27738), .X(n27736) );
  nand_x4_sg U65834 ( .A(n28010), .B(n46235), .X(n28009) );
  nor_x1_sg U65835 ( .A(n28011), .B(n28012), .X(n28010) );
  nand_x4_sg U65836 ( .A(n28015), .B(n46235), .X(n28014) );
  nor_x1_sg U65837 ( .A(n28016), .B(n28017), .X(n28015) );
  nand_x4_sg U65838 ( .A(n28290), .B(n46235), .X(n28289) );
  nor_x1_sg U65839 ( .A(n28291), .B(n28292), .X(n28290) );
  nand_x4_sg U65840 ( .A(n28295), .B(n46235), .X(n28294) );
  nor_x1_sg U65841 ( .A(n28296), .B(n28297), .X(n28295) );
  nand_x4_sg U65842 ( .A(n28568), .B(n46235), .X(n28567) );
  nor_x1_sg U65843 ( .A(n28569), .B(n28570), .X(n28568) );
  nand_x4_sg U65844 ( .A(n28573), .B(n46235), .X(n28572) );
  nor_x1_sg U65845 ( .A(n28574), .B(n28575), .X(n28573) );
  nand_x4_sg U65846 ( .A(n28848), .B(n46235), .X(n28847) );
  nor_x1_sg U65847 ( .A(n28849), .B(n28850), .X(n28848) );
  nand_x4_sg U65848 ( .A(n28853), .B(n46235), .X(n28852) );
  nor_x1_sg U65849 ( .A(n28854), .B(n28855), .X(n28853) );
  nand_x4_sg U65850 ( .A(n29127), .B(n46235), .X(n29126) );
  nor_x1_sg U65851 ( .A(n29128), .B(n29129), .X(n29127) );
  nand_x4_sg U65852 ( .A(n29132), .B(n46235), .X(n29131) );
  nor_x1_sg U65853 ( .A(n29133), .B(n29134), .X(n29132) );
  nand_x4_sg U65854 ( .A(n29409), .B(n46235), .X(n29408) );
  nor_x1_sg U65855 ( .A(n29410), .B(n29411), .X(n29409) );
  nand_x4_sg U65856 ( .A(n29414), .B(n46235), .X(n29413) );
  nor_x1_sg U65857 ( .A(n29415), .B(n29416), .X(n29414) );
  nand_x2_sg U65858 ( .A(n46232), .B(n25485), .X(n25494) );
  nand_x2_sg U65859 ( .A(n46230), .B(n25763), .X(n25772) );
  nand_x2_sg U65860 ( .A(n46228), .B(n26041), .X(n26051) );
  nand_x2_sg U65861 ( .A(n46226), .B(n26322), .X(n26332) );
  nand_x2_sg U65862 ( .A(n46224), .B(n26601), .X(n26611) );
  nand_x2_sg U65863 ( .A(n46222), .B(n26879), .X(n26888) );
  nand_x2_sg U65864 ( .A(n46220), .B(n27158), .X(n27168) );
  nand_x2_sg U65865 ( .A(n46218), .B(n27438), .X(n27447) );
  nand_x2_sg U65866 ( .A(n46216), .B(n27718), .X(n27728) );
  nand_x2_sg U65867 ( .A(n46214), .B(n27998), .X(n28007) );
  nand_x2_sg U65868 ( .A(n46212), .B(n28278), .X(n28287) );
  nand_x2_sg U65869 ( .A(n46210), .B(n28556), .X(n28565) );
  nand_x2_sg U65870 ( .A(n46208), .B(n28836), .X(n28845) );
  nand_x2_sg U65871 ( .A(n46206), .B(n29115), .X(n29124) );
  nand_x1_sg U65872 ( .A(n46598), .B(n50872), .X(n9451) );
  nand_x1_sg U65873 ( .A(n46598), .B(n50828), .X(n9500) );
  nand_x1_sg U65874 ( .A(n46598), .B(n50784), .X(n9549) );
  nand_x1_sg U65875 ( .A(n46598), .B(n50738), .X(n9597) );
  nand_x1_sg U65876 ( .A(n46598), .B(n50692), .X(n9645) );
  nand_x1_sg U65877 ( .A(n46598), .B(n50601), .X(n9740) );
  nand_x1_sg U65878 ( .A(n46598), .B(n50555), .X(n9788) );
  nand_x1_sg U65879 ( .A(n50013), .B(n46598), .X(n24559) );
  nand_x1_sg U65880 ( .A(n49969), .B(n46598), .X(n24608) );
  nand_x1_sg U65881 ( .A(n49925), .B(n46598), .X(n24657) );
  nand_x1_sg U65882 ( .A(n49879), .B(n46598), .X(n24705) );
  nand_x1_sg U65883 ( .A(n49833), .B(n46598), .X(n24753) );
  nand_x1_sg U65884 ( .A(n49742), .B(n46598), .X(n24848) );
  nand_x1_sg U65885 ( .A(n49696), .B(n46598), .X(n24896) );
  nand_x4_sg U65886 ( .A(n11567), .B(n11568), .X(n11565) );
  nand_x1_sg U65887 ( .A(n11575), .B(n11573), .X(n11567) );
  nor_x1_sg U65888 ( .A(n51616), .B(n46543), .X(n11569) );
  nand_x4_sg U65889 ( .A(n13128), .B(n13129), .X(n13126) );
  nand_x1_sg U65890 ( .A(n13136), .B(n13134), .X(n13128) );
  nor_x1_sg U65891 ( .A(n52174), .B(n46499), .X(n13130) );
  nand_x4_sg U65892 ( .A(n15461), .B(n15462), .X(n15459) );
  nand_x1_sg U65893 ( .A(n15469), .B(n15467), .X(n15461) );
  nor_x1_sg U65894 ( .A(n53008), .B(n46431), .X(n15463) );
  nand_x4_sg U65895 ( .A(n17027), .B(n17028), .X(n17025) );
  nand_x1_sg U65896 ( .A(n17035), .B(n17033), .X(n17027) );
  nor_x1_sg U65897 ( .A(n53566), .B(n46387), .X(n17029) );
  nand_x4_sg U65898 ( .A(n26614), .B(n46235), .X(n26613) );
  nor_x1_sg U65899 ( .A(n26615), .B(n26616), .X(n26614) );
  nand_x4_sg U65900 ( .A(n26619), .B(n46235), .X(n26618) );
  nor_x1_sg U65901 ( .A(n26620), .B(n26621), .X(n26619) );
  nand_x4_sg U65902 ( .A(n26896), .B(n46235), .X(n26895) );
  nor_x1_sg U65903 ( .A(n26897), .B(n26898), .X(n26896) );
  nand_x4_sg U65904 ( .A(n14408), .B(n52714), .X(n14373) );
  nand_x1_sg U65905 ( .A(n14403), .B(n52690), .X(n14408) );
  nor_x1_sg U65906 ( .A(n52690), .B(n14403), .X(n14409) );
  nand_x4_sg U65907 ( .A(n17828), .B(n17866), .X(n17864) );
  nand_x4_sg U65908 ( .A(n19373), .B(n19411), .X(n19409) );
  nand_x4_sg U65909 ( .A(n20917), .B(n20955), .X(n20953) );
  nor_x1_sg U65910 ( .A(n46561), .B(n25428), .X(n25437) );
  nor_x1_sg U65911 ( .A(n46533), .B(n25707), .X(n25716) );
  nor_x1_sg U65912 ( .A(n46514), .B(n25985), .X(n25994) );
  nor_x1_sg U65913 ( .A(n46489), .B(n26266), .X(n26275) );
  nor_x1_sg U65914 ( .A(n46469), .B(n26545), .X(n26554) );
  nor_x1_sg U65915 ( .A(n46445), .B(n26823), .X(n26832) );
  nor_x1_sg U65916 ( .A(n46421), .B(n27102), .X(n27111) );
  nor_x1_sg U65917 ( .A(n46402), .B(n27382), .X(n27391) );
  nor_x1_sg U65918 ( .A(n46377), .B(n27662), .X(n27671) );
  nor_x1_sg U65919 ( .A(n53814), .B(n27942), .X(n27951) );
  nor_x1_sg U65920 ( .A(n54097), .B(n28221), .X(n28230) );
  nor_x1_sg U65921 ( .A(n54379), .B(n28500), .X(n28509) );
  nor_x1_sg U65922 ( .A(n46289), .B(n28779), .X(n28788) );
  nor_x1_sg U65923 ( .A(n54947), .B(n29059), .X(n29068) );
  nor_x1_sg U65924 ( .A(n46244), .B(n29340), .X(n29349) );
  nand_x4_sg U65925 ( .A(n13729), .B(n13730), .X(n13665) );
  nand_x1_sg U65926 ( .A(n13732), .B(n13733), .X(n13729) );
  nand_x4_sg U65927 ( .A(n12348), .B(n12349), .X(n12346) );
  nand_x1_sg U65928 ( .A(n12356), .B(n12354), .X(n12348) );
  nor_x1_sg U65929 ( .A(n12214), .B(n46518), .X(n12356) );
  nand_x4_sg U65930 ( .A(n13908), .B(n13909), .X(n13906) );
  nand_x1_sg U65931 ( .A(n13916), .B(n13914), .X(n13908) );
  nor_x1_sg U65932 ( .A(n46475), .B(n13775), .X(n13916) );
  nor_x1_sg U65933 ( .A(n24524), .B(n24473), .X(\L1_0/n4819 ) );
  nor_x1_sg U65934 ( .A(n24573), .B(n46234), .X(\L1_0/n4815 ) );
  nor_x1_sg U65935 ( .A(n24671), .B(n24473), .X(\L1_0/n4807 ) );
  nor_x1_sg U65936 ( .A(n24719), .B(n46234), .X(\L1_0/n4803 ) );
  nor_x1_sg U65937 ( .A(n24814), .B(n24473), .X(\L1_0/n4795 ) );
  nor_x1_sg U65938 ( .A(n24862), .B(n46234), .X(\L1_0/n4791 ) );
  nor_x1_sg U65939 ( .A(n24958), .B(n24473), .X(\L1_0/n4783 ) );
  nor_x1_sg U65940 ( .A(n25006), .B(n46234), .X(\L1_0/n4779 ) );
  nor_x1_sg U65941 ( .A(n25103), .B(n24473), .X(\L1_0/n4771 ) );
  nor_x1_sg U65942 ( .A(n25151), .B(n46234), .X(\L1_0/n4767 ) );
  nor_x1_sg U65943 ( .A(n25249), .B(n24473), .X(\L1_0/n4759 ) );
  nor_x1_sg U65944 ( .A(n25296), .B(n46234), .X(\L1_0/n4755 ) );
  nand_x4_sg U65945 ( .A(n14351), .B(n14352), .X(n14349) );
  nand_x1_sg U65946 ( .A(n14354), .B(n14355), .X(n14351) );
  nand_x4_sg U65947 ( .A(n18241), .B(n18242), .X(n18235) );
  nand_x1_sg U65948 ( .A(n18244), .B(n18245), .X(n18241) );
  nand_x4_sg U65949 ( .A(n19786), .B(n19787), .X(n19781) );
  nand_x1_sg U65950 ( .A(n19789), .B(n19790), .X(n19786) );
  nand_x4_sg U65951 ( .A(n21331), .B(n21332), .X(n21326) );
  nand_x1_sg U65952 ( .A(n21334), .B(n21335), .X(n21331) );
  nand_x4_sg U65953 ( .A(n10947), .B(n10948), .X(n10932) );
  nand_x1_sg U65954 ( .A(n43798), .B(n10950), .X(n10948) );
  nand_x1_sg U65955 ( .A(n10952), .B(n10951), .X(n10947) );
  nand_x1_sg U65956 ( .A(n10951), .B(n10282), .X(n10950) );
  nand_x4_sg U65957 ( .A(n16405), .B(n16406), .X(n16390) );
  nand_x1_sg U65958 ( .A(n43051), .B(n16408), .X(n16406) );
  nand_x1_sg U65959 ( .A(n16410), .B(n16409), .X(n16405) );
  nand_x1_sg U65960 ( .A(n16409), .B(n46413), .X(n16408) );
  nand_x4_sg U65961 ( .A(n25490), .B(n25491), .X(n25489) );
  nor_x1_sg U65962 ( .A(n42489), .B(n25493), .X(n25491) );
  nor_x1_sg U65963 ( .A(n25495), .B(n46236), .X(n25490) );
  nand_x4_sg U65964 ( .A(n19615), .B(n19616), .X(n9181) );
  nand_x4_sg U65965 ( .A(n21160), .B(n21161), .X(n9101) );
  nand_x4_sg U65966 ( .A(n17802), .B(n17803), .X(n17714) );
  nand_x1_sg U65967 ( .A(n17805), .B(n17806), .X(n17802) );
  nor_x1_sg U65968 ( .A(n17805), .B(n46362), .X(n17804) );
  nand_x4_sg U65969 ( .A(n19347), .B(n19348), .X(n19259) );
  nand_x1_sg U65970 ( .A(n19350), .B(n19351), .X(n19347) );
  nor_x1_sg U65971 ( .A(n19350), .B(n46315), .X(n19349) );
  nand_x4_sg U65972 ( .A(n20891), .B(n20892), .X(n20803) );
  nand_x1_sg U65973 ( .A(n20894), .B(n20895), .X(n20891) );
  nor_x1_sg U65974 ( .A(n20894), .B(n46270), .X(n20893) );
  nor_x1_sg U65975 ( .A(n46480), .B(n46471), .X(n13594) );
  nand_x4_sg U65976 ( .A(n16351), .B(n16352), .X(n16350) );
  nand_x1_sg U65977 ( .A(n16353), .B(n53424), .X(n16352) );
  nand_x1_sg U65978 ( .A(n16355), .B(n53340), .X(n16351) );
  nor_x1_sg U65979 ( .A(n16354), .B(n53446), .X(n16353) );
  nand_x4_sg U65980 ( .A(n51880), .B(n12075), .X(n12034) );
  nand_x1_sg U65981 ( .A(n12069), .B(n12076), .X(n12075) );
  nor_x1_sg U65982 ( .A(n12076), .B(n12069), .X(n12077) );
  nand_x4_sg U65983 ( .A(n53267), .B(n15970), .X(n15929) );
  nand_x1_sg U65984 ( .A(n15964), .B(n15971), .X(n15970) );
  nor_x1_sg U65985 ( .A(n15971), .B(n15964), .X(n15972) );
  nand_x4_sg U65986 ( .A(n12551), .B(n12552), .X(n12540) );
  nand_x1_sg U65987 ( .A(n12555), .B(n51945), .X(n12551) );
  nand_x1_sg U65988 ( .A(n12553), .B(n12554), .X(n12552) );
  nand_x4_sg U65989 ( .A(n51599), .B(n11295), .X(n11257) );
  nand_x1_sg U65990 ( .A(n11289), .B(n11296), .X(n11295) );
  nor_x1_sg U65991 ( .A(n11296), .B(n11289), .X(n11297) );
  nand_x4_sg U65992 ( .A(n25390), .B(n25391), .X(n25389) );
  nor_x1_sg U65993 ( .A(n51256), .B(n25392), .X(n25391) );
  nor_x1_sg U65994 ( .A(n25393), .B(n46236), .X(n25390) );
  nand_x4_sg U65995 ( .A(n25670), .B(n25671), .X(n25669) );
  nor_x1_sg U65996 ( .A(n51532), .B(n25672), .X(n25671) );
  nor_x1_sg U65997 ( .A(n25673), .B(n46236), .X(n25670) );
  nand_x4_sg U65998 ( .A(n25948), .B(n25949), .X(n25947) );
  nor_x1_sg U65999 ( .A(n51814), .B(n25950), .X(n25949) );
  nor_x1_sg U66000 ( .A(n25951), .B(n46236), .X(n25948) );
  nand_x4_sg U66001 ( .A(n26229), .B(n26230), .X(n26228) );
  nor_x1_sg U66002 ( .A(n52090), .B(n26231), .X(n26230) );
  nor_x1_sg U66003 ( .A(n26232), .B(n46236), .X(n26229) );
  nand_x4_sg U66004 ( .A(n26786), .B(n26787), .X(n26785) );
  nor_x1_sg U66005 ( .A(n52643), .B(n26788), .X(n26787) );
  nor_x1_sg U66006 ( .A(n26789), .B(n46236), .X(n26786) );
  nand_x4_sg U66007 ( .A(n27065), .B(n27066), .X(n27064) );
  nor_x1_sg U66008 ( .A(n52924), .B(n27067), .X(n27066) );
  nor_x1_sg U66009 ( .A(n27068), .B(n46236), .X(n27065) );
  nand_x4_sg U66010 ( .A(n27345), .B(n27346), .X(n27344) );
  nor_x1_sg U66011 ( .A(n53202), .B(n27347), .X(n27346) );
  nor_x1_sg U66012 ( .A(n27348), .B(n46236), .X(n27345) );
  nand_x4_sg U66013 ( .A(n27625), .B(n27626), .X(n27624) );
  nor_x1_sg U66014 ( .A(n53482), .B(n27627), .X(n27626) );
  nor_x1_sg U66015 ( .A(n27628), .B(n46236), .X(n27625) );
  nand_x4_sg U66016 ( .A(n27905), .B(n27906), .X(n27904) );
  nor_x1_sg U66017 ( .A(n53760), .B(n27907), .X(n27906) );
  nor_x1_sg U66018 ( .A(n27908), .B(n46236), .X(n27905) );
  nand_x4_sg U66019 ( .A(n28184), .B(n28185), .X(n28183) );
  nor_x1_sg U66020 ( .A(n54044), .B(n28186), .X(n28185) );
  nor_x1_sg U66021 ( .A(n28187), .B(n46236), .X(n28184) );
  nand_x4_sg U66022 ( .A(n28463), .B(n28464), .X(n28462) );
  nor_x1_sg U66023 ( .A(n54325), .B(n28465), .X(n28464) );
  nor_x1_sg U66024 ( .A(n28466), .B(n46236), .X(n28463) );
  nand_x4_sg U66025 ( .A(n12949), .B(n12950), .X(n12885) );
  nand_x1_sg U66026 ( .A(n12952), .B(n12953), .X(n12949) );
  nor_x1_sg U66027 ( .A(n46508), .B(n12952), .X(n12951) );
  nand_x4_sg U66028 ( .A(n15282), .B(n15283), .X(n15218) );
  nand_x1_sg U66029 ( .A(n15285), .B(n15286), .X(n15282) );
  nor_x1_sg U66030 ( .A(n46440), .B(n15285), .X(n15284) );
  nand_x4_sg U66031 ( .A(n16848), .B(n16849), .X(n16784) );
  nand_x1_sg U66032 ( .A(n16851), .B(n16852), .X(n16848) );
  nor_x1_sg U66033 ( .A(n46396), .B(n16851), .X(n16850) );
  nand_x4_sg U66034 ( .A(n28742), .B(n28743), .X(n28741) );
  nor_x1_sg U66035 ( .A(n54609), .B(n28744), .X(n28743) );
  nor_x1_sg U66036 ( .A(n28745), .B(n46236), .X(n28742) );
  nand_x4_sg U66037 ( .A(n29022), .B(n29023), .X(n29021) );
  nor_x1_sg U66038 ( .A(n54893), .B(n29024), .X(n29023) );
  nor_x1_sg U66039 ( .A(n29025), .B(n46236), .X(n29022) );
  nand_x4_sg U66040 ( .A(n29303), .B(n29304), .X(n29302) );
  nor_x1_sg U66041 ( .A(n55177), .B(n29305), .X(n29304) );
  nor_x1_sg U66042 ( .A(n29306), .B(n46236), .X(n29303) );
  nand_x4_sg U66043 ( .A(n14112), .B(n14113), .X(n14101) );
  nand_x1_sg U66044 ( .A(n14116), .B(n52497), .X(n14112) );
  nand_x1_sg U66045 ( .A(n14114), .B(n14115), .X(n14113) );
  nand_x4_sg U66046 ( .A(n52157), .B(n12856), .X(n12818) );
  nand_x1_sg U66047 ( .A(n12850), .B(n12857), .X(n12856) );
  nor_x1_sg U66048 ( .A(n12857), .B(n12850), .X(n12858) );
  nand_x4_sg U66049 ( .A(n52991), .B(n15189), .X(n15151) );
  nand_x1_sg U66050 ( .A(n15183), .B(n15190), .X(n15189) );
  nor_x1_sg U66051 ( .A(n15190), .B(n15183), .X(n15191) );
  nand_x4_sg U66052 ( .A(n53549), .B(n16755), .X(n16717) );
  nand_x1_sg U66053 ( .A(n16749), .B(n16756), .X(n16755) );
  nor_x1_sg U66054 ( .A(n16756), .B(n16749), .X(n16757) );
  nand_x4_sg U66055 ( .A(n11388), .B(n11389), .X(n11324) );
  nand_x1_sg U66056 ( .A(n11391), .B(n11392), .X(n11388) );
  nor_x1_sg U66057 ( .A(n46552), .B(n11391), .X(n11390) );
  nand_x2_sg U66058 ( .A(n41521), .B(n28201), .X(n28200) );
  nand_x4_sg U66059 ( .A(n10786), .B(n10787), .X(n10784) );
  nand_x1_sg U66060 ( .A(n10794), .B(n10792), .X(n10786) );
  nor_x1_sg U66061 ( .A(n41277), .B(n46568), .X(n10788) );
  nand_x4_sg U66062 ( .A(n20112), .B(n20113), .X(n20110) );
  nand_x1_sg U66063 ( .A(n20120), .B(n20118), .X(n20112) );
  nor_x1_sg U66064 ( .A(n41574), .B(n46297), .X(n20114) );
  nand_x4_sg U66065 ( .A(n21657), .B(n21658), .X(n21655) );
  nand_x1_sg U66066 ( .A(n21665), .B(n21663), .X(n21657) );
  nor_x1_sg U66067 ( .A(n41572), .B(n46252), .X(n21659) );
  nand_x4_sg U66068 ( .A(n11259), .B(n11260), .X(n11248) );
  nor_x1_sg U66069 ( .A(n11261), .B(n46546), .X(n11260) );
  nor_x1_sg U66070 ( .A(n11267), .B(n11238), .X(n11259) );
  nand_x4_sg U66071 ( .A(n11570), .B(n11571), .X(n11482) );
  nand_x1_sg U66072 ( .A(n11573), .B(n11574), .X(n11570) );
  nor_x1_sg U66073 ( .A(n11573), .B(n46541), .X(n11572) );
  nand_x4_sg U66074 ( .A(n13131), .B(n13132), .X(n13043) );
  nand_x1_sg U66075 ( .A(n13134), .B(n13135), .X(n13131) );
  nor_x1_sg U66076 ( .A(n13134), .B(n46497), .X(n13133) );
  nand_x4_sg U66077 ( .A(n15464), .B(n15465), .X(n15376) );
  nand_x1_sg U66078 ( .A(n15467), .B(n15468), .X(n15464) );
  nor_x1_sg U66079 ( .A(n15467), .B(n46429), .X(n15466) );
  nand_x4_sg U66080 ( .A(n17030), .B(n17031), .X(n16942) );
  nand_x1_sg U66081 ( .A(n17033), .B(n17034), .X(n17030) );
  nor_x1_sg U66082 ( .A(n17033), .B(n46385), .X(n17032) );
  nand_x4_sg U66083 ( .A(n12604), .B(n12605), .X(n12440) );
  nand_x1_sg U66084 ( .A(n12214), .B(n12606), .X(n12604) );
  nand_x4_sg U66085 ( .A(n17981), .B(n17982), .X(n17979) );
  nand_x1_sg U66086 ( .A(n53999), .B(n17984), .X(n17981) );
  nand_x1_sg U66087 ( .A(n53827), .B(n53862), .X(n17984) );
  nand_x4_sg U66088 ( .A(n19526), .B(n19527), .X(n19524) );
  nand_x1_sg U66089 ( .A(n54564), .B(n19529), .X(n19526) );
  nand_x1_sg U66090 ( .A(n54392), .B(n54427), .X(n19529) );
  nand_x4_sg U66091 ( .A(n21070), .B(n21071), .X(n21068) );
  nand_x1_sg U66092 ( .A(n55132), .B(n21073), .X(n21070) );
  nand_x1_sg U66093 ( .A(n54960), .B(n54995), .X(n21073) );
  nand_x4_sg U66094 ( .A(n11411), .B(n11465), .X(n11463) );
  nand_x1_sg U66095 ( .A(n51696), .B(n11466), .X(n11465) );
  nand_x4_sg U66096 ( .A(n12972), .B(n13026), .X(n13024) );
  nand_x1_sg U66097 ( .A(n52252), .B(n13027), .X(n13026) );
  nand_x4_sg U66098 ( .A(n15305), .B(n15359), .X(n15357) );
  nand_x1_sg U66099 ( .A(n53086), .B(n15360), .X(n15359) );
  nand_x4_sg U66100 ( .A(n16871), .B(n16925), .X(n16923) );
  nand_x1_sg U66101 ( .A(n53644), .B(n16926), .X(n16925) );
  nand_x4_sg U66102 ( .A(n12102), .B(n51912), .X(n12094) );
  nor_x1_sg U66103 ( .A(n12104), .B(n12105), .X(n12103) );
  nand_x4_sg U66104 ( .A(n15997), .B(n53299), .X(n15989) );
  nor_x1_sg U66105 ( .A(n15999), .B(n16000), .X(n15998) );
  nand_x4_sg U66106 ( .A(n11990), .B(n11991), .X(n11979) );
  nand_x1_sg U66107 ( .A(n51849), .B(n11986), .X(n11990) );
  nand_x1_sg U66108 ( .A(n11985), .B(n51855), .X(n11991) );
  nand_x4_sg U66109 ( .A(n15885), .B(n15886), .X(n15874) );
  nand_x1_sg U66110 ( .A(n53235), .B(n15881), .X(n15885) );
  nand_x1_sg U66111 ( .A(n15880), .B(n53241), .X(n15886) );
  nand_x4_sg U66112 ( .A(n51367), .B(n10581), .X(n10566) );
  nand_x1_sg U66113 ( .A(n51366), .B(n10582), .X(n10581) );
  nor_x1_sg U66114 ( .A(n10582), .B(n51366), .X(n10583) );
  nand_x4_sg U66115 ( .A(n10577), .B(n10578), .X(n10570) );
  nand_x1_sg U66116 ( .A(n10580), .B(n51346), .X(n10577) );
  nand_x1_sg U66117 ( .A(n10579), .B(n51301), .X(n10578) );
  nand_x4_sg U66118 ( .A(n10438), .B(n10439), .X(n10427) );
  nand_x1_sg U66119 ( .A(n51289), .B(n10434), .X(n10438) );
  nand_x1_sg U66120 ( .A(n10433), .B(n51294), .X(n10439) );
  nand_x4_sg U66121 ( .A(n14330), .B(n14331), .X(n14319) );
  nand_x1_sg U66122 ( .A(n52679), .B(n14326), .X(n14330) );
  nand_x1_sg U66123 ( .A(n14325), .B(n52684), .X(n14331) );
  nand_x4_sg U66124 ( .A(n19765), .B(n19766), .X(n19754) );
  nand_x1_sg U66125 ( .A(n54643), .B(n19761), .X(n19765) );
  nand_x1_sg U66126 ( .A(n19760), .B(n54648), .X(n19766) );
  nand_x4_sg U66127 ( .A(n21310), .B(n21311), .X(n21299) );
  nand_x1_sg U66128 ( .A(n55211), .B(n21306), .X(n21310) );
  nand_x1_sg U66129 ( .A(n21305), .B(n55216), .X(n21311) );
  nand_x4_sg U66130 ( .A(n18302), .B(n18303), .X(n18286) );
  nand_x1_sg U66131 ( .A(n54092), .B(n54130), .X(n18303) );
  nand_x4_sg U66132 ( .A(n17453), .B(n17454), .X(n17442) );
  nand_x1_sg U66133 ( .A(n53798), .B(n17449), .X(n17453) );
  nand_x1_sg U66134 ( .A(n17448), .B(n53803), .X(n17454) );
  nand_x4_sg U66135 ( .A(n18219), .B(n18220), .X(n18208) );
  nand_x1_sg U66136 ( .A(n54079), .B(n18215), .X(n18219) );
  nand_x1_sg U66137 ( .A(n18214), .B(n54085), .X(n18220) );
  nand_x4_sg U66138 ( .A(n18998), .B(n18999), .X(n18987) );
  nand_x1_sg U66139 ( .A(n54363), .B(n18994), .X(n18998) );
  nand_x1_sg U66140 ( .A(n18993), .B(n54368), .X(n18999) );
  nand_x4_sg U66141 ( .A(n20542), .B(n20543), .X(n20531) );
  nand_x1_sg U66142 ( .A(n54931), .B(n20538), .X(n20542) );
  nand_x1_sg U66143 ( .A(n20537), .B(n54936), .X(n20543) );
  nand_x4_sg U66144 ( .A(n17589), .B(n17590), .X(n17582) );
  nand_x1_sg U66145 ( .A(n17592), .B(n53856), .X(n17589) );
  nand_x1_sg U66146 ( .A(n17591), .B(n53810), .X(n17590) );
  nand_x4_sg U66147 ( .A(n19134), .B(n19135), .X(n19127) );
  nand_x1_sg U66148 ( .A(n19137), .B(n54421), .X(n19134) );
  nand_x1_sg U66149 ( .A(n19136), .B(n54375), .X(n19135) );
  nand_x4_sg U66150 ( .A(n20678), .B(n20679), .X(n20671) );
  nand_x1_sg U66151 ( .A(n20681), .B(n54989), .X(n20678) );
  nand_x1_sg U66152 ( .A(n20680), .B(n54943), .X(n20679) );
  nor_x1_sg U66153 ( .A(n46615), .B(n29578), .X(n29581) );
  nor_x1_sg U66154 ( .A(n46615), .B(n24474), .X(n24478) );
  nor_x1_sg U66155 ( .A(n46615), .B(n24623), .X(n24626) );
  nor_x1_sg U66156 ( .A(n46615), .B(n24768), .X(n24771) );
  nor_x1_sg U66157 ( .A(n46615), .B(n24911), .X(n24914) );
  nor_x1_sg U66158 ( .A(n46615), .B(n25055), .X(n25058) );
  nor_x1_sg U66159 ( .A(n46615), .B(n25201), .X(n25204) );
  nand_x4_sg U66160 ( .A(n14681), .B(n14682), .X(n14593) );
  nand_x1_sg U66161 ( .A(n14684), .B(n14685), .X(n14681) );
  nor_x1_sg U66162 ( .A(n14684), .B(n46451), .X(n14683) );
  nand_x4_sg U66163 ( .A(n12590), .B(n12591), .X(n12409) );
  nand_x1_sg U66164 ( .A(n52025), .B(n12587), .X(n12591) );
  nand_x1_sg U66165 ( .A(n51890), .B(n12586), .X(n12590) );
  nand_x4_sg U66166 ( .A(n12820), .B(n12821), .X(n12809) );
  nor_x1_sg U66167 ( .A(n12828), .B(n12799), .X(n12820) );
  nor_x1_sg U66168 ( .A(n12822), .B(n46502), .X(n12821) );
  nand_x4_sg U66169 ( .A(n15153), .B(n15154), .X(n15142) );
  nor_x1_sg U66170 ( .A(n15161), .B(n15132), .X(n15153) );
  nor_x1_sg U66171 ( .A(n15155), .B(n46434), .X(n15154) );
  nand_x4_sg U66172 ( .A(n16719), .B(n16720), .X(n16708) );
  nor_x1_sg U66173 ( .A(n16727), .B(n16698), .X(n16719) );
  nor_x1_sg U66174 ( .A(n16721), .B(n46390), .X(n16720) );
  nand_x4_sg U66175 ( .A(n51919), .B(n12135), .X(n12116) );
  nand_x1_sg U66176 ( .A(n51918), .B(n12136), .X(n12135) );
  nor_x1_sg U66177 ( .A(n12136), .B(n51918), .X(n12137) );
  nand_x4_sg U66178 ( .A(n53306), .B(n16030), .X(n16011) );
  nand_x1_sg U66179 ( .A(n53305), .B(n16031), .X(n16030) );
  nor_x1_sg U66180 ( .A(n16031), .B(n53305), .X(n16032) );
  nand_x4_sg U66181 ( .A(n10789), .B(n10790), .X(n10701) );
  nand_x1_sg U66182 ( .A(n10792), .B(n10793), .X(n10789) );
  nor_x1_sg U66183 ( .A(n10792), .B(n10655), .X(n10791) );
  nand_x4_sg U66184 ( .A(n20115), .B(n20116), .X(n20028) );
  nand_x1_sg U66185 ( .A(n20118), .B(n20119), .X(n20115) );
  nor_x1_sg U66186 ( .A(n20118), .B(n19982), .X(n20117) );
  nand_x4_sg U66187 ( .A(n21660), .B(n21661), .X(n21573) );
  nand_x1_sg U66188 ( .A(n21663), .B(n21664), .X(n21660) );
  nor_x1_sg U66189 ( .A(n21663), .B(n21527), .X(n21662) );
  nand_x4_sg U66190 ( .A(n12351), .B(n12352), .X(n12262) );
  nand_x1_sg U66191 ( .A(n12354), .B(n12355), .X(n12351) );
  nor_x1_sg U66192 ( .A(n12354), .B(n12214), .X(n12353) );
  nand_x4_sg U66193 ( .A(n16246), .B(n16247), .X(n16157) );
  nand_x1_sg U66194 ( .A(n16249), .B(n16250), .X(n16246) );
  nor_x1_sg U66195 ( .A(n16249), .B(n16109), .X(n16248) );
  nand_x4_sg U66196 ( .A(n12603), .B(n52016), .X(n26050) );
  nand_x4_sg U66197 ( .A(n13385), .B(n52292), .X(n26331) );
  nand_x4_sg U66198 ( .A(n14165), .B(n52567), .X(n26610) );
  nand_x4_sg U66199 ( .A(n15718), .B(n53126), .X(n27167) );
  nand_x4_sg U66200 ( .A(n17284), .B(n53684), .X(n27727) );
  nand_x4_sg U66201 ( .A(n10920), .B(n10921), .X(n10913) );
  nand_x1_sg U66202 ( .A(n10744), .B(n10924), .X(n10920) );
  nor_x1_sg U66203 ( .A(n10744), .B(n10923), .X(n10922) );
  nand_x4_sg U66204 ( .A(n51466), .B(n10839), .X(n10827) );
  nand_x4_sg U66205 ( .A(n14707), .B(n14745), .X(n14743) );
  nand_x4_sg U66206 ( .A(n51382), .B(n11035), .X(n11000) );
  nand_x1_sg U66207 ( .A(n10998), .B(n11036), .X(n11035) );
  nor_x1_sg U66208 ( .A(n11036), .B(n10998), .X(n11037) );
  nand_x4_sg U66209 ( .A(n10995), .B(n10996), .X(n10976) );
  nand_x1_sg U66210 ( .A(n10999), .B(n11000), .X(n10995) );
  nand_x1_sg U66211 ( .A(n10997), .B(n10998), .X(n10996) );
  nor_x1_sg U66212 ( .A(n10660), .B(n46563), .X(n10997) );
  nand_x4_sg U66213 ( .A(n18782), .B(n18783), .X(n18762) );
  nand_x1_sg U66214 ( .A(n18786), .B(n18787), .X(n18782) );
  nand_x1_sg U66215 ( .A(n18784), .B(n18785), .X(n18783) );
  nor_x1_sg U66216 ( .A(n46337), .B(n18442), .X(n18784) );
  nand_x4_sg U66217 ( .A(n20328), .B(n20329), .X(n20308) );
  nand_x1_sg U66218 ( .A(n20332), .B(n20333), .X(n20328) );
  nand_x1_sg U66219 ( .A(n20330), .B(n20331), .X(n20329) );
  nor_x1_sg U66220 ( .A(n46293), .B(n19987), .X(n20330) );
  nand_x4_sg U66221 ( .A(n21873), .B(n21874), .X(n21853) );
  nand_x1_sg U66222 ( .A(n21877), .B(n21878), .X(n21873) );
  nand_x1_sg U66223 ( .A(n21875), .B(n21876), .X(n21874) );
  nor_x1_sg U66224 ( .A(n46248), .B(n21532), .X(n21875) );
  nand_x4_sg U66225 ( .A(n10751), .B(n51436), .X(n10747) );
  nand_x1_sg U66226 ( .A(n10754), .B(n10753), .X(n10751) );
  nor_x1_sg U66227 ( .A(n10753), .B(n10754), .X(n10752) );
  nand_x4_sg U66228 ( .A(n18532), .B(n54230), .X(n18528) );
  nand_x1_sg U66229 ( .A(n18535), .B(n18534), .X(n18532) );
  nor_x1_sg U66230 ( .A(n18534), .B(n18535), .X(n18533) );
  nand_x4_sg U66231 ( .A(n20363), .B(n20364), .X(n20174) );
  nand_x1_sg U66232 ( .A(n54677), .B(n20359), .X(n20363) );
  nand_x1_sg U66233 ( .A(n54823), .B(n20360), .X(n20364) );
  nand_x4_sg U66234 ( .A(n21908), .B(n21909), .X(n21719) );
  nand_x1_sg U66235 ( .A(n55245), .B(n21904), .X(n21908) );
  nand_x1_sg U66236 ( .A(n55391), .B(n21905), .X(n21909) );
  nand_x4_sg U66237 ( .A(n16454), .B(n16455), .X(n16434) );
  nand_x1_sg U66238 ( .A(n16458), .B(n53333), .X(n16454) );
  nand_x1_sg U66239 ( .A(n16456), .B(n16457), .X(n16455) );
  nand_x4_sg U66240 ( .A(n53864), .B(n17593), .X(n17578) );
  nand_x1_sg U66241 ( .A(n53863), .B(n17594), .X(n17593) );
  nor_x1_sg U66242 ( .A(n17594), .B(n53863), .X(n17595) );
  nand_x4_sg U66243 ( .A(n54429), .B(n19138), .X(n19123) );
  nand_x1_sg U66244 ( .A(n54428), .B(n19139), .X(n19138) );
  nor_x1_sg U66245 ( .A(n19139), .B(n54428), .X(n19140) );
  nand_x4_sg U66246 ( .A(n54997), .B(n20682), .X(n20667) );
  nand_x1_sg U66247 ( .A(n54996), .B(n20683), .X(n20682) );
  nor_x1_sg U66248 ( .A(n20683), .B(n54996), .X(n20684) );
  nand_x4_sg U66249 ( .A(n19719), .B(n19720), .X(n19622) );
  nand_x1_sg U66250 ( .A(n19722), .B(n19723), .X(n19719) );
  nand_x4_sg U66251 ( .A(n21264), .B(n21265), .X(n21167) );
  nand_x1_sg U66252 ( .A(n21267), .B(n21268), .X(n21264) );
  nand_x4_sg U66253 ( .A(n11316), .B(n11317), .X(n11285) );
  nand_x1_sg U66254 ( .A(n11319), .B(n11320), .X(n11316) );
  nand_x4_sg U66255 ( .A(n12096), .B(n12097), .X(n12065) );
  nand_x1_sg U66256 ( .A(n12099), .B(n12100), .X(n12096) );
  nand_x4_sg U66257 ( .A(n12877), .B(n12878), .X(n12846) );
  nand_x1_sg U66258 ( .A(n12880), .B(n12881), .X(n12877) );
  nand_x4_sg U66259 ( .A(n15210), .B(n15211), .X(n15179) );
  nand_x1_sg U66260 ( .A(n15213), .B(n15214), .X(n15210) );
  nand_x4_sg U66261 ( .A(n15991), .B(n15992), .X(n15960) );
  nand_x1_sg U66262 ( .A(n15994), .B(n15995), .X(n15991) );
  nand_x4_sg U66263 ( .A(n16776), .B(n16777), .X(n16745) );
  nand_x1_sg U66264 ( .A(n16779), .B(n16780), .X(n16776) );
  nand_x4_sg U66265 ( .A(n9374), .B(n9375), .X(n9356) );
  nor_x1_sg U66266 ( .A(n9376), .B(n9377), .X(n9375) );
  nor_x1_sg U66267 ( .A(n9395), .B(n9396), .X(n9374) );
  nand_x2_sg U66268 ( .A(n9386), .B(n9387), .X(n9376) );
  nand_x4_sg U66269 ( .A(n9674), .B(n9675), .X(n9660) );
  nor_x1_sg U66270 ( .A(n9676), .B(n9677), .X(n9675) );
  nor_x1_sg U66271 ( .A(n9690), .B(n9691), .X(n9674) );
  nand_x2_sg U66272 ( .A(n9684), .B(n9685), .X(n9676) );
  nand_x4_sg U66273 ( .A(n24489), .B(n24490), .X(n24474) );
  nor_x1_sg U66274 ( .A(n24491), .B(n24492), .X(n24490) );
  nor_x1_sg U66275 ( .A(n24507), .B(n24508), .X(n24489) );
  nand_x2_sg U66276 ( .A(n24500), .B(n24501), .X(n24491) );
  nand_x4_sg U66277 ( .A(n24782), .B(n24783), .X(n24768) );
  nor_x1_sg U66278 ( .A(n24784), .B(n24785), .X(n24783) );
  nor_x1_sg U66279 ( .A(n24798), .B(n24799), .X(n24782) );
  nand_x2_sg U66280 ( .A(n24792), .B(n24793), .X(n24784) );
  nand_x4_sg U66281 ( .A(n9431), .B(n9432), .X(n9417) );
  nor_x1_sg U66282 ( .A(n9448), .B(n9449), .X(n9431) );
  nor_x1_sg U66283 ( .A(n9433), .B(n9434), .X(n9432) );
  nand_x2_sg U66284 ( .A(n9450), .B(n9451), .X(n9449) );
  nand_x4_sg U66285 ( .A(n9480), .B(n9481), .X(n9466) );
  nor_x1_sg U66286 ( .A(n9497), .B(n9498), .X(n9480) );
  nor_x1_sg U66287 ( .A(n9482), .B(n9483), .X(n9481) );
  nand_x2_sg U66288 ( .A(n9499), .B(n9500), .X(n9498) );
  nand_x4_sg U66289 ( .A(n9529), .B(n9530), .X(n9515) );
  nor_x1_sg U66290 ( .A(n9546), .B(n9547), .X(n9529) );
  nor_x1_sg U66291 ( .A(n9531), .B(n9532), .X(n9530) );
  nand_x2_sg U66292 ( .A(n9548), .B(n9549), .X(n9547) );
  nand_x4_sg U66293 ( .A(n24539), .B(n24540), .X(n24525) );
  nor_x1_sg U66294 ( .A(n24556), .B(n24557), .X(n24539) );
  nor_x1_sg U66295 ( .A(n24541), .B(n24542), .X(n24540) );
  nand_x2_sg U66296 ( .A(n24558), .B(n24559), .X(n24557) );
  nand_x4_sg U66297 ( .A(n24588), .B(n24589), .X(n24574) );
  nor_x1_sg U66298 ( .A(n24605), .B(n24606), .X(n24588) );
  nor_x1_sg U66299 ( .A(n24590), .B(n24591), .X(n24589) );
  nand_x2_sg U66300 ( .A(n24607), .B(n24608), .X(n24606) );
  nand_x4_sg U66301 ( .A(n24637), .B(n24638), .X(n24623) );
  nor_x1_sg U66302 ( .A(n24654), .B(n24655), .X(n24637) );
  nor_x1_sg U66303 ( .A(n24639), .B(n24640), .X(n24638) );
  nand_x2_sg U66304 ( .A(n24656), .B(n24657), .X(n24655) );
  nand_x4_sg U66305 ( .A(n10058), .B(n10059), .X(n10044) );
  nor_x1_sg U66306 ( .A(n10060), .B(n10061), .X(n10059) );
  nor_x1_sg U66307 ( .A(n10074), .B(n10075), .X(n10058) );
  nand_x2_sg U66308 ( .A(n10068), .B(n10069), .X(n10060) );
  nand_x4_sg U66309 ( .A(n10107), .B(n10108), .X(n10093) );
  nor_x1_sg U66310 ( .A(n10109), .B(n10110), .X(n10108) );
  nor_x1_sg U66311 ( .A(n10123), .B(n10124), .X(n10107) );
  nand_x2_sg U66312 ( .A(n10117), .B(n10118), .X(n10109) );
  nand_x4_sg U66313 ( .A(n25166), .B(n25167), .X(n25152) );
  nor_x1_sg U66314 ( .A(n25168), .B(n25169), .X(n25167) );
  nor_x1_sg U66315 ( .A(n25182), .B(n25183), .X(n25166) );
  nand_x2_sg U66316 ( .A(n25176), .B(n25177), .X(n25168) );
  nand_x4_sg U66317 ( .A(n25215), .B(n25216), .X(n25201) );
  nor_x1_sg U66318 ( .A(n25217), .B(n25218), .X(n25216) );
  nor_x1_sg U66319 ( .A(n25231), .B(n25232), .X(n25215) );
  nand_x2_sg U66320 ( .A(n25225), .B(n25226), .X(n25217) );
  nand_x4_sg U66321 ( .A(n9961), .B(n9962), .X(n9947) );
  nor_x1_sg U66322 ( .A(n9963), .B(n9964), .X(n9962) );
  nor_x1_sg U66323 ( .A(n9977), .B(n9978), .X(n9961) );
  nand_x2_sg U66324 ( .A(n9971), .B(n9972), .X(n9963) );
  nand_x4_sg U66325 ( .A(n25069), .B(n25070), .X(n25055) );
  nor_x1_sg U66326 ( .A(n25071), .B(n25072), .X(n25070) );
  nor_x1_sg U66327 ( .A(n25085), .B(n25086), .X(n25069) );
  nand_x2_sg U66328 ( .A(n25079), .B(n25080), .X(n25071) );
  nand_x4_sg U66329 ( .A(n9578), .B(n9579), .X(n9564) );
  nor_x1_sg U66330 ( .A(n9594), .B(n9595), .X(n9578) );
  nor_x1_sg U66331 ( .A(n9580), .B(n9581), .X(n9579) );
  nand_x2_sg U66332 ( .A(n9596), .B(n9597), .X(n9595) );
  nand_x4_sg U66333 ( .A(n9626), .B(n9627), .X(n9612) );
  nor_x1_sg U66334 ( .A(n9642), .B(n9643), .X(n9626) );
  nor_x1_sg U66335 ( .A(n9628), .B(n9629), .X(n9627) );
  nand_x2_sg U66336 ( .A(n9644), .B(n9645), .X(n9643) );
  nand_x4_sg U66337 ( .A(n9721), .B(n9722), .X(n9707) );
  nor_x1_sg U66338 ( .A(n9737), .B(n9738), .X(n9721) );
  nor_x1_sg U66339 ( .A(n9723), .B(n9724), .X(n9722) );
  nand_x2_sg U66340 ( .A(n9739), .B(n9740), .X(n9738) );
  nand_x4_sg U66341 ( .A(n9769), .B(n9770), .X(n9755) );
  nor_x1_sg U66342 ( .A(n9785), .B(n9786), .X(n9769) );
  nor_x1_sg U66343 ( .A(n9771), .B(n9772), .X(n9770) );
  nand_x2_sg U66344 ( .A(n9787), .B(n9788), .X(n9786) );
  nand_x4_sg U66345 ( .A(n9817), .B(n9818), .X(n9803) );
  nor_x1_sg U66346 ( .A(n9833), .B(n9834), .X(n9817) );
  nor_x1_sg U66347 ( .A(n9819), .B(n9820), .X(n9818) );
  nand_x2_sg U66348 ( .A(n9835), .B(n9836), .X(n9834) );
  nand_x4_sg U66349 ( .A(n9865), .B(n9866), .X(n9851) );
  nor_x1_sg U66350 ( .A(n9881), .B(n9882), .X(n9865) );
  nor_x1_sg U66351 ( .A(n9867), .B(n9868), .X(n9866) );
  nand_x2_sg U66352 ( .A(n9883), .B(n9884), .X(n9882) );
  nand_x4_sg U66353 ( .A(n9913), .B(n9914), .X(n9899) );
  nor_x1_sg U66354 ( .A(n9929), .B(n9930), .X(n9913) );
  nor_x1_sg U66355 ( .A(n9915), .B(n9916), .X(n9914) );
  nand_x2_sg U66356 ( .A(n9931), .B(n9932), .X(n9930) );
  nand_x4_sg U66357 ( .A(n10010), .B(n10011), .X(n9996) );
  nor_x1_sg U66358 ( .A(n10026), .B(n10027), .X(n10010) );
  nor_x1_sg U66359 ( .A(n10012), .B(n10013), .X(n10011) );
  nand_x2_sg U66360 ( .A(n10028), .B(n10029), .X(n10027) );
  nand_x4_sg U66361 ( .A(n10156), .B(n10157), .X(n10142) );
  nor_x1_sg U66362 ( .A(n10172), .B(n10173), .X(n10156) );
  nor_x1_sg U66363 ( .A(n10158), .B(n10159), .X(n10157) );
  nand_x2_sg U66364 ( .A(n10174), .B(n10175), .X(n10173) );
  nand_x4_sg U66365 ( .A(n24686), .B(n24687), .X(n24672) );
  nor_x1_sg U66366 ( .A(n24702), .B(n24703), .X(n24686) );
  nor_x1_sg U66367 ( .A(n24688), .B(n24689), .X(n24687) );
  nand_x2_sg U66368 ( .A(n24704), .B(n24705), .X(n24703) );
  nand_x4_sg U66369 ( .A(n24734), .B(n24735), .X(n24720) );
  nor_x1_sg U66370 ( .A(n24750), .B(n24751), .X(n24734) );
  nor_x1_sg U66371 ( .A(n24736), .B(n24737), .X(n24735) );
  nand_x2_sg U66372 ( .A(n24752), .B(n24753), .X(n24751) );
  nand_x4_sg U66373 ( .A(n24829), .B(n24830), .X(n24815) );
  nor_x1_sg U66374 ( .A(n24845), .B(n24846), .X(n24829) );
  nor_x1_sg U66375 ( .A(n24831), .B(n24832), .X(n24830) );
  nand_x2_sg U66376 ( .A(n24847), .B(n24848), .X(n24846) );
  nand_x4_sg U66377 ( .A(n24877), .B(n24878), .X(n24863) );
  nor_x1_sg U66378 ( .A(n24893), .B(n24894), .X(n24877) );
  nor_x1_sg U66379 ( .A(n24879), .B(n24880), .X(n24878) );
  nand_x2_sg U66380 ( .A(n24895), .B(n24896), .X(n24894) );
  nand_x4_sg U66381 ( .A(n24925), .B(n24926), .X(n24911) );
  nor_x1_sg U66382 ( .A(n24941), .B(n24942), .X(n24925) );
  nor_x1_sg U66383 ( .A(n24927), .B(n24928), .X(n24926) );
  nand_x2_sg U66384 ( .A(n24943), .B(n24944), .X(n24942) );
  nand_x4_sg U66385 ( .A(n24973), .B(n24974), .X(n24959) );
  nor_x1_sg U66386 ( .A(n24989), .B(n24990), .X(n24973) );
  nor_x1_sg U66387 ( .A(n24975), .B(n24976), .X(n24974) );
  nand_x2_sg U66388 ( .A(n24991), .B(n24992), .X(n24990) );
  nand_x4_sg U66389 ( .A(n25021), .B(n25022), .X(n25007) );
  nor_x1_sg U66390 ( .A(n25037), .B(n25038), .X(n25021) );
  nor_x1_sg U66391 ( .A(n25023), .B(n25024), .X(n25022) );
  nand_x2_sg U66392 ( .A(n25039), .B(n25040), .X(n25038) );
  nand_x4_sg U66393 ( .A(n25118), .B(n25119), .X(n25104) );
  nor_x1_sg U66394 ( .A(n25134), .B(n25135), .X(n25118) );
  nor_x1_sg U66395 ( .A(n25120), .B(n25121), .X(n25119) );
  nand_x2_sg U66396 ( .A(n25136), .B(n25137), .X(n25135) );
  nand_x4_sg U66397 ( .A(n25264), .B(n25265), .X(n25250) );
  nor_x1_sg U66398 ( .A(n25280), .B(n25281), .X(n25264) );
  nor_x1_sg U66399 ( .A(n25266), .B(n25267), .X(n25265) );
  nand_x2_sg U66400 ( .A(n25282), .B(n25283), .X(n25281) );
  nand_x4_sg U66401 ( .A(n21942), .B(n21943), .X(n21928) );
  nor_x1_sg U66402 ( .A(n21960), .B(n21961), .X(n21942) );
  nor_x1_sg U66403 ( .A(n21944), .B(n21945), .X(n21943) );
  nand_x2_sg U66404 ( .A(n21966), .B(n21967), .X(n21960) );
  nand_x4_sg U66405 ( .A(n29596), .B(n29597), .X(n29578) );
  nor_x1_sg U66406 ( .A(n29621), .B(n29622), .X(n29596) );
  nor_x1_sg U66407 ( .A(n29598), .B(n29599), .X(n29597) );
  nand_x2_sg U66408 ( .A(n29629), .B(n29630), .X(n29621) );
  nand_x4_sg U66409 ( .A(n10201), .B(n10202), .X(n10189) );
  nor_x1_sg U66410 ( .A(n10203), .B(n10204), .X(n10202) );
  nor_x1_sg U66411 ( .A(n10214), .B(n10215), .X(n10201) );
  nand_x2_sg U66412 ( .A(n10209), .B(n10210), .X(n10203) );
  nand_x4_sg U66413 ( .A(n25309), .B(n25310), .X(n25297) );
  nor_x1_sg U66414 ( .A(n25311), .B(n25312), .X(n25310) );
  nor_x1_sg U66415 ( .A(n25322), .B(n25323), .X(n25309) );
  nand_x2_sg U66416 ( .A(n25317), .B(n25318), .X(n25311) );
  nor_x1_sg U66417 ( .A(n46575), .B(n9356), .X(n9359) );
  nor_x1_sg U66418 ( .A(n46575), .B(n9417), .X(n9420) );
  nor_x1_sg U66419 ( .A(n46575), .B(n9466), .X(n9469) );
  nor_x1_sg U66420 ( .A(n46575), .B(n9515), .X(n9518) );
  nor_x1_sg U66421 ( .A(n46575), .B(n9564), .X(n9567) );
  nor_x1_sg U66422 ( .A(n46575), .B(n9612), .X(n9615) );
  nor_x1_sg U66423 ( .A(n46575), .B(n9660), .X(n9663) );
  nor_x1_sg U66424 ( .A(n46575), .B(n9707), .X(n9710) );
  nor_x1_sg U66425 ( .A(n46575), .B(n9755), .X(n9758) );
  nor_x1_sg U66426 ( .A(n46575), .B(n9803), .X(n9806) );
  nor_x1_sg U66427 ( .A(n46575), .B(n9851), .X(n9854) );
  nor_x1_sg U66428 ( .A(n46575), .B(n9899), .X(n9902) );
  nor_x1_sg U66429 ( .A(n46575), .B(n9947), .X(n9950) );
  nand_x4_sg U66430 ( .A(n18013), .B(n18014), .X(n17993) );
  nand_x1_sg U66431 ( .A(n18017), .B(n53890), .X(n18013) );
  nand_x1_sg U66432 ( .A(n18015), .B(n18016), .X(n18014) );
  nand_x4_sg U66433 ( .A(n19558), .B(n19559), .X(n19538) );
  nand_x1_sg U66434 ( .A(n19562), .B(n54455), .X(n19558) );
  nand_x1_sg U66435 ( .A(n19560), .B(n19561), .X(n19559) );
  nand_x4_sg U66436 ( .A(n21102), .B(n21103), .X(n21082) );
  nand_x1_sg U66437 ( .A(n21106), .B(n55023), .X(n21102) );
  nand_x1_sg U66438 ( .A(n21104), .B(n21105), .X(n21103) );
  nand_x4_sg U66439 ( .A(n17529), .B(n17530), .X(n17495) );
  nand_x4_sg U66440 ( .A(n19074), .B(n19075), .X(n19040) );
  nand_x4_sg U66441 ( .A(n20618), .B(n20619), .X(n20584) );
  nand_x4_sg U66442 ( .A(n12818), .B(n12817), .X(n12819) );
  nand_x4_sg U66443 ( .A(n15151), .B(n15150), .X(n15152) );
  nand_x4_sg U66444 ( .A(n16717), .B(n16716), .X(n16718) );
  nand_x2_sg U66445 ( .A(n46478), .B(n26518), .X(n26517) );
  nand_x4_sg U66446 ( .A(n52788), .B(n14553), .X(n14535) );
  nand_x1_sg U66447 ( .A(n52787), .B(n14554), .X(n14553) );
  nor_x1_sg U66448 ( .A(n52787), .B(n14554), .X(n14555) );
  nand_x4_sg U66449 ( .A(n53908), .B(n17674), .X(n17656) );
  nand_x1_sg U66450 ( .A(n53907), .B(n17675), .X(n17674) );
  nor_x1_sg U66451 ( .A(n53907), .B(n17675), .X(n17676) );
  nand_x4_sg U66452 ( .A(n54473), .B(n19219), .X(n19201) );
  nand_x1_sg U66453 ( .A(n54472), .B(n19220), .X(n19219) );
  nor_x1_sg U66454 ( .A(n54472), .B(n19220), .X(n19221) );
  nand_x4_sg U66455 ( .A(n55041), .B(n20763), .X(n20745) );
  nand_x1_sg U66456 ( .A(n55040), .B(n20764), .X(n20763) );
  nor_x1_sg U66457 ( .A(n55040), .B(n20764), .X(n20765) );
  nand_x4_sg U66458 ( .A(n18818), .B(n18819), .X(n18628) );
  nand_x1_sg U66459 ( .A(n54256), .B(n18815), .X(n18819) );
  nand_x1_sg U66460 ( .A(n54114), .B(n18814), .X(n18818) );
  nand_x4_sg U66461 ( .A(n10893), .B(n51518), .X(n10891) );
  nand_x1_sg U66462 ( .A(n41586), .B(n10895), .X(n10893) );
  nor_x1_sg U66463 ( .A(n10895), .B(n51517), .X(n10894) );
  nand_x4_sg U66464 ( .A(n16348), .B(n53467), .X(n16346) );
  nand_x1_sg U66465 ( .A(n41428), .B(n16350), .X(n16348) );
  nor_x1_sg U66466 ( .A(n16350), .B(n53466), .X(n16349) );
  nand_x4_sg U66467 ( .A(n11031), .B(n11032), .X(n10848) );
  nand_x1_sg U66468 ( .A(n51323), .B(n11027), .X(n11031) );
  nand_x1_sg U66469 ( .A(n51463), .B(n11028), .X(n11032) );
  nand_x4_sg U66470 ( .A(n20077), .B(n54795), .X(n20073) );
  nor_x1_sg U66471 ( .A(n20079), .B(n20080), .X(n20078) );
  nand_x4_sg U66472 ( .A(n21622), .B(n55363), .X(n21618) );
  nor_x1_sg U66473 ( .A(n21624), .B(n21625), .X(n21623) );
  nand_x4_sg U66474 ( .A(n14643), .B(n52825), .X(n14639) );
  nor_x1_sg U66475 ( .A(n14645), .B(n14646), .X(n14644) );
  nand_x4_sg U66476 ( .A(n17764), .B(n53945), .X(n17760) );
  nor_x1_sg U66477 ( .A(n17766), .B(n17767), .X(n17765) );
  nand_x4_sg U66478 ( .A(n19309), .B(n54510), .X(n19305) );
  nor_x1_sg U66479 ( .A(n19311), .B(n19312), .X(n19310) );
  nand_x4_sg U66480 ( .A(n20853), .B(n55078), .X(n20849) );
  nor_x1_sg U66481 ( .A(n20855), .B(n20856), .X(n20854) );
  nor_x1_sg U66482 ( .A(n46615), .B(n24525), .X(n24528) );
  nor_x1_sg U66483 ( .A(n46615), .B(n24574), .X(n24577) );
  nor_x1_sg U66484 ( .A(n46615), .B(n24672), .X(n24675) );
  nor_x1_sg U66485 ( .A(n46615), .B(n24720), .X(n24723) );
  nor_x1_sg U66486 ( .A(n46615), .B(n24815), .X(n24818) );
  nor_x1_sg U66487 ( .A(n46615), .B(n24863), .X(n24866) );
  nor_x1_sg U66488 ( .A(n46615), .B(n24959), .X(n24962) );
  nor_x1_sg U66489 ( .A(n46615), .B(n25007), .X(n25010) );
  nor_x1_sg U66490 ( .A(n46615), .B(n25104), .X(n25107) );
  nor_x1_sg U66491 ( .A(n46615), .B(n25152), .X(n25155) );
  nor_x1_sg U66492 ( .A(n46615), .B(n25250), .X(n25253) );
  nor_x1_sg U66493 ( .A(n46615), .B(n25297), .X(n25300) );
  nand_x4_sg U66494 ( .A(n12616), .B(n12617), .X(n8846) );
  nand_x4_sg U66495 ( .A(n13400), .B(n13401), .X(n8805) );
  nand_x4_sg U66496 ( .A(n14949), .B(n14950), .X(n8988) );
  nand_x4_sg U66497 ( .A(n16515), .B(n16516), .X(n9313) );
  nor_x1_sg U66498 ( .A(n53792), .B(n42166), .X(n17427) );
  nor_x1_sg U66499 ( .A(n54073), .B(n44195), .X(n18194) );
  nor_x1_sg U66500 ( .A(n54357), .B(n42164), .X(n18972) );
  nor_x1_sg U66501 ( .A(n54925), .B(n42162), .X(n20516) );
  nor_x1_sg U66502 ( .A(n52673), .B(n44199), .X(n14306) );
  nor_x1_sg U66503 ( .A(n51845), .B(n44203), .X(n11964) );
  nor_x1_sg U66504 ( .A(n53231), .B(n44197), .X(n15859) );
  nor_x1_sg U66505 ( .A(n51567), .B(n42160), .X(n11186) );
  nor_x1_sg U66506 ( .A(n52124), .B(n42158), .X(n12747) );
  nor_x1_sg U66507 ( .A(n52958), .B(n42156), .X(n15080) );
  nor_x1_sg U66508 ( .A(n53516), .B(n42154), .X(n16646) );
  nor_x1_sg U66509 ( .A(n51283), .B(n42152), .X(n10414) );
  nor_x1_sg U66510 ( .A(n54637), .B(n41964), .X(n19741) );
  nor_x1_sg U66511 ( .A(n55205), .B(n41962), .X(n21286) );
  nand_x4_sg U66512 ( .A(n20296), .B(n20297), .X(n20294) );
  nand_x1_sg U66513 ( .A(n54849), .B(n20299), .X(n20296) );
  nor_x1_sg U66514 ( .A(n54849), .B(n46287), .X(n20298) );
  nand_x4_sg U66515 ( .A(n21841), .B(n21842), .X(n21839) );
  nand_x1_sg U66516 ( .A(n55417), .B(n21844), .X(n21841) );
  nor_x1_sg U66517 ( .A(n55417), .B(n46242), .X(n21843) );
  nand_x4_sg U66518 ( .A(n17471), .B(n17472), .X(n17462) );
  nand_x4_sg U66519 ( .A(n19016), .B(n19017), .X(n19007) );
  nand_x4_sg U66520 ( .A(n20560), .B(n20561), .X(n20551) );
  nand_x4_sg U66521 ( .A(n14860), .B(n14861), .X(n14858) );
  nand_x1_sg U66522 ( .A(n52879), .B(n14863), .X(n14860) );
  nand_x1_sg U66523 ( .A(n52707), .B(n52742), .X(n14863) );
  nand_x4_sg U66524 ( .A(n18070), .B(n18071), .X(n9071) );
  nand_x4_sg U66525 ( .A(n18237), .B(n18238), .X(n18228) );
  nand_x1_sg U66526 ( .A(n41711), .B(n54099), .X(n18238) );
  nand_x4_sg U66527 ( .A(n14345), .B(n14346), .X(n14339) );
  nand_x1_sg U66528 ( .A(n46450), .B(n52698), .X(n14346) );
  nand_x4_sg U66529 ( .A(n11212), .B(n11213), .X(n11201) );
  nand_x1_sg U66530 ( .A(n51572), .B(n51576), .X(n11213) );
  nand_x4_sg U66531 ( .A(n12773), .B(n12774), .X(n12762) );
  nand_x1_sg U66532 ( .A(n52129), .B(n52134), .X(n12774) );
  nand_x4_sg U66533 ( .A(n15106), .B(n15107), .X(n15095) );
  nand_x1_sg U66534 ( .A(n52963), .B(n52968), .X(n15107) );
  nand_x4_sg U66535 ( .A(n16672), .B(n16673), .X(n16661) );
  nand_x1_sg U66536 ( .A(n53521), .B(n53526), .X(n16673) );
  nand_x4_sg U66537 ( .A(n10456), .B(n10457), .X(n10447) );
  nand_x1_sg U66538 ( .A(n46564), .B(n51309), .X(n10457) );
  nand_x4_sg U66539 ( .A(n19783), .B(n19784), .X(n19774) );
  nand_x1_sg U66540 ( .A(n46294), .B(n54663), .X(n19784) );
  nand_x4_sg U66541 ( .A(n21328), .B(n21329), .X(n21319) );
  nand_x1_sg U66542 ( .A(n46249), .B(n55231), .X(n21329) );
  nand_x4_sg U66543 ( .A(n10392), .B(n10393), .X(n10294) );
  nand_x1_sg U66544 ( .A(n10395), .B(n10396), .X(n10392) );
  nor_x1_sg U66545 ( .A(n10395), .B(n46570), .X(n10394) );
  nor_x1_sg U66546 ( .A(n46575), .B(n21928), .X(n21931) );
  nor_x1_sg U66547 ( .A(n46575), .B(n9996), .X(n9999) );
  nor_x1_sg U66548 ( .A(n46575), .B(n10044), .X(n10047) );
  nor_x1_sg U66549 ( .A(n46575), .B(n10093), .X(n10096) );
  nor_x1_sg U66550 ( .A(n46575), .B(n10142), .X(n10145) );
  nor_x1_sg U66551 ( .A(n46575), .B(n10189), .X(n10192) );
  nand_x4_sg U66552 ( .A(n18750), .B(n18751), .X(n18748) );
  nand_x1_sg U66553 ( .A(n54282), .B(n18753), .X(n18750) );
  nor_x1_sg U66554 ( .A(n54282), .B(n46331), .X(n18752) );
  nor_x1_sg U66555 ( .A(n25794), .B(n25795), .X(\L1_0/n4591 ) );
  nand_x2_sg U66556 ( .A(n25796), .B(n46235), .X(n25794) );
  nor_x1_sg U66557 ( .A(n46611), .B(n51804), .X(n25796) );
  nor_x1_sg U66558 ( .A(n26910), .B(n26911), .X(\L1_0/n4271 ) );
  nand_x2_sg U66559 ( .A(n26912), .B(n46235), .X(n26910) );
  nor_x1_sg U66560 ( .A(n46625), .B(n52914), .X(n26912) );
  nor_x1_sg U66561 ( .A(n27469), .B(n27470), .X(\L1_0/n4111 ) );
  nand_x2_sg U66562 ( .A(n27471), .B(n46235), .X(n27469) );
  nor_x1_sg U66563 ( .A(n55786), .B(n53472), .X(n27471) );
  nor_x1_sg U66564 ( .A(n28029), .B(n28030), .X(\L1_0/n3951 ) );
  nand_x2_sg U66565 ( .A(n28031), .B(n46592), .X(n28029) );
  nor_x1_sg U66566 ( .A(n54034), .B(n46236), .X(n28031) );
  nor_x1_sg U66567 ( .A(n28309), .B(n28310), .X(\L1_0/n3871 ) );
  nand_x2_sg U66568 ( .A(n28311), .B(n46594), .X(n28309) );
  nor_x1_sg U66569 ( .A(n54315), .B(n46236), .X(n28311) );
  nor_x1_sg U66570 ( .A(n28587), .B(n28588), .X(\L1_0/n3791 ) );
  nand_x2_sg U66571 ( .A(n28589), .B(n46595), .X(n28587) );
  nor_x1_sg U66572 ( .A(n54599), .B(n46236), .X(n28589) );
  nor_x1_sg U66573 ( .A(n28867), .B(n28868), .X(\L1_0/n3711 ) );
  nand_x2_sg U66574 ( .A(n28869), .B(n46235), .X(n28867) );
  nor_x1_sg U66575 ( .A(n55784), .B(n54883), .X(n28869) );
  nor_x1_sg U66576 ( .A(n29428), .B(n29429), .X(\L1_0/n3551 ) );
  nand_x2_sg U66577 ( .A(n29430), .B(n46597), .X(n29428) );
  nor_x1_sg U66578 ( .A(n55451), .B(n46236), .X(n29430) );
  nand_x4_sg U66579 ( .A(n11257), .B(n11256), .X(n11258) );
  nand_x4_sg U66580 ( .A(n12202), .B(n12215), .X(n12198) );
  nand_x1_sg U66581 ( .A(n51867), .B(n51889), .X(n12216) );
  nand_x4_sg U66582 ( .A(n16097), .B(n16110), .X(n16093) );
  nand_x1_sg U66583 ( .A(n53254), .B(n53276), .X(n16111) );
  nand_x4_sg U66584 ( .A(n11422), .B(n11435), .X(n11418) );
  nand_x1_sg U66585 ( .A(n51595), .B(n51608), .X(n11436) );
  nand_x4_sg U66586 ( .A(n12983), .B(n12996), .X(n12979) );
  nand_x1_sg U66587 ( .A(n52153), .B(n52166), .X(n12997) );
  nand_x4_sg U66588 ( .A(n15316), .B(n15329), .X(n15312) );
  nand_x1_sg U66589 ( .A(n52987), .B(n53000), .X(n15330) );
  nand_x4_sg U66590 ( .A(n16882), .B(n16895), .X(n16878) );
  nand_x1_sg U66591 ( .A(n53545), .B(n53558), .X(n16896) );
  nor_x1_sg U66592 ( .A(n26073), .B(n26074), .X(\L1_0/n4511 ) );
  nor_x1_sg U66593 ( .A(n52080), .B(n46236), .X(n26075) );
  nor_x1_sg U66594 ( .A(n26354), .B(n26355), .X(\L1_0/n4431 ) );
  nand_x2_sg U66595 ( .A(n26356), .B(n46586), .X(n26354) );
  nor_x1_sg U66596 ( .A(n52358), .B(n46236), .X(n26356) );
  nor_x1_sg U66597 ( .A(n26633), .B(n26634), .X(\L1_0/n4351 ) );
  nand_x2_sg U66598 ( .A(n26635), .B(n46588), .X(n26633) );
  nor_x1_sg U66599 ( .A(n52633), .B(n46236), .X(n26635) );
  nor_x1_sg U66600 ( .A(n27190), .B(n27191), .X(\L1_0/n4191 ) );
  nand_x2_sg U66601 ( .A(n27192), .B(n46590), .X(n27190) );
  nor_x1_sg U66602 ( .A(n53192), .B(n46236), .X(n27192) );
  nor_x1_sg U66603 ( .A(n27750), .B(n27751), .X(\L1_0/n4031 ) );
  nand_x2_sg U66604 ( .A(n27752), .B(n46235), .X(n27750) );
  nor_x1_sg U66605 ( .A(n55785), .B(n53750), .X(n27752) );
  nor_x1_sg U66606 ( .A(n46611), .B(n55527), .X(\L1_0/n4594 ) );
  nand_x2_sg U66607 ( .A(n46339), .B(n28208), .X(n28207) );
  nand_x4_sg U66608 ( .A(n13386), .B(n13387), .X(n13221) );
  nand_x1_sg U66609 ( .A(n12995), .B(n13388), .X(n13386) );
  nand_x4_sg U66610 ( .A(n15719), .B(n15720), .X(n15554) );
  nand_x1_sg U66611 ( .A(n15328), .B(n15721), .X(n15719) );
  nand_x4_sg U66612 ( .A(n17285), .B(n17286), .X(n17120) );
  nand_x1_sg U66613 ( .A(n16894), .B(n17287), .X(n17285) );
  nand_x4_sg U66614 ( .A(n13504), .B(n13505), .X(n13407) );
  nand_x1_sg U66615 ( .A(n13507), .B(n13508), .X(n13504) );
  nor_x1_sg U66616 ( .A(n13507), .B(n46480), .X(n13506) );
  nand_x4_sg U66617 ( .A(n12006), .B(n12007), .X(n11999) );
  nand_x1_sg U66618 ( .A(n46517), .B(n51868), .X(n12007) );
  nand_x4_sg U66619 ( .A(n13567), .B(n13568), .X(n13560) );
  nand_x1_sg U66620 ( .A(n46474), .B(n52420), .X(n13568) );
  nand_x4_sg U66621 ( .A(n12573), .B(n12581), .X(n12380) );
  nand_x1_sg U66622 ( .A(n12582), .B(n12583), .X(n12581) );
  nor_x1_sg U66623 ( .A(n44677), .B(n40880), .X(n12582) );
  nor_x1_sg U66624 ( .A(n12586), .B(n12587), .X(n12585) );
  nand_x1_sg U66625 ( .A(n11204), .B(n11205), .X(n11203) );
  nor_x1_sg U66626 ( .A(n51577), .B(n11206), .X(n11204) );
  nand_x1_sg U66627 ( .A(n12765), .B(n12766), .X(n12764) );
  nor_x1_sg U66628 ( .A(n52135), .B(n12767), .X(n12765) );
  nand_x1_sg U66629 ( .A(n15098), .B(n15099), .X(n15097) );
  nor_x1_sg U66630 ( .A(n52969), .B(n15100), .X(n15098) );
  nand_x1_sg U66631 ( .A(n16664), .B(n16665), .X(n16663) );
  nor_x1_sg U66632 ( .A(n53527), .B(n16666), .X(n16664) );
  nand_x4_sg U66633 ( .A(n10827), .B(n10833), .X(n10758) );
  nand_x1_sg U66634 ( .A(n10834), .B(n10835), .X(n10833) );
  nor_x1_sg U66635 ( .A(n10836), .B(n10837), .X(n10834) );
  nand_x4_sg U66636 ( .A(n18607), .B(n18613), .X(n18539) );
  nand_x1_sg U66637 ( .A(n18614), .B(n18615), .X(n18613) );
  nor_x1_sg U66638 ( .A(n43848), .B(n18617), .X(n18614) );
  nand_x4_sg U66639 ( .A(n17840), .B(n17846), .X(n17771) );
  nand_x1_sg U66640 ( .A(n17847), .B(n17848), .X(n17846) );
  nor_x1_sg U66641 ( .A(n43978), .B(n17850), .X(n17847) );
  nand_x4_sg U66642 ( .A(n19385), .B(n19391), .X(n19316) );
  nand_x1_sg U66643 ( .A(n19392), .B(n19393), .X(n19391) );
  nor_x1_sg U66644 ( .A(n43977), .B(n19395), .X(n19392) );
  nand_x4_sg U66645 ( .A(n20929), .B(n20935), .X(n20860) );
  nand_x1_sg U66646 ( .A(n20936), .B(n20937), .X(n20935) );
  nor_x1_sg U66647 ( .A(n43976), .B(n20939), .X(n20936) );
  nand_x4_sg U66648 ( .A(n16283), .B(n16289), .X(n16215) );
  nand_x1_sg U66649 ( .A(n16290), .B(n16291), .X(n16289) );
  nor_x1_sg U66650 ( .A(n44358), .B(n16293), .X(n16290) );
  nand_x4_sg U66651 ( .A(n20153), .B(n20159), .X(n20084) );
  nand_x1_sg U66652 ( .A(n20160), .B(n20161), .X(n20159) );
  nor_x1_sg U66653 ( .A(n43803), .B(n20163), .X(n20160) );
  nand_x4_sg U66654 ( .A(n21698), .B(n21704), .X(n21629) );
  nand_x1_sg U66655 ( .A(n21705), .B(n21706), .X(n21704) );
  nor_x1_sg U66656 ( .A(n43782), .B(n21708), .X(n21705) );
  nand_x4_sg U66657 ( .A(n12388), .B(n12394), .X(n12320) );
  nand_x1_sg U66658 ( .A(n12395), .B(n12396), .X(n12394) );
  nor_x1_sg U66659 ( .A(n44361), .B(n12398), .X(n12395) );
  nand_x1_sg U66660 ( .A(n15877), .B(n15878), .X(n15876) );
  nor_x1_sg U66661 ( .A(n53242), .B(n15879), .X(n15877) );
  nand_x1_sg U66662 ( .A(n11982), .B(n11983), .X(n11981) );
  nor_x1_sg U66663 ( .A(n51856), .B(n11984), .X(n11982) );
  nand_x4_sg U66664 ( .A(n14719), .B(n14725), .X(n14650) );
  nand_x1_sg U66665 ( .A(n14726), .B(n14727), .X(n14725) );
  nor_x1_sg U66666 ( .A(n43783), .B(n14729), .X(n14726) );
  nand_x4_sg U66667 ( .A(n11607), .B(n11613), .X(n11540) );
  nand_x1_sg U66668 ( .A(n11614), .B(n11615), .X(n11613) );
  nor_x1_sg U66669 ( .A(n43980), .B(n11617), .X(n11614) );
  nand_x4_sg U66670 ( .A(n13168), .B(n13174), .X(n13101) );
  nand_x1_sg U66671 ( .A(n13175), .B(n13176), .X(n13174) );
  nor_x1_sg U66672 ( .A(n44360), .B(n13178), .X(n13175) );
  nand_x4_sg U66673 ( .A(n15501), .B(n15507), .X(n15434) );
  nand_x1_sg U66674 ( .A(n15508), .B(n15509), .X(n15507) );
  nor_x1_sg U66675 ( .A(n44359), .B(n15511), .X(n15508) );
  nand_x4_sg U66676 ( .A(n17067), .B(n17073), .X(n17000) );
  nand_x1_sg U66677 ( .A(n17074), .B(n17075), .X(n17073) );
  nor_x1_sg U66678 ( .A(n44357), .B(n17077), .X(n17074) );
  nand_x4_sg U66679 ( .A(n15901), .B(n15902), .X(n15894) );
  nand_x1_sg U66680 ( .A(n46405), .B(n53255), .X(n15902) );
  nand_x4_sg U66681 ( .A(n12198), .B(n12200), .X(n12152) );
  nor_x1_sg U66682 ( .A(n12203), .B(n12204), .X(n12201) );
  nand_x4_sg U66683 ( .A(n16093), .B(n16095), .X(n16047) );
  nor_x1_sg U66684 ( .A(n16098), .B(n16099), .X(n16096) );
  nand_x4_sg U66685 ( .A(n11418), .B(n11420), .X(n11372) );
  nor_x1_sg U66686 ( .A(n11423), .B(n11424), .X(n11421) );
  nand_x4_sg U66687 ( .A(n12979), .B(n12981), .X(n12933) );
  nor_x1_sg U66688 ( .A(n12984), .B(n12985), .X(n12982) );
  nand_x4_sg U66689 ( .A(n15312), .B(n15314), .X(n15266) );
  nor_x1_sg U66690 ( .A(n15317), .B(n15318), .X(n15315) );
  nand_x4_sg U66691 ( .A(n16878), .B(n16880), .X(n16832) );
  nor_x1_sg U66692 ( .A(n16883), .B(n16884), .X(n16881) );
  nor_x1_sg U66693 ( .A(n54086), .B(n18213), .X(n18211) );
  nor_x1_sg U66694 ( .A(n51295), .B(n10432), .X(n10430) );
  nor_x1_sg U66695 ( .A(n52685), .B(n14324), .X(n14322) );
  nor_x1_sg U66696 ( .A(n54649), .B(n19759), .X(n19757) );
  nor_x1_sg U66697 ( .A(n55217), .B(n21304), .X(n21302) );
  nor_x1_sg U66698 ( .A(n21927), .B(n9355), .X(\L2_0/n2904 ) );
  nand_x2_sg U66699 ( .A(n10205), .B(n10206), .X(n10204) );
  nor_x1_sg U66700 ( .A(n10207), .B(n10208), .X(n10205) );
  nand_x1_sg U66701 ( .A(n46602), .B(n50153), .X(n10206) );
  nand_x2_sg U66702 ( .A(n25313), .B(n25314), .X(n25312) );
  nor_x1_sg U66703 ( .A(n25315), .B(n25316), .X(n25313) );
  nand_x1_sg U66704 ( .A(n49294), .B(n46602), .X(n25314) );
  nor_x1_sg U66705 ( .A(n55621), .B(n46618), .X(\L1_0/n3634 ) );
  nor_x1_sg U66706 ( .A(n46616), .B(n29140), .X(\L1_0/n3635 ) );
  nor_x1_sg U66707 ( .A(n46614), .B(n26067), .X(\L1_0/n4515 ) );
  nor_x1_sg U66708 ( .A(n55534), .B(n46612), .X(\L1_0/n4514 ) );
  nor_x1_sg U66709 ( .A(n46625), .B(n55558), .X(\L1_0/n4274 ) );
  nor_x1_sg U66710 ( .A(n46621), .B(n55581), .X(\L1_0/n4034 ) );
  nor_x1_sg U66711 ( .A(n46623), .B(n55573), .X(\L1_0/n4114 ) );
  nor_x1_sg U66712 ( .A(n46619), .B(n55613), .X(\L1_0/n3714 ) );
  nor_x1_sg U66713 ( .A(n46615), .B(n55520), .X(\L1_0/n4674 ) );
  nand_x2_sg U66714 ( .A(n10216), .B(n10217), .X(n10215) );
  nand_x1_sg U66715 ( .A(n46598), .B(n50143), .X(n10217) );
  nand_x1_sg U66716 ( .A(n50141), .B(n46608), .X(n10216) );
  nand_x2_sg U66717 ( .A(n25324), .B(n25325), .X(n25323) );
  nand_x1_sg U66718 ( .A(n49284), .B(n46598), .X(n25325) );
  nand_x1_sg U66719 ( .A(n49282), .B(n46608), .X(n25324) );
  nand_x2_sg U66720 ( .A(n24800), .B(n24801), .X(n24799) );
  nand_x1_sg U66721 ( .A(n49788), .B(n46598), .X(n24801) );
  nand_x2_sg U66722 ( .A(n9692), .B(n9693), .X(n9691) );
  nand_x1_sg U66723 ( .A(n46598), .B(n50647), .X(n9693) );
  inv_x4_sg U66724 ( .A(n46660), .X(n46659) );
  inv_x4_sg U66725 ( .A(n43784), .X(n46640) );
  nand_x1_sg U66726 ( .A(n44088), .B(n46355), .X(n9055) );
  nand_x1_sg U66727 ( .A(n46355), .B(n44108), .X(n9051) );
  nand_x1_sg U66728 ( .A(n42865), .B(n46355), .X(n9078) );
  nand_x1_sg U66729 ( .A(n44395), .B(n46355), .X(n9058) );
  nand_x1_sg U66730 ( .A(n44086), .B(n46308), .X(n9167) );
  nand_x1_sg U66731 ( .A(n41970), .B(n46308), .X(n9174) );
  nand_x1_sg U66732 ( .A(n42861), .B(n46308), .X(n9188) );
  nand_x1_sg U66733 ( .A(n44391), .B(n46308), .X(n9184) );
  nand_x2_sg U66734 ( .A(n25821), .B(n25820), .X(n25818) );
  nor_x1_sg U66735 ( .A(n25820), .B(n25821), .X(n25819) );
  nand_x2_sg U66736 ( .A(n26937), .B(n26936), .X(n26934) );
  nor_x1_sg U66737 ( .A(n26936), .B(n26937), .X(n26935) );
  nand_x2_sg U66738 ( .A(n27508), .B(n27507), .X(n27505) );
  nor_x1_sg U66739 ( .A(n27507), .B(n27508), .X(n27506) );
  nand_x2_sg U66740 ( .A(n27496), .B(n27495), .X(n27493) );
  nor_x1_sg U66741 ( .A(n27495), .B(n27496), .X(n27494) );
  nand_x4_sg U66742 ( .A(n12826), .B(n46496), .X(n12987) );
  nand_x4_sg U66743 ( .A(n15159), .B(n46428), .X(n15320) );
  nand_x4_sg U66744 ( .A(n16725), .B(n46384), .X(n16886) );
  nand_x2_sg U66745 ( .A(n25833), .B(n25832), .X(n25830) );
  nor_x1_sg U66746 ( .A(n25832), .B(n25833), .X(n25831) );
  nand_x2_sg U66747 ( .A(n26392), .B(n26391), .X(n26389) );
  nor_x1_sg U66748 ( .A(n26391), .B(n26392), .X(n26390) );
  nand_x2_sg U66749 ( .A(n27229), .B(n27228), .X(n27226) );
  nor_x1_sg U66750 ( .A(n27228), .B(n27229), .X(n27227) );
  nand_x2_sg U66751 ( .A(n27787), .B(n27786), .X(n27784) );
  nor_x1_sg U66752 ( .A(n27786), .B(n27787), .X(n27785) );
  nand_x4_sg U66753 ( .A(n54818), .B(n46305), .X(n20359) );
  nand_x4_sg U66754 ( .A(n55386), .B(n46260), .X(n21904) );
  nand_x4_sg U66755 ( .A(n51738), .B(n46551), .X(n11811) );
  nand_x4_sg U66756 ( .A(n52848), .B(n46462), .X(n14922) );
  nand_x4_sg U66757 ( .A(n53408), .B(n46417), .X(n16486) );
  nand_x4_sg U66758 ( .A(n53968), .B(n46372), .X(n18043) );
  nand_x4_sg U66759 ( .A(n54250), .B(n46352), .X(n18814) );
  nand_x4_sg U66760 ( .A(n54533), .B(n46325), .X(n19588) );
  nand_x4_sg U66761 ( .A(n55101), .B(n46280), .X(n21132) );
  nand_x4_sg U66762 ( .A(n13268), .B(n46507), .X(n13368) );
  nand_x4_sg U66763 ( .A(n15601), .B(n46439), .X(n15701) );
  nand_x4_sg U66764 ( .A(n17167), .B(n46395), .X(n17267) );
  nand_x4_sg U66765 ( .A(n12487), .B(n46529), .X(n12586) );
  nand_x2_sg U66766 ( .A(n28910), .B(n28909), .X(n28907) );
  nor_x1_sg U66767 ( .A(n28909), .B(n28910), .X(n28908) );
  nand_x2_sg U66768 ( .A(n29471), .B(n29470), .X(n29468) );
  nor_x1_sg U66769 ( .A(n29470), .B(n29471), .X(n29469) );
  nand_x2_sg U66770 ( .A(n25536), .B(n25535), .X(n25533) );
  nor_x1_sg U66771 ( .A(n25535), .B(n25536), .X(n25534) );
  nand_x2_sg U66772 ( .A(n26095), .B(n26094), .X(n26092) );
  nor_x1_sg U66773 ( .A(n26094), .B(n26095), .X(n26093) );
  nand_x2_sg U66774 ( .A(n27490), .B(n27489), .X(n27487) );
  nor_x1_sg U66775 ( .A(n27489), .B(n27490), .X(n27488) );
  nand_x2_sg U66776 ( .A(n26119), .B(n26118), .X(n26116) );
  nor_x1_sg U66777 ( .A(n26118), .B(n26119), .X(n26117) );
  nand_x2_sg U66778 ( .A(n26113), .B(n26112), .X(n26110) );
  nor_x1_sg U66779 ( .A(n26112), .B(n26113), .X(n26111) );
  nand_x2_sg U66780 ( .A(n26670), .B(n26669), .X(n26667) );
  nor_x1_sg U66781 ( .A(n26669), .B(n26670), .X(n26668) );
  nand_x2_sg U66782 ( .A(n26101), .B(n26100), .X(n26098) );
  nor_x1_sg U66783 ( .A(n26100), .B(n26101), .X(n26099) );
  nand_x2_sg U66784 ( .A(n26380), .B(n26379), .X(n26377) );
  nor_x1_sg U66785 ( .A(n26379), .B(n26380), .X(n26378) );
  nand_x2_sg U66786 ( .A(n26658), .B(n26657), .X(n26655) );
  nor_x1_sg U66787 ( .A(n26657), .B(n26658), .X(n26656) );
  nand_x2_sg U66788 ( .A(n26949), .B(n26948), .X(n26946) );
  nor_x1_sg U66789 ( .A(n26948), .B(n26949), .X(n26947) );
  nand_x2_sg U66790 ( .A(n27217), .B(n27216), .X(n27214) );
  nor_x1_sg U66791 ( .A(n27216), .B(n27217), .X(n27215) );
  nand_x2_sg U66792 ( .A(n27775), .B(n27774), .X(n27772) );
  nor_x1_sg U66793 ( .A(n27774), .B(n27775), .X(n27773) );
  nand_x2_sg U66794 ( .A(n28068), .B(n28067), .X(n28065) );
  nor_x1_sg U66795 ( .A(n28067), .B(n28068), .X(n28066) );
  nand_x2_sg U66796 ( .A(n28056), .B(n28055), .X(n28053) );
  nor_x1_sg U66797 ( .A(n28055), .B(n28056), .X(n28054) );
  nand_x2_sg U66798 ( .A(n28337), .B(n28336), .X(n28334) );
  nor_x1_sg U66799 ( .A(n28336), .B(n28337), .X(n28335) );
  nand_x2_sg U66800 ( .A(n28626), .B(n28625), .X(n28623) );
  nor_x1_sg U66801 ( .A(n28625), .B(n28626), .X(n28624) );
  nand_x2_sg U66802 ( .A(n28614), .B(n28613), .X(n28611) );
  nor_x1_sg U66803 ( .A(n28613), .B(n28614), .X(n28612) );
  nand_x2_sg U66804 ( .A(n29187), .B(n29186), .X(n29184) );
  nor_x1_sg U66805 ( .A(n29186), .B(n29187), .X(n29185) );
  nand_x2_sg U66806 ( .A(n29175), .B(n29174), .X(n29172) );
  nor_x1_sg U66807 ( .A(n29174), .B(n29175), .X(n29173) );
  nand_x2_sg U66808 ( .A(n46582), .B(n26358), .X(n32136) );
  nand_x4_sg U66809 ( .A(n54751), .B(n46305), .X(n20059) );
  nand_x4_sg U66810 ( .A(n55319), .B(n46260), .X(n21604) );
  nand_x2_sg U66811 ( .A(n25558), .B(n25557), .X(n25555) );
  nor_x1_sg U66812 ( .A(n25557), .B(n25558), .X(n25556) );
  nand_x2_sg U66813 ( .A(n28353), .B(n28352), .X(n28350) );
  nor_x1_sg U66814 ( .A(n28352), .B(n28353), .X(n28351) );
  nand_x2_sg U66815 ( .A(n28343), .B(n28342), .X(n28340) );
  nor_x1_sg U66816 ( .A(n28342), .B(n28343), .X(n28341) );
  nand_x2_sg U66817 ( .A(n28900), .B(n28899), .X(n28897) );
  nor_x1_sg U66818 ( .A(n28899), .B(n28900), .X(n28898) );
  nand_x2_sg U66819 ( .A(n29461), .B(n29460), .X(n29458) );
  nor_x1_sg U66820 ( .A(n29460), .B(n29461), .X(n29459) );
  nand_x2_sg U66821 ( .A(n26676), .B(n26675), .X(n26673) );
  nor_x1_sg U66822 ( .A(n26675), .B(n26676), .X(n26674) );
  nand_x2_sg U66823 ( .A(n27514), .B(n27513), .X(n27511) );
  nor_x1_sg U66824 ( .A(n27513), .B(n27514), .X(n27512) );
  nand_x4_sg U66825 ( .A(n51458), .B(n46574), .X(n11027) );
  nand_x2_sg U66826 ( .A(n14768), .B(n46443), .X(n14851) );
  nand_x2_sg U66827 ( .A(n17889), .B(n46356), .X(n17972) );
  nand_x2_sg U66828 ( .A(n19434), .B(n46309), .X(n19517) );
  nand_x2_sg U66829 ( .A(n20978), .B(n46264), .X(n21061) );
  nand_x1_sg U66830 ( .A(n10907), .B(n46574), .X(n10909) );
  nand_x2_sg U66831 ( .A(n25548), .B(n25547), .X(n25545) );
  nor_x1_sg U66832 ( .A(n25547), .B(n25548), .X(n25546) );
  nand_x2_sg U66833 ( .A(n25827), .B(n25826), .X(n25824) );
  nor_x1_sg U66834 ( .A(n25826), .B(n25827), .X(n25825) );
  nand_x2_sg U66835 ( .A(n25815), .B(n25814), .X(n25812) );
  nor_x1_sg U66836 ( .A(n25814), .B(n25815), .X(n25813) );
  nand_x2_sg U66837 ( .A(n26107), .B(n26106), .X(n26104) );
  nor_x1_sg U66838 ( .A(n26106), .B(n26107), .X(n26105) );
  nand_x2_sg U66839 ( .A(n26386), .B(n26385), .X(n26383) );
  nor_x1_sg U66840 ( .A(n26385), .B(n26386), .X(n26384) );
  nand_x2_sg U66841 ( .A(n26664), .B(n26663), .X(n26661) );
  nor_x1_sg U66842 ( .A(n26663), .B(n26664), .X(n26662) );
  nand_x2_sg U66843 ( .A(n26943), .B(n26942), .X(n26940) );
  nor_x1_sg U66844 ( .A(n26942), .B(n26943), .X(n26941) );
  nand_x2_sg U66845 ( .A(n27223), .B(n27222), .X(n27220) );
  nor_x1_sg U66846 ( .A(n27222), .B(n27223), .X(n27221) );
  nand_x2_sg U66847 ( .A(n27502), .B(n27501), .X(n27499) );
  nor_x1_sg U66848 ( .A(n27501), .B(n27502), .X(n27500) );
  nand_x2_sg U66849 ( .A(n27781), .B(n27780), .X(n27778) );
  nor_x1_sg U66850 ( .A(n27780), .B(n27781), .X(n27779) );
  nand_x2_sg U66851 ( .A(n28062), .B(n28061), .X(n28059) );
  nor_x1_sg U66852 ( .A(n28061), .B(n28062), .X(n28060) );
  nand_x2_sg U66853 ( .A(n28620), .B(n28619), .X(n28617) );
  nor_x1_sg U66854 ( .A(n28619), .B(n28620), .X(n28618) );
  nand_x2_sg U66855 ( .A(n28888), .B(n28887), .X(n28885) );
  nor_x1_sg U66856 ( .A(n28887), .B(n28888), .X(n28886) );
  nand_x2_sg U66857 ( .A(n29181), .B(n29180), .X(n29178) );
  nor_x1_sg U66858 ( .A(n29180), .B(n29181), .X(n29179) );
  nand_x2_sg U66859 ( .A(n29449), .B(n29448), .X(n29446) );
  nor_x1_sg U66860 ( .A(n29448), .B(n29449), .X(n29447) );
  nand_x1_sg U66861 ( .A(n10907), .B(n25513), .X(n25514) );
  nand_x2_sg U66862 ( .A(n46529), .B(n12316), .X(n12403) );
  nand_x2_sg U66863 ( .A(n12725), .B(n13096), .X(n13183) );
  nand_x2_sg U66864 ( .A(n46462), .B(n14646), .X(n14734) );
  nand_x2_sg U66865 ( .A(n15058), .B(n15429), .X(n15516) );
  nand_x2_sg U66866 ( .A(n16624), .B(n16995), .X(n17082) );
  nand_x2_sg U66867 ( .A(n46372), .B(n17767), .X(n17855) );
  nand_x2_sg U66868 ( .A(n46325), .B(n19312), .X(n19400) );
  nand_x2_sg U66869 ( .A(n46280), .B(n20856), .X(n20944) );
  nand_x2_sg U66870 ( .A(n26089), .B(n26088), .X(n26086) );
  nor_x1_sg U66871 ( .A(n26088), .B(n26089), .X(n26087) );
  nand_x2_sg U66872 ( .A(n26368), .B(n26367), .X(n26365) );
  nor_x1_sg U66873 ( .A(n26367), .B(n26368), .X(n26366) );
  nand_x2_sg U66874 ( .A(n26646), .B(n26645), .X(n26643) );
  nor_x1_sg U66875 ( .A(n26645), .B(n26646), .X(n26644) );
  nand_x2_sg U66876 ( .A(n26925), .B(n26924), .X(n26922) );
  nor_x1_sg U66877 ( .A(n26924), .B(n26925), .X(n26923) );
  nand_x2_sg U66878 ( .A(n27205), .B(n27204), .X(n27202) );
  nor_x1_sg U66879 ( .A(n27204), .B(n27205), .X(n27203) );
  nand_x2_sg U66880 ( .A(n27763), .B(n27762), .X(n27760) );
  nor_x1_sg U66881 ( .A(n27762), .B(n27763), .X(n27761) );
  nand_x2_sg U66882 ( .A(n28044), .B(n28043), .X(n28041) );
  nor_x1_sg U66883 ( .A(n28043), .B(n28044), .X(n28042) );
  nand_x2_sg U66884 ( .A(n28602), .B(n28601), .X(n28599) );
  nor_x1_sg U66885 ( .A(n28601), .B(n28602), .X(n28600) );
  nand_x2_sg U66886 ( .A(n28894), .B(n28893), .X(n28891) );
  nor_x1_sg U66887 ( .A(n28893), .B(n28894), .X(n28892) );
  nand_x2_sg U66888 ( .A(n29163), .B(n29162), .X(n29160) );
  nor_x1_sg U66889 ( .A(n29162), .B(n29163), .X(n29161) );
  nand_x2_sg U66890 ( .A(n29455), .B(n29454), .X(n29452) );
  nor_x1_sg U66891 ( .A(n29454), .B(n29455), .X(n29453) );
  nand_x2_sg U66892 ( .A(n11164), .B(n11535), .X(n11622) );
  nand_x2_sg U66893 ( .A(n46417), .B(n16211), .X(n16298) );
  nand_x2_sg U66894 ( .A(n46305), .B(n20080), .X(n20168) );
  nand_x2_sg U66895 ( .A(n46260), .B(n21625), .X(n21713) );
  nand_x2_sg U66896 ( .A(n14025), .B(n14026), .X(n14024) );
  nand_x1_sg U66897 ( .A(n14029), .B(n14030), .X(n14025) );
  nand_x2_sg U66898 ( .A(n18687), .B(n18688), .X(n18686) );
  nand_x1_sg U66899 ( .A(n18691), .B(n18692), .X(n18687) );
  nand_x2_sg U66900 ( .A(n17496), .B(n17522), .X(n17521) );
  nand_x1_sg U66901 ( .A(n17523), .B(n53808), .X(n17522) );
  nor_x1_sg U66902 ( .A(n46373), .B(n17524), .X(n17523) );
  nand_x2_sg U66903 ( .A(n19041), .B(n19067), .X(n19066) );
  nand_x1_sg U66904 ( .A(n19068), .B(n54373), .X(n19067) );
  nor_x1_sg U66905 ( .A(n46326), .B(n19069), .X(n19068) );
  nand_x2_sg U66906 ( .A(n20585), .B(n20611), .X(n20610) );
  nand_x1_sg U66907 ( .A(n20612), .B(n54941), .X(n20611) );
  nor_x1_sg U66908 ( .A(n46281), .B(n20613), .X(n20612) );
  nand_x2_sg U66909 ( .A(n14797), .B(n14798), .X(n14796) );
  nand_x1_sg U66910 ( .A(n14801), .B(n14802), .X(n14797) );
  nand_x2_sg U66911 ( .A(n20233), .B(n20234), .X(n20232) );
  nand_x1_sg U66912 ( .A(n20237), .B(n20238), .X(n20233) );
  nand_x2_sg U66913 ( .A(n21778), .B(n21779), .X(n21777) );
  nand_x1_sg U66914 ( .A(n21782), .B(n21783), .X(n21778) );
  nand_x1_sg U66915 ( .A(n16363), .B(n16364), .X(n16359) );
  nand_x2_sg U66916 ( .A(n12464), .B(n12465), .X(n12463) );
  nand_x1_sg U66917 ( .A(n12468), .B(n12469), .X(n12464) );
  nand_x2_sg U66918 ( .A(n46352), .B(n18535), .X(n18622) );
  nand_x1_sg U66919 ( .A(n10908), .B(n10909), .X(n10904) );
  nand_x1_sg U66920 ( .A(n10906), .B(n10907), .X(n10905) );
  nand_x2_sg U66921 ( .A(n11685), .B(n11686), .X(n11684) );
  nand_x1_sg U66922 ( .A(n11689), .B(n11690), .X(n11685) );
  nand_x2_sg U66923 ( .A(n13245), .B(n13246), .X(n13244) );
  nand_x1_sg U66924 ( .A(n13249), .B(n13250), .X(n13245) );
  nand_x2_sg U66925 ( .A(n15578), .B(n15579), .X(n15577) );
  nand_x1_sg U66926 ( .A(n15582), .B(n15583), .X(n15578) );
  nand_x2_sg U66927 ( .A(n17144), .B(n17145), .X(n17143) );
  nand_x1_sg U66928 ( .A(n17148), .B(n17149), .X(n17144) );
  nand_x2_sg U66929 ( .A(n17918), .B(n17919), .X(n17917) );
  nand_x1_sg U66930 ( .A(n17922), .B(n17923), .X(n17918) );
  nand_x2_sg U66931 ( .A(n19463), .B(n19464), .X(n19462) );
  nand_x1_sg U66932 ( .A(n19467), .B(n19468), .X(n19463) );
  nand_x2_sg U66933 ( .A(n21007), .B(n21008), .X(n21006) );
  nand_x1_sg U66934 ( .A(n21011), .B(n21012), .X(n21007) );
  nand_x4_sg U66935 ( .A(n53282), .B(n46417), .X(n16020) );
  nand_x2_sg U66936 ( .A(n13589), .B(n13628), .X(n13627) );
  nand_x1_sg U66937 ( .A(n13629), .B(n13630), .X(n13628) );
  nor_x1_sg U66938 ( .A(n46485), .B(n46467), .X(n13629) );
  nand_x1_sg U66939 ( .A(n13734), .B(n13732), .X(n13728) );
  nor_x1_sg U66940 ( .A(n46485), .B(n13735), .X(n13734) );
  nand_x4_sg U66941 ( .A(n51819), .B(n46529), .X(n11837) );
  nand_x4_sg U66942 ( .A(n53207), .B(n46417), .X(n15732) );
  nand_x4_sg U66943 ( .A(n54124), .B(n46352), .X(n18305) );
  nand_x2_sg U66944 ( .A(n26840), .B(n46235), .X(n26835) );
  nand_x2_sg U66945 ( .A(n26837), .B(n52918), .X(n26836) );
  nand_x2_sg U66946 ( .A(n27959), .B(n46235), .X(n27954) );
  nand_x2_sg U66947 ( .A(n27956), .B(n54038), .X(n27955) );
  nand_x2_sg U66948 ( .A(n28517), .B(n46235), .X(n28512) );
  nand_x2_sg U66949 ( .A(n28514), .B(n54603), .X(n28513) );
  nand_x2_sg U66950 ( .A(n29076), .B(n46235), .X(n29071) );
  nand_x2_sg U66951 ( .A(n29073), .B(n55171), .X(n29072) );
  nand_x2_sg U66952 ( .A(n25839), .B(n25838), .X(n25836) );
  nor_x1_sg U66953 ( .A(n25838), .B(n25839), .X(n25837) );
  nand_x2_sg U66954 ( .A(n26955), .B(n26954), .X(n26952) );
  nor_x1_sg U66955 ( .A(n26954), .B(n26955), .X(n26953) );
  nand_x2_sg U66956 ( .A(n28074), .B(n28073), .X(n28071) );
  nor_x1_sg U66957 ( .A(n28073), .B(n28074), .X(n28072) );
  nand_x2_sg U66958 ( .A(n28632), .B(n28631), .X(n28629) );
  nor_x1_sg U66959 ( .A(n28631), .B(n28632), .X(n28630) );
  nand_x2_sg U66960 ( .A(n29193), .B(n29192), .X(n29190) );
  nor_x1_sg U66961 ( .A(n29192), .B(n29193), .X(n29191) );
  nand_x2_sg U66962 ( .A(n26374), .B(n26373), .X(n26371) );
  nor_x1_sg U66963 ( .A(n26373), .B(n26374), .X(n26372) );
  nand_x2_sg U66964 ( .A(n26652), .B(n26651), .X(n26649) );
  nor_x1_sg U66965 ( .A(n26651), .B(n26652), .X(n26650) );
  nand_x2_sg U66966 ( .A(n26931), .B(n26930), .X(n26928) );
  nor_x1_sg U66967 ( .A(n26930), .B(n26931), .X(n26929) );
  nand_x2_sg U66968 ( .A(n27211), .B(n27210), .X(n27208) );
  nor_x1_sg U66969 ( .A(n27210), .B(n27211), .X(n27209) );
  nand_x2_sg U66970 ( .A(n27769), .B(n27768), .X(n27766) );
  nor_x1_sg U66971 ( .A(n27768), .B(n27769), .X(n27767) );
  nand_x2_sg U66972 ( .A(n28050), .B(n28049), .X(n28047) );
  nor_x1_sg U66973 ( .A(n28049), .B(n28050), .X(n28048) );
  nand_x2_sg U66974 ( .A(n28331), .B(n28330), .X(n28328) );
  nor_x1_sg U66975 ( .A(n28330), .B(n28331), .X(n28329) );
  nand_x2_sg U66976 ( .A(n28608), .B(n28607), .X(n28605) );
  nor_x1_sg U66977 ( .A(n28607), .B(n28608), .X(n28606) );
  nand_x2_sg U66978 ( .A(n29169), .B(n29168), .X(n29166) );
  nor_x1_sg U66979 ( .A(n29168), .B(n29169), .X(n29167) );
  nand_x2_sg U66980 ( .A(n26398), .B(n26397), .X(n26395) );
  nor_x1_sg U66981 ( .A(n26397), .B(n26398), .X(n26396) );
  nand_x2_sg U66982 ( .A(n27235), .B(n27234), .X(n27232) );
  nor_x1_sg U66983 ( .A(n27234), .B(n27235), .X(n27233) );
  nand_x2_sg U66984 ( .A(n27793), .B(n27792), .X(n27790) );
  nor_x1_sg U66985 ( .A(n27792), .B(n27793), .X(n27791) );
  nand_x2_sg U66986 ( .A(n25617), .B(n25616), .X(n25614) );
  nor_x1_sg U66987 ( .A(n25616), .B(n25617), .X(n25615) );
  nand_x2_sg U66988 ( .A(n25898), .B(n25897), .X(n25895) );
  nor_x1_sg U66989 ( .A(n25897), .B(n25898), .X(n25896) );
  nand_x2_sg U66990 ( .A(n26178), .B(n26177), .X(n26175) );
  nor_x1_sg U66991 ( .A(n26177), .B(n26178), .X(n26176) );
  nand_x2_sg U66992 ( .A(n26457), .B(n26456), .X(n26454) );
  nor_x1_sg U66993 ( .A(n26456), .B(n26457), .X(n26455) );
  nand_x2_sg U66994 ( .A(n26735), .B(n26734), .X(n26732) );
  nor_x1_sg U66995 ( .A(n26734), .B(n26735), .X(n26733) );
  nand_x2_sg U66996 ( .A(n27014), .B(n27013), .X(n27011) );
  nor_x1_sg U66997 ( .A(n27013), .B(n27014), .X(n27012) );
  nand_x2_sg U66998 ( .A(n27294), .B(n27293), .X(n27291) );
  nor_x1_sg U66999 ( .A(n27293), .B(n27294), .X(n27292) );
  nand_x2_sg U67000 ( .A(n27573), .B(n27572), .X(n27570) );
  nor_x1_sg U67001 ( .A(n27572), .B(n27573), .X(n27571) );
  nand_x2_sg U67002 ( .A(n27852), .B(n27851), .X(n27849) );
  nor_x1_sg U67003 ( .A(n27851), .B(n27852), .X(n27850) );
  nand_x2_sg U67004 ( .A(n28133), .B(n28132), .X(n28130) );
  nor_x1_sg U67005 ( .A(n28132), .B(n28133), .X(n28131) );
  nand_x2_sg U67006 ( .A(n28412), .B(n28411), .X(n28409) );
  nor_x1_sg U67007 ( .A(n28411), .B(n28412), .X(n28410) );
  nand_x2_sg U67008 ( .A(n28691), .B(n28690), .X(n28688) );
  nor_x1_sg U67009 ( .A(n28690), .B(n28691), .X(n28689) );
  nand_x2_sg U67010 ( .A(n28969), .B(n28968), .X(n28966) );
  nor_x1_sg U67011 ( .A(n28968), .B(n28969), .X(n28967) );
  nand_x2_sg U67012 ( .A(n29252), .B(n29251), .X(n29249) );
  nor_x1_sg U67013 ( .A(n29251), .B(n29252), .X(n29250) );
  nand_x2_sg U67014 ( .A(n29530), .B(n29529), .X(n29527) );
  nor_x1_sg U67015 ( .A(n29529), .B(n29530), .X(n29528) );
  nand_x2_sg U67016 ( .A(n25809), .B(n25808), .X(n25806) );
  nor_x1_sg U67017 ( .A(n25808), .B(n25809), .X(n25807) );
  nand_x2_sg U67018 ( .A(n27484), .B(n27483), .X(n27481) );
  nor_x1_sg U67019 ( .A(n27483), .B(n27484), .X(n27482) );
  nand_x2_sg U67020 ( .A(n28882), .B(n28881), .X(n28879) );
  nor_x1_sg U67021 ( .A(n28881), .B(n28882), .X(n28880) );
  nand_x2_sg U67022 ( .A(n29443), .B(n29442), .X(n29440) );
  nor_x1_sg U67023 ( .A(n29442), .B(n29443), .X(n29441) );
  nand_x4_sg U67024 ( .A(n55462), .B(n46576), .X(n18836) );
  nand_x4_sg U67025 ( .A(n10951), .B(n46574), .X(n11043) );
  nand_x4_sg U67026 ( .A(n11735), .B(n46551), .X(n11827) );
  nand_x4_sg U67027 ( .A(n14847), .B(n46462), .X(n14939) );
  nand_x4_sg U67028 ( .A(n17968), .B(n46372), .X(n18060) );
  nand_x4_sg U67029 ( .A(n18737), .B(n46352), .X(n18832) );
  nand_x4_sg U67030 ( .A(n19513), .B(n46325), .X(n19605) );
  nand_x4_sg U67031 ( .A(n20283), .B(n46305), .X(n20377) );
  nand_x4_sg U67032 ( .A(n21057), .B(n46280), .X(n21149) );
  nand_x4_sg U67033 ( .A(n21828), .B(n46260), .X(n21922) );
  nor_x1_sg U67034 ( .A(n21937), .B(n9367), .X(n21934) );
  nor_x1_sg U67035 ( .A(n29588), .B(n9367), .X(n29584) );
  nand_x2_sg U67036 ( .A(n16409), .B(n46417), .X(n16504) );
  nand_x2_sg U67037 ( .A(n12515), .B(n46529), .X(n12606) );
  nand_x2_sg U67038 ( .A(n13296), .B(n46507), .X(n13388) );
  nand_x2_sg U67039 ( .A(n15629), .B(n46439), .X(n15721) );
  nand_x2_sg U67040 ( .A(n17195), .B(n46395), .X(n17287) );
  nand_x4_sg U67041 ( .A(n51896), .B(n46529), .X(n12125) );
  nand_x1_sg U67042 ( .A(n12826), .B(n46507), .X(n12825) );
  nand_x1_sg U67043 ( .A(n15159), .B(n46439), .X(n15158) );
  nand_x1_sg U67044 ( .A(n16725), .B(n46395), .X(n16724) );
  nand_x4_sg U67045 ( .A(n51839), .B(n46529), .X(n11977) );
  nand_x4_sg U67046 ( .A(n53227), .B(n46417), .X(n15872) );
  nand_x4_sg U67047 ( .A(n51598), .B(n46551), .X(n11296) );
  nand_x4_sg U67048 ( .A(n51879), .B(n46529), .X(n12076) );
  nand_x4_sg U67049 ( .A(n52156), .B(n46507), .X(n12857) );
  nand_x4_sg U67050 ( .A(n52990), .B(n46439), .X(n15190) );
  nand_x4_sg U67051 ( .A(n53266), .B(n46417), .X(n15971) );
  nand_x4_sg U67052 ( .A(n53548), .B(n46395), .X(n16756) );
  nand_x4_sg U67053 ( .A(n54614), .B(n46305), .X(n19614) );
  nand_x4_sg U67054 ( .A(n55182), .B(n46260), .X(n21159) );
  nand_x2_sg U67055 ( .A(n25524), .B(n25523), .X(n25521) );
  nor_x1_sg U67056 ( .A(n25523), .B(n25524), .X(n25522) );
  nor_x1_sg U67057 ( .A(n46485), .B(n13732), .X(n13731) );
  nand_x2_sg U67058 ( .A(n25530), .B(n25529), .X(n25527) );
  nor_x1_sg U67059 ( .A(n25529), .B(n25530), .X(n25528) );
  nand_x2_sg U67060 ( .A(n28325), .B(n28324), .X(n28322) );
  nor_x1_sg U67061 ( .A(n28324), .B(n28325), .X(n28323) );
  nand_x4_sg U67062 ( .A(n13393), .B(n15725), .X(n14942) );
  nand_x2_sg U67063 ( .A(n11266), .B(n11265), .X(n11262) );
  nor_x1_sg U67064 ( .A(n46552), .B(n11180), .X(n11266) );
  nor_x1_sg U67065 ( .A(n53446), .B(n16357), .X(n16356) );
  nor_x1_sg U67066 ( .A(n52057), .B(n12462), .X(n12461) );
  nor_x1_sg U67067 ( .A(n25238), .B(n49356), .X(n31422) );
  nor_x1_sg U67068 ( .A(n10130), .B(n50215), .X(n23756) );
  nand_x4_sg U67069 ( .A(n16063), .B(n16064), .X(n15999) );
  nand_x1_sg U67070 ( .A(n16066), .B(n16067), .X(n16063) );
  nand_x1_sg U67071 ( .A(n16065), .B(n53298), .X(n16064) );
  nand_x1_sg U67072 ( .A(n53298), .B(n46417), .X(n16067) );
  nand_x4_sg U67073 ( .A(n52670), .B(n46462), .X(n14313) );
  nor_x1_sg U67074 ( .A(n46485), .B(n14029), .X(n14027) );
  nand_x4_sg U67075 ( .A(n54634), .B(n46305), .X(n19748) );
  nand_x4_sg U67076 ( .A(n55202), .B(n46260), .X(n21293) );
  nand_x4_sg U67077 ( .A(n51280), .B(n46574), .X(n10421) );
  nand_x4_sg U67078 ( .A(n54070), .B(n46352), .X(n18201) );
  nor_x1_sg U67079 ( .A(n10518), .B(n10782), .X(n10858) );
  nand_x4_sg U67080 ( .A(n12852), .B(n12853), .X(n12817) );
  nand_x1_sg U67081 ( .A(n12752), .B(n12855), .X(n12852) );
  nand_x1_sg U67082 ( .A(n12854), .B(n12826), .X(n12853) );
  nand_x1_sg U67083 ( .A(n12826), .B(n46503), .X(n12855) );
  nand_x4_sg U67084 ( .A(n15185), .B(n15186), .X(n15150) );
  nand_x1_sg U67085 ( .A(n15085), .B(n15188), .X(n15185) );
  nand_x1_sg U67086 ( .A(n15187), .B(n15159), .X(n15186) );
  nand_x1_sg U67087 ( .A(n15159), .B(n46435), .X(n15188) );
  nand_x4_sg U67088 ( .A(n16751), .B(n16752), .X(n16716) );
  nand_x1_sg U67089 ( .A(n16651), .B(n16754), .X(n16751) );
  nand_x1_sg U67090 ( .A(n16753), .B(n16725), .X(n16752) );
  nand_x1_sg U67091 ( .A(n16725), .B(n46391), .X(n16754) );
  nand_x1_sg U67092 ( .A(n49401), .B(n25189), .X(n31419) );
  nand_x1_sg U67093 ( .A(n50260), .B(n10081), .X(n23753) );
  nand_x1_sg U67094 ( .A(n49822), .B(n24756), .X(n31391) );
  nand_x1_sg U67095 ( .A(n50681), .B(n9648), .X(n23725) );
  nand_x1_sg U67096 ( .A(n50004), .B(n24562), .X(n30515) );
  nand_x1_sg U67097 ( .A(n49916), .B(n24660), .X(n30996) );
  nand_x1_sg U67098 ( .A(n50863), .B(n9454), .X(n22849) );
  nand_x1_sg U67099 ( .A(n50775), .B(n9552), .X(n23330) );
  nand_x4_sg U67100 ( .A(n17871), .B(n53838), .X(n17828) );
  nor_x1_sg U67101 ( .A(n17596), .B(n17795), .X(n17871) );
  nand_x4_sg U67102 ( .A(n19416), .B(n54403), .X(n19373) );
  nor_x1_sg U67103 ( .A(n19141), .B(n19340), .X(n19416) );
  nand_x4_sg U67104 ( .A(n20960), .B(n54971), .X(n20917) );
  nor_x1_sg U67105 ( .A(n20685), .B(n20884), .X(n20960) );
  nand_x2_sg U67106 ( .A(n21972), .B(n50966), .X(n21971) );
  nand_x2_sg U67107 ( .A(n29637), .B(n50107), .X(n29636) );
  nand_x4_sg U67108 ( .A(n46539), .B(n46551), .X(n11198) );
  nand_x4_sg U67109 ( .A(n46495), .B(n46507), .X(n12759) );
  nand_x4_sg U67110 ( .A(n46427), .B(n46439), .X(n15092) );
  nand_x4_sg U67111 ( .A(n46383), .B(n46395), .X(n16658) );
  nand_x4_sg U67112 ( .A(n46532), .B(n46551), .X(n11345) );
  nand_x4_sg U67113 ( .A(n46488), .B(n46507), .X(n12906) );
  nand_x4_sg U67114 ( .A(n46420), .B(n46439), .X(n15239) );
  nand_x4_sg U67115 ( .A(n46376), .B(n46395), .X(n16805) );
  nand_x4_sg U67116 ( .A(n29141), .B(n46235), .X(n29140) );
  nor_x1_sg U67117 ( .A(n29142), .B(n29143), .X(n29141) );
  nand_x4_sg U67118 ( .A(n46480), .B(n46485), .X(n26518) );
  nand_x4_sg U67119 ( .A(n46360), .B(n46372), .X(n17435) );
  nand_x4_sg U67120 ( .A(n46313), .B(n46325), .X(n18980) );
  nand_x4_sg U67121 ( .A(n46268), .B(n46280), .X(n20524) );
  nand_x2_sg U67122 ( .A(n29437), .B(n29436), .X(n29434) );
  nor_x1_sg U67123 ( .A(n29436), .B(n29437), .X(n29435) );
  nand_x2_sg U67124 ( .A(n25803), .B(n25802), .X(n25800) );
  nor_x1_sg U67125 ( .A(n25802), .B(n25803), .X(n25801) );
  nand_x2_sg U67126 ( .A(n26919), .B(n26918), .X(n26916) );
  nor_x1_sg U67127 ( .A(n26918), .B(n26919), .X(n26917) );
  nand_x2_sg U67128 ( .A(n27478), .B(n27477), .X(n27475) );
  nor_x1_sg U67129 ( .A(n27477), .B(n27478), .X(n27476) );
  nand_x2_sg U67130 ( .A(n28038), .B(n28037), .X(n28035) );
  nor_x1_sg U67131 ( .A(n28037), .B(n28038), .X(n28036) );
  nand_x2_sg U67132 ( .A(n28319), .B(n28318), .X(n28316) );
  nor_x1_sg U67133 ( .A(n28318), .B(n28319), .X(n28317) );
  nand_x2_sg U67134 ( .A(n28596), .B(n28595), .X(n28593) );
  nor_x1_sg U67135 ( .A(n28595), .B(n28596), .X(n28594) );
  nand_x2_sg U67136 ( .A(n28876), .B(n28875), .X(n28873) );
  nor_x1_sg U67137 ( .A(n28875), .B(n28876), .X(n28874) );
  nand_x2_sg U67138 ( .A(n29157), .B(n29156), .X(n29154) );
  nor_x1_sg U67139 ( .A(n29156), .B(n29157), .X(n29155) );
  nor_x1_sg U67140 ( .A(n46236), .B(n25666), .X(\L1_0/n4667 ) );
  nand_x2_sg U67141 ( .A(n25667), .B(n46551), .X(n25666) );
  nor_x1_sg U67142 ( .A(n46236), .B(n26782), .X(\L1_0/n4347 ) );
  nand_x2_sg U67143 ( .A(n26783), .B(n14295), .X(n26782) );
  nor_x1_sg U67144 ( .A(n46236), .B(n27341), .X(\L1_0/n4187 ) );
  nand_x2_sg U67145 ( .A(n27342), .B(n46417), .X(n27341) );
  nor_x1_sg U67146 ( .A(n46236), .B(n27621), .X(\L1_0/n4107 ) );
  nand_x2_sg U67147 ( .A(n27622), .B(n46395), .X(n27621) );
  nor_x1_sg U67148 ( .A(n46236), .B(n28738), .X(\L1_0/n3787 ) );
  nand_x2_sg U67149 ( .A(n28739), .B(n46305), .X(n28738) );
  nand_x4_sg U67150 ( .A(n46576), .B(n32137), .X(n25667) );
  nand_x4_sg U67151 ( .A(n46576), .B(n27620), .X(n27342) );
  nor_x1_sg U67152 ( .A(n10231), .B(n9355), .X(\L2_0/n4148 ) );
  nand_x4_sg U67153 ( .A(n11291), .B(n11292), .X(n11256) );
  nand_x1_sg U67154 ( .A(n11191), .B(n11294), .X(n11291) );
  nor_x1_sg U67155 ( .A(n11191), .B(n46546), .X(n11293) );
  nor_x1_sg U67156 ( .A(n26357), .B(n46585), .X(\L1_0/n4430 ) );
  nand_x2_sg U67157 ( .A(n46235), .B(n26353), .X(n26359) );
  nor_x1_sg U67158 ( .A(n26636), .B(n46587), .X(\L1_0/n4350 ) );
  nand_x2_sg U67159 ( .A(n46235), .B(n26632), .X(n26637) );
  nor_x1_sg U67160 ( .A(n28032), .B(n46591), .X(\L1_0/n3950 ) );
  nand_x2_sg U67161 ( .A(n46235), .B(n28028), .X(n28033) );
  nor_x1_sg U67162 ( .A(n28590), .B(n28459), .X(\L1_0/n3790 ) );
  nand_x2_sg U67163 ( .A(n46235), .B(n28586), .X(n28591) );
  nor_x1_sg U67164 ( .A(n29431), .B(n46596), .X(\L1_0/n3550 ) );
  nand_x2_sg U67165 ( .A(n46235), .B(n29427), .X(n29432) );
  nand_x4_sg U67166 ( .A(n29593), .B(n15726), .X(n29589) );
  nor_x1_sg U67167 ( .A(n27193), .B(n46589), .X(\L1_0/n4190 ) );
  nand_x2_sg U67168 ( .A(n46235), .B(n27189), .X(n27196) );
  nor_x1_sg U67169 ( .A(n28312), .B(n46593), .X(\L1_0/n3870 ) );
  nand_x2_sg U67170 ( .A(n46235), .B(n28308), .X(n28314) );
  nor_x1_sg U67171 ( .A(n46616), .B(n29019), .X(\L1_0/n3707 ) );
  nand_x2_sg U67172 ( .A(n46235), .B(n46280), .X(n29019) );
  nor_x1_sg U67173 ( .A(n46612), .B(n25945), .X(\L1_0/n4587 ) );
  nand_x2_sg U67174 ( .A(n46235), .B(n46529), .X(n25945) );
  inv_x4_sg U67175 ( .A(n46606), .X(n46605) );
  nor_x1_sg U67176 ( .A(n25339), .B(n46233), .X(\L1_0/n4751 ) );
  nand_x4_sg U67177 ( .A(n25511), .B(n46235), .X(n25510) );
  nor_x1_sg U67178 ( .A(n51525), .B(n25512), .X(n25511) );
  nand_x4_sg U67179 ( .A(n25789), .B(n46235), .X(n25788) );
  nor_x1_sg U67180 ( .A(n25790), .B(n25791), .X(n25789) );
  nand_x4_sg U67181 ( .A(n26068), .B(n46235), .X(n26067) );
  nor_x1_sg U67182 ( .A(n26069), .B(n26070), .X(n26068) );
  nand_x4_sg U67183 ( .A(n26349), .B(n46235), .X(n26348) );
  nor_x1_sg U67184 ( .A(n26350), .B(n26351), .X(n26349) );
  nand_x4_sg U67185 ( .A(n27185), .B(n46235), .X(n27184) );
  nor_x1_sg U67186 ( .A(n27186), .B(n27187), .X(n27185) );
  nand_x4_sg U67187 ( .A(n27464), .B(n46235), .X(n27463) );
  nor_x1_sg U67188 ( .A(n27465), .B(n27466), .X(n27464) );
  nand_x4_sg U67189 ( .A(n27745), .B(n46235), .X(n27744) );
  nor_x1_sg U67190 ( .A(n27746), .B(n27747), .X(n27745) );
  nand_x4_sg U67191 ( .A(n28024), .B(n46235), .X(n28023) );
  nor_x1_sg U67192 ( .A(n28025), .B(n28026), .X(n28024) );
  nand_x4_sg U67193 ( .A(n28304), .B(n46235), .X(n28303) );
  nor_x1_sg U67194 ( .A(n28305), .B(n28306), .X(n28304) );
  nand_x4_sg U67195 ( .A(n28582), .B(n46235), .X(n28581) );
  nor_x1_sg U67196 ( .A(n28583), .B(n28584), .X(n28582) );
  nand_x4_sg U67197 ( .A(n28862), .B(n46235), .X(n28861) );
  nor_x1_sg U67198 ( .A(n28863), .B(n28864), .X(n28862) );
  nand_x4_sg U67199 ( .A(n29423), .B(n46235), .X(n29422) );
  nor_x1_sg U67200 ( .A(n29424), .B(n29425), .X(n29423) );
  nor_x1_sg U67201 ( .A(n46519), .B(n12030), .X(n12029) );
  nor_x1_sg U67202 ( .A(n46407), .B(n15925), .X(n15924) );
  nand_x4_sg U67203 ( .A(n26905), .B(n46235), .X(n26904) );
  nor_x1_sg U67204 ( .A(n26906), .B(n26907), .X(n26905) );
  nand_x4_sg U67205 ( .A(n12168), .B(n12169), .X(n12104) );
  nand_x1_sg U67206 ( .A(n12171), .B(n12172), .X(n12168) );
  nand_x4_sg U67207 ( .A(n26628), .B(n46235), .X(n26627) );
  nor_x1_sg U67208 ( .A(n26629), .B(n26630), .X(n26628) );
  nor_x1_sg U67209 ( .A(n46485), .B(n46483), .X(\L2_0/n3824 ) );
  nor_x1_sg U67210 ( .A(n14411), .B(n26839), .X(n26838) );
  nand_x2_sg U67211 ( .A(n46222), .B(n26830), .X(n26839) );
  nor_x1_sg U67212 ( .A(n17524), .B(n27958), .X(n27957) );
  nand_x2_sg U67213 ( .A(n46214), .B(n27949), .X(n27958) );
  nor_x1_sg U67214 ( .A(n19069), .B(n28516), .X(n28515) );
  nand_x2_sg U67215 ( .A(n46210), .B(n28507), .X(n28516) );
  nor_x1_sg U67216 ( .A(n20613), .B(n29075), .X(n29074) );
  nand_x2_sg U67217 ( .A(n46206), .B(n29066), .X(n29075) );
  nor_x1_sg U67218 ( .A(n25541), .B(n25542), .X(n25540) );
  nor_x1_sg U67219 ( .A(n46615), .B(n25340), .X(n25343) );
  nand_x4_sg U67220 ( .A(n9951), .B(n9952), .X(n9948) );
  nor_x1_sg U67221 ( .A(n9953), .B(n9954), .X(n9952) );
  nor_x1_sg U67222 ( .A(n9957), .B(n9958), .X(n9951) );
  nand_x4_sg U67223 ( .A(n10048), .B(n10049), .X(n10045) );
  nor_x1_sg U67224 ( .A(n10050), .B(n10051), .X(n10049) );
  nor_x1_sg U67225 ( .A(n10054), .B(n10055), .X(n10048) );
  nand_x4_sg U67226 ( .A(n10097), .B(n10098), .X(n10094) );
  nor_x1_sg U67227 ( .A(n10099), .B(n10100), .X(n10098) );
  nor_x1_sg U67228 ( .A(n10103), .B(n10104), .X(n10097) );
  nand_x4_sg U67229 ( .A(n25059), .B(n25060), .X(n25056) );
  nor_x1_sg U67230 ( .A(n25065), .B(n25066), .X(n25059) );
  nor_x1_sg U67231 ( .A(n25061), .B(n25062), .X(n25060) );
  nand_x4_sg U67232 ( .A(n25156), .B(n25157), .X(n25153) );
  nor_x1_sg U67233 ( .A(n25162), .B(n25163), .X(n25156) );
  nor_x1_sg U67234 ( .A(n25158), .B(n25159), .X(n25157) );
  nand_x4_sg U67235 ( .A(n25205), .B(n25206), .X(n25202) );
  nor_x1_sg U67236 ( .A(n25211), .B(n25212), .X(n25205) );
  nor_x1_sg U67237 ( .A(n25207), .B(n25208), .X(n25206) );
  nand_x4_sg U67238 ( .A(n9360), .B(n9361), .X(n9357) );
  nor_x1_sg U67239 ( .A(n9362), .B(n9363), .X(n9361) );
  nor_x1_sg U67240 ( .A(n9368), .B(n9369), .X(n9360) );
  nand_x4_sg U67241 ( .A(n24479), .B(n24480), .X(n24475) );
  nor_x1_sg U67242 ( .A(n24485), .B(n24486), .X(n24479) );
  nor_x1_sg U67243 ( .A(n24481), .B(n24482), .X(n24480) );
  nand_x4_sg U67244 ( .A(n9807), .B(n9808), .X(n9804) );
  nor_x1_sg U67245 ( .A(n9813), .B(n9814), .X(n9807) );
  nor_x1_sg U67246 ( .A(n9809), .B(n9810), .X(n9808) );
  nand_x4_sg U67247 ( .A(n9855), .B(n9856), .X(n9852) );
  nor_x1_sg U67248 ( .A(n9861), .B(n9862), .X(n9855) );
  nor_x1_sg U67249 ( .A(n9857), .B(n9858), .X(n9856) );
  nand_x4_sg U67250 ( .A(n9903), .B(n9904), .X(n9900) );
  nor_x1_sg U67251 ( .A(n9909), .B(n9910), .X(n9903) );
  nor_x1_sg U67252 ( .A(n9905), .B(n9906), .X(n9904) );
  nand_x4_sg U67253 ( .A(n10000), .B(n10001), .X(n9997) );
  nor_x1_sg U67254 ( .A(n10006), .B(n10007), .X(n10000) );
  nor_x1_sg U67255 ( .A(n10002), .B(n10003), .X(n10001) );
  nand_x4_sg U67256 ( .A(n10146), .B(n10147), .X(n10143) );
  nor_x1_sg U67257 ( .A(n10152), .B(n10153), .X(n10146) );
  nor_x1_sg U67258 ( .A(n10148), .B(n10149), .X(n10147) );
  nand_x4_sg U67259 ( .A(n24915), .B(n24916), .X(n24912) );
  nor_x1_sg U67260 ( .A(n24921), .B(n24922), .X(n24915) );
  nor_x1_sg U67261 ( .A(n24917), .B(n24918), .X(n24916) );
  nand_x4_sg U67262 ( .A(n24963), .B(n24964), .X(n24960) );
  nor_x1_sg U67263 ( .A(n24969), .B(n24970), .X(n24963) );
  nor_x1_sg U67264 ( .A(n24965), .B(n24966), .X(n24964) );
  nand_x4_sg U67265 ( .A(n25011), .B(n25012), .X(n25008) );
  nor_x1_sg U67266 ( .A(n25017), .B(n25018), .X(n25011) );
  nor_x1_sg U67267 ( .A(n25013), .B(n25014), .X(n25012) );
  nand_x4_sg U67268 ( .A(n25108), .B(n25109), .X(n25105) );
  nor_x1_sg U67269 ( .A(n25114), .B(n25115), .X(n25108) );
  nor_x1_sg U67270 ( .A(n25110), .B(n25111), .X(n25109) );
  nand_x4_sg U67271 ( .A(n25254), .B(n25255), .X(n25251) );
  nor_x1_sg U67272 ( .A(n25260), .B(n25261), .X(n25254) );
  nor_x1_sg U67273 ( .A(n25256), .B(n25257), .X(n25255) );
  nand_x4_sg U67274 ( .A(n9421), .B(n9422), .X(n9418) );
  nor_x1_sg U67275 ( .A(n9423), .B(n9424), .X(n9422) );
  nor_x1_sg U67276 ( .A(n9427), .B(n9428), .X(n9421) );
  nand_x4_sg U67277 ( .A(n9470), .B(n9471), .X(n9467) );
  nor_x1_sg U67278 ( .A(n9472), .B(n9473), .X(n9471) );
  nor_x1_sg U67279 ( .A(n9476), .B(n9477), .X(n9470) );
  nand_x4_sg U67280 ( .A(n9519), .B(n9520), .X(n9516) );
  nor_x1_sg U67281 ( .A(n9521), .B(n9522), .X(n9520) );
  nor_x1_sg U67282 ( .A(n9525), .B(n9526), .X(n9519) );
  nand_x4_sg U67283 ( .A(n9568), .B(n9569), .X(n9565) );
  nor_x1_sg U67284 ( .A(n9570), .B(n9571), .X(n9569) );
  nor_x1_sg U67285 ( .A(n9574), .B(n9575), .X(n9568) );
  nand_x4_sg U67286 ( .A(n9616), .B(n9617), .X(n9613) );
  nor_x1_sg U67287 ( .A(n9618), .B(n9619), .X(n9617) );
  nor_x1_sg U67288 ( .A(n9622), .B(n9623), .X(n9616) );
  nand_x4_sg U67289 ( .A(n9664), .B(n9665), .X(n9661) );
  nor_x1_sg U67290 ( .A(n9666), .B(n9667), .X(n9665) );
  nor_x1_sg U67291 ( .A(n9670), .B(n9671), .X(n9664) );
  nand_x4_sg U67292 ( .A(n9711), .B(n9712), .X(n9708) );
  nor_x1_sg U67293 ( .A(n9713), .B(n9714), .X(n9712) );
  nor_x1_sg U67294 ( .A(n9717), .B(n9718), .X(n9711) );
  nand_x4_sg U67295 ( .A(n9759), .B(n9760), .X(n9756) );
  nor_x1_sg U67296 ( .A(n9761), .B(n9762), .X(n9760) );
  nor_x1_sg U67297 ( .A(n9765), .B(n9766), .X(n9759) );
  nand_x4_sg U67298 ( .A(n24529), .B(n24530), .X(n24526) );
  nor_x1_sg U67299 ( .A(n24535), .B(n24536), .X(n24529) );
  nor_x1_sg U67300 ( .A(n24531), .B(n24532), .X(n24530) );
  nand_x4_sg U67301 ( .A(n24578), .B(n24579), .X(n24575) );
  nor_x1_sg U67302 ( .A(n24584), .B(n24585), .X(n24578) );
  nor_x1_sg U67303 ( .A(n24580), .B(n24581), .X(n24579) );
  nand_x4_sg U67304 ( .A(n24627), .B(n24628), .X(n24624) );
  nor_x1_sg U67305 ( .A(n24633), .B(n24634), .X(n24627) );
  nor_x1_sg U67306 ( .A(n24629), .B(n24630), .X(n24628) );
  nand_x4_sg U67307 ( .A(n24676), .B(n24677), .X(n24673) );
  nor_x1_sg U67308 ( .A(n24682), .B(n24683), .X(n24676) );
  nor_x1_sg U67309 ( .A(n24678), .B(n24679), .X(n24677) );
  nand_x4_sg U67310 ( .A(n24724), .B(n24725), .X(n24721) );
  nor_x1_sg U67311 ( .A(n24730), .B(n24731), .X(n24724) );
  nor_x1_sg U67312 ( .A(n24726), .B(n24727), .X(n24725) );
  nand_x4_sg U67313 ( .A(n24772), .B(n24773), .X(n24769) );
  nor_x1_sg U67314 ( .A(n24778), .B(n24779), .X(n24772) );
  nor_x1_sg U67315 ( .A(n24774), .B(n24775), .X(n24773) );
  nand_x4_sg U67316 ( .A(n24819), .B(n24820), .X(n24816) );
  nor_x1_sg U67317 ( .A(n24825), .B(n24826), .X(n24819) );
  nor_x1_sg U67318 ( .A(n24821), .B(n24822), .X(n24820) );
  nand_x4_sg U67319 ( .A(n24867), .B(n24868), .X(n24864) );
  nor_x1_sg U67320 ( .A(n24873), .B(n24874), .X(n24867) );
  nor_x1_sg U67321 ( .A(n24869), .B(n24870), .X(n24868) );
  nand_x4_sg U67322 ( .A(n25552), .B(n25551), .X(n11039) );
  nand_x4_sg U67323 ( .A(n28347), .B(n28346), .X(n18826) );
  nand_x4_sg U67324 ( .A(n28904), .B(n28903), .X(n20371) );
  nand_x4_sg U67325 ( .A(n29465), .B(n29464), .X(n21916) );
  nand_x4_sg U67326 ( .A(n25611), .B(n25610), .X(n11045) );
  nand_x4_sg U67327 ( .A(n27567), .B(n27566), .X(n16506) );
  nand_x4_sg U67328 ( .A(n25892), .B(n25891), .X(n11829) );
  nand_x4_sg U67329 ( .A(n26172), .B(n26171), .X(n12608) );
  nand_x4_sg U67330 ( .A(n26083), .B(n26082), .X(n12603) );
  nand_x4_sg U67331 ( .A(n26451), .B(n26450), .X(n13390) );
  nand_x4_sg U67332 ( .A(n26362), .B(n26361), .X(n13385) );
  nand_x4_sg U67333 ( .A(n26729), .B(n26728), .X(n14170) );
  nand_x4_sg U67334 ( .A(n26640), .B(n26639), .X(n14165) );
  nand_x4_sg U67335 ( .A(n27008), .B(n27007), .X(n14941) );
  nand_x4_sg U67336 ( .A(n27288), .B(n27287), .X(n15723) );
  nand_x4_sg U67337 ( .A(n27199), .B(n27198), .X(n15718) );
  nand_x4_sg U67338 ( .A(n27846), .B(n27845), .X(n17289) );
  nand_x4_sg U67339 ( .A(n27757), .B(n27756), .X(n17284) );
  nand_x4_sg U67340 ( .A(n28127), .B(n28126), .X(n18062) );
  nand_x4_sg U67341 ( .A(n28406), .B(n28405), .X(n18834) );
  nand_x4_sg U67342 ( .A(n28685), .B(n28684), .X(n19607) );
  nand_x4_sg U67343 ( .A(n28963), .B(n28962), .X(n20379) );
  nand_x4_sg U67344 ( .A(n29246), .B(n29245), .X(n21151) );
  nand_x4_sg U67345 ( .A(n29524), .B(n29523), .X(n21924) );
  nand_x4_sg U67346 ( .A(n10246), .B(n10247), .X(n10232) );
  nor_x1_sg U67347 ( .A(n10268), .B(n10269), .X(n10246) );
  nor_x1_sg U67348 ( .A(n10248), .B(n10249), .X(n10247) );
  nand_x2_sg U67349 ( .A(n10270), .B(n10271), .X(n10269) );
  nand_x4_sg U67350 ( .A(n25354), .B(n25355), .X(n25340) );
  nor_x1_sg U67351 ( .A(n25374), .B(n25375), .X(n25354) );
  nor_x1_sg U67352 ( .A(n25356), .B(n25357), .X(n25355) );
  nand_x2_sg U67353 ( .A(n25376), .B(n25377), .X(n25375) );
  nand_x4_sg U67354 ( .A(n21932), .B(n21933), .X(n21929) );
  nor_x1_sg U67355 ( .A(n21938), .B(n21939), .X(n21932) );
  nor_x1_sg U67356 ( .A(n40882), .B(n21935), .X(n21933) );
  nand_x4_sg U67357 ( .A(n29582), .B(n29583), .X(n29579) );
  nor_x1_sg U67358 ( .A(n29590), .B(n29591), .X(n29582) );
  nor_x1_sg U67359 ( .A(n40884), .B(n29585), .X(n29583) );
  nand_x4_sg U67360 ( .A(n10193), .B(n10194), .X(n10190) );
  nor_x1_sg U67361 ( .A(n10195), .B(n10196), .X(n10194) );
  nor_x1_sg U67362 ( .A(n10198), .B(n10199), .X(n10193) );
  nand_x4_sg U67363 ( .A(n25301), .B(n25302), .X(n25298) );
  nor_x1_sg U67364 ( .A(n25305), .B(n25306), .X(n25301) );
  nor_x1_sg U67365 ( .A(n25303), .B(n25304), .X(n25302) );
  nand_x1_sg U67366 ( .A(n25519), .B(n25508), .X(n25518) );
  nor_x1_sg U67367 ( .A(n10907), .B(n46231), .X(n25519) );
  nor_x1_sg U67368 ( .A(n46575), .B(n10232), .X(n10235) );
  nor_x1_sg U67369 ( .A(n55782), .B(n25515), .X(\L1_0/n4671 ) );
  nor_x1_sg U67370 ( .A(n46234), .B(n10907), .X(n25516) );
  nor_x1_sg U67371 ( .A(n29146), .B(n29147), .X(\L1_0/n3631 ) );
  nor_x1_sg U67372 ( .A(n55167), .B(n46236), .X(n29148) );
  nor_x1_sg U67373 ( .A(n46611), .B(n25797), .X(\L1_0/n4590 ) );
  nand_x2_sg U67374 ( .A(n46235), .B(n25793), .X(n25798) );
  nand_x2_sg U67375 ( .A(n9401), .B(n9402), .X(n9395) );
  nor_x1_sg U67376 ( .A(n9404), .B(n9405), .X(n9401) );
  nand_x1_sg U67377 ( .A(n46600), .B(n50925), .X(n9402) );
  nand_x2_sg U67378 ( .A(n9694), .B(n9695), .X(n9690) );
  nor_x1_sg U67379 ( .A(n9696), .B(n9697), .X(n9694) );
  nand_x1_sg U67380 ( .A(n46600), .B(n50655), .X(n9695) );
  nand_x2_sg U67381 ( .A(n24512), .B(n24513), .X(n24507) );
  nor_x1_sg U67382 ( .A(n24514), .B(n24515), .X(n24512) );
  nand_x1_sg U67383 ( .A(n46600), .B(n50066), .X(n24513) );
  nand_x2_sg U67384 ( .A(n24802), .B(n24803), .X(n24798) );
  nor_x1_sg U67385 ( .A(n24804), .B(n24805), .X(n24802) );
  nand_x1_sg U67386 ( .A(n46600), .B(n49796), .X(n24803) );
  nor_x1_sg U67387 ( .A(n28459), .B(n28460), .X(\L1_0/n3867 ) );
  nand_x2_sg U67388 ( .A(n46235), .B(n46325), .X(n28460) );
  nand_x2_sg U67389 ( .A(n9441), .B(n9442), .X(n9433) );
  nor_x1_sg U67390 ( .A(n9444), .B(n9445), .X(n9441) );
  nand_x1_sg U67391 ( .A(n46607), .B(n9443), .X(n9442) );
  nand_x2_sg U67392 ( .A(n9490), .B(n9491), .X(n9482) );
  nor_x1_sg U67393 ( .A(n9493), .B(n9494), .X(n9490) );
  nand_x1_sg U67394 ( .A(n46607), .B(n9492), .X(n9491) );
  nand_x2_sg U67395 ( .A(n9539), .B(n9540), .X(n9531) );
  nor_x1_sg U67396 ( .A(n9542), .B(n9543), .X(n9539) );
  nand_x1_sg U67397 ( .A(n46607), .B(n9541), .X(n9540) );
  nand_x2_sg U67398 ( .A(n24549), .B(n24550), .X(n24541) );
  nor_x1_sg U67399 ( .A(n24552), .B(n24553), .X(n24549) );
  nand_x1_sg U67400 ( .A(n24551), .B(n46607), .X(n24550) );
  nand_x2_sg U67401 ( .A(n24598), .B(n24599), .X(n24590) );
  nor_x1_sg U67402 ( .A(n24601), .B(n24602), .X(n24598) );
  nand_x1_sg U67403 ( .A(n24600), .B(n46607), .X(n24599) );
  nand_x2_sg U67404 ( .A(n24647), .B(n24648), .X(n24639) );
  nor_x1_sg U67405 ( .A(n24650), .B(n24651), .X(n24647) );
  nand_x1_sg U67406 ( .A(n24649), .B(n46607), .X(n24648) );
  nand_x2_sg U67407 ( .A(n10125), .B(n10126), .X(n10124) );
  nand_x1_sg U67408 ( .A(n46598), .B(n50229), .X(n10126) );
  nand_x1_sg U67409 ( .A(n10127), .B(n46608), .X(n10125) );
  nand_x2_sg U67410 ( .A(n25233), .B(n25234), .X(n25232) );
  nand_x1_sg U67411 ( .A(n49370), .B(n46598), .X(n25234) );
  nand_x1_sg U67412 ( .A(n25235), .B(n46608), .X(n25233) );
  nand_x2_sg U67413 ( .A(n10076), .B(n10077), .X(n10075) );
  nand_x1_sg U67414 ( .A(n46598), .B(n50275), .X(n10077) );
  nand_x1_sg U67415 ( .A(n10078), .B(n46608), .X(n10076) );
  nand_x2_sg U67416 ( .A(n25184), .B(n25185), .X(n25183) );
  nand_x1_sg U67417 ( .A(n49416), .B(n46598), .X(n25185) );
  nand_x1_sg U67418 ( .A(n25186), .B(n46608), .X(n25184) );
  nor_x1_sg U67419 ( .A(n26506), .B(n46587), .X(\L1_0/n4426 ) );
  nand_x2_sg U67420 ( .A(n9979), .B(n9980), .X(n9978) );
  nand_x1_sg U67421 ( .A(n46598), .B(n50368), .X(n9980) );
  nand_x1_sg U67422 ( .A(n9981), .B(n46608), .X(n9979) );
  nand_x2_sg U67423 ( .A(n25087), .B(n25088), .X(n25086) );
  nand_x1_sg U67424 ( .A(n49509), .B(n46598), .X(n25088) );
  nand_x1_sg U67425 ( .A(n25089), .B(n46608), .X(n25087) );
  nand_x2_sg U67426 ( .A(n9378), .B(n9379), .X(n9377) );
  nand_x1_sg U67427 ( .A(n46602), .B(n9380), .X(n9379) );
  nor_x1_sg U67428 ( .A(n9381), .B(n9382), .X(n9378) );
  nand_x2_sg U67429 ( .A(n24493), .B(n24494), .X(n24492) );
  nand_x1_sg U67430 ( .A(n24495), .B(n46602), .X(n24494) );
  nor_x1_sg U67431 ( .A(n24496), .B(n24497), .X(n24493) );
  nand_x2_sg U67432 ( .A(n9484), .B(n9485), .X(n9483) );
  nand_x1_sg U67433 ( .A(n46602), .B(n50849), .X(n9485) );
  nor_x1_sg U67434 ( .A(n9486), .B(n9487), .X(n9484) );
  nand_x2_sg U67435 ( .A(n9533), .B(n9534), .X(n9532) );
  nand_x1_sg U67436 ( .A(n46602), .B(n50804), .X(n9534) );
  nor_x1_sg U67437 ( .A(n9535), .B(n9536), .X(n9533) );
  nand_x2_sg U67438 ( .A(n9582), .B(n9583), .X(n9581) );
  nand_x1_sg U67439 ( .A(n46602), .B(n50756), .X(n9583) );
  nor_x1_sg U67440 ( .A(n9584), .B(n9585), .X(n9582) );
  nand_x2_sg U67441 ( .A(n9588), .B(n9589), .X(n9580) );
  nand_x1_sg U67442 ( .A(n46607), .B(n50752), .X(n9589) );
  nor_x1_sg U67443 ( .A(n9590), .B(n9591), .X(n9588) );
  nand_x2_sg U67444 ( .A(n9630), .B(n9631), .X(n9629) );
  nand_x1_sg U67445 ( .A(n46602), .B(n50709), .X(n9631) );
  nor_x1_sg U67446 ( .A(n9632), .B(n9633), .X(n9630) );
  nand_x2_sg U67447 ( .A(n9636), .B(n9637), .X(n9628) );
  nand_x1_sg U67448 ( .A(n46607), .B(n50705), .X(n9637) );
  nor_x1_sg U67449 ( .A(n9638), .B(n9639), .X(n9636) );
  nand_x2_sg U67450 ( .A(n9678), .B(n9679), .X(n9677) );
  nand_x1_sg U67451 ( .A(n46602), .B(n50661), .X(n9679) );
  nor_x1_sg U67452 ( .A(n9680), .B(n9681), .X(n9678) );
  nand_x2_sg U67453 ( .A(n9725), .B(n9726), .X(n9724) );
  nand_x1_sg U67454 ( .A(n46602), .B(n50614), .X(n9726) );
  nor_x1_sg U67455 ( .A(n9727), .B(n9728), .X(n9725) );
  nand_x2_sg U67456 ( .A(n9731), .B(n9732), .X(n9723) );
  nand_x1_sg U67457 ( .A(n46607), .B(n50610), .X(n9732) );
  nor_x1_sg U67458 ( .A(n9733), .B(n9734), .X(n9731) );
  nand_x2_sg U67459 ( .A(n9773), .B(n9774), .X(n9772) );
  nand_x1_sg U67460 ( .A(n46602), .B(n50565), .X(n9774) );
  nor_x1_sg U67461 ( .A(n9775), .B(n9776), .X(n9773) );
  nand_x2_sg U67462 ( .A(n9779), .B(n9780), .X(n9771) );
  nand_x1_sg U67463 ( .A(n46607), .B(n50561), .X(n9780) );
  nor_x1_sg U67464 ( .A(n9781), .B(n9782), .X(n9779) );
  nand_x2_sg U67465 ( .A(n9821), .B(n9822), .X(n9820) );
  nand_x1_sg U67466 ( .A(n46602), .B(n50518), .X(n9822) );
  nor_x1_sg U67467 ( .A(n9823), .B(n9824), .X(n9821) );
  nand_x2_sg U67468 ( .A(n9827), .B(n9828), .X(n9819) );
  nand_x1_sg U67469 ( .A(n46607), .B(n50514), .X(n9828) );
  nor_x1_sg U67470 ( .A(n9829), .B(n9830), .X(n9827) );
  nand_x2_sg U67471 ( .A(n9869), .B(n9870), .X(n9868) );
  nand_x1_sg U67472 ( .A(n46602), .B(n50471), .X(n9870) );
  nor_x1_sg U67473 ( .A(n9871), .B(n9872), .X(n9869) );
  nand_x2_sg U67474 ( .A(n9875), .B(n9876), .X(n9867) );
  nand_x1_sg U67475 ( .A(n46607), .B(n50467), .X(n9876) );
  nor_x1_sg U67476 ( .A(n9877), .B(n9878), .X(n9875) );
  nand_x2_sg U67477 ( .A(n9917), .B(n9918), .X(n9916) );
  nand_x1_sg U67478 ( .A(n46602), .B(n50425), .X(n9918) );
  nor_x1_sg U67479 ( .A(n9919), .B(n9920), .X(n9917) );
  nand_x2_sg U67480 ( .A(n9923), .B(n9924), .X(n9915) );
  nand_x1_sg U67481 ( .A(n46607), .B(n50421), .X(n9924) );
  nor_x1_sg U67482 ( .A(n9925), .B(n9926), .X(n9923) );
  nand_x2_sg U67483 ( .A(n9965), .B(n9966), .X(n9964) );
  nand_x1_sg U67484 ( .A(n46602), .B(n50378), .X(n9966) );
  nor_x1_sg U67485 ( .A(n9967), .B(n9968), .X(n9965) );
  nand_x2_sg U67486 ( .A(n10014), .B(n10015), .X(n10013) );
  nand_x1_sg U67487 ( .A(n46602), .B(n50331), .X(n10015) );
  nor_x1_sg U67488 ( .A(n10016), .B(n10017), .X(n10014) );
  nand_x2_sg U67489 ( .A(n10020), .B(n10021), .X(n10012) );
  nand_x1_sg U67490 ( .A(n46607), .B(n50327), .X(n10021) );
  nor_x1_sg U67491 ( .A(n10022), .B(n10023), .X(n10020) );
  nand_x2_sg U67492 ( .A(n10062), .B(n10063), .X(n10061) );
  nand_x1_sg U67493 ( .A(n46602), .B(n50285), .X(n10063) );
  nor_x1_sg U67494 ( .A(n10064), .B(n10065), .X(n10062) );
  nand_x2_sg U67495 ( .A(n10111), .B(n10112), .X(n10110) );
  nand_x1_sg U67496 ( .A(n46602), .B(n50239), .X(n10112) );
  nor_x1_sg U67497 ( .A(n10113), .B(n10114), .X(n10111) );
  nand_x2_sg U67498 ( .A(n10160), .B(n10161), .X(n10159) );
  nand_x1_sg U67499 ( .A(n46602), .B(n50195), .X(n10161) );
  nor_x1_sg U67500 ( .A(n10162), .B(n10163), .X(n10160) );
  nand_x2_sg U67501 ( .A(n10166), .B(n10167), .X(n10158) );
  nand_x1_sg U67502 ( .A(n46607), .B(n50191), .X(n10167) );
  nor_x1_sg U67503 ( .A(n10168), .B(n10169), .X(n10166) );
  nand_x2_sg U67504 ( .A(n24592), .B(n24593), .X(n24591) );
  nand_x1_sg U67505 ( .A(n49990), .B(n46602), .X(n24593) );
  nor_x1_sg U67506 ( .A(n24594), .B(n24595), .X(n24592) );
  nand_x2_sg U67507 ( .A(n24641), .B(n24642), .X(n24640) );
  nand_x1_sg U67508 ( .A(n49945), .B(n46602), .X(n24642) );
  nor_x1_sg U67509 ( .A(n24643), .B(n24644), .X(n24641) );
  nand_x2_sg U67510 ( .A(n24690), .B(n24691), .X(n24689) );
  nand_x1_sg U67511 ( .A(n49897), .B(n46602), .X(n24691) );
  nor_x1_sg U67512 ( .A(n24692), .B(n24693), .X(n24690) );
  nand_x2_sg U67513 ( .A(n24696), .B(n24697), .X(n24688) );
  nand_x1_sg U67514 ( .A(n49893), .B(n46607), .X(n24697) );
  nor_x1_sg U67515 ( .A(n24698), .B(n24699), .X(n24696) );
  nand_x2_sg U67516 ( .A(n24738), .B(n24739), .X(n24737) );
  nand_x1_sg U67517 ( .A(n49850), .B(n46602), .X(n24739) );
  nor_x1_sg U67518 ( .A(n24740), .B(n24741), .X(n24738) );
  nand_x2_sg U67519 ( .A(n24744), .B(n24745), .X(n24736) );
  nand_x1_sg U67520 ( .A(n49846), .B(n46607), .X(n24745) );
  nor_x1_sg U67521 ( .A(n24746), .B(n24747), .X(n24744) );
  nand_x2_sg U67522 ( .A(n24786), .B(n24787), .X(n24785) );
  nand_x1_sg U67523 ( .A(n49802), .B(n46602), .X(n24787) );
  nor_x1_sg U67524 ( .A(n24788), .B(n24789), .X(n24786) );
  nand_x2_sg U67525 ( .A(n24833), .B(n24834), .X(n24832) );
  nand_x1_sg U67526 ( .A(n49755), .B(n46602), .X(n24834) );
  nor_x1_sg U67527 ( .A(n24835), .B(n24836), .X(n24833) );
  nand_x2_sg U67528 ( .A(n24839), .B(n24840), .X(n24831) );
  nand_x1_sg U67529 ( .A(n49751), .B(n46607), .X(n24840) );
  nor_x1_sg U67530 ( .A(n24841), .B(n24842), .X(n24839) );
  nand_x2_sg U67531 ( .A(n24881), .B(n24882), .X(n24880) );
  nand_x1_sg U67532 ( .A(n49706), .B(n46602), .X(n24882) );
  nor_x1_sg U67533 ( .A(n24883), .B(n24884), .X(n24881) );
  nand_x2_sg U67534 ( .A(n24887), .B(n24888), .X(n24879) );
  nand_x1_sg U67535 ( .A(n49702), .B(n46607), .X(n24888) );
  nor_x1_sg U67536 ( .A(n24889), .B(n24890), .X(n24887) );
  nand_x2_sg U67537 ( .A(n24929), .B(n24930), .X(n24928) );
  nand_x1_sg U67538 ( .A(n49659), .B(n46602), .X(n24930) );
  nor_x1_sg U67539 ( .A(n24931), .B(n24932), .X(n24929) );
  nand_x2_sg U67540 ( .A(n24935), .B(n24936), .X(n24927) );
  nand_x1_sg U67541 ( .A(n49655), .B(n46607), .X(n24936) );
  nor_x1_sg U67542 ( .A(n24937), .B(n24938), .X(n24935) );
  nand_x2_sg U67543 ( .A(n24977), .B(n24978), .X(n24976) );
  nand_x1_sg U67544 ( .A(n49612), .B(n46602), .X(n24978) );
  nor_x1_sg U67545 ( .A(n24979), .B(n24980), .X(n24977) );
  nand_x2_sg U67546 ( .A(n24983), .B(n24984), .X(n24975) );
  nand_x1_sg U67547 ( .A(n49608), .B(n46607), .X(n24984) );
  nor_x1_sg U67548 ( .A(n24985), .B(n24986), .X(n24983) );
  nand_x2_sg U67549 ( .A(n25025), .B(n25026), .X(n25024) );
  nand_x1_sg U67550 ( .A(n49566), .B(n46602), .X(n25026) );
  nor_x1_sg U67551 ( .A(n25027), .B(n25028), .X(n25025) );
  nand_x2_sg U67552 ( .A(n25031), .B(n25032), .X(n25023) );
  nand_x1_sg U67553 ( .A(n49562), .B(n46607), .X(n25032) );
  nor_x1_sg U67554 ( .A(n25033), .B(n25034), .X(n25031) );
  nand_x2_sg U67555 ( .A(n25073), .B(n25074), .X(n25072) );
  nand_x1_sg U67556 ( .A(n49519), .B(n46602), .X(n25074) );
  nor_x1_sg U67557 ( .A(n25075), .B(n25076), .X(n25073) );
  nand_x2_sg U67558 ( .A(n25122), .B(n25123), .X(n25121) );
  nand_x1_sg U67559 ( .A(n49472), .B(n46602), .X(n25123) );
  nor_x1_sg U67560 ( .A(n25124), .B(n25125), .X(n25122) );
  nand_x2_sg U67561 ( .A(n25128), .B(n25129), .X(n25120) );
  nand_x1_sg U67562 ( .A(n49468), .B(n46607), .X(n25129) );
  nor_x1_sg U67563 ( .A(n25130), .B(n25131), .X(n25128) );
  nand_x2_sg U67564 ( .A(n25170), .B(n25171), .X(n25169) );
  nand_x1_sg U67565 ( .A(n49426), .B(n46602), .X(n25171) );
  nor_x1_sg U67566 ( .A(n25172), .B(n25173), .X(n25170) );
  nand_x2_sg U67567 ( .A(n25219), .B(n25220), .X(n25218) );
  nand_x1_sg U67568 ( .A(n49380), .B(n46602), .X(n25220) );
  nor_x1_sg U67569 ( .A(n25221), .B(n25222), .X(n25219) );
  nand_x2_sg U67570 ( .A(n25268), .B(n25269), .X(n25267) );
  nand_x1_sg U67571 ( .A(n49336), .B(n46602), .X(n25269) );
  nor_x1_sg U67572 ( .A(n25270), .B(n25271), .X(n25268) );
  nand_x2_sg U67573 ( .A(n25274), .B(n25275), .X(n25266) );
  nand_x1_sg U67574 ( .A(n49332), .B(n46607), .X(n25275) );
  nor_x1_sg U67575 ( .A(n25276), .B(n25277), .X(n25274) );
  nand_x2_sg U67576 ( .A(n9435), .B(n9436), .X(n9434) );
  nand_x1_sg U67577 ( .A(n46602), .B(n50898), .X(n9436) );
  nor_x1_sg U67578 ( .A(n9437), .B(n9438), .X(n9435) );
  nand_x2_sg U67579 ( .A(n9452), .B(n9453), .X(n9448) );
  nor_x1_sg U67580 ( .A(n9455), .B(n9456), .X(n9452) );
  nand_x2_sg U67581 ( .A(n9501), .B(n9502), .X(n9497) );
  nor_x1_sg U67582 ( .A(n9504), .B(n9505), .X(n9501) );
  nand_x2_sg U67583 ( .A(n9550), .B(n9551), .X(n9546) );
  nor_x1_sg U67584 ( .A(n9553), .B(n9554), .X(n9550) );
  nand_x2_sg U67585 ( .A(n9598), .B(n9599), .X(n9594) );
  nor_x1_sg U67586 ( .A(n9601), .B(n9602), .X(n9598) );
  nand_x2_sg U67587 ( .A(n9646), .B(n9647), .X(n9642) );
  nor_x1_sg U67588 ( .A(n9649), .B(n9650), .X(n9646) );
  nand_x2_sg U67589 ( .A(n9741), .B(n9742), .X(n9737) );
  nor_x1_sg U67590 ( .A(n9744), .B(n9745), .X(n9741) );
  nand_x2_sg U67591 ( .A(n9789), .B(n9790), .X(n9785) );
  nor_x1_sg U67592 ( .A(n9792), .B(n9793), .X(n9789) );
  nand_x2_sg U67593 ( .A(n9837), .B(n9838), .X(n9833) );
  nor_x1_sg U67594 ( .A(n9840), .B(n9841), .X(n9837) );
  nand_x2_sg U67595 ( .A(n9885), .B(n9886), .X(n9881) );
  nor_x1_sg U67596 ( .A(n9888), .B(n9889), .X(n9885) );
  nand_x2_sg U67597 ( .A(n9933), .B(n9934), .X(n9929) );
  nor_x1_sg U67598 ( .A(n9936), .B(n9937), .X(n9933) );
  nand_x2_sg U67599 ( .A(n9982), .B(n9983), .X(n9977) );
  nor_x1_sg U67600 ( .A(n9985), .B(n9986), .X(n9982) );
  nand_x2_sg U67601 ( .A(n10030), .B(n10031), .X(n10026) );
  nor_x1_sg U67602 ( .A(n10033), .B(n10034), .X(n10030) );
  nand_x2_sg U67603 ( .A(n10079), .B(n10080), .X(n10074) );
  nor_x1_sg U67604 ( .A(n10082), .B(n10083), .X(n10079) );
  nand_x2_sg U67605 ( .A(n10128), .B(n10129), .X(n10123) );
  nor_x1_sg U67606 ( .A(n10131), .B(n10132), .X(n10128) );
  nand_x2_sg U67607 ( .A(n10176), .B(n10177), .X(n10172) );
  nand_x1_sg U67608 ( .A(n46600), .B(n50188), .X(n10177) );
  nor_x1_sg U67609 ( .A(n10178), .B(n10179), .X(n10176) );
  nand_x2_sg U67610 ( .A(n24543), .B(n24544), .X(n24542) );
  nand_x1_sg U67611 ( .A(n50039), .B(n46602), .X(n24544) );
  nor_x1_sg U67612 ( .A(n24545), .B(n24546), .X(n24543) );
  nand_x2_sg U67613 ( .A(n24560), .B(n24561), .X(n24556) );
  nor_x1_sg U67614 ( .A(n24563), .B(n24564), .X(n24560) );
  nand_x2_sg U67615 ( .A(n24609), .B(n24610), .X(n24605) );
  nor_x1_sg U67616 ( .A(n24612), .B(n24613), .X(n24609) );
  nand_x2_sg U67617 ( .A(n24658), .B(n24659), .X(n24654) );
  nor_x1_sg U67618 ( .A(n24661), .B(n24662), .X(n24658) );
  nand_x2_sg U67619 ( .A(n24706), .B(n24707), .X(n24702) );
  nor_x1_sg U67620 ( .A(n24709), .B(n24710), .X(n24706) );
  nand_x2_sg U67621 ( .A(n24754), .B(n24755), .X(n24750) );
  nor_x1_sg U67622 ( .A(n24757), .B(n24758), .X(n24754) );
  nand_x2_sg U67623 ( .A(n24849), .B(n24850), .X(n24845) );
  nor_x1_sg U67624 ( .A(n24852), .B(n24853), .X(n24849) );
  nand_x2_sg U67625 ( .A(n24897), .B(n24898), .X(n24893) );
  nor_x1_sg U67626 ( .A(n24900), .B(n24901), .X(n24897) );
  nand_x2_sg U67627 ( .A(n24945), .B(n24946), .X(n24941) );
  nor_x1_sg U67628 ( .A(n24948), .B(n24949), .X(n24945) );
  nand_x2_sg U67629 ( .A(n24993), .B(n24994), .X(n24989) );
  nor_x1_sg U67630 ( .A(n24996), .B(n24997), .X(n24993) );
  nand_x2_sg U67631 ( .A(n25041), .B(n25042), .X(n25037) );
  nor_x1_sg U67632 ( .A(n25044), .B(n25045), .X(n25041) );
  nand_x2_sg U67633 ( .A(n25090), .B(n25091), .X(n25085) );
  nor_x1_sg U67634 ( .A(n25093), .B(n25094), .X(n25090) );
  nand_x2_sg U67635 ( .A(n25138), .B(n25139), .X(n25134) );
  nor_x1_sg U67636 ( .A(n25141), .B(n25142), .X(n25138) );
  nand_x2_sg U67637 ( .A(n25187), .B(n25188), .X(n25182) );
  nor_x1_sg U67638 ( .A(n25190), .B(n25191), .X(n25187) );
  nand_x2_sg U67639 ( .A(n25236), .B(n25237), .X(n25231) );
  nor_x1_sg U67640 ( .A(n25239), .B(n25240), .X(n25236) );
  nand_x2_sg U67641 ( .A(n25284), .B(n25285), .X(n25280) );
  nand_x1_sg U67642 ( .A(n46600), .B(n49329), .X(n25285) );
  nor_x1_sg U67643 ( .A(n25286), .B(n25287), .X(n25284) );
  nor_x1_sg U67644 ( .A(n46585), .B(n26226), .X(\L1_0/n4507 ) );
  nand_x2_sg U67645 ( .A(n46235), .B(n46507), .X(n26226) );
  nor_x1_sg U67646 ( .A(n46591), .B(n27902), .X(\L1_0/n4027 ) );
  nand_x2_sg U67647 ( .A(n46235), .B(n46372), .X(n27902) );
  nor_x1_sg U67648 ( .A(n46596), .B(n29300), .X(\L1_0/n3627 ) );
  nand_x2_sg U67649 ( .A(n46235), .B(n46260), .X(n29300) );
  nor_x1_sg U67650 ( .A(n46625), .B(n26913), .X(\L1_0/n4270 ) );
  nand_x2_sg U67651 ( .A(n46235), .B(n26909), .X(n26914) );
  nor_x1_sg U67652 ( .A(n46623), .B(n27472), .X(\L1_0/n4110 ) );
  nand_x2_sg U67653 ( .A(n46235), .B(n27468), .X(n27473) );
  nor_x1_sg U67654 ( .A(n46619), .B(n28870), .X(\L1_0/n3710 ) );
  nand_x2_sg U67655 ( .A(n46235), .B(n28866), .X(n28871) );
  nor_x1_sg U67656 ( .A(n29150), .B(n46616), .X(\L1_0/n3630 ) );
  nand_x2_sg U67657 ( .A(n46235), .B(n29145), .X(n29152) );
  nor_x1_sg U67658 ( .A(n26077), .B(n46612), .X(\L1_0/n4510 ) );
  nand_x2_sg U67659 ( .A(n46235), .B(n26072), .X(n26080) );
  nor_x1_sg U67660 ( .A(n46621), .B(n27753), .X(\L1_0/n4030 ) );
  nand_x2_sg U67661 ( .A(n46235), .B(n27749), .X(n27754) );
  nand_x2_sg U67662 ( .A(n21962), .B(n21963), .X(n21961) );
  nand_x1_sg U67663 ( .A(n21965), .B(n46608), .X(n21962) );
  nand_x1_sg U67664 ( .A(n21964), .B(n46598), .X(n21963) );
  nand_x2_sg U67665 ( .A(n29623), .B(n29624), .X(n29622) );
  nand_x1_sg U67666 ( .A(n29628), .B(n46608), .X(n29623) );
  nand_x1_sg U67667 ( .A(n29625), .B(n46598), .X(n29624) );
  nand_x2_sg U67668 ( .A(n21946), .B(n21947), .X(n21945) );
  nor_x1_sg U67669 ( .A(n21949), .B(n21950), .X(n21946) );
  nand_x1_sg U67670 ( .A(n21948), .B(n46602), .X(n21947) );
  nand_x2_sg U67671 ( .A(n21953), .B(n21954), .X(n21944) );
  nor_x1_sg U67672 ( .A(n21956), .B(n21957), .X(n21953) );
  nand_x1_sg U67673 ( .A(n21955), .B(n46607), .X(n21954) );
  nand_x2_sg U67674 ( .A(n29600), .B(n29601), .X(n29599) );
  nor_x1_sg U67675 ( .A(n29604), .B(n29605), .X(n29600) );
  nand_x1_sg U67676 ( .A(n29602), .B(n46602), .X(n29601) );
  nand_x2_sg U67677 ( .A(n29609), .B(n29610), .X(n29598) );
  nor_x1_sg U67678 ( .A(n29613), .B(n29614), .X(n29609) );
  nand_x1_sg U67679 ( .A(n29611), .B(n46607), .X(n29610) );
  nor_x1_sg U67680 ( .A(n46589), .B(n27062), .X(\L1_0/n4267 ) );
  nand_x2_sg U67681 ( .A(n46235), .B(n46439), .X(n27062) );
  nor_x1_sg U67682 ( .A(n46593), .B(n28181), .X(\L1_0/n3947 ) );
  nand_x2_sg U67683 ( .A(n46235), .B(n46352), .X(n28181) );
  nand_x2_sg U67684 ( .A(n9397), .B(n9398), .X(n9396) );
  nand_x1_sg U67685 ( .A(n46598), .B(n50916), .X(n9398) );
  nand_x1_sg U67686 ( .A(n9400), .B(n46608), .X(n9397) );
  nand_x2_sg U67687 ( .A(n24509), .B(n24510), .X(n24508) );
  nand_x1_sg U67688 ( .A(n50057), .B(n46598), .X(n24510) );
  nand_x1_sg U67689 ( .A(n24511), .B(n46608), .X(n24509) );
  nand_x2_sg U67690 ( .A(n10218), .B(n10219), .X(n10214) );
  nor_x1_sg U67691 ( .A(n10221), .B(n10222), .X(n10218) );
  nand_x2_sg U67692 ( .A(n25326), .B(n25327), .X(n25322) );
  nor_x1_sg U67693 ( .A(n25329), .B(n25330), .X(n25326) );
  nor_x1_sg U67694 ( .A(n10078), .B(n41141), .X(n24331) );
  nor_x1_sg U67695 ( .A(n25186), .B(n41140), .X(n31997) );
  nor_x1_sg U67696 ( .A(n9981), .B(n41609), .X(n24344) );
  nor_x1_sg U67697 ( .A(n25089), .B(n41613), .X(n32010) );
  nor_x1_sg U67698 ( .A(n9388), .B(n50892), .X(n22778) );
  nor_x1_sg U67699 ( .A(n24502), .B(n50033), .X(n30444) );
  nor_x1_sg U67700 ( .A(n9380), .B(n50904), .X(n22174) );
  nor_x1_sg U67701 ( .A(n24495), .B(n50045), .X(n29839) );
  nor_x1_sg U67702 ( .A(n9400), .B(n50868), .X(n22802) );
  nor_x1_sg U67703 ( .A(n24511), .B(n50009), .X(n30468) );
  nor_x1_sg U67704 ( .A(n45493), .B(n24352), .X(n24349) );
  nor_x1_sg U67705 ( .A(n45491), .B(n32018), .X(n32015) );
  nor_x1_sg U67706 ( .A(n42761), .B(n41181), .X(n22510) );
  nor_x1_sg U67707 ( .A(n42759), .B(n41145), .X(n22498) );
  nor_x1_sg U67708 ( .A(n42689), .B(n41179), .X(n30176) );
  nor_x1_sg U67709 ( .A(n42687), .B(n41143), .X(n30164) );
  nor_x1_sg U67710 ( .A(n41350), .B(n22526), .X(n22525) );
  nor_x1_sg U67711 ( .A(n41348), .B(n30192), .X(n30191) );
  nor_x1_sg U67712 ( .A(n41486), .B(n21980), .X(n21978) );
  nor_x1_sg U67713 ( .A(n41488), .B(n22508), .X(n22507) );
  nor_x1_sg U67714 ( .A(n41482), .B(n29645), .X(n29643) );
  nor_x1_sg U67715 ( .A(n41484), .B(n30174), .X(n30173) );
  nand_x2_sg U67716 ( .A(n22533), .B(n22532), .X(n22534) );
  nand_x2_sg U67717 ( .A(n30199), .B(n30198), .X(n30200) );
  nand_x2_sg U67718 ( .A(n25575), .B(n25576), .X(n25573) );
  nor_x1_sg U67719 ( .A(n25575), .B(n25576), .X(n25574) );
  nand_x2_sg U67720 ( .A(n27531), .B(n27532), .X(n27529) );
  nor_x1_sg U67721 ( .A(n27531), .B(n27532), .X(n27530) );
  nand_x2_sg U67722 ( .A(n26136), .B(n26137), .X(n26134) );
  nor_x1_sg U67723 ( .A(n26136), .B(n26137), .X(n26135) );
  nand_x2_sg U67724 ( .A(n28091), .B(n28092), .X(n28089) );
  nor_x1_sg U67725 ( .A(n28091), .B(n28092), .X(n28090) );
  nand_x2_sg U67726 ( .A(n28649), .B(n28650), .X(n28647) );
  nor_x1_sg U67727 ( .A(n28649), .B(n28650), .X(n28648) );
  nand_x2_sg U67728 ( .A(n29210), .B(n29211), .X(n29208) );
  nor_x1_sg U67729 ( .A(n29210), .B(n29211), .X(n29209) );
  inv_x8_sg U67730 ( .A(n46201), .X(n11265) );
  nor_x1_sg U67731 ( .A(n22806), .B(n41213), .X(n22805) );
  nor_x1_sg U67732 ( .A(n30472), .B(n41212), .X(n30471) );
  nand_x2_sg U67733 ( .A(n52692), .B(n52706), .X(n26959) );
  nand_x2_sg U67734 ( .A(n26960), .B(n26961), .X(n26958) );
  nand_x2_sg U67735 ( .A(n53811), .B(n53826), .X(n28078) );
  nand_x2_sg U67736 ( .A(n28079), .B(n28080), .X(n28077) );
  nand_x2_sg U67737 ( .A(n54376), .B(n54391), .X(n28636) );
  nand_x2_sg U67738 ( .A(n28637), .B(n28638), .X(n28635) );
  nand_x2_sg U67739 ( .A(n54944), .B(n54959), .X(n29197) );
  nand_x2_sg U67740 ( .A(n29198), .B(n29199), .X(n29196) );
  nor_x1_sg U67741 ( .A(n41958), .B(n10154), .X(n23770) );
  nor_x1_sg U67742 ( .A(n41956), .B(n25262), .X(n31436) );
  nand_x4_sg U67743 ( .A(n55468), .B(n55458), .X(n29627) );
  nor_x1_sg U67744 ( .A(n16367), .B(n41622), .X(n16366) );
  nor_x1_sg U67745 ( .A(n11693), .B(n41648), .X(n11692) );
  nor_x1_sg U67746 ( .A(n12472), .B(n41646), .X(n12471) );
  nor_x1_sg U67747 ( .A(n13253), .B(n41644), .X(n13252) );
  nor_x1_sg U67748 ( .A(n14033), .B(n41642), .X(n14032) );
  nor_x1_sg U67749 ( .A(n14805), .B(n41640), .X(n14804) );
  nor_x1_sg U67750 ( .A(n15586), .B(n41638), .X(n15585) );
  nor_x1_sg U67751 ( .A(n17152), .B(n41636), .X(n17151) );
  nor_x1_sg U67752 ( .A(n17926), .B(n41634), .X(n17925) );
  nor_x1_sg U67753 ( .A(n18695), .B(n41632), .X(n18694) );
  nor_x1_sg U67754 ( .A(n19471), .B(n41630), .X(n19470) );
  nor_x1_sg U67755 ( .A(n20241), .B(n41628), .X(n20240) );
  nor_x1_sg U67756 ( .A(n21015), .B(n41626), .X(n21014) );
  nor_x1_sg U67757 ( .A(n21786), .B(n41624), .X(n21785) );
  nor_x1_sg U67758 ( .A(n22772), .B(n9447), .X(n22872) );
  nor_x1_sg U67759 ( .A(n30438), .B(n24555), .X(n30538) );
  nor_x1_sg U67760 ( .A(n22766), .B(n9496), .X(n22875) );
  nor_x1_sg U67761 ( .A(n22760), .B(n9545), .X(n22878) );
  nor_x1_sg U67762 ( .A(n30432), .B(n24604), .X(n30541) );
  nor_x1_sg U67763 ( .A(n30426), .B(n24653), .X(n30544) );
  nor_x1_sg U67764 ( .A(n24226), .B(n10057), .X(n24299) );
  nor_x1_sg U67765 ( .A(n24220), .B(n10106), .X(n24302) );
  nor_x1_sg U67766 ( .A(n31892), .B(n25160), .X(n31965) );
  nor_x1_sg U67767 ( .A(n31886), .B(n25209), .X(n31968) );
  nor_x1_sg U67768 ( .A(n24238), .B(n9960), .X(n24293) );
  nor_x1_sg U67769 ( .A(n31904), .B(n25063), .X(n31959) );
  nor_x1_sg U67770 ( .A(n22612), .B(n9393), .X(n22611) );
  nor_x1_sg U67771 ( .A(n9412), .B(n9383), .X(n22001) );
  nor_x1_sg U67772 ( .A(n30278), .B(n24506), .X(n30277) );
  nor_x1_sg U67773 ( .A(n24521), .B(n24498), .X(n29666) );
  nor_x1_sg U67774 ( .A(n22554), .B(n9372), .X(n22553) );
  nor_x1_sg U67775 ( .A(n30220), .B(n24483), .X(n30219) );
  nor_x1_sg U67776 ( .A(n22682), .B(n10171), .X(n22917) );
  nor_x1_sg U67777 ( .A(n30348), .B(n25279), .X(n30583) );
  nor_x1_sg U67778 ( .A(n22736), .B(n9736), .X(n22890) );
  nor_x1_sg U67779 ( .A(n23978), .B(n9812), .X(n24043) );
  nor_x1_sg U67780 ( .A(n22700), .B(n10025), .X(n22908) );
  nor_x1_sg U67781 ( .A(n22688), .B(n10122), .X(n22914) );
  nor_x1_sg U67782 ( .A(n23936), .B(n10151), .X(n24064) );
  nor_x1_sg U67783 ( .A(n30402), .B(n24844), .X(n30556) );
  nor_x1_sg U67784 ( .A(n30366), .B(n25133), .X(n30574) );
  nor_x1_sg U67785 ( .A(n30354), .B(n25230), .X(n30580) );
  nor_x1_sg U67786 ( .A(n9511), .B(n9488), .X(n22007) );
  nor_x1_sg U67787 ( .A(n9560), .B(n9537), .X(n22010) );
  nor_x1_sg U67788 ( .A(n22754), .B(n9593), .X(n22881) );
  nor_x1_sg U67789 ( .A(n9608), .B(n9586), .X(n22013) );
  nor_x1_sg U67790 ( .A(n22748), .B(n9641), .X(n22884) );
  nor_x1_sg U67791 ( .A(n9656), .B(n9634), .X(n22016) );
  nor_x1_sg U67792 ( .A(n22742), .B(n9689), .X(n22887) );
  nor_x1_sg U67793 ( .A(n9703), .B(n9682), .X(n22019) );
  nor_x1_sg U67794 ( .A(n9751), .B(n9729), .X(n22022) );
  nor_x1_sg U67795 ( .A(n22730), .B(n9784), .X(n22893) );
  nor_x1_sg U67796 ( .A(n9799), .B(n9777), .X(n22025) );
  nor_x1_sg U67797 ( .A(n22724), .B(n9832), .X(n22896) );
  nor_x1_sg U67798 ( .A(n9847), .B(n9825), .X(n22028) );
  nor_x1_sg U67799 ( .A(n22718), .B(n9880), .X(n22899) );
  nor_x1_sg U67800 ( .A(n9895), .B(n9873), .X(n22031) );
  nor_x1_sg U67801 ( .A(n22712), .B(n9928), .X(n22902) );
  nor_x1_sg U67802 ( .A(n9943), .B(n9921), .X(n22034) );
  nor_x1_sg U67803 ( .A(n23954), .B(n10005), .X(n24055) );
  nor_x1_sg U67804 ( .A(n22706), .B(n9976), .X(n22905) );
  nor_x1_sg U67805 ( .A(n9992), .B(n9969), .X(n22037) );
  nor_x1_sg U67806 ( .A(n10040), .B(n10018), .X(n22040) );
  nor_x1_sg U67807 ( .A(n23942), .B(n10102), .X(n24061) );
  nor_x1_sg U67808 ( .A(n22694), .B(n10073), .X(n22911) );
  nor_x1_sg U67809 ( .A(n10089), .B(n10066), .X(n22043) );
  nor_x1_sg U67810 ( .A(n10138), .B(n10115), .X(n22046) );
  nor_x1_sg U67811 ( .A(n10185), .B(n10164), .X(n22049) );
  nor_x1_sg U67812 ( .A(n24619), .B(n24596), .X(n29672) );
  nor_x1_sg U67813 ( .A(n24668), .B(n24645), .X(n29675) );
  nor_x1_sg U67814 ( .A(n30420), .B(n24701), .X(n30547) );
  nor_x1_sg U67815 ( .A(n24716), .B(n24694), .X(n29678) );
  nor_x1_sg U67816 ( .A(n30414), .B(n24749), .X(n30550) );
  nor_x1_sg U67817 ( .A(n24764), .B(n24742), .X(n29681) );
  nor_x1_sg U67818 ( .A(n30408), .B(n24797), .X(n30553) );
  nor_x1_sg U67819 ( .A(n24811), .B(n24790), .X(n29684) );
  nor_x1_sg U67820 ( .A(n24859), .B(n24837), .X(n29687) );
  nor_x1_sg U67821 ( .A(n30396), .B(n24892), .X(n30559) );
  nor_x1_sg U67822 ( .A(n24907), .B(n24885), .X(n29690) );
  nor_x1_sg U67823 ( .A(n30390), .B(n24940), .X(n30562) );
  nor_x1_sg U67824 ( .A(n24955), .B(n24933), .X(n29693) );
  nor_x1_sg U67825 ( .A(n30384), .B(n24988), .X(n30565) );
  nor_x1_sg U67826 ( .A(n25003), .B(n24981), .X(n29696) );
  nor_x1_sg U67827 ( .A(n30378), .B(n25036), .X(n30568) );
  nor_x1_sg U67828 ( .A(n25051), .B(n25029), .X(n29699) );
  nor_x1_sg U67829 ( .A(n30372), .B(n25084), .X(n30571) );
  nor_x1_sg U67830 ( .A(n25100), .B(n25077), .X(n29702) );
  nor_x1_sg U67831 ( .A(n25148), .B(n25126), .X(n29705) );
  nor_x1_sg U67832 ( .A(n30360), .B(n25181), .X(n30577) );
  nor_x1_sg U67833 ( .A(n25197), .B(n25174), .X(n29708) );
  nor_x1_sg U67834 ( .A(n25246), .B(n25223), .X(n29711) );
  nor_x1_sg U67835 ( .A(n25293), .B(n25272), .X(n29714) );
  nor_x1_sg U67836 ( .A(n23972), .B(n9860), .X(n24046) );
  nor_x1_sg U67837 ( .A(n23966), .B(n9908), .X(n24049) );
  nor_x1_sg U67838 ( .A(n23960), .B(n9956), .X(n24052) );
  nor_x1_sg U67839 ( .A(n23948), .B(n10053), .X(n24058) );
  nor_x1_sg U67840 ( .A(n31644), .B(n24920), .X(n31709) );
  nor_x1_sg U67841 ( .A(n31638), .B(n24968), .X(n31712) );
  nor_x1_sg U67842 ( .A(n31632), .B(n25016), .X(n31715) );
  nor_x1_sg U67843 ( .A(n31626), .B(n25064), .X(n31718) );
  nor_x1_sg U67844 ( .A(n31620), .B(n25113), .X(n31721) );
  nor_x1_sg U67845 ( .A(n31614), .B(n25161), .X(n31724) );
  nor_x1_sg U67846 ( .A(n31608), .B(n25210), .X(n31727) );
  nor_x1_sg U67847 ( .A(n31602), .B(n25259), .X(n31730) );
  nor_x1_sg U67848 ( .A(n24232), .B(n10009), .X(n24296) );
  nor_x1_sg U67849 ( .A(n31898), .B(n25112), .X(n31962) );
  nor_x1_sg U67850 ( .A(n24214), .B(n10155), .X(n24305) );
  nor_x1_sg U67851 ( .A(n24244), .B(n9912), .X(n24290) );
  nor_x1_sg U67852 ( .A(n31910), .B(n25015), .X(n31956) );
  nor_x1_sg U67853 ( .A(n31880), .B(n25258), .X(n31971) );
  nor_x1_sg U67854 ( .A(n23319), .B(n9524), .X(n23318) );
  nor_x1_sg U67855 ( .A(n23714), .B(n9621), .X(n23713) );
  nor_x1_sg U67856 ( .A(n23990), .B(n9716), .X(n24037) );
  nor_x1_sg U67857 ( .A(n23093), .B(n9475), .X(n23092) );
  nor_x1_sg U67858 ( .A(n23524), .B(n9573), .X(n23523) );
  nor_x1_sg U67859 ( .A(n23885), .B(n9669), .X(n23884) );
  nor_x1_sg U67860 ( .A(n23984), .B(n9764), .X(n24040) );
  nor_x1_sg U67861 ( .A(n22838), .B(n9426), .X(n22837) );
  nor_x1_sg U67862 ( .A(n9462), .B(n9439), .X(n22004) );
  nor_x1_sg U67863 ( .A(n24570), .B(n24547), .X(n29669) );
  nor_x1_sg U67864 ( .A(n22569), .B(n9366), .X(n22568) );
  nor_x1_sg U67865 ( .A(n30235), .B(n24484), .X(n30234) );
  nor_x1_sg U67866 ( .A(n30504), .B(n24534), .X(n30503) );
  nor_x1_sg U67867 ( .A(n30759), .B(n24583), .X(n30758) );
  nor_x1_sg U67868 ( .A(n30985), .B(n24632), .X(n30984) );
  nor_x1_sg U67869 ( .A(n31190), .B(n24681), .X(n31189) );
  nor_x1_sg U67870 ( .A(n31380), .B(n24729), .X(n31379) );
  nor_x1_sg U67871 ( .A(n31551), .B(n24777), .X(n31550) );
  nor_x1_sg U67872 ( .A(n31656), .B(n24824), .X(n31703) );
  nor_x1_sg U67873 ( .A(n31650), .B(n24872), .X(n31706) );
  nor_x1_sg U67874 ( .A(n24250), .B(n9864), .X(n24287) );
  nor_x1_sg U67875 ( .A(n23701), .B(n9625), .X(n23700) );
  nor_x1_sg U67876 ( .A(n24025), .B(n9720), .X(n24024) );
  nor_x1_sg U67877 ( .A(n24256), .B(n9816), .X(n24284) );
  nor_x1_sg U67878 ( .A(n23306), .B(n9528), .X(n23305) );
  nor_x1_sg U67879 ( .A(n23511), .B(n9577), .X(n23510) );
  nor_x1_sg U67880 ( .A(n23872), .B(n9673), .X(n23871) );
  nor_x1_sg U67881 ( .A(n24169), .B(n9768), .X(n24168) );
  nor_x1_sg U67882 ( .A(n31916), .B(n24967), .X(n31953) );
  nor_x1_sg U67883 ( .A(n23080), .B(n9479), .X(n23079) );
  nor_x1_sg U67884 ( .A(n31922), .B(n24919), .X(n31950) );
  nor_x1_sg U67885 ( .A(n22825), .B(n9430), .X(n22824) );
  nor_x1_sg U67886 ( .A(n30491), .B(n24533), .X(n30490) );
  nor_x1_sg U67887 ( .A(n30746), .B(n24582), .X(n30745) );
  nor_x1_sg U67888 ( .A(n30972), .B(n24631), .X(n30971) );
  nor_x1_sg U67889 ( .A(n31177), .B(n24680), .X(n31176) );
  nor_x1_sg U67890 ( .A(n31367), .B(n24728), .X(n31366) );
  nor_x1_sg U67891 ( .A(n31538), .B(n24776), .X(n31537) );
  nor_x1_sg U67892 ( .A(n31691), .B(n24823), .X(n31690) );
  nor_x1_sg U67893 ( .A(n31835), .B(n24871), .X(n31834) );
  nor_x1_sg U67894 ( .A(n23193), .B(n10067), .X(n23374) );
  nor_x1_sg U67895 ( .A(n23181), .B(n10165), .X(n23380) );
  nor_x1_sg U67896 ( .A(n30859), .B(n25175), .X(n31040) );
  nor_x1_sg U67897 ( .A(n30847), .B(n25273), .X(n31046) );
  nor_x1_sg U67898 ( .A(n22322), .B(n9658), .X(n22364) );
  nor_x1_sg U67899 ( .A(n22316), .B(n9705), .X(n22367) );
  nor_x1_sg U67900 ( .A(n22310), .B(n9753), .X(n22370) );
  nor_x1_sg U67901 ( .A(n22304), .B(n9801), .X(n22373) );
  nor_x1_sg U67902 ( .A(n23223), .B(n9826), .X(n23359) );
  nor_x1_sg U67903 ( .A(n22298), .B(n9849), .X(n22376) );
  nor_x1_sg U67904 ( .A(n23217), .B(n9874), .X(n23362) );
  nor_x1_sg U67905 ( .A(n22292), .B(n9897), .X(n22379) );
  nor_x1_sg U67906 ( .A(n23211), .B(n9922), .X(n23365) );
  nor_x1_sg U67907 ( .A(n22286), .B(n9945), .X(n22382) );
  nor_x1_sg U67908 ( .A(n23205), .B(n9970), .X(n23368) );
  nor_x1_sg U67909 ( .A(n22280), .B(n9994), .X(n22385) );
  nor_x1_sg U67910 ( .A(n23199), .B(n10019), .X(n23371) );
  nor_x1_sg U67911 ( .A(n22274), .B(n10042), .X(n22388) );
  nor_x1_sg U67912 ( .A(n22268), .B(n10091), .X(n22391) );
  nor_x1_sg U67913 ( .A(n23187), .B(n10116), .X(n23377) );
  nor_x1_sg U67914 ( .A(n22262), .B(n10140), .X(n22394) );
  nor_x1_sg U67915 ( .A(n22256), .B(n10187), .X(n22397) );
  nor_x1_sg U67916 ( .A(n29987), .B(n24766), .X(n30029) );
  nor_x1_sg U67917 ( .A(n29981), .B(n24813), .X(n30032) );
  nor_x1_sg U67918 ( .A(n29975), .B(n24861), .X(n30035) );
  nor_x1_sg U67919 ( .A(n29969), .B(n24909), .X(n30038) );
  nor_x1_sg U67920 ( .A(n30889), .B(n24934), .X(n31025) );
  nor_x1_sg U67921 ( .A(n29963), .B(n24957), .X(n30041) );
  nor_x1_sg U67922 ( .A(n30883), .B(n24982), .X(n31028) );
  nor_x1_sg U67923 ( .A(n29957), .B(n25005), .X(n30044) );
  nor_x1_sg U67924 ( .A(n30877), .B(n25030), .X(n31031) );
  nor_x1_sg U67925 ( .A(n29951), .B(n25053), .X(n30047) );
  nor_x1_sg U67926 ( .A(n30871), .B(n25078), .X(n31034) );
  nor_x1_sg U67927 ( .A(n29945), .B(n25102), .X(n30050) );
  nor_x1_sg U67928 ( .A(n30865), .B(n25127), .X(n31037) );
  nor_x1_sg U67929 ( .A(n29939), .B(n25150), .X(n30053) );
  nor_x1_sg U67930 ( .A(n29933), .B(n25199), .X(n30056) );
  nor_x1_sg U67931 ( .A(n30853), .B(n25224), .X(n31043) );
  nor_x1_sg U67932 ( .A(n29927), .B(n25248), .X(n30059) );
  nor_x1_sg U67933 ( .A(n29921), .B(n25295), .X(n30062) );
  nor_x1_sg U67934 ( .A(n22328), .B(n9610), .X(n22361) );
  nor_x1_sg U67935 ( .A(n23229), .B(n9778), .X(n23356) );
  nor_x1_sg U67936 ( .A(n29993), .B(n24718), .X(n30026) );
  nor_x1_sg U67937 ( .A(n30895), .B(n24886), .X(n31022) );
  nor_x1_sg U67938 ( .A(n22334), .B(n9562), .X(n22358) );
  nor_x1_sg U67939 ( .A(n23235), .B(n9730), .X(n23353) );
  nor_x1_sg U67940 ( .A(n29999), .B(n24670), .X(n30023) );
  nor_x1_sg U67941 ( .A(n30901), .B(n24838), .X(n31019) );
  nor_x1_sg U67942 ( .A(n22340), .B(n9513), .X(n22355) );
  nor_x1_sg U67943 ( .A(n23241), .B(n9683), .X(n23350) );
  nor_x1_sg U67944 ( .A(n30005), .B(n24621), .X(n30020) );
  nor_x1_sg U67945 ( .A(n30907), .B(n24791), .X(n31016) );
  nor_x1_sg U67946 ( .A(n22190), .B(n9464), .X(n22189) );
  nor_x1_sg U67947 ( .A(n22861), .B(n9440), .X(n22860) );
  nor_x1_sg U67948 ( .A(n23247), .B(n9635), .X(n23347) );
  nor_x1_sg U67949 ( .A(n29855), .B(n24572), .X(n29854) );
  nor_x1_sg U67950 ( .A(n30527), .B(n24548), .X(n30526) );
  nor_x1_sg U67951 ( .A(n30913), .B(n24743), .X(n31013) );
  nor_x1_sg U67952 ( .A(n21988), .B(n9414), .X(n21987) );
  nor_x1_sg U67953 ( .A(n22598), .B(n9384), .X(n22597) );
  nor_x1_sg U67954 ( .A(n23118), .B(n9489), .X(n23117) );
  nor_x1_sg U67955 ( .A(n23259), .B(n9538), .X(n23341) );
  nor_x1_sg U67956 ( .A(n23253), .B(n9587), .X(n23344) );
  nor_x1_sg U67957 ( .A(n29653), .B(n24523), .X(n29652) );
  nor_x1_sg U67958 ( .A(n30264), .B(n24499), .X(n30263) );
  nor_x1_sg U67959 ( .A(n30784), .B(n24597), .X(n30783) );
  nor_x1_sg U67960 ( .A(n30925), .B(n24646), .X(n31007) );
  nor_x1_sg U67961 ( .A(n30919), .B(n24695), .X(n31010) );
  nor_x1_sg U67962 ( .A(n41923), .B(n24780), .X(n31496) );
  nand_x1_sg U67963 ( .A(n24780), .B(n41923), .X(n31497) );
  nor_x1_sg U67964 ( .A(n41931), .B(n9370), .X(n22789) );
  nand_x1_sg U67965 ( .A(n9370), .B(n41931), .X(n22790) );
  nor_x1_sg U67966 ( .A(n41929), .B(n24487), .X(n30455) );
  nand_x1_sg U67967 ( .A(n24487), .B(n41929), .X(n30456) );
  nor_x1_sg U67968 ( .A(n41933), .B(n9672), .X(n23830) );
  nand_x1_sg U67969 ( .A(n9672), .B(n41933), .X(n23831) );
  nor_x1_sg U67970 ( .A(n9447), .B(n22770), .X(n22769) );
  nor_x1_sg U67971 ( .A(n9496), .B(n22764), .X(n22763) );
  nor_x1_sg U67972 ( .A(n9545), .B(n22758), .X(n22757) );
  nor_x1_sg U67973 ( .A(n24555), .B(n30436), .X(n30435) );
  nor_x1_sg U67974 ( .A(n24604), .B(n30430), .X(n30429) );
  nor_x1_sg U67975 ( .A(n24653), .B(n30424), .X(n30423) );
  nor_x1_sg U67976 ( .A(n9393), .B(n22776), .X(n22775) );
  nor_x1_sg U67977 ( .A(n24506), .B(n30442), .X(n30441) );
  nor_x1_sg U67978 ( .A(n9689), .B(n22740), .X(n22739) );
  nor_x1_sg U67979 ( .A(n9976), .B(n22704), .X(n22703) );
  nor_x1_sg U67980 ( .A(n10073), .B(n22692), .X(n22691) );
  nor_x1_sg U67981 ( .A(n10122), .B(n22686), .X(n22685) );
  nor_x1_sg U67982 ( .A(n24797), .B(n30406), .X(n30405) );
  nor_x1_sg U67983 ( .A(n25084), .B(n30370), .X(n30369) );
  nor_x1_sg U67984 ( .A(n25181), .B(n30358), .X(n30357) );
  nor_x1_sg U67985 ( .A(n25230), .B(n30352), .X(n30351) );
  nor_x1_sg U67986 ( .A(n9956), .B(n23958), .X(n23957) );
  nor_x1_sg U67987 ( .A(n10053), .B(n23946), .X(n23945) );
  nor_x1_sg U67988 ( .A(n10102), .B(n23940), .X(n23939) );
  nor_x1_sg U67989 ( .A(n25259), .B(n31600), .X(n31599) );
  nor_x1_sg U67990 ( .A(n9593), .B(n22752), .X(n22751) );
  nor_x1_sg U67991 ( .A(n9641), .B(n22746), .X(n22745) );
  nor_x1_sg U67992 ( .A(n9736), .B(n22734), .X(n22733) );
  nor_x1_sg U67993 ( .A(n9784), .B(n22728), .X(n22727) );
  nor_x1_sg U67994 ( .A(n9832), .B(n22722), .X(n22721) );
  nor_x1_sg U67995 ( .A(n9880), .B(n22716), .X(n22715) );
  nor_x1_sg U67996 ( .A(n9928), .B(n22710), .X(n22709) );
  nor_x1_sg U67997 ( .A(n10025), .B(n22698), .X(n22697) );
  nor_x1_sg U67998 ( .A(n10171), .B(n22680), .X(n22679) );
  nor_x1_sg U67999 ( .A(n24701), .B(n30418), .X(n30417) );
  nor_x1_sg U68000 ( .A(n24749), .B(n30412), .X(n30411) );
  nor_x1_sg U68001 ( .A(n24844), .B(n30400), .X(n30399) );
  nor_x1_sg U68002 ( .A(n24892), .B(n30394), .X(n30393) );
  nor_x1_sg U68003 ( .A(n24940), .B(n30388), .X(n30387) );
  nor_x1_sg U68004 ( .A(n24988), .B(n30382), .X(n30381) );
  nor_x1_sg U68005 ( .A(n25036), .B(n30376), .X(n30375) );
  nor_x1_sg U68006 ( .A(n25133), .B(n30364), .X(n30363) );
  nor_x1_sg U68007 ( .A(n25279), .B(n30346), .X(n30345) );
  nor_x1_sg U68008 ( .A(n9812), .B(n23976), .X(n23975) );
  nor_x1_sg U68009 ( .A(n9860), .B(n23970), .X(n23969) );
  nor_x1_sg U68010 ( .A(n9908), .B(n23964), .X(n23963) );
  nor_x1_sg U68011 ( .A(n10005), .B(n23952), .X(n23951) );
  nor_x1_sg U68012 ( .A(n10151), .B(n23934), .X(n23933) );
  nor_x1_sg U68013 ( .A(n24920), .B(n31642), .X(n31641) );
  nor_x1_sg U68014 ( .A(n24968), .B(n31636), .X(n31635) );
  nor_x1_sg U68015 ( .A(n25016), .B(n31630), .X(n31629) );
  nor_x1_sg U68016 ( .A(n25064), .B(n31624), .X(n31623) );
  nor_x1_sg U68017 ( .A(n25113), .B(n31618), .X(n31617) );
  nor_x1_sg U68018 ( .A(n25161), .B(n31612), .X(n31611) );
  nor_x1_sg U68019 ( .A(n25210), .B(n31606), .X(n31605) );
  nor_x1_sg U68020 ( .A(n9366), .B(n22794), .X(n22793) );
  nor_x1_sg U68021 ( .A(n9475), .B(n23275), .X(n23274) );
  nor_x1_sg U68022 ( .A(n9573), .B(n23670), .X(n23669) );
  nor_x1_sg U68023 ( .A(n9669), .B(n23994), .X(n23993) );
  nor_x1_sg U68024 ( .A(n9426), .B(n23049), .X(n23048) );
  nor_x1_sg U68025 ( .A(n9524), .B(n23480), .X(n23479) );
  nor_x1_sg U68026 ( .A(n9621), .B(n23841), .X(n23840) );
  nor_x1_sg U68027 ( .A(n9716), .B(n23988), .X(n23987) );
  nor_x1_sg U68028 ( .A(n9764), .B(n23982), .X(n23981) );
  nor_x1_sg U68029 ( .A(n24484), .B(n30460), .X(n30459) );
  nor_x1_sg U68030 ( .A(n24534), .B(n30715), .X(n30714) );
  nor_x1_sg U68031 ( .A(n24583), .B(n30941), .X(n30940) );
  nor_x1_sg U68032 ( .A(n24632), .B(n31146), .X(n31145) );
  nor_x1_sg U68033 ( .A(n24681), .B(n31336), .X(n31335) );
  nor_x1_sg U68034 ( .A(n24729), .B(n31507), .X(n31506) );
  nor_x1_sg U68035 ( .A(n24777), .B(n31660), .X(n31659) );
  nor_x1_sg U68036 ( .A(n24824), .B(n31654), .X(n31653) );
  nor_x1_sg U68037 ( .A(n24872), .B(n31648), .X(n31647) );
  nor_x1_sg U68038 ( .A(n44257), .B(n42829), .X(n25597) );
  nor_x1_sg U68039 ( .A(n44263), .B(n42833), .X(n28949) );
  nor_x1_sg U68040 ( .A(n44267), .B(n42831), .X(n29510) );
  nor_x1_sg U68041 ( .A(n42949), .B(n50066), .X(n30454) );
  nor_x1_sg U68042 ( .A(n41667), .B(n49796), .X(n31318) );
  nor_x1_sg U68043 ( .A(n43013), .B(n50925), .X(n22788) );
  nor_x1_sg U68044 ( .A(n41677), .B(n50655), .X(n23652) );
  nand_x2_sg U68045 ( .A(n50169), .B(n23592), .X(n23589) );
  nand_x2_sg U68046 ( .A(n49310), .B(n31258), .X(n31255) );
  nand_x2_sg U68047 ( .A(n30935), .B(n49979), .X(n30933) );
  nor_x1_sg U68048 ( .A(n49979), .B(n30935), .X(n30934) );
  nand_x2_sg U68049 ( .A(n31330), .B(n49889), .X(n31328) );
  nor_x1_sg U68050 ( .A(n49889), .B(n31330), .X(n31329) );
  nand_x2_sg U68051 ( .A(n23269), .B(n50838), .X(n23267) );
  nor_x1_sg U68052 ( .A(n50838), .B(n23269), .X(n23268) );
  nand_x2_sg U68053 ( .A(n23664), .B(n50748), .X(n23662) );
  nor_x1_sg U68054 ( .A(n50748), .B(n23664), .X(n23663) );
  nand_x1_sg U68055 ( .A(n41233), .B(n28389), .X(n28387) );
  nand_x2_sg U68056 ( .A(n9839), .B(n43022), .X(n23632) );
  nor_x1_sg U68057 ( .A(n43022), .B(n9839), .X(n23634) );
  nand_x2_sg U68058 ( .A(n9887), .B(n41445), .X(n23626) );
  nor_x1_sg U68059 ( .A(n41445), .B(n9887), .X(n23628) );
  nand_x2_sg U68060 ( .A(n9935), .B(n41443), .X(n23620) );
  nor_x1_sg U68061 ( .A(n41443), .B(n9935), .X(n23622) );
  nand_x2_sg U68062 ( .A(n10032), .B(n41441), .X(n23608) );
  nor_x1_sg U68063 ( .A(n41441), .B(n10032), .X(n23610) );
  nand_x2_sg U68064 ( .A(n24851), .B(n41618), .X(n31310) );
  nor_x1_sg U68065 ( .A(n41618), .B(n24851), .X(n31312) );
  nand_x2_sg U68066 ( .A(n24899), .B(n41439), .X(n31304) );
  nor_x1_sg U68067 ( .A(n41439), .B(n24899), .X(n31306) );
  nand_x2_sg U68068 ( .A(n24947), .B(n42940), .X(n31298) );
  nor_x1_sg U68069 ( .A(n42940), .B(n24947), .X(n31300) );
  nand_x2_sg U68070 ( .A(n24995), .B(n41437), .X(n31292) );
  nor_x1_sg U68071 ( .A(n41437), .B(n24995), .X(n31294) );
  nand_x2_sg U68072 ( .A(n25043), .B(n41435), .X(n31286) );
  nor_x1_sg U68073 ( .A(n41435), .B(n25043), .X(n31288) );
  nand_x2_sg U68074 ( .A(n25092), .B(n42935), .X(n31280) );
  nor_x1_sg U68075 ( .A(n42935), .B(n25092), .X(n31282) );
  nand_x2_sg U68076 ( .A(n25140), .B(n41433), .X(n31274) );
  nor_x1_sg U68077 ( .A(n41433), .B(n25140), .X(n31276) );
  nand_x2_sg U68078 ( .A(n9743), .B(n41620), .X(n23644) );
  nor_x1_sg U68079 ( .A(n41620), .B(n9743), .X(n23646) );
  nand_x2_sg U68080 ( .A(n9791), .B(n41447), .X(n23638) );
  nor_x1_sg U68081 ( .A(n41447), .B(n9791), .X(n23640) );
  nand_x2_sg U68082 ( .A(n9984), .B(n43017), .X(n23614) );
  nor_x1_sg U68083 ( .A(n43017), .B(n9984), .X(n23616) );
  nand_x2_sg U68084 ( .A(n24562), .B(n42947), .X(n30707) );
  nor_x1_sg U68085 ( .A(n42947), .B(n24562), .X(n30709) );
  nand_x2_sg U68086 ( .A(n24660), .B(n42945), .X(n31138) );
  nor_x1_sg U68087 ( .A(n42945), .B(n24660), .X(n31140) );
  nand_x2_sg U68088 ( .A(n24756), .B(n41671), .X(n31322) );
  nor_x1_sg U68089 ( .A(n41671), .B(n24756), .X(n31324) );
  nand_x2_sg U68090 ( .A(n25189), .B(n41663), .X(n31268) );
  nor_x1_sg U68091 ( .A(n41663), .B(n25189), .X(n31270) );
  nand_x2_sg U68092 ( .A(n25238), .B(n44371), .X(n31262) );
  nor_x1_sg U68093 ( .A(n44371), .B(n25238), .X(n31264) );
  nand_x2_sg U68094 ( .A(n9454), .B(n43029), .X(n23041) );
  nor_x1_sg U68095 ( .A(n43029), .B(n9454), .X(n23043) );
  nand_x2_sg U68096 ( .A(n9552), .B(n43027), .X(n23472) );
  nor_x1_sg U68097 ( .A(n43027), .B(n9552), .X(n23474) );
  nand_x2_sg U68098 ( .A(n9648), .B(n41681), .X(n23656) );
  nor_x1_sg U68099 ( .A(n41681), .B(n9648), .X(n23658) );
  nand_x2_sg U68100 ( .A(n10081), .B(n41673), .X(n23602) );
  nor_x1_sg U68101 ( .A(n41673), .B(n10081), .X(n23604) );
  nand_x2_sg U68102 ( .A(n10130), .B(n44373), .X(n23596) );
  nor_x1_sg U68103 ( .A(n44373), .B(n10130), .X(n23598) );
  nor_x1_sg U68104 ( .A(n42172), .B(n25569), .X(n25570) );
  nor_x1_sg U68105 ( .A(n42184), .B(n26130), .X(n26131) );
  nor_x1_sg U68106 ( .A(n42168), .B(n27525), .X(n27526) );
  nor_x1_sg U68107 ( .A(n42180), .B(n28921), .X(n28922) );
  nor_x1_sg U68108 ( .A(n42176), .B(n29482), .X(n29483) );
  nor_x1_sg U68109 ( .A(n42148), .B(n26687), .X(n26688) );
  nand_x2_sg U68110 ( .A(n10264), .B(n40789), .X(n10267) );
  nand_x2_sg U68111 ( .A(n9815), .B(n45369), .X(n23812) );
  nor_x1_sg U68112 ( .A(n45369), .B(n9815), .X(n23814) );
  nand_x2_sg U68113 ( .A(n9863), .B(n45367), .X(n23806) );
  nor_x1_sg U68114 ( .A(n45367), .B(n9863), .X(n23808) );
  nand_x2_sg U68115 ( .A(n9911), .B(n45365), .X(n23800) );
  nor_x1_sg U68116 ( .A(n45365), .B(n9911), .X(n23802) );
  nand_x2_sg U68117 ( .A(n10008), .B(n45363), .X(n23788) );
  nor_x1_sg U68118 ( .A(n45363), .B(n10008), .X(n23790) );
  nand_x2_sg U68119 ( .A(n24537), .B(n45359), .X(n30710) );
  nor_x1_sg U68120 ( .A(n45359), .B(n24537), .X(n30712) );
  nand_x2_sg U68121 ( .A(n24635), .B(n45357), .X(n31141) );
  nor_x1_sg U68122 ( .A(n45357), .B(n24635), .X(n31143) );
  nand_x2_sg U68123 ( .A(n24732), .B(n45355), .X(n31502) );
  nor_x1_sg U68124 ( .A(n45355), .B(n24732), .X(n31504) );
  nand_x2_sg U68125 ( .A(n24827), .B(n45353), .X(n31490) );
  nor_x1_sg U68126 ( .A(n45353), .B(n24827), .X(n31492) );
  nand_x2_sg U68127 ( .A(n24875), .B(n45351), .X(n31484) );
  nor_x1_sg U68128 ( .A(n45351), .B(n24875), .X(n31486) );
  nand_x2_sg U68129 ( .A(n24923), .B(n45349), .X(n31478) );
  nor_x1_sg U68130 ( .A(n45349), .B(n24923), .X(n31480) );
  nand_x2_sg U68131 ( .A(n24971), .B(n45347), .X(n31472) );
  nor_x1_sg U68132 ( .A(n45347), .B(n24971), .X(n31474) );
  nand_x2_sg U68133 ( .A(n25019), .B(n45345), .X(n31466) );
  nor_x1_sg U68134 ( .A(n45345), .B(n25019), .X(n31468) );
  nand_x2_sg U68135 ( .A(n25067), .B(n45343), .X(n31460) );
  nor_x1_sg U68136 ( .A(n45343), .B(n25067), .X(n31462) );
  nand_x2_sg U68137 ( .A(n25116), .B(n45341), .X(n31454) );
  nor_x1_sg U68138 ( .A(n45341), .B(n25116), .X(n31456) );
  nand_x2_sg U68139 ( .A(n25164), .B(n45339), .X(n31448) );
  nor_x1_sg U68140 ( .A(n45339), .B(n25164), .X(n31450) );
  nand_x2_sg U68141 ( .A(n25213), .B(n45337), .X(n31442) );
  nor_x1_sg U68142 ( .A(n45337), .B(n25213), .X(n31444) );
  nand_x2_sg U68143 ( .A(n9429), .B(n45387), .X(n23044) );
  nor_x1_sg U68144 ( .A(n45387), .B(n9429), .X(n23046) );
  nand_x2_sg U68145 ( .A(n9527), .B(n45385), .X(n23475) );
  nor_x1_sg U68146 ( .A(n45385), .B(n9527), .X(n23477) );
  nand_x2_sg U68147 ( .A(n9624), .B(n45383), .X(n23836) );
  nor_x1_sg U68148 ( .A(n45383), .B(n9624), .X(n23838) );
  nand_x2_sg U68149 ( .A(n9719), .B(n45381), .X(n23824) );
  nor_x1_sg U68150 ( .A(n45381), .B(n9719), .X(n23826) );
  nand_x2_sg U68151 ( .A(n9767), .B(n45379), .X(n23818) );
  nor_x1_sg U68152 ( .A(n45379), .B(n9767), .X(n23820) );
  nand_x2_sg U68153 ( .A(n9959), .B(n45377), .X(n23794) );
  nor_x1_sg U68154 ( .A(n45377), .B(n9959), .X(n23796) );
  nand_x2_sg U68155 ( .A(n10056), .B(n45375), .X(n23782) );
  nor_x1_sg U68156 ( .A(n45375), .B(n10056), .X(n23784) );
  nand_x2_sg U68157 ( .A(n10105), .B(n45373), .X(n23776) );
  nor_x1_sg U68158 ( .A(n45373), .B(n10105), .X(n23778) );
  nor_x1_sg U68159 ( .A(n43163), .B(n44321), .X(n26967) );
  nand_x2_sg U68160 ( .A(n25371), .B(n40790), .X(n25373) );
  nand_x1_sg U68161 ( .A(n24417), .B(n40721), .X(n24461) );
  nand_x1_sg U68162 ( .A(n32083), .B(n40722), .X(n32127) );
  nand_x1_sg U68163 ( .A(n23625), .B(n9935), .X(n23744) );
  nand_x1_sg U68164 ( .A(n31315), .B(n24851), .X(n31398) );
  nand_x1_sg U68165 ( .A(n31309), .B(n24899), .X(n31401) );
  nand_x1_sg U68166 ( .A(n31303), .B(n24947), .X(n31404) );
  nand_x1_sg U68167 ( .A(n31297), .B(n24995), .X(n31407) );
  nand_x1_sg U68168 ( .A(n31291), .B(n25043), .X(n31410) );
  nand_x1_sg U68169 ( .A(n23631), .B(n9887), .X(n23741) );
  nand_x1_sg U68170 ( .A(n23649), .B(n9743), .X(n23732) );
  nand_x1_sg U68171 ( .A(n23643), .B(n9791), .X(n23735) );
  nand_x1_sg U68172 ( .A(n23637), .B(n9839), .X(n23738) );
  nand_x1_sg U68173 ( .A(n23619), .B(n9984), .X(n23747) );
  nand_x1_sg U68174 ( .A(n31285), .B(n25092), .X(n31413) );
  nand_x1_sg U68175 ( .A(n31279), .B(n25140), .X(n31416) );
  nand_x1_sg U68176 ( .A(n23613), .B(n10032), .X(n23750) );
  nand_x1_sg U68177 ( .A(n43161), .B(n28383), .X(n28381) );
  nor_x1_sg U68178 ( .A(n9372), .B(n22800), .X(n22799) );
  nor_x1_sg U68179 ( .A(n24483), .B(n30466), .X(n30465) );
  nor_x1_sg U68180 ( .A(n9479), .B(n23281), .X(n23280) );
  nor_x1_sg U68181 ( .A(n9577), .B(n23676), .X(n23675) );
  nor_x1_sg U68182 ( .A(n9673), .B(n24000), .X(n23999) );
  nor_x1_sg U68183 ( .A(n9768), .B(n24260), .X(n24259) );
  nor_x1_sg U68184 ( .A(n9430), .B(n23055), .X(n23054) );
  nor_x1_sg U68185 ( .A(n9528), .B(n23486), .X(n23485) );
  nor_x1_sg U68186 ( .A(n9625), .B(n23847), .X(n23846) );
  nor_x1_sg U68187 ( .A(n9720), .B(n24144), .X(n24143) );
  nor_x1_sg U68188 ( .A(n24871), .B(n31926), .X(n31925) );
  nor_x1_sg U68189 ( .A(n24533), .B(n30721), .X(n30720) );
  nor_x1_sg U68190 ( .A(n24582), .B(n30947), .X(n30946) );
  nor_x1_sg U68191 ( .A(n24631), .B(n31152), .X(n31151) );
  nor_x1_sg U68192 ( .A(n24680), .B(n31342), .X(n31341) );
  nor_x1_sg U68193 ( .A(n24728), .B(n31513), .X(n31512) );
  nor_x1_sg U68194 ( .A(n24776), .B(n31666), .X(n31665) );
  nor_x1_sg U68195 ( .A(n24823), .B(n31810), .X(n31809) );
  nor_x1_sg U68196 ( .A(n9464), .B(n22344), .X(n22343) );
  nor_x1_sg U68197 ( .A(n24572), .B(n30009), .X(n30008) );
  nand_x4_sg U68198 ( .A(n26444), .B(n26445), .X(n12611) );
  nand_x1_sg U68199 ( .A(n52089), .B(n26446), .X(n26445) );
  nand_x1_sg U68200 ( .A(n26447), .B(n52087), .X(n26444) );
  nand_x4_sg U68201 ( .A(n27281), .B(n27282), .X(n14944) );
  nand_x1_sg U68202 ( .A(n52923), .B(n27283), .X(n27282) );
  nand_x1_sg U68203 ( .A(n27284), .B(n52921), .X(n27281) );
  nand_x4_sg U68204 ( .A(n27839), .B(n27840), .X(n16510) );
  nand_x1_sg U68205 ( .A(n53481), .B(n27841), .X(n27840) );
  nand_x1_sg U68206 ( .A(n27842), .B(n53479), .X(n27839) );
  nand_x4_sg U68207 ( .A(n25885), .B(n25886), .X(n11050) );
  nand_x1_sg U68208 ( .A(n51531), .B(n25887), .X(n25886) );
  nand_x1_sg U68209 ( .A(n25888), .B(n51529), .X(n25885) );
  nand_x4_sg U68210 ( .A(n25604), .B(n25605), .X(n10282) );
  nand_x1_sg U68211 ( .A(n51255), .B(n25606), .X(n25605) );
  nand_x1_sg U68212 ( .A(n25607), .B(n51253), .X(n25604) );
  nand_x1_sg U68213 ( .A(n24428), .B(n40795), .X(n24455) );
  nand_x1_sg U68214 ( .A(n32094), .B(n40796), .X(n32121) );
  nand_x4_sg U68215 ( .A(n26722), .B(n26723), .X(n13395) );
  nand_x1_sg U68216 ( .A(n52366), .B(n52364), .X(n26723) );
  nand_x4_sg U68217 ( .A(n25585), .B(n25586), .X(n10408) );
  nand_x1_sg U68218 ( .A(n25587), .B(n51264), .X(n25586) );
  nand_x4_sg U68219 ( .A(n28937), .B(n28938), .X(n19735) );
  nand_x1_sg U68220 ( .A(n28939), .B(n54618), .X(n28938) );
  nand_x4_sg U68221 ( .A(n29498), .B(n29499), .X(n21280) );
  nand_x1_sg U68222 ( .A(n29500), .B(n55186), .X(n29499) );
  nand_x4_sg U68223 ( .A(n25866), .B(n25867), .X(n11173) );
  nand_x4_sg U68224 ( .A(n26425), .B(n26426), .X(n12734) );
  nand_x4_sg U68225 ( .A(n27262), .B(n27263), .X(n15067) );
  nand_x4_sg U68226 ( .A(n27820), .B(n27821), .X(n16633) );
  nand_x4_sg U68227 ( .A(n26152), .B(n26153), .X(n11947) );
  nand_x4_sg U68228 ( .A(n26988), .B(n26989), .X(n14289) );
  nand_x4_sg U68229 ( .A(n27547), .B(n27548), .X(n15842) );
  nor_x1_sg U68230 ( .A(n50933), .B(n22605), .X(n22604) );
  nor_x1_sg U68231 ( .A(n50943), .B(n21995), .X(n21994) );
  nor_x1_sg U68232 ( .A(n50074), .B(n30271), .X(n30270) );
  nor_x1_sg U68233 ( .A(n50084), .B(n29660), .X(n29659) );
  nor_x1_sg U68234 ( .A(n50910), .B(n22547), .X(n22546) );
  nor_x1_sg U68235 ( .A(n50051), .B(n30213), .X(n30212) );
  nand_x4_sg U68236 ( .A(n46576), .B(n29151), .X(n21153) );
  nor_x1_sg U68237 ( .A(n50990), .B(n25862), .X(n25930) );
  nor_x1_sg U68238 ( .A(n51028), .B(n26421), .X(n26489) );
  nor_x1_sg U68239 ( .A(n51086), .B(n27258), .X(n27326) );
  nor_x1_sg U68240 ( .A(n51124), .B(n27816), .X(n27884) );
  nor_x1_sg U68241 ( .A(n50992), .B(n25850), .X(n25924) );
  nor_x1_sg U68242 ( .A(n51030), .B(n26409), .X(n26483) );
  nor_x1_sg U68243 ( .A(n51088), .B(n27246), .X(n27320) );
  nor_x1_sg U68244 ( .A(n51126), .B(n27804), .X(n27878) );
  nor_x1_sg U68245 ( .A(n51143), .B(n28097), .X(n28165) );
  nor_x1_sg U68246 ( .A(n51180), .B(n28655), .X(n28723) );
  nor_x1_sg U68247 ( .A(n51218), .B(n29216), .X(n29284) );
  nor_x1_sg U68248 ( .A(n51145), .B(n28085), .X(n28159) );
  nor_x1_sg U68249 ( .A(n51182), .B(n28643), .X(n28717) );
  nor_x1_sg U68250 ( .A(n51220), .B(n29204), .X(n29278) );
  nand_x2_sg U68251 ( .A(n25891), .B(n25893), .X(n25912) );
  nand_x2_sg U68252 ( .A(n26171), .B(n26173), .X(n26192) );
  nand_x2_sg U68253 ( .A(n26450), .B(n26452), .X(n26471) );
  nand_x2_sg U68254 ( .A(n26728), .B(n26730), .X(n26749) );
  nand_x2_sg U68255 ( .A(n27007), .B(n27009), .X(n27028) );
  nand_x2_sg U68256 ( .A(n27287), .B(n27289), .X(n27308) );
  nand_x2_sg U68257 ( .A(n27566), .B(n27568), .X(n27587) );
  nand_x2_sg U68258 ( .A(n27845), .B(n27847), .X(n27866) );
  nand_x2_sg U68259 ( .A(n28126), .B(n28128), .X(n28147) );
  nand_x2_sg U68260 ( .A(n28405), .B(n28407), .X(n28426) );
  nand_x2_sg U68261 ( .A(n28684), .B(n28686), .X(n28705) );
  nand_x2_sg U68262 ( .A(n28962), .B(n28964), .X(n28983) );
  nand_x2_sg U68263 ( .A(n29245), .B(n29247), .X(n29266) );
  nand_x2_sg U68264 ( .A(n29523), .B(n29525), .X(n29544) );
  nor_x1_sg U68265 ( .A(n41233), .B(n28389), .X(n28386) );
  nor_x1_sg U68266 ( .A(n44265), .B(n42835), .X(n26994) );
  nor_x1_sg U68267 ( .A(n44261), .B(n42827), .X(n27553) );
  nor_x1_sg U68268 ( .A(n44259), .B(n42823), .X(n25878) );
  nor_x1_sg U68269 ( .A(n44255), .B(n42841), .X(n28113) );
  nor_x1_sg U68270 ( .A(n44253), .B(n42839), .X(n28671) );
  nor_x1_sg U68271 ( .A(n44251), .B(n42837), .X(n29232) );
  nor_x1_sg U68272 ( .A(n44269), .B(n42805), .X(n26715) );
  nor_x1_sg U68273 ( .A(n44277), .B(n42825), .X(n26158) );
  nor_x1_sg U68274 ( .A(n44275), .B(n42821), .X(n26437) );
  nor_x1_sg U68275 ( .A(n44273), .B(n42819), .X(n27274) );
  nor_x1_sg U68276 ( .A(n44271), .B(n42817), .X(n27832) );
  nor_x1_sg U68277 ( .A(n10265), .B(n10266), .X(n10263) );
  nor_x1_sg U68278 ( .A(n25372), .B(n10266), .X(n25370) );
  nand_x2_sg U68279 ( .A(n23287), .B(n50776), .X(n23285) );
  nand_x2_sg U68280 ( .A(n50822), .B(n23065), .X(n23286) );
  nand_x2_sg U68281 ( .A(n23682), .B(n50684), .X(n23680) );
  nand_x2_sg U68282 ( .A(n50732), .B(n23496), .X(n23681) );
  nand_x2_sg U68283 ( .A(n24006), .B(n50593), .X(n24004) );
  nand_x2_sg U68284 ( .A(n50641), .B(n23857), .X(n24005) );
  nand_x2_sg U68285 ( .A(n30953), .B(n49917), .X(n30951) );
  nand_x2_sg U68286 ( .A(n49963), .B(n30731), .X(n30952) );
  nand_x2_sg U68287 ( .A(n31348), .B(n49825), .X(n31346) );
  nand_x2_sg U68288 ( .A(n49873), .B(n31162), .X(n31347) );
  nand_x2_sg U68289 ( .A(n31672), .B(n49734), .X(n31670) );
  nand_x2_sg U68290 ( .A(n49782), .B(n31523), .X(n31671) );
  nand_x2_sg U68291 ( .A(n24266), .B(n50502), .X(n24264) );
  nand_x2_sg U68292 ( .A(n50549), .B(n24154), .X(n24265) );
  nand_x2_sg U68293 ( .A(n31932), .B(n49643), .X(n31930) );
  nand_x2_sg U68294 ( .A(n49690), .B(n31820), .X(n31931) );
  nand_x2_sg U68295 ( .A(n22673), .B(n50130), .X(n22672) );
  nand_x2_sg U68296 ( .A(n22674), .B(n50150), .X(n22671) );
  nand_x2_sg U68297 ( .A(n30339), .B(n49271), .X(n30338) );
  nand_x2_sg U68298 ( .A(n30340), .B(n49291), .X(n30337) );
  nand_x2_sg U68299 ( .A(n23927), .B(n50136), .X(n23926) );
  nand_x2_sg U68300 ( .A(n23928), .B(n50144), .X(n23925) );
  nand_x2_sg U68301 ( .A(n31593), .B(n49277), .X(n31592) );
  nand_x2_sg U68302 ( .A(n31594), .B(n49285), .X(n31591) );
  nand_x4_sg U68303 ( .A(n24216), .B(n50228), .X(n24086) );
  nand_x1_sg U68304 ( .A(n24218), .B(n10106), .X(n24216) );
  nor_x1_sg U68305 ( .A(n10106), .B(n24218), .X(n24217) );
  nand_x4_sg U68306 ( .A(n24222), .B(n50274), .X(n24093) );
  nand_x1_sg U68307 ( .A(n24224), .B(n10057), .X(n24222) );
  nor_x1_sg U68308 ( .A(n10057), .B(n24224), .X(n24223) );
  nand_x4_sg U68309 ( .A(n31888), .B(n49415), .X(n31759) );
  nand_x1_sg U68310 ( .A(n31890), .B(n25160), .X(n31888) );
  nor_x1_sg U68311 ( .A(n25160), .B(n31890), .X(n31889) );
  nand_x4_sg U68312 ( .A(n31882), .B(n49369), .X(n31752) );
  nand_x1_sg U68313 ( .A(n31884), .B(n25209), .X(n31882) );
  nor_x1_sg U68314 ( .A(n25209), .B(n31884), .X(n31883) );
  nand_x4_sg U68315 ( .A(n24234), .B(n50367), .X(n24107) );
  nand_x1_sg U68316 ( .A(n24236), .B(n9960), .X(n24234) );
  nor_x1_sg U68317 ( .A(n9960), .B(n24236), .X(n24235) );
  nand_x4_sg U68318 ( .A(n31900), .B(n49508), .X(n31773) );
  nand_x1_sg U68319 ( .A(n31902), .B(n25063), .X(n31900) );
  nor_x1_sg U68320 ( .A(n25063), .B(n31902), .X(n31901) );
  nand_x4_sg U68321 ( .A(n24228), .B(n50320), .X(n24100) );
  nand_x1_sg U68322 ( .A(n24230), .B(n10009), .X(n24228) );
  nor_x1_sg U68323 ( .A(n10009), .B(n24230), .X(n24229) );
  nand_x4_sg U68324 ( .A(n31894), .B(n49461), .X(n31766) );
  nand_x1_sg U68325 ( .A(n31896), .B(n25112), .X(n31894) );
  nor_x1_sg U68326 ( .A(n25112), .B(n31896), .X(n31895) );
  nand_x4_sg U68327 ( .A(n24210), .B(n50184), .X(n24079) );
  nand_x1_sg U68328 ( .A(n24212), .B(n10155), .X(n24210) );
  nor_x1_sg U68329 ( .A(n10155), .B(n24212), .X(n24211) );
  nand_x4_sg U68330 ( .A(n31876), .B(n49325), .X(n31745) );
  nand_x1_sg U68331 ( .A(n31878), .B(n25258), .X(n31876) );
  nor_x1_sg U68332 ( .A(n25258), .B(n31878), .X(n31877) );
  nand_x4_sg U68333 ( .A(n24240), .B(n50414), .X(n24114) );
  nand_x1_sg U68334 ( .A(n24242), .B(n9912), .X(n24240) );
  nor_x1_sg U68335 ( .A(n9912), .B(n24242), .X(n24241) );
  nand_x4_sg U68336 ( .A(n31906), .B(n49555), .X(n31780) );
  nand_x1_sg U68337 ( .A(n31908), .B(n25015), .X(n31906) );
  nor_x1_sg U68338 ( .A(n25015), .B(n31908), .X(n31907) );
  nand_x4_sg U68339 ( .A(n24252), .B(n50507), .X(n24128) );
  nand_x1_sg U68340 ( .A(n24254), .B(n9816), .X(n24252) );
  nor_x1_sg U68341 ( .A(n9816), .B(n24254), .X(n24253) );
  nand_x4_sg U68342 ( .A(n24246), .B(n50460), .X(n24121) );
  nand_x1_sg U68343 ( .A(n24248), .B(n9864), .X(n24246) );
  nor_x1_sg U68344 ( .A(n9864), .B(n24248), .X(n24247) );
  nand_x4_sg U68345 ( .A(n31918), .B(n49648), .X(n31794) );
  nand_x1_sg U68346 ( .A(n31920), .B(n24919), .X(n31918) );
  nor_x1_sg U68347 ( .A(n24919), .B(n31920), .X(n31919) );
  nand_x4_sg U68348 ( .A(n31912), .B(n49601), .X(n31787) );
  nand_x1_sg U68349 ( .A(n31914), .B(n24967), .X(n31912) );
  nor_x1_sg U68350 ( .A(n24967), .B(n31914), .X(n31913) );
  nand_x4_sg U68351 ( .A(n23177), .B(n50190), .X(n22932) );
  nand_x1_sg U68352 ( .A(n23179), .B(n10165), .X(n23177) );
  nor_x1_sg U68353 ( .A(n10165), .B(n23179), .X(n23178) );
  nand_x4_sg U68354 ( .A(n30843), .B(n49331), .X(n30598) );
  nand_x1_sg U68355 ( .A(n30845), .B(n25273), .X(n30843) );
  nor_x1_sg U68356 ( .A(n25273), .B(n30845), .X(n30844) );
  nand_x4_sg U68357 ( .A(n23231), .B(n50609), .X(n22995) );
  nand_x1_sg U68358 ( .A(n23233), .B(n9730), .X(n23231) );
  nor_x1_sg U68359 ( .A(n9730), .B(n23233), .X(n23232) );
  nand_x4_sg U68360 ( .A(n23195), .B(n50326), .X(n22953) );
  nand_x1_sg U68361 ( .A(n23197), .B(n10019), .X(n23195) );
  nor_x1_sg U68362 ( .A(n10019), .B(n23197), .X(n23196) );
  nand_x4_sg U68363 ( .A(n23183), .B(n50234), .X(n22939) );
  nand_x1_sg U68364 ( .A(n23185), .B(n10116), .X(n23183) );
  nor_x1_sg U68365 ( .A(n10116), .B(n23185), .X(n23184) );
  nand_x4_sg U68366 ( .A(n30897), .B(n49750), .X(n30661) );
  nand_x1_sg U68367 ( .A(n30899), .B(n24838), .X(n30897) );
  nor_x1_sg U68368 ( .A(n24838), .B(n30899), .X(n30898) );
  nand_x4_sg U68369 ( .A(n30861), .B(n49467), .X(n30619) );
  nand_x1_sg U68370 ( .A(n30863), .B(n25127), .X(n30861) );
  nor_x1_sg U68371 ( .A(n25127), .B(n30863), .X(n30862) );
  nand_x4_sg U68372 ( .A(n30849), .B(n49375), .X(n30605) );
  nand_x1_sg U68373 ( .A(n30851), .B(n25224), .X(n30849) );
  nor_x1_sg U68374 ( .A(n25224), .B(n30851), .X(n30850) );
  nand_x4_sg U68375 ( .A(n22336), .B(n50848), .X(n22162) );
  nand_x1_sg U68376 ( .A(n22338), .B(n9513), .X(n22336) );
  nor_x1_sg U68377 ( .A(n9513), .B(n22338), .X(n22337) );
  nand_x4_sg U68378 ( .A(n22330), .B(n50803), .X(n22155) );
  nand_x1_sg U68379 ( .A(n22332), .B(n9562), .X(n22330) );
  nor_x1_sg U68380 ( .A(n9562), .B(n22332), .X(n22331) );
  nand_x4_sg U68381 ( .A(n23249), .B(n50751), .X(n23016) );
  nand_x1_sg U68382 ( .A(n23251), .B(n9587), .X(n23249) );
  nor_x1_sg U68383 ( .A(n9587), .B(n23251), .X(n23250) );
  nand_x4_sg U68384 ( .A(n22324), .B(n50755), .X(n22148) );
  nand_x1_sg U68385 ( .A(n22326), .B(n9610), .X(n22324) );
  nor_x1_sg U68386 ( .A(n9610), .B(n22326), .X(n22325) );
  nand_x4_sg U68387 ( .A(n23243), .B(n50704), .X(n23009) );
  nand_x1_sg U68388 ( .A(n23245), .B(n9635), .X(n23243) );
  nor_x1_sg U68389 ( .A(n9635), .B(n23245), .X(n23244) );
  nand_x4_sg U68390 ( .A(n22318), .B(n50708), .X(n22141) );
  nand_x1_sg U68391 ( .A(n22320), .B(n9658), .X(n22318) );
  nor_x1_sg U68392 ( .A(n9658), .B(n22320), .X(n22319) );
  nand_x4_sg U68393 ( .A(n23237), .B(n50657), .X(n23002) );
  nand_x1_sg U68394 ( .A(n23239), .B(n9683), .X(n23237) );
  nor_x1_sg U68395 ( .A(n9683), .B(n23239), .X(n23238) );
  nand_x4_sg U68396 ( .A(n22312), .B(n50660), .X(n22134) );
  nand_x1_sg U68397 ( .A(n22314), .B(n9705), .X(n22312) );
  nor_x1_sg U68398 ( .A(n9705), .B(n22314), .X(n22313) );
  nand_x4_sg U68399 ( .A(n22306), .B(n50613), .X(n22127) );
  nand_x1_sg U68400 ( .A(n22308), .B(n9753), .X(n22306) );
  nor_x1_sg U68401 ( .A(n9753), .B(n22308), .X(n22307) );
  nand_x4_sg U68402 ( .A(n23225), .B(n50560), .X(n22988) );
  nand_x1_sg U68403 ( .A(n23227), .B(n9778), .X(n23225) );
  nor_x1_sg U68404 ( .A(n9778), .B(n23227), .X(n23226) );
  nand_x4_sg U68405 ( .A(n22300), .B(n50564), .X(n22120) );
  nand_x1_sg U68406 ( .A(n22302), .B(n9801), .X(n22300) );
  nor_x1_sg U68407 ( .A(n9801), .B(n22302), .X(n22301) );
  nand_x4_sg U68408 ( .A(n23219), .B(n50513), .X(n22981) );
  nand_x1_sg U68409 ( .A(n23221), .B(n9826), .X(n23219) );
  nor_x1_sg U68410 ( .A(n9826), .B(n23221), .X(n23220) );
  nand_x4_sg U68411 ( .A(n22294), .B(n50517), .X(n22113) );
  nand_x1_sg U68412 ( .A(n22296), .B(n9849), .X(n22294) );
  nor_x1_sg U68413 ( .A(n9849), .B(n22296), .X(n22295) );
  nand_x4_sg U68414 ( .A(n23213), .B(n50466), .X(n22974) );
  nand_x1_sg U68415 ( .A(n23215), .B(n9874), .X(n23213) );
  nor_x1_sg U68416 ( .A(n9874), .B(n23215), .X(n23214) );
  nand_x4_sg U68417 ( .A(n22288), .B(n50470), .X(n22106) );
  nand_x1_sg U68418 ( .A(n22290), .B(n9897), .X(n22288) );
  nor_x1_sg U68419 ( .A(n9897), .B(n22290), .X(n22289) );
  nand_x4_sg U68420 ( .A(n23207), .B(n50420), .X(n22967) );
  nand_x1_sg U68421 ( .A(n23209), .B(n9922), .X(n23207) );
  nor_x1_sg U68422 ( .A(n9922), .B(n23209), .X(n23208) );
  nand_x4_sg U68423 ( .A(n22282), .B(n50424), .X(n22099) );
  nand_x1_sg U68424 ( .A(n22284), .B(n9945), .X(n22282) );
  nor_x1_sg U68425 ( .A(n9945), .B(n22284), .X(n22283) );
  nand_x4_sg U68426 ( .A(n23201), .B(n50373), .X(n22960) );
  nand_x1_sg U68427 ( .A(n23203), .B(n9970), .X(n23201) );
  nor_x1_sg U68428 ( .A(n9970), .B(n23203), .X(n23202) );
  nand_x4_sg U68429 ( .A(n22276), .B(n50377), .X(n22092) );
  nand_x1_sg U68430 ( .A(n22278), .B(n9994), .X(n22276) );
  nor_x1_sg U68431 ( .A(n9994), .B(n22278), .X(n22277) );
  nand_x4_sg U68432 ( .A(n22270), .B(n50330), .X(n22085) );
  nand_x1_sg U68433 ( .A(n22272), .B(n10042), .X(n22270) );
  nor_x1_sg U68434 ( .A(n10042), .B(n22272), .X(n22271) );
  nand_x4_sg U68435 ( .A(n23189), .B(n50280), .X(n22946) );
  nand_x1_sg U68436 ( .A(n23191), .B(n10067), .X(n23189) );
  nor_x1_sg U68437 ( .A(n10067), .B(n23191), .X(n23190) );
  nand_x4_sg U68438 ( .A(n22264), .B(n50284), .X(n22078) );
  nand_x1_sg U68439 ( .A(n22266), .B(n10091), .X(n22264) );
  nor_x1_sg U68440 ( .A(n10091), .B(n22266), .X(n22265) );
  nand_x4_sg U68441 ( .A(n22258), .B(n50238), .X(n22071) );
  nand_x1_sg U68442 ( .A(n22260), .B(n10140), .X(n22258) );
  nor_x1_sg U68443 ( .A(n10140), .B(n22260), .X(n22259) );
  nand_x4_sg U68444 ( .A(n22252), .B(n50194), .X(n22064) );
  nand_x1_sg U68445 ( .A(n22254), .B(n10187), .X(n22252) );
  nor_x1_sg U68446 ( .A(n10187), .B(n22254), .X(n22253) );
  nand_x4_sg U68447 ( .A(n30001), .B(n49989), .X(n29827) );
  nand_x1_sg U68448 ( .A(n30003), .B(n24621), .X(n30001) );
  nor_x1_sg U68449 ( .A(n24621), .B(n30003), .X(n30002) );
  nand_x4_sg U68450 ( .A(n29995), .B(n49944), .X(n29820) );
  nand_x1_sg U68451 ( .A(n29997), .B(n24670), .X(n29995) );
  nor_x1_sg U68452 ( .A(n24670), .B(n29997), .X(n29996) );
  nand_x4_sg U68453 ( .A(n30915), .B(n49892), .X(n30682) );
  nand_x1_sg U68454 ( .A(n30917), .B(n24695), .X(n30915) );
  nor_x1_sg U68455 ( .A(n24695), .B(n30917), .X(n30916) );
  nand_x4_sg U68456 ( .A(n29989), .B(n49896), .X(n29813) );
  nand_x1_sg U68457 ( .A(n29991), .B(n24718), .X(n29989) );
  nor_x1_sg U68458 ( .A(n24718), .B(n29991), .X(n29990) );
  nand_x4_sg U68459 ( .A(n30909), .B(n49845), .X(n30675) );
  nand_x1_sg U68460 ( .A(n30911), .B(n24743), .X(n30909) );
  nor_x1_sg U68461 ( .A(n24743), .B(n30911), .X(n30910) );
  nand_x4_sg U68462 ( .A(n29983), .B(n49849), .X(n29806) );
  nand_x1_sg U68463 ( .A(n29985), .B(n24766), .X(n29983) );
  nor_x1_sg U68464 ( .A(n24766), .B(n29985), .X(n29984) );
  nand_x4_sg U68465 ( .A(n30903), .B(n49798), .X(n30668) );
  nand_x1_sg U68466 ( .A(n30905), .B(n24791), .X(n30903) );
  nor_x1_sg U68467 ( .A(n24791), .B(n30905), .X(n30904) );
  nand_x4_sg U68468 ( .A(n29977), .B(n49801), .X(n29799) );
  nand_x1_sg U68469 ( .A(n29979), .B(n24813), .X(n29977) );
  nor_x1_sg U68470 ( .A(n24813), .B(n29979), .X(n29978) );
  nand_x4_sg U68471 ( .A(n29971), .B(n49754), .X(n29792) );
  nand_x1_sg U68472 ( .A(n29973), .B(n24861), .X(n29971) );
  nor_x1_sg U68473 ( .A(n24861), .B(n29973), .X(n29972) );
  nand_x4_sg U68474 ( .A(n30891), .B(n49701), .X(n30654) );
  nand_x1_sg U68475 ( .A(n30893), .B(n24886), .X(n30891) );
  nor_x1_sg U68476 ( .A(n24886), .B(n30893), .X(n30892) );
  nand_x4_sg U68477 ( .A(n29965), .B(n49705), .X(n29785) );
  nand_x1_sg U68478 ( .A(n29967), .B(n24909), .X(n29965) );
  nor_x1_sg U68479 ( .A(n24909), .B(n29967), .X(n29966) );
  nand_x4_sg U68480 ( .A(n30885), .B(n49654), .X(n30647) );
  nand_x1_sg U68481 ( .A(n30887), .B(n24934), .X(n30885) );
  nor_x1_sg U68482 ( .A(n24934), .B(n30887), .X(n30886) );
  nand_x4_sg U68483 ( .A(n29959), .B(n49658), .X(n29778) );
  nand_x1_sg U68484 ( .A(n29961), .B(n24957), .X(n29959) );
  nor_x1_sg U68485 ( .A(n24957), .B(n29961), .X(n29960) );
  nand_x4_sg U68486 ( .A(n30879), .B(n49607), .X(n30640) );
  nand_x1_sg U68487 ( .A(n30881), .B(n24982), .X(n30879) );
  nor_x1_sg U68488 ( .A(n24982), .B(n30881), .X(n30880) );
  nand_x4_sg U68489 ( .A(n29953), .B(n49611), .X(n29771) );
  nand_x1_sg U68490 ( .A(n29955), .B(n25005), .X(n29953) );
  nor_x1_sg U68491 ( .A(n25005), .B(n29955), .X(n29954) );
  nand_x4_sg U68492 ( .A(n30873), .B(n49561), .X(n30633) );
  nand_x1_sg U68493 ( .A(n30875), .B(n25030), .X(n30873) );
  nor_x1_sg U68494 ( .A(n25030), .B(n30875), .X(n30874) );
  nand_x4_sg U68495 ( .A(n29947), .B(n49565), .X(n29764) );
  nand_x1_sg U68496 ( .A(n29949), .B(n25053), .X(n29947) );
  nor_x1_sg U68497 ( .A(n25053), .B(n29949), .X(n29948) );
  nand_x4_sg U68498 ( .A(n30867), .B(n49514), .X(n30626) );
  nand_x1_sg U68499 ( .A(n30869), .B(n25078), .X(n30867) );
  nor_x1_sg U68500 ( .A(n25078), .B(n30869), .X(n30868) );
  nand_x4_sg U68501 ( .A(n29941), .B(n49518), .X(n29757) );
  nand_x1_sg U68502 ( .A(n29943), .B(n25102), .X(n29941) );
  nor_x1_sg U68503 ( .A(n25102), .B(n29943), .X(n29942) );
  nand_x4_sg U68504 ( .A(n29935), .B(n49471), .X(n29750) );
  nand_x1_sg U68505 ( .A(n29937), .B(n25150), .X(n29935) );
  nor_x1_sg U68506 ( .A(n25150), .B(n29937), .X(n29936) );
  nand_x4_sg U68507 ( .A(n30855), .B(n49421), .X(n30612) );
  nand_x1_sg U68508 ( .A(n30857), .B(n25175), .X(n30855) );
  nor_x1_sg U68509 ( .A(n25175), .B(n30857), .X(n30856) );
  nand_x4_sg U68510 ( .A(n29929), .B(n49425), .X(n29743) );
  nand_x1_sg U68511 ( .A(n29931), .B(n25199), .X(n29929) );
  nor_x1_sg U68512 ( .A(n25199), .B(n29931), .X(n29930) );
  nand_x4_sg U68513 ( .A(n29923), .B(n49379), .X(n29736) );
  nand_x1_sg U68514 ( .A(n29925), .B(n25248), .X(n29923) );
  nor_x1_sg U68515 ( .A(n25248), .B(n29925), .X(n29924) );
  nand_x4_sg U68516 ( .A(n29917), .B(n49335), .X(n29729) );
  nand_x1_sg U68517 ( .A(n29919), .B(n25295), .X(n29917) );
  nor_x1_sg U68518 ( .A(n25295), .B(n29919), .X(n29918) );
  nand_x2_sg U68519 ( .A(n23061), .B(n22809), .X(n23059) );
  nor_x1_sg U68520 ( .A(n23061), .B(n22809), .X(n23060) );
  nand_x2_sg U68521 ( .A(n23492), .B(n23290), .X(n23490) );
  nor_x1_sg U68522 ( .A(n23492), .B(n23290), .X(n23491) );
  nand_x2_sg U68523 ( .A(n23853), .B(n23685), .X(n23851) );
  nor_x1_sg U68524 ( .A(n23853), .B(n23685), .X(n23852) );
  nand_x2_sg U68525 ( .A(n24150), .B(n24009), .X(n24148) );
  nor_x1_sg U68526 ( .A(n24150), .B(n24009), .X(n24149) );
  nand_x2_sg U68527 ( .A(n24446), .B(n24372), .X(n24444) );
  nor_x1_sg U68528 ( .A(n24446), .B(n24372), .X(n24445) );
  nand_x2_sg U68529 ( .A(n32112), .B(n32038), .X(n32110) );
  nor_x1_sg U68530 ( .A(n32112), .B(n32038), .X(n32111) );
  nand_x2_sg U68531 ( .A(n30727), .B(n30475), .X(n30725) );
  nor_x1_sg U68532 ( .A(n30727), .B(n30475), .X(n30726) );
  nand_x2_sg U68533 ( .A(n31158), .B(n30956), .X(n31156) );
  nor_x1_sg U68534 ( .A(n31158), .B(n30956), .X(n31157) );
  nand_x2_sg U68535 ( .A(n31519), .B(n31351), .X(n31517) );
  nor_x1_sg U68536 ( .A(n31519), .B(n31351), .X(n31518) );
  nand_x2_sg U68537 ( .A(n31816), .B(n31675), .X(n31814) );
  nor_x1_sg U68538 ( .A(n31816), .B(n31675), .X(n31815) );
  nand_x2_sg U68539 ( .A(n24368), .B(n24269), .X(n24366) );
  nor_x1_sg U68540 ( .A(n24368), .B(n24269), .X(n24367) );
  nand_x2_sg U68541 ( .A(n32034), .B(n31935), .X(n32032) );
  nor_x1_sg U68542 ( .A(n32034), .B(n31935), .X(n32033) );
  nand_x2_sg U68543 ( .A(n25328), .B(n49275), .X(n31250) );
  nand_x2_sg U68544 ( .A(n31251), .B(n49287), .X(n31249) );
  nand_x2_sg U68545 ( .A(n10220), .B(n50134), .X(n23584) );
  nand_x2_sg U68546 ( .A(n23585), .B(n50146), .X(n23583) );
  nand_x2_sg U68547 ( .A(n25557), .B(n25559), .X(n25641) );
  nand_x2_sg U68548 ( .A(n28352), .B(n28354), .X(n28434) );
  nand_x2_sg U68549 ( .A(n28909), .B(n28911), .X(n28991) );
  nand_x2_sg U68550 ( .A(n29470), .B(n29472), .X(n29552) );
  nand_x2_sg U68551 ( .A(n25616), .B(n25618), .X(n25634) );
  nand_x2_sg U68552 ( .A(n27572), .B(n27574), .X(n27588) );
  nand_x2_sg U68553 ( .A(n25897), .B(n25899), .X(n25913) );
  nand_x2_sg U68554 ( .A(n26177), .B(n26179), .X(n26193) );
  nand_x2_sg U68555 ( .A(n26456), .B(n26458), .X(n26472) );
  nand_x2_sg U68556 ( .A(n26734), .B(n26736), .X(n26750) );
  nand_x2_sg U68557 ( .A(n27013), .B(n27015), .X(n27029) );
  nand_x2_sg U68558 ( .A(n27293), .B(n27295), .X(n27309) );
  nand_x2_sg U68559 ( .A(n27851), .B(n27853), .X(n27867) );
  nand_x2_sg U68560 ( .A(n28132), .B(n28134), .X(n28148) );
  nand_x2_sg U68561 ( .A(n28411), .B(n28413), .X(n28427) );
  nand_x2_sg U68562 ( .A(n28690), .B(n28692), .X(n28706) );
  nand_x2_sg U68563 ( .A(n28968), .B(n28970), .X(n28984) );
  nand_x2_sg U68564 ( .A(n29251), .B(n29253), .X(n29267) );
  nand_x2_sg U68565 ( .A(n29529), .B(n29531), .X(n29545) );
  nor_x1_sg U68566 ( .A(n21959), .B(n22503), .X(n22502) );
  nor_x1_sg U68567 ( .A(n29618), .B(n30169), .X(n30168) );
  nor_x1_sg U68568 ( .A(n21937), .B(n22521), .X(n22520) );
  nor_x1_sg U68569 ( .A(n29588), .B(n30187), .X(n30186) );
  nand_x4_sg U68570 ( .A(n50318), .B(n24426), .X(n24339) );
  nand_x1_sg U68571 ( .A(n41927), .B(n24428), .X(n24426) );
  nor_x1_sg U68572 ( .A(n41927), .B(n24428), .X(n24429) );
  nand_x4_sg U68573 ( .A(n49459), .B(n32092), .X(n32005) );
  nand_x1_sg U68574 ( .A(n41935), .B(n32094), .X(n32092) );
  nor_x1_sg U68575 ( .A(n41935), .B(n32094), .X(n32095) );
  nor_x1_sg U68576 ( .A(n44100), .B(n21968), .X(n22515) );
  nor_x1_sg U68577 ( .A(n44098), .B(n29631), .X(n30181) );
  nand_x2_sg U68578 ( .A(n41648), .B(n11693), .X(n25910) );
  nand_x2_sg U68579 ( .A(n41646), .B(n12472), .X(n26190) );
  nand_x2_sg U68580 ( .A(n41644), .B(n13253), .X(n26469) );
  nand_x2_sg U68581 ( .A(n41642), .B(n14033), .X(n26747) );
  nand_x2_sg U68582 ( .A(n41640), .B(n14805), .X(n27026) );
  nand_x2_sg U68583 ( .A(n41638), .B(n15586), .X(n27306) );
  nand_x2_sg U68584 ( .A(n41622), .B(n16367), .X(n27585) );
  nand_x2_sg U68585 ( .A(n41636), .B(n17152), .X(n27864) );
  nand_x2_sg U68586 ( .A(n41634), .B(n17926), .X(n28145) );
  nand_x2_sg U68587 ( .A(n41632), .B(n18695), .X(n28424) );
  nand_x2_sg U68588 ( .A(n41630), .B(n19471), .X(n28703) );
  nand_x2_sg U68589 ( .A(n41628), .B(n20241), .X(n28981) );
  nand_x2_sg U68590 ( .A(n41626), .B(n21015), .X(n29264) );
  nand_x2_sg U68591 ( .A(n41624), .B(n21786), .X(n29542) );
  nor_x1_sg U68592 ( .A(n45371), .B(n21940), .X(n22518) );
  nor_x1_sg U68593 ( .A(n45361), .B(n29592), .X(n30184) );
  nand_x4_sg U68594 ( .A(n24402), .B(n24403), .X(n24312) );
  nand_x1_sg U68595 ( .A(n50140), .B(n24404), .X(n24403) );
  nand_x1_sg U68596 ( .A(n24405), .B(n50108), .X(n24402) );
  nand_x4_sg U68597 ( .A(n32068), .B(n32069), .X(n31978) );
  nand_x1_sg U68598 ( .A(n49281), .B(n32070), .X(n32069) );
  nand_x1_sg U68599 ( .A(n32071), .B(n49249), .X(n32068) );
  nand_x4_sg U68600 ( .A(n24438), .B(n24439), .X(n24352) );
  nand_x1_sg U68601 ( .A(n24440), .B(n24441), .X(n24439) );
  nand_x4_sg U68602 ( .A(n32104), .B(n32105), .X(n32018) );
  nand_x1_sg U68603 ( .A(n32106), .B(n32107), .X(n32105) );
  nand_x4_sg U68604 ( .A(n51305), .B(n25567), .X(n10490) );
  nand_x1_sg U68605 ( .A(n42172), .B(n25569), .X(n25567) );
  nand_x4_sg U68606 ( .A(n51866), .B(n26128), .X(n12043) );
  nand_x1_sg U68607 ( .A(n42184), .B(n26130), .X(n26128) );
  nand_x4_sg U68608 ( .A(n53252), .B(n27523), .X(n15938) );
  nand_x1_sg U68609 ( .A(n42168), .B(n27525), .X(n27523) );
  nand_x4_sg U68610 ( .A(n54659), .B(n28919), .X(n19817) );
  nand_x1_sg U68611 ( .A(n42180), .B(n28921), .X(n28919) );
  nand_x4_sg U68612 ( .A(n55227), .B(n29480), .X(n21362) );
  nand_x1_sg U68613 ( .A(n42176), .B(n29482), .X(n29480) );
  nand_x4_sg U68614 ( .A(n52418), .B(n26685), .X(n13604) );
  nand_x1_sg U68615 ( .A(n42148), .B(n26687), .X(n26685) );
  nand_x4_sg U68616 ( .A(n46576), .B(n29016), .X(n28739) );
  nand_x1_sg U68617 ( .A(n29017), .B(n55460), .X(n29016) );
  nor_x1_sg U68618 ( .A(n55780), .B(n29018), .X(n29017) );
  nand_x1_sg U68619 ( .A(n43163), .B(n44321), .X(n26964) );
  nand_x4_sg U68620 ( .A(n28956), .B(n28957), .X(n19610) );
  nand_x1_sg U68621 ( .A(n54608), .B(n28958), .X(n28957) );
  nand_x1_sg U68622 ( .A(n28959), .B(n54606), .X(n28956) );
  nand_x4_sg U68623 ( .A(n29517), .B(n29518), .X(n21155) );
  nand_x1_sg U68624 ( .A(n55176), .B(n29519), .X(n29518) );
  nand_x1_sg U68625 ( .A(n29520), .B(n55174), .X(n29517) );
  nand_x4_sg U68626 ( .A(n27001), .B(n27002), .X(n14174) );
  nand_x1_sg U68627 ( .A(n52642), .B(n27003), .X(n27002) );
  nand_x1_sg U68628 ( .A(n27004), .B(n52640), .X(n27001) );
  nand_x4_sg U68629 ( .A(n28120), .B(n28121), .X(n17293) );
  nand_x1_sg U68630 ( .A(n53759), .B(n28122), .X(n28121) );
  nand_x1_sg U68631 ( .A(n28123), .B(n53757), .X(n28120) );
  nand_x4_sg U68632 ( .A(n28399), .B(n28400), .X(n18065) );
  nand_x1_sg U68633 ( .A(n54043), .B(n28401), .X(n28400) );
  nand_x1_sg U68634 ( .A(n28402), .B(n54041), .X(n28399) );
  nand_x4_sg U68635 ( .A(n28678), .B(n28679), .X(n18838) );
  nand_x1_sg U68636 ( .A(n54324), .B(n28680), .X(n28679) );
  nand_x1_sg U68637 ( .A(n28681), .B(n54322), .X(n28678) );
  nand_x4_sg U68638 ( .A(n29239), .B(n29240), .X(n20382) );
  nand_x1_sg U68639 ( .A(n54892), .B(n29241), .X(n29240) );
  nand_x1_sg U68640 ( .A(n29242), .B(n54890), .X(n29239) );
  nand_x4_sg U68641 ( .A(n26165), .B(n26166), .X(n11833) );
  nand_x1_sg U68642 ( .A(n51813), .B(n26167), .X(n26166) );
  nand_x1_sg U68643 ( .A(n26168), .B(n51811), .X(n26165) );
  nand_x4_sg U68644 ( .A(n27560), .B(n27561), .X(n15728) );
  nand_x1_sg U68645 ( .A(n53201), .B(n27562), .X(n27561) );
  nand_x1_sg U68646 ( .A(n27563), .B(n53199), .X(n27560) );
  nor_x1_sg U68647 ( .A(n22491), .B(n9544), .X(n22627) );
  nor_x1_sg U68648 ( .A(n30156), .B(n24652), .X(n30293) );
  nor_x1_sg U68649 ( .A(n22497), .B(n9495), .X(n22624) );
  nor_x1_sg U68650 ( .A(n30162), .B(n24603), .X(n30290) );
  nor_x1_sg U68651 ( .A(n22350), .B(n9446), .X(n22621) );
  nor_x1_sg U68652 ( .A(n30015), .B(n24554), .X(n30287) );
  nor_x1_sg U68653 ( .A(n22184), .B(n9391), .X(n22618) );
  nor_x1_sg U68654 ( .A(n29849), .B(n24505), .X(n30284) );
  nor_x1_sg U68655 ( .A(n22473), .B(n9688), .X(n22636) );
  nor_x1_sg U68656 ( .A(n22467), .B(n9735), .X(n22639) );
  nor_x1_sg U68657 ( .A(n22461), .B(n9783), .X(n22642) );
  nor_x1_sg U68658 ( .A(n22455), .B(n9831), .X(n22645) );
  nor_x1_sg U68659 ( .A(n22449), .B(n9879), .X(n22648) );
  nor_x1_sg U68660 ( .A(n22443), .B(n9927), .X(n22651) );
  nor_x1_sg U68661 ( .A(n22437), .B(n9975), .X(n22654) );
  nor_x1_sg U68662 ( .A(n22431), .B(n10024), .X(n22657) );
  nor_x1_sg U68663 ( .A(n22425), .B(n10072), .X(n22660) );
  nor_x1_sg U68664 ( .A(n22419), .B(n10121), .X(n22663) );
  nor_x1_sg U68665 ( .A(n22413), .B(n10170), .X(n22666) );
  nor_x1_sg U68666 ( .A(n30138), .B(n24796), .X(n30302) );
  nor_x1_sg U68667 ( .A(n30132), .B(n24843), .X(n30305) );
  nor_x1_sg U68668 ( .A(n30126), .B(n24891), .X(n30308) );
  nor_x1_sg U68669 ( .A(n30120), .B(n24939), .X(n30311) );
  nor_x1_sg U68670 ( .A(n30114), .B(n24987), .X(n30314) );
  nor_x1_sg U68671 ( .A(n30108), .B(n25035), .X(n30317) );
  nor_x1_sg U68672 ( .A(n30102), .B(n25083), .X(n30320) );
  nor_x1_sg U68673 ( .A(n30096), .B(n25132), .X(n30323) );
  nor_x1_sg U68674 ( .A(n30090), .B(n25180), .X(n30326) );
  nor_x1_sg U68675 ( .A(n30084), .B(n25229), .X(n30329) );
  nor_x1_sg U68676 ( .A(n30078), .B(n25278), .X(n30332) );
  nor_x1_sg U68677 ( .A(n22479), .B(n9640), .X(n22633) );
  nor_x1_sg U68678 ( .A(n30144), .B(n24748), .X(n30299) );
  nor_x1_sg U68679 ( .A(n22485), .B(n9592), .X(n22630) );
  nor_x1_sg U68680 ( .A(n30150), .B(n24700), .X(n30296) );
  nor_x1_sg U68681 ( .A(n23805), .B(n9911), .X(n23905) );
  nor_x1_sg U68682 ( .A(n23799), .B(n9959), .X(n23908) );
  nor_x1_sg U68683 ( .A(n31483), .B(n24923), .X(n31565) );
  nor_x1_sg U68684 ( .A(n31477), .B(n24971), .X(n31568) );
  nor_x1_sg U68685 ( .A(n31471), .B(n25019), .X(n31571) );
  nor_x1_sg U68686 ( .A(n31465), .B(n25067), .X(n31574) );
  nor_x1_sg U68687 ( .A(n31459), .B(n25116), .X(n31577) );
  nor_x1_sg U68688 ( .A(n31453), .B(n25164), .X(n31580) );
  nor_x1_sg U68689 ( .A(n31447), .B(n25213), .X(n31583) );
  nor_x1_sg U68690 ( .A(n31441), .B(n25262), .X(n31586) );
  nor_x1_sg U68691 ( .A(n23811), .B(n9863), .X(n23902) );
  nor_x1_sg U68692 ( .A(n23787), .B(n10056), .X(n23914) );
  nor_x1_sg U68693 ( .A(n23817), .B(n9815), .X(n23899) );
  nor_x1_sg U68694 ( .A(n23793), .B(n10008), .X(n23911) );
  nor_x1_sg U68695 ( .A(n23781), .B(n10105), .X(n23917) );
  nor_x1_sg U68696 ( .A(n23775), .B(n10154), .X(n23920) );
  nor_x1_sg U68697 ( .A(n22844), .B(n9429), .X(n22843) );
  nor_x1_sg U68698 ( .A(n30510), .B(n24537), .X(n30509) );
  nor_x1_sg U68699 ( .A(n30991), .B(n24635), .X(n30990) );
  nor_x1_sg U68700 ( .A(n31386), .B(n24732), .X(n31385) );
  nor_x1_sg U68701 ( .A(n31495), .B(n24827), .X(n31559) );
  nor_x1_sg U68702 ( .A(n9370), .B(n22576), .X(n22575) );
  nor_x1_sg U68703 ( .A(n24487), .B(n30242), .X(n30241) );
  nor_x1_sg U68704 ( .A(n30765), .B(n24586), .X(n30764) );
  nor_x1_sg U68705 ( .A(n31196), .B(n24684), .X(n31195) );
  nor_x1_sg U68706 ( .A(n31501), .B(n24780), .X(n31556) );
  nor_x1_sg U68707 ( .A(n31489), .B(n24875), .X(n31562) );
  nor_x1_sg U68708 ( .A(n23325), .B(n9527), .X(n23324) );
  nor_x1_sg U68709 ( .A(n23720), .B(n9624), .X(n23719) );
  nor_x1_sg U68710 ( .A(n23829), .B(n9719), .X(n23893) );
  nor_x1_sg U68711 ( .A(n23099), .B(n9478), .X(n23098) );
  nor_x1_sg U68712 ( .A(n23530), .B(n9576), .X(n23529) );
  nor_x1_sg U68713 ( .A(n23835), .B(n9672), .X(n23890) );
  nor_x1_sg U68714 ( .A(n23823), .B(n9767), .X(n23896) );
  nand_x4_sg U68715 ( .A(n25854), .B(n51575), .X(n11240) );
  nand_x1_sg U68716 ( .A(n28370), .B(n54067), .X(n28369) );
  nand_x4_sg U68717 ( .A(n26976), .B(n26977), .X(n14356) );
  nand_x1_sg U68718 ( .A(n26978), .B(n52660), .X(n26977) );
  nand_x4_sg U68719 ( .A(n26982), .B(n26983), .X(n14300) );
  nand_x1_sg U68720 ( .A(n26984), .B(n52652), .X(n26983) );
  nand_x4_sg U68721 ( .A(n26140), .B(n26141), .X(n12061) );
  nand_x1_sg U68722 ( .A(n26142), .B(n51831), .X(n26141) );
  nand_x4_sg U68723 ( .A(n26697), .B(n26698), .X(n13622) );
  nand_x1_sg U68724 ( .A(n26699), .B(n52383), .X(n26698) );
  nand_x4_sg U68725 ( .A(n26703), .B(n26704), .X(n13518) );
  nand_x1_sg U68726 ( .A(n26705), .B(n52375), .X(n26704) );
  nand_x4_sg U68727 ( .A(n27541), .B(n27542), .X(n15852) );
  nand_x1_sg U68728 ( .A(n27543), .B(n53211), .X(n27542) );
  nand_x4_sg U68729 ( .A(n26146), .B(n26147), .X(n11957) );
  nand_x1_sg U68730 ( .A(n26148), .B(n51823), .X(n26147) );
  nand_x4_sg U68731 ( .A(n25579), .B(n25580), .X(n10464) );
  nand_x1_sg U68732 ( .A(n25581), .B(n51271), .X(n25580) );
  nand_x4_sg U68733 ( .A(n28931), .B(n28932), .X(n19791) );
  nand_x1_sg U68734 ( .A(n28933), .B(n54625), .X(n28932) );
  nand_x4_sg U68735 ( .A(n29492), .B(n29493), .X(n21336) );
  nand_x1_sg U68736 ( .A(n29494), .B(n55193), .X(n29493) );
  nand_x4_sg U68737 ( .A(n27535), .B(n27536), .X(n15956) );
  nand_x1_sg U68738 ( .A(n27537), .B(n53219), .X(n27536) );
  nand_x4_sg U68739 ( .A(n28101), .B(n28102), .X(n17417) );
  nand_x4_sg U68740 ( .A(n28659), .B(n28660), .X(n18962) );
  nand_x4_sg U68741 ( .A(n29220), .B(n29221), .X(n20506) );
  nand_x4_sg U68742 ( .A(n28107), .B(n28108), .X(n17408) );
  nand_x4_sg U68743 ( .A(n28665), .B(n28666), .X(n18953) );
  nand_x4_sg U68744 ( .A(n28943), .B(n28944), .X(n19724) );
  nand_x4_sg U68745 ( .A(n29226), .B(n29227), .X(n20497) );
  nand_x4_sg U68746 ( .A(n29504), .B(n29505), .X(n21269) );
  nand_x4_sg U68747 ( .A(n25591), .B(n25592), .X(n10397) );
  nand_x4_sg U68748 ( .A(n28374), .B(n28375), .X(n18246) );
  nand_x4_sg U68749 ( .A(n23170), .B(n23171), .X(n22924) );
  nand_x1_sg U68750 ( .A(n23173), .B(n50148), .X(n23170) );
  nand_x4_sg U68751 ( .A(n30836), .B(n30837), .X(n30590) );
  nand_x1_sg U68752 ( .A(n30839), .B(n49289), .X(n30836) );
  nand_x4_sg U68753 ( .A(n22245), .B(n22246), .X(n22056) );
  nand_x1_sg U68754 ( .A(n22248), .B(n50152), .X(n22245) );
  nand_x4_sg U68755 ( .A(n29910), .B(n29911), .X(n29721) );
  nand_x1_sg U68756 ( .A(n29913), .B(n49293), .X(n29910) );
  nand_x4_sg U68757 ( .A(n24408), .B(n24409), .X(n24320) );
  nand_x1_sg U68758 ( .A(n50182), .B(n50179), .X(n24409) );
  nand_x4_sg U68759 ( .A(n32074), .B(n32075), .X(n31986) );
  nand_x1_sg U68760 ( .A(n49323), .B(n49320), .X(n32075) );
  nand_x4_sg U68761 ( .A(n26122), .B(n26123), .X(n12070) );
  nand_x4_sg U68762 ( .A(n26679), .B(n26680), .X(n13631) );
  nand_x4_sg U68763 ( .A(n27517), .B(n27518), .X(n15965) );
  nand_x4_sg U68764 ( .A(n25561), .B(n25562), .X(n10519) );
  nand_x4_sg U68765 ( .A(n28913), .B(n28914), .X(n19846) );
  nand_x4_sg U68766 ( .A(n29474), .B(n29475), .X(n21391) );
  nand_x4_sg U68767 ( .A(n24203), .B(n24204), .X(n24071) );
  nand_x1_sg U68768 ( .A(n24206), .B(n50142), .X(n24203) );
  nand_x4_sg U68769 ( .A(n31869), .B(n31870), .X(n31737) );
  nand_x1_sg U68770 ( .A(n31872), .B(n49283), .X(n31869) );
  nand_x4_sg U68771 ( .A(n28356), .B(n28357), .X(n18301) );
  nand_x4_sg U68772 ( .A(n25842), .B(n25843), .X(n11290) );
  nand_x4_sg U68773 ( .A(n26401), .B(n26402), .X(n12851) );
  nand_x4_sg U68774 ( .A(n27238), .B(n27239), .X(n15184) );
  nand_x4_sg U68775 ( .A(n27796), .B(n27797), .X(n16750) );
  nand_x4_sg U68776 ( .A(n25543), .B(n25544), .X(n25542) );
  nand_x4_sg U68777 ( .A(n25553), .B(n25554), .X(n25552) );
  nand_x4_sg U68778 ( .A(n28348), .B(n28349), .X(n28347) );
  nand_x4_sg U68779 ( .A(n28905), .B(n28906), .X(n28904) );
  nand_x4_sg U68780 ( .A(n29466), .B(n29467), .X(n29465) );
  nand_x4_sg U68781 ( .A(n25840), .B(n25841), .X(n25839) );
  nand_x4_sg U68782 ( .A(n26399), .B(n26400), .X(n26398) );
  nand_x4_sg U68783 ( .A(n26956), .B(n26957), .X(n26955) );
  nand_x4_sg U68784 ( .A(n27236), .B(n27237), .X(n27235) );
  nand_x4_sg U68785 ( .A(n27794), .B(n27795), .X(n27793) );
  nand_x4_sg U68786 ( .A(n28075), .B(n28076), .X(n28074) );
  nand_x4_sg U68787 ( .A(n28633), .B(n28634), .X(n28632) );
  nand_x4_sg U68788 ( .A(n29194), .B(n29195), .X(n29193) );
  nand_x4_sg U68789 ( .A(n25612), .B(n25613), .X(n25611) );
  nand_x4_sg U68790 ( .A(n27568), .B(n27569), .X(n27567) );
  nand_x4_sg U68791 ( .A(n25893), .B(n25894), .X(n25892) );
  nand_x4_sg U68792 ( .A(n26173), .B(n26174), .X(n26172) );
  nand_x4_sg U68793 ( .A(n26084), .B(n26085), .X(n26083) );
  nand_x4_sg U68794 ( .A(n26452), .B(n26453), .X(n26451) );
  nand_x4_sg U68795 ( .A(n26363), .B(n26364), .X(n26362) );
  nand_x4_sg U68796 ( .A(n26730), .B(n26731), .X(n26729) );
  nand_x4_sg U68797 ( .A(n26641), .B(n26642), .X(n26640) );
  nand_x4_sg U68798 ( .A(n27009), .B(n27010), .X(n27008) );
  nand_x4_sg U68799 ( .A(n27289), .B(n27290), .X(n27288) );
  nand_x4_sg U68800 ( .A(n27200), .B(n27201), .X(n27199) );
  nand_x4_sg U68801 ( .A(n27847), .B(n27848), .X(n27846) );
  nand_x4_sg U68802 ( .A(n27758), .B(n27759), .X(n27757) );
  nand_x4_sg U68803 ( .A(n28128), .B(n28129), .X(n28127) );
  nand_x4_sg U68804 ( .A(n28407), .B(n28408), .X(n28406) );
  nand_x4_sg U68805 ( .A(n28686), .B(n28687), .X(n28685) );
  nand_x4_sg U68806 ( .A(n28964), .B(n28965), .X(n28963) );
  nand_x4_sg U68807 ( .A(n29247), .B(n29248), .X(n29246) );
  nand_x4_sg U68808 ( .A(n29525), .B(n29526), .X(n29524) );
  nand_x4_sg U68809 ( .A(n25559), .B(n25560), .X(n25558) );
  nand_x4_sg U68810 ( .A(n25549), .B(n25550), .X(n25548) );
  nand_x4_sg U68811 ( .A(n25537), .B(n25538), .X(n25536) );
  nand_x4_sg U68812 ( .A(n25531), .B(n25532), .X(n25530) );
  nand_x4_sg U68813 ( .A(n25834), .B(n25835), .X(n25833) );
  nand_x4_sg U68814 ( .A(n25828), .B(n25829), .X(n25827) );
  nand_x4_sg U68815 ( .A(n25822), .B(n25823), .X(n25821) );
  nand_x4_sg U68816 ( .A(n25816), .B(n25817), .X(n25815) );
  nand_x4_sg U68817 ( .A(n25810), .B(n25811), .X(n25809) );
  nand_x4_sg U68818 ( .A(n26120), .B(n26121), .X(n26119) );
  nand_x4_sg U68819 ( .A(n26114), .B(n26115), .X(n26113) );
  nand_x4_sg U68820 ( .A(n26108), .B(n26109), .X(n26107) );
  nand_x4_sg U68821 ( .A(n26102), .B(n26103), .X(n26101) );
  nand_x4_sg U68822 ( .A(n26096), .B(n26097), .X(n26095) );
  nand_x4_sg U68823 ( .A(n26090), .B(n26091), .X(n26089) );
  nand_x4_sg U68824 ( .A(n26393), .B(n26394), .X(n26392) );
  nand_x4_sg U68825 ( .A(n26387), .B(n26388), .X(n26386) );
  nand_x4_sg U68826 ( .A(n26381), .B(n26382), .X(n26380) );
  nand_x4_sg U68827 ( .A(n26375), .B(n26376), .X(n26374) );
  nand_x4_sg U68828 ( .A(n26369), .B(n26370), .X(n26368) );
  nand_x4_sg U68829 ( .A(n26677), .B(n26678), .X(n26676) );
  nand_x4_sg U68830 ( .A(n26671), .B(n26672), .X(n26670) );
  nand_x4_sg U68831 ( .A(n26665), .B(n26666), .X(n26664) );
  nand_x4_sg U68832 ( .A(n26659), .B(n26660), .X(n26658) );
  nand_x4_sg U68833 ( .A(n26653), .B(n26654), .X(n26652) );
  nand_x4_sg U68834 ( .A(n26647), .B(n26648), .X(n26646) );
  nand_x4_sg U68835 ( .A(n26950), .B(n26951), .X(n26949) );
  nand_x4_sg U68836 ( .A(n26944), .B(n26945), .X(n26943) );
  nand_x4_sg U68837 ( .A(n26938), .B(n26939), .X(n26937) );
  nand_x4_sg U68838 ( .A(n26932), .B(n26933), .X(n26931) );
  nand_x4_sg U68839 ( .A(n26926), .B(n26927), .X(n26925) );
  nand_x4_sg U68840 ( .A(n27230), .B(n27231), .X(n27229) );
  nand_x4_sg U68841 ( .A(n27224), .B(n27225), .X(n27223) );
  nand_x4_sg U68842 ( .A(n27218), .B(n27219), .X(n27217) );
  nand_x4_sg U68843 ( .A(n27212), .B(n27213), .X(n27211) );
  nand_x4_sg U68844 ( .A(n27206), .B(n27207), .X(n27205) );
  nand_x4_sg U68845 ( .A(n27515), .B(n27516), .X(n27514) );
  nand_x4_sg U68846 ( .A(n27509), .B(n27510), .X(n27508) );
  nand_x4_sg U68847 ( .A(n27503), .B(n27504), .X(n27502) );
  nand_x4_sg U68848 ( .A(n27497), .B(n27498), .X(n27496) );
  nand_x4_sg U68849 ( .A(n27491), .B(n27492), .X(n27490) );
  nand_x4_sg U68850 ( .A(n27485), .B(n27486), .X(n27484) );
  nand_x4_sg U68851 ( .A(n27788), .B(n27789), .X(n27787) );
  nand_x4_sg U68852 ( .A(n27782), .B(n27783), .X(n27781) );
  nand_x4_sg U68853 ( .A(n27776), .B(n27777), .X(n27775) );
  nand_x4_sg U68854 ( .A(n27770), .B(n27771), .X(n27769) );
  nand_x4_sg U68855 ( .A(n27764), .B(n27765), .X(n27763) );
  nand_x4_sg U68856 ( .A(n28069), .B(n28070), .X(n28068) );
  nand_x4_sg U68857 ( .A(n28063), .B(n28064), .X(n28062) );
  nand_x4_sg U68858 ( .A(n28057), .B(n28058), .X(n28056) );
  nand_x4_sg U68859 ( .A(n28051), .B(n28052), .X(n28050) );
  nand_x4_sg U68860 ( .A(n28045), .B(n28046), .X(n28044) );
  nand_x4_sg U68861 ( .A(n28354), .B(n28355), .X(n28353) );
  nand_x4_sg U68862 ( .A(n28344), .B(n28345), .X(n28343) );
  nand_x4_sg U68863 ( .A(n28338), .B(n28339), .X(n28337) );
  nand_x4_sg U68864 ( .A(n28332), .B(n28333), .X(n28331) );
  nand_x4_sg U68865 ( .A(n28326), .B(n28327), .X(n28325) );
  nand_x4_sg U68866 ( .A(n28627), .B(n28628), .X(n28626) );
  nand_x4_sg U68867 ( .A(n28621), .B(n28622), .X(n28620) );
  nand_x4_sg U68868 ( .A(n28615), .B(n28616), .X(n28614) );
  nand_x4_sg U68869 ( .A(n28609), .B(n28610), .X(n28608) );
  nand_x4_sg U68870 ( .A(n28603), .B(n28604), .X(n28602) );
  nand_x4_sg U68871 ( .A(n28911), .B(n28912), .X(n28910) );
  nand_x4_sg U68872 ( .A(n28901), .B(n28902), .X(n28900) );
  nand_x4_sg U68873 ( .A(n28895), .B(n28896), .X(n28894) );
  nand_x4_sg U68874 ( .A(n28889), .B(n28890), .X(n28888) );
  nand_x4_sg U68875 ( .A(n28883), .B(n28884), .X(n28882) );
  nand_x4_sg U68876 ( .A(n29188), .B(n29189), .X(n29187) );
  nand_x4_sg U68877 ( .A(n29182), .B(n29183), .X(n29181) );
  nand_x4_sg U68878 ( .A(n29176), .B(n29177), .X(n29175) );
  nand_x4_sg U68879 ( .A(n29170), .B(n29171), .X(n29169) );
  nand_x4_sg U68880 ( .A(n29164), .B(n29165), .X(n29163) );
  nand_x4_sg U68881 ( .A(n29472), .B(n29473), .X(n29471) );
  nand_x4_sg U68882 ( .A(n29462), .B(n29463), .X(n29461) );
  nand_x4_sg U68883 ( .A(n29456), .B(n29457), .X(n29455) );
  nand_x4_sg U68884 ( .A(n29450), .B(n29451), .X(n29449) );
  nand_x4_sg U68885 ( .A(n29444), .B(n29445), .X(n29443) );
  nand_x4_sg U68886 ( .A(n29438), .B(n29439), .X(n29437) );
  nand_x4_sg U68887 ( .A(n25525), .B(n25526), .X(n25524) );
  nand_x4_sg U68888 ( .A(n25618), .B(n25619), .X(n25617) );
  nand_x4_sg U68889 ( .A(n25804), .B(n25805), .X(n25803) );
  nand_x4_sg U68890 ( .A(n25899), .B(n25900), .X(n25898) );
  nand_x4_sg U68891 ( .A(n26179), .B(n26180), .X(n26178) );
  nand_x4_sg U68892 ( .A(n26458), .B(n26459), .X(n26457) );
  nand_x4_sg U68893 ( .A(n26736), .B(n26737), .X(n26735) );
  nand_x4_sg U68894 ( .A(n26920), .B(n26921), .X(n26919) );
  nand_x4_sg U68895 ( .A(n27015), .B(n27016), .X(n27014) );
  nand_x4_sg U68896 ( .A(n27295), .B(n27296), .X(n27294) );
  nand_x4_sg U68897 ( .A(n27479), .B(n27480), .X(n27478) );
  nand_x4_sg U68898 ( .A(n27574), .B(n27575), .X(n27573) );
  nand_x4_sg U68899 ( .A(n27853), .B(n27854), .X(n27852) );
  nand_x4_sg U68900 ( .A(n28039), .B(n28040), .X(n28038) );
  nand_x4_sg U68901 ( .A(n28134), .B(n28135), .X(n28133) );
  nand_x4_sg U68902 ( .A(n28320), .B(n28321), .X(n28319) );
  nand_x4_sg U68903 ( .A(n28413), .B(n28414), .X(n28412) );
  nand_x4_sg U68904 ( .A(n28597), .B(n28598), .X(n28596) );
  nand_x4_sg U68905 ( .A(n28692), .B(n28693), .X(n28691) );
  nand_x4_sg U68906 ( .A(n28877), .B(n28878), .X(n28876) );
  nand_x4_sg U68907 ( .A(n28970), .B(n28971), .X(n28969) );
  nand_x4_sg U68908 ( .A(n29158), .B(n29159), .X(n29157) );
  nand_x4_sg U68909 ( .A(n29253), .B(n29254), .X(n29252) );
  nand_x4_sg U68910 ( .A(n29531), .B(n29532), .X(n29530) );
  nand_x4_sg U68911 ( .A(n49978), .B(n30936), .X(n24611) );
  nand_x1_sg U68912 ( .A(n24586), .B(n45331), .X(n30936) );
  nor_x1_sg U68913 ( .A(n45331), .B(n24586), .X(n30938) );
  nand_x4_sg U68914 ( .A(n49888), .B(n31331), .X(n24708) );
  nand_x1_sg U68915 ( .A(n24684), .B(n45329), .X(n31331) );
  nor_x1_sg U68916 ( .A(n45329), .B(n24684), .X(n31333) );
  nand_x4_sg U68917 ( .A(n50837), .B(n23270), .X(n9503) );
  nand_x1_sg U68918 ( .A(n9478), .B(n45335), .X(n23270) );
  nor_x1_sg U68919 ( .A(n45335), .B(n9478), .X(n23272) );
  nand_x4_sg U68920 ( .A(n50747), .B(n23665), .X(n9600) );
  nand_x1_sg U68921 ( .A(n9576), .B(n45333), .X(n23665) );
  nor_x1_sg U68922 ( .A(n45333), .B(n9576), .X(n23667) );
  nor_x1_sg U68923 ( .A(n28927), .B(n28928), .X(n28926) );
  nor_x1_sg U68924 ( .A(n29488), .B(n29489), .X(n29487) );
  nor_x1_sg U68925 ( .A(n26693), .B(n26694), .X(n26692) );
  nand_x4_sg U68926 ( .A(n24310), .B(n24311), .X(n24205) );
  nand_x1_sg U68927 ( .A(n24313), .B(n50141), .X(n24310) );
  nand_x4_sg U68928 ( .A(n31976), .B(n31977), .X(n31871) );
  nand_x1_sg U68929 ( .A(n31979), .B(n49282), .X(n31976) );
  nand_x4_sg U68930 ( .A(n24069), .B(n24070), .X(n23927) );
  nand_x1_sg U68931 ( .A(n24072), .B(n50143), .X(n24069) );
  nand_x4_sg U68932 ( .A(n31735), .B(n31736), .X(n31593) );
  nand_x1_sg U68933 ( .A(n31738), .B(n49284), .X(n31735) );
  nand_x4_sg U68934 ( .A(n22922), .B(n22923), .X(n22673) );
  nand_x1_sg U68935 ( .A(n22925), .B(n50149), .X(n22922) );
  nand_x4_sg U68936 ( .A(n30588), .B(n30589), .X(n30339) );
  nand_x1_sg U68937 ( .A(n30591), .B(n49290), .X(n30588) );
  nand_x4_sg U68938 ( .A(n22054), .B(n22055), .X(n10226) );
  nand_x1_sg U68939 ( .A(n22057), .B(n50153), .X(n22054) );
  nand_x4_sg U68940 ( .A(n29719), .B(n29720), .X(n25334) );
  nand_x1_sg U68941 ( .A(n29722), .B(n49294), .X(n29719) );
  nor_x1_sg U68942 ( .A(n22591), .B(n9364), .X(n22590) );
  nor_x1_sg U68943 ( .A(n23456), .B(n9668), .X(n23548) );
  nor_x1_sg U68944 ( .A(n30257), .B(n24488), .X(n30256) );
  nor_x1_sg U68945 ( .A(n31122), .B(n24781), .X(n31214) );
  nor_x1_sg U68946 ( .A(n26972), .B(n26973), .X(n26971) );
  nor_x1_sg U68947 ( .A(n23396), .B(n10150), .X(n23578) );
  nor_x1_sg U68948 ( .A(n31062), .B(n25263), .X(n31244) );
  nor_x1_sg U68949 ( .A(n25856), .B(n25857), .X(n25855) );
  nor_x1_sg U68950 ( .A(n26415), .B(n26416), .X(n26414) );
  nor_x1_sg U68951 ( .A(n27252), .B(n27253), .X(n27251) );
  nor_x1_sg U68952 ( .A(n27810), .B(n27811), .X(n27809) );
  nor_x1_sg U68953 ( .A(n23112), .B(n9474), .X(n23111) );
  nor_x1_sg U68954 ( .A(n23468), .B(n9572), .X(n23542) );
  nor_x1_sg U68955 ( .A(n30778), .B(n24587), .X(n30777) );
  nor_x1_sg U68956 ( .A(n31134), .B(n24685), .X(n31208) );
  nor_x1_sg U68957 ( .A(n21951), .B(n21974), .X(n21973) );
  nor_x1_sg U68958 ( .A(n29606), .B(n29639), .X(n29638) );
  nand_x4_sg U68959 ( .A(n22402), .B(n22403), .X(n22247) );
  nand_x4_sg U68960 ( .A(n30067), .B(n30068), .X(n29912) );
  nand_x4_sg U68961 ( .A(n23385), .B(n23386), .X(n23172) );
  nand_x4_sg U68962 ( .A(n31051), .B(n31052), .X(n30838) );
  nor_x1_sg U68963 ( .A(n23450), .B(n9715), .X(n23551) );
  nor_x1_sg U68964 ( .A(n23444), .B(n9763), .X(n23554) );
  nor_x1_sg U68965 ( .A(n23438), .B(n9811), .X(n23557) );
  nor_x1_sg U68966 ( .A(n23432), .B(n9859), .X(n23560) );
  nor_x1_sg U68967 ( .A(n23426), .B(n9907), .X(n23563) );
  nor_x1_sg U68968 ( .A(n23420), .B(n9955), .X(n23566) );
  nor_x1_sg U68969 ( .A(n31116), .B(n24828), .X(n31217) );
  nor_x1_sg U68970 ( .A(n31110), .B(n24876), .X(n31220) );
  nor_x1_sg U68971 ( .A(n31104), .B(n24924), .X(n31223) );
  nor_x1_sg U68972 ( .A(n31098), .B(n24972), .X(n31226) );
  nor_x1_sg U68973 ( .A(n31092), .B(n25020), .X(n31229) );
  nor_x1_sg U68974 ( .A(n31086), .B(n25068), .X(n31232) );
  nor_x1_sg U68975 ( .A(n23414), .B(n10004), .X(n23569) );
  nor_x1_sg U68976 ( .A(n31080), .B(n25117), .X(n31235) );
  nor_x1_sg U68977 ( .A(n22855), .B(n9425), .X(n22854) );
  nor_x1_sg U68978 ( .A(n23336), .B(n9523), .X(n23335) );
  nor_x1_sg U68979 ( .A(n23462), .B(n9620), .X(n23545) );
  nor_x1_sg U68980 ( .A(n23408), .B(n10052), .X(n23572) );
  nor_x1_sg U68981 ( .A(n23402), .B(n10101), .X(n23575) );
  nor_x1_sg U68982 ( .A(n30521), .B(n24538), .X(n30520) );
  nor_x1_sg U68983 ( .A(n31002), .B(n24636), .X(n31001) );
  nor_x1_sg U68984 ( .A(n31128), .B(n24733), .X(n31211) );
  nor_x1_sg U68985 ( .A(n31074), .B(n25165), .X(n31238) );
  nor_x1_sg U68986 ( .A(n31068), .B(n25214), .X(n31241) );
  nor_x1_sg U68987 ( .A(n22561), .B(n22562), .X(n22560) );
  nor_x1_sg U68988 ( .A(n30227), .B(n30228), .X(n30226) );
  nor_x1_sg U68989 ( .A(n23312), .B(n23313), .X(n23311) );
  nor_x1_sg U68990 ( .A(n23707), .B(n23708), .X(n23706) );
  nor_x1_sg U68991 ( .A(n24031), .B(n24032), .X(n24030) );
  nor_x1_sg U68992 ( .A(n23086), .B(n23087), .X(n23085) );
  nor_x1_sg U68993 ( .A(n23517), .B(n23518), .X(n23516) );
  nor_x1_sg U68994 ( .A(n23878), .B(n23879), .X(n23877) );
  nor_x1_sg U68995 ( .A(n24138), .B(n24135), .X(n24174) );
  nor_x1_sg U68996 ( .A(n22831), .B(n22832), .X(n22830) );
  nor_x1_sg U68997 ( .A(n22172), .B(n22169), .X(n22195) );
  nor_x1_sg U68998 ( .A(n29837), .B(n29834), .X(n29860) );
  nor_x1_sg U68999 ( .A(n30497), .B(n30498), .X(n30496) );
  nor_x1_sg U69000 ( .A(n30752), .B(n30753), .X(n30751) );
  nor_x1_sg U69001 ( .A(n30978), .B(n30979), .X(n30977) );
  nor_x1_sg U69002 ( .A(n31183), .B(n31184), .X(n31182) );
  nor_x1_sg U69003 ( .A(n31373), .B(n31374), .X(n31372) );
  nor_x1_sg U69004 ( .A(n31544), .B(n31545), .X(n31543) );
  nor_x1_sg U69005 ( .A(n31697), .B(n31698), .X(n31696) );
  nor_x1_sg U69006 ( .A(n31804), .B(n31801), .X(n31840) );
  nand_x2_sg U69007 ( .A(n9408), .B(n50946), .X(n9407) );
  nand_x1_sg U69008 ( .A(n9410), .B(n9383), .X(n9408) );
  nor_x1_sg U69009 ( .A(n9383), .B(n9410), .X(n9409) );
  nand_x2_sg U69010 ( .A(n24517), .B(n50087), .X(n24516) );
  nand_x1_sg U69011 ( .A(n24519), .B(n24498), .X(n24517) );
  nor_x1_sg U69012 ( .A(n24498), .B(n24519), .X(n24518) );
  nand_x2_sg U69013 ( .A(n9507), .B(n50850), .X(n9506) );
  nand_x1_sg U69014 ( .A(n9509), .B(n9488), .X(n9507) );
  nor_x1_sg U69015 ( .A(n9488), .B(n9509), .X(n9508) );
  nand_x2_sg U69016 ( .A(n9556), .B(n50805), .X(n9555) );
  nand_x1_sg U69017 ( .A(n9558), .B(n9537), .X(n9556) );
  nor_x1_sg U69018 ( .A(n9537), .B(n9558), .X(n9557) );
  nand_x2_sg U69019 ( .A(n9604), .B(n50757), .X(n9603) );
  nand_x1_sg U69020 ( .A(n9606), .B(n9586), .X(n9604) );
  nor_x1_sg U69021 ( .A(n9586), .B(n9606), .X(n9605) );
  nand_x2_sg U69022 ( .A(n9652), .B(n50710), .X(n9651) );
  nand_x1_sg U69023 ( .A(n9654), .B(n9634), .X(n9652) );
  nor_x1_sg U69024 ( .A(n9634), .B(n9654), .X(n9653) );
  nand_x2_sg U69025 ( .A(n9699), .B(n50662), .X(n9698) );
  nand_x1_sg U69026 ( .A(n9701), .B(n9682), .X(n9699) );
  nor_x1_sg U69027 ( .A(n9682), .B(n9701), .X(n9700) );
  nand_x2_sg U69028 ( .A(n9747), .B(n50615), .X(n9746) );
  nand_x1_sg U69029 ( .A(n9749), .B(n9729), .X(n9747) );
  nor_x1_sg U69030 ( .A(n9729), .B(n9749), .X(n9748) );
  nand_x2_sg U69031 ( .A(n9795), .B(n50566), .X(n9794) );
  nand_x1_sg U69032 ( .A(n9797), .B(n9777), .X(n9795) );
  nor_x1_sg U69033 ( .A(n9777), .B(n9797), .X(n9796) );
  nand_x2_sg U69034 ( .A(n9843), .B(n50519), .X(n9842) );
  nand_x1_sg U69035 ( .A(n9845), .B(n9825), .X(n9843) );
  nor_x1_sg U69036 ( .A(n9825), .B(n9845), .X(n9844) );
  nand_x2_sg U69037 ( .A(n9891), .B(n50472), .X(n9890) );
  nand_x1_sg U69038 ( .A(n9893), .B(n9873), .X(n9891) );
  nor_x1_sg U69039 ( .A(n9873), .B(n9893), .X(n9892) );
  nand_x2_sg U69040 ( .A(n9939), .B(n50426), .X(n9938) );
  nand_x1_sg U69041 ( .A(n9941), .B(n9921), .X(n9939) );
  nor_x1_sg U69042 ( .A(n9921), .B(n9941), .X(n9940) );
  nand_x2_sg U69043 ( .A(n9988), .B(n50379), .X(n9987) );
  nand_x1_sg U69044 ( .A(n9990), .B(n9969), .X(n9988) );
  nor_x1_sg U69045 ( .A(n9969), .B(n9990), .X(n9989) );
  nand_x2_sg U69046 ( .A(n10036), .B(n50332), .X(n10035) );
  nand_x1_sg U69047 ( .A(n10038), .B(n10018), .X(n10036) );
  nor_x1_sg U69048 ( .A(n10018), .B(n10038), .X(n10037) );
  nand_x2_sg U69049 ( .A(n10085), .B(n50286), .X(n10084) );
  nand_x1_sg U69050 ( .A(n10087), .B(n10066), .X(n10085) );
  nor_x1_sg U69051 ( .A(n10066), .B(n10087), .X(n10086) );
  nand_x2_sg U69052 ( .A(n10134), .B(n50240), .X(n10133) );
  nand_x1_sg U69053 ( .A(n10136), .B(n10115), .X(n10134) );
  nor_x1_sg U69054 ( .A(n10115), .B(n10136), .X(n10135) );
  nand_x2_sg U69055 ( .A(n10181), .B(n50196), .X(n10180) );
  nand_x1_sg U69056 ( .A(n10183), .B(n10164), .X(n10181) );
  nor_x1_sg U69057 ( .A(n10164), .B(n10183), .X(n10182) );
  nand_x2_sg U69058 ( .A(n24615), .B(n49991), .X(n24614) );
  nand_x1_sg U69059 ( .A(n24617), .B(n24596), .X(n24615) );
  nor_x1_sg U69060 ( .A(n24596), .B(n24617), .X(n24616) );
  nand_x2_sg U69061 ( .A(n24664), .B(n49946), .X(n24663) );
  nand_x1_sg U69062 ( .A(n24666), .B(n24645), .X(n24664) );
  nor_x1_sg U69063 ( .A(n24645), .B(n24666), .X(n24665) );
  nand_x2_sg U69064 ( .A(n24712), .B(n49898), .X(n24711) );
  nand_x1_sg U69065 ( .A(n24714), .B(n24694), .X(n24712) );
  nor_x1_sg U69066 ( .A(n24694), .B(n24714), .X(n24713) );
  nand_x2_sg U69067 ( .A(n24760), .B(n49851), .X(n24759) );
  nand_x1_sg U69068 ( .A(n24762), .B(n24742), .X(n24760) );
  nor_x1_sg U69069 ( .A(n24742), .B(n24762), .X(n24761) );
  nand_x2_sg U69070 ( .A(n24807), .B(n49803), .X(n24806) );
  nand_x1_sg U69071 ( .A(n24809), .B(n24790), .X(n24807) );
  nor_x1_sg U69072 ( .A(n24790), .B(n24809), .X(n24808) );
  nand_x2_sg U69073 ( .A(n24855), .B(n49756), .X(n24854) );
  nand_x1_sg U69074 ( .A(n24857), .B(n24837), .X(n24855) );
  nor_x1_sg U69075 ( .A(n24837), .B(n24857), .X(n24856) );
  nand_x2_sg U69076 ( .A(n24903), .B(n49707), .X(n24902) );
  nand_x1_sg U69077 ( .A(n24905), .B(n24885), .X(n24903) );
  nor_x1_sg U69078 ( .A(n24885), .B(n24905), .X(n24904) );
  nand_x2_sg U69079 ( .A(n24951), .B(n49660), .X(n24950) );
  nand_x1_sg U69080 ( .A(n24953), .B(n24933), .X(n24951) );
  nor_x1_sg U69081 ( .A(n24933), .B(n24953), .X(n24952) );
  nand_x2_sg U69082 ( .A(n24999), .B(n49613), .X(n24998) );
  nand_x1_sg U69083 ( .A(n25001), .B(n24981), .X(n24999) );
  nor_x1_sg U69084 ( .A(n24981), .B(n25001), .X(n25000) );
  nand_x2_sg U69085 ( .A(n25047), .B(n49567), .X(n25046) );
  nand_x1_sg U69086 ( .A(n25049), .B(n25029), .X(n25047) );
  nor_x1_sg U69087 ( .A(n25029), .B(n25049), .X(n25048) );
  nand_x2_sg U69088 ( .A(n25096), .B(n49520), .X(n25095) );
  nand_x1_sg U69089 ( .A(n25098), .B(n25077), .X(n25096) );
  nor_x1_sg U69090 ( .A(n25077), .B(n25098), .X(n25097) );
  nand_x2_sg U69091 ( .A(n25144), .B(n49473), .X(n25143) );
  nand_x1_sg U69092 ( .A(n25146), .B(n25126), .X(n25144) );
  nor_x1_sg U69093 ( .A(n25126), .B(n25146), .X(n25145) );
  nand_x2_sg U69094 ( .A(n25193), .B(n49427), .X(n25192) );
  nand_x1_sg U69095 ( .A(n25195), .B(n25174), .X(n25193) );
  nor_x1_sg U69096 ( .A(n25174), .B(n25195), .X(n25194) );
  nand_x2_sg U69097 ( .A(n25242), .B(n49381), .X(n25241) );
  nand_x1_sg U69098 ( .A(n25244), .B(n25223), .X(n25242) );
  nor_x1_sg U69099 ( .A(n25223), .B(n25244), .X(n25243) );
  nand_x2_sg U69100 ( .A(n25289), .B(n49337), .X(n25288) );
  nand_x1_sg U69101 ( .A(n25291), .B(n25272), .X(n25289) );
  nor_x1_sg U69102 ( .A(n25272), .B(n25291), .X(n25290) );
  nand_x2_sg U69103 ( .A(n9458), .B(n50899), .X(n9457) );
  nand_x1_sg U69104 ( .A(n9460), .B(n9439), .X(n9458) );
  nor_x1_sg U69105 ( .A(n9439), .B(n9460), .X(n9459) );
  nand_x2_sg U69106 ( .A(n24566), .B(n50040), .X(n24565) );
  nand_x1_sg U69107 ( .A(n24568), .B(n24547), .X(n24566) );
  nor_x1_sg U69108 ( .A(n24547), .B(n24568), .X(n24567) );
  nand_x4_sg U69109 ( .A(n10236), .B(n10237), .X(n10233) );
  nor_x1_sg U69110 ( .A(n10238), .B(n10239), .X(n10237) );
  nor_x1_sg U69111 ( .A(n10242), .B(n10243), .X(n10236) );
  nand_x4_sg U69112 ( .A(n25344), .B(n25345), .X(n25341) );
  nor_x1_sg U69113 ( .A(n25346), .B(n25347), .X(n25345) );
  nor_x1_sg U69114 ( .A(n25350), .B(n25351), .X(n25344) );
  nand_x2_sg U69115 ( .A(n10258), .B(n55463), .X(n10248) );
  nor_x1_sg U69116 ( .A(n10261), .B(n10262), .X(n10258) );
  nor_x1_sg U69117 ( .A(n10260), .B(n9394), .X(n10259) );
  nand_x2_sg U69118 ( .A(n10274), .B(n10275), .X(n10268) );
  nor_x1_sg U69119 ( .A(n10277), .B(n10278), .X(n10274) );
  nand_x2_sg U69120 ( .A(n10250), .B(n55466), .X(n10249) );
  nor_x1_sg U69121 ( .A(n10253), .B(n10254), .X(n10250) );
  nor_x1_sg U69122 ( .A(n9385), .B(n10252), .X(n10251) );
  nand_x2_sg U69123 ( .A(n25365), .B(n55464), .X(n25356) );
  nor_x1_sg U69124 ( .A(n25368), .B(n25369), .X(n25365) );
  nor_x1_sg U69125 ( .A(n25367), .B(n9394), .X(n25366) );
  nand_x2_sg U69126 ( .A(n25380), .B(n25381), .X(n25374) );
  nor_x1_sg U69127 ( .A(n25383), .B(n25384), .X(n25380) );
  nand_x2_sg U69128 ( .A(n25358), .B(n55467), .X(n25357) );
  nor_x1_sg U69129 ( .A(n25361), .B(n25362), .X(n25358) );
  nor_x1_sg U69130 ( .A(n25360), .B(n9385), .X(n25359) );
  nand_x2_sg U69131 ( .A(n10224), .B(n10225), .X(n10223) );
  nand_x1_sg U69132 ( .A(n10227), .B(n50154), .X(n10224) );
  nand_x2_sg U69133 ( .A(n25332), .B(n25333), .X(n25331) );
  nand_x1_sg U69134 ( .A(n25335), .B(n49295), .X(n25332) );
  nand_x2_sg U69135 ( .A(n32139), .B(output_taken), .X(n32138) );
  nor_x1_sg U69136 ( .A(state[0]), .B(n55796), .X(n32139) );
  nand_x1_sg U69137 ( .A(n46657), .B(n46085), .X(n39915) );
  nand_x1_sg U69138 ( .A(n46643), .B(n45237), .X(n39923) );
  nand_x1_sg U69139 ( .A(n46654), .B(n46063), .X(n39955) );
  nand_x1_sg U69140 ( .A(n46654), .B(n46077), .X(n39957) );
  nand_x1_sg U69141 ( .A(n46655), .B(n46035), .X(n39961) );
  nand_x1_sg U69142 ( .A(n46652), .B(n46073), .X(n39995) );
  nand_x1_sg U69143 ( .A(n46655), .B(n45235), .X(n40003) );
  nand_x1_sg U69144 ( .A(n46653), .B(n46055), .X(n40035) );
  nand_x1_sg U69145 ( .A(n46651), .B(n46049), .X(n40037) );
  nand_x1_sg U69146 ( .A(n46652), .B(n45225), .X(n40041) );
  nand_x1_sg U69147 ( .A(n46652), .B(n46071), .X(n40075) );
  nand_x1_sg U69148 ( .A(n46657), .B(n45227), .X(n40083) );
  nand_x1_sg U69149 ( .A(n46646), .B(n46083), .X(n40115) );
  nand_x1_sg U69150 ( .A(n46642), .B(n46033), .X(n40123) );
  nand_x1_sg U69151 ( .A(n46650), .B(n46053), .X(n40155) );
  nand_x1_sg U69152 ( .A(n46650), .B(n46047), .X(n40157) );
  nand_x1_sg U69153 ( .A(n46655), .B(n45223), .X(n40161) );
  nand_x1_sg U69154 ( .A(n46642), .B(n46075), .X(n40195) );
  nand_x1_sg U69155 ( .A(n46648), .B(n45233), .X(n40203) );
  nand_x1_sg U69156 ( .A(n46648), .B(n46051), .X(n40235) );
  nand_x1_sg U69157 ( .A(n46651), .B(n46045), .X(n40237) );
  nand_x1_sg U69158 ( .A(n46643), .B(n45221), .X(n40241) );
  nand_x1_sg U69159 ( .A(n46655), .B(n46067), .X(n40275) );
  nand_x1_sg U69160 ( .A(n46647), .B(n46059), .X(n40277) );
  nand_x1_sg U69161 ( .A(n46651), .B(n46041), .X(n40281) );
  nand_x1_sg U69162 ( .A(n46646), .B(n46043), .X(n40321) );
  nand_x1_sg U69163 ( .A(n46653), .B(n46091), .X(n39825) );
  nand_x1_sg U69164 ( .A(n46650), .B(n46155), .X(n39833) );
  nand_x1_sg U69165 ( .A(n46646), .B(n46097), .X(n39865) );
  nand_x1_sg U69166 ( .A(n46650), .B(n46175), .X(n39873) );
  nand_x1_sg U69167 ( .A(n46657), .B(n46145), .X(n39877) );
  nand_x1_sg U69168 ( .A(n46651), .B(n46135), .X(n39879) );
  nand_x1_sg U69169 ( .A(n46647), .B(n46121), .X(n39883) );
  nand_x1_sg U69170 ( .A(n46655), .B(n46089), .X(n39905) );
  nand_x1_sg U69171 ( .A(n46653), .B(n45303), .X(n39913) );
  nand_x1_sg U69172 ( .A(n46657), .B(n45275), .X(n39917) );
  nand_x1_sg U69173 ( .A(n46654), .B(n45327), .X(n39919) );
  nand_x1_sg U69174 ( .A(n46655), .B(n45241), .X(n39945) );
  nand_x1_sg U69175 ( .A(n46647), .B(n45305), .X(n39953) );
  nand_x1_sg U69176 ( .A(n46646), .B(n45259), .X(n39985) );
  nand_x1_sg U69177 ( .A(n46653), .B(n45325), .X(n39993) );
  nand_x1_sg U69178 ( .A(n46647), .B(n45281), .X(n39997) );
  nand_x1_sg U69179 ( .A(n46645), .B(n45293), .X(n39999) );
  nand_x1_sg U69180 ( .A(n46642), .B(n45263), .X(n40025) );
  nand_x1_sg U69181 ( .A(n46643), .B(n45323), .X(n40033) );
  nand_x1_sg U69182 ( .A(n46646), .B(n45269), .X(n40065) );
  nand_x1_sg U69183 ( .A(n46654), .B(n45317), .X(n40073) );
  nand_x1_sg U69184 ( .A(n46643), .B(n45291), .X(n40077) );
  nand_x1_sg U69185 ( .A(n46652), .B(n45273), .X(n40079) );
  nand_x1_sg U69186 ( .A(n46650), .B(n45261), .X(n40105) );
  nand_x1_sg U69187 ( .A(n46652), .B(n45313), .X(n40113) );
  nand_x1_sg U69188 ( .A(n46653), .B(n45309), .X(n40117) );
  nand_x1_sg U69189 ( .A(n46654), .B(n45283), .X(n40119) );
  nand_x1_sg U69190 ( .A(n46654), .B(n45249), .X(n40145) );
  nand_x1_sg U69191 ( .A(n46653), .B(n45321), .X(n40153) );
  nand_x1_sg U69192 ( .A(n46651), .B(n45267), .X(n40185) );
  nand_x1_sg U69193 ( .A(n46652), .B(n45307), .X(n40193) );
  nand_x1_sg U69194 ( .A(n46652), .B(n45285), .X(n40197) );
  nand_x1_sg U69195 ( .A(n46657), .B(n45301), .X(n40199) );
  nand_x1_sg U69196 ( .A(n46655), .B(n45257), .X(n40225) );
  nand_x1_sg U69197 ( .A(n46652), .B(n45319), .X(n40233) );
  nand_x1_sg U69198 ( .A(n46646), .B(n45265), .X(n40265) );
  nand_x1_sg U69199 ( .A(n46643), .B(n45299), .X(n40273) );
  nand_x1_sg U69200 ( .A(n46652), .B(n45255), .X(n40305) );
  nand_x1_sg U69201 ( .A(n46642), .B(n45271), .X(n40317) );
  nand_x1_sg U69202 ( .A(n46653), .B(n46001), .X(n39831) );
  nand_x1_sg U69203 ( .A(n46645), .B(n46025), .X(n39871) );
  nand_x1_sg U69204 ( .A(n46647), .B(n46031), .X(n39959) );
  nand_x1_sg U69205 ( .A(n46648), .B(n46029), .X(n39963) );
  nand_x1_sg U69206 ( .A(n46643), .B(n45999), .X(n40039) );
  nand_x1_sg U69207 ( .A(n46650), .B(n45217), .X(n40043) );
  nand_x1_sg U69208 ( .A(n46645), .B(n45997), .X(n40159) );
  nand_x1_sg U69209 ( .A(n46652), .B(n45215), .X(n40163) );
  nand_x1_sg U69210 ( .A(n46655), .B(n45995), .X(n40239) );
  nand_x1_sg U69211 ( .A(n46652), .B(n45213), .X(n40243) );
  nand_x1_sg U69212 ( .A(n46657), .B(n45993), .X(n40279) );
  nand_x1_sg U69213 ( .A(n46652), .B(n45981), .X(n40283) );
  nand_x1_sg U69214 ( .A(n46650), .B(n45219), .X(n40319) );
  nand_x1_sg U69215 ( .A(n46650), .B(n45211), .X(n40323) );
  nand_x1_sg U69216 ( .A(n46642), .B(n45953), .X(n39829) );
  nand_x1_sg U69217 ( .A(n46654), .B(n45973), .X(n39869) );
  nand_x1_sg U69218 ( .A(n46654), .B(n45947), .X(n40069) );
  nand_x1_sg U69219 ( .A(n46646), .B(n45209), .X(n40315) );
  nand_x1_sg U69220 ( .A(n46655), .B(n44943), .X(n39813) );
  nand_x1_sg U69221 ( .A(n46657), .B(n45151), .X(n39815) );
  nand_x1_sg U69222 ( .A(n46648), .B(n45157), .X(n39817) );
  nand_x1_sg U69223 ( .A(n46641), .B(n44941), .X(n39819) );
  nand_x1_sg U69224 ( .A(n46657), .B(n44939), .X(n39821) );
  nand_x1_sg U69225 ( .A(n46647), .B(n44937), .X(n39823) );
  nand_x1_sg U69226 ( .A(n44763), .B(n46652), .X(n39827) );
  nand_x1_sg U69227 ( .A(n46648), .B(n44893), .X(n39835) );
  nand_x1_sg U69228 ( .A(n46647), .B(n44883), .X(n39837) );
  nand_x1_sg U69229 ( .A(n46655), .B(n44803), .X(n39839) );
  nand_x1_sg U69230 ( .A(n46646), .B(n44809), .X(n39841) );
  nand_x1_sg U69231 ( .A(n46644), .B(n44797), .X(n39843) );
  nand_x1_sg U69232 ( .A(n46653), .B(n44935), .X(n39845) );
  nand_x1_sg U69233 ( .A(n46647), .B(n45193), .X(n39847) );
  nand_x1_sg U69234 ( .A(n46654), .B(n44933), .X(n39849) );
  nand_x1_sg U69235 ( .A(n46648), .B(n44931), .X(n39851) );
  nand_x1_sg U69236 ( .A(n46651), .B(n45187), .X(n39853) );
  nand_x1_sg U69237 ( .A(n46646), .B(n44929), .X(n39855) );
  nand_x1_sg U69238 ( .A(n46652), .B(n45131), .X(n39857) );
  nand_x1_sg U69239 ( .A(n46642), .B(n44927), .X(n39859) );
  nand_x1_sg U69240 ( .A(n46647), .B(n44925), .X(n39861) );
  nand_x1_sg U69241 ( .A(n46648), .B(n44923), .X(n39863) );
  nand_x1_sg U69242 ( .A(n44761), .B(n46646), .X(n39867) );
  nand_x1_sg U69243 ( .A(n46643), .B(n44899), .X(n39875) );
  nand_x1_sg U69244 ( .A(n46651), .B(n45643), .X(n39881) );
  nand_x1_sg U69245 ( .A(n46652), .B(n44921), .X(n39885) );
  nand_x1_sg U69246 ( .A(n46657), .B(n45203), .X(n39887) );
  nand_x1_sg U69247 ( .A(n46643), .B(n44919), .X(n39889) );
  nand_x1_sg U69248 ( .A(n46650), .B(n44917), .X(n39891) );
  nand_x1_sg U69249 ( .A(n46655), .B(n44915), .X(n39893) );
  nand_x1_sg U69250 ( .A(n46652), .B(n45149), .X(n39895) );
  nand_x1_sg U69251 ( .A(n46643), .B(n45155), .X(n39897) );
  nand_x1_sg U69252 ( .A(n46651), .B(n44913), .X(n39899) );
  nand_x1_sg U69253 ( .A(n46655), .B(n44911), .X(n39901) );
  nand_x1_sg U69254 ( .A(n46657), .B(n44909), .X(n39903) );
  nand_x1_sg U69255 ( .A(n44759), .B(n46654), .X(n39907) );
  nand_x1_sg U69256 ( .A(n46648), .B(n44865), .X(n39911) );
  nand_x1_sg U69257 ( .A(n46650), .B(n44789), .X(n39921) );
  nand_x1_sg U69258 ( .A(n46641), .B(n45863), .X(n39925) );
  nand_x1_sg U69259 ( .A(n46650), .B(n45945), .X(n39927) );
  nand_x1_sg U69260 ( .A(n46653), .B(n45861), .X(n39929) );
  nand_x1_sg U69261 ( .A(n46654), .B(n45859), .X(n39931) );
  nand_x1_sg U69262 ( .A(n46651), .B(n45857), .X(n39933) );
  nand_x1_sg U69263 ( .A(n46652), .B(n45921), .X(n39935) );
  nand_x1_sg U69264 ( .A(n46655), .B(n45855), .X(n39937) );
  nand_x1_sg U69265 ( .A(n46657), .B(n45853), .X(n39939) );
  nand_x1_sg U69266 ( .A(n46648), .B(n45883), .X(n39941) );
  nand_x1_sg U69267 ( .A(n46654), .B(n45865), .X(n39943) );
  nand_x1_sg U69268 ( .A(n45631), .B(n46646), .X(n39947) );
  nand_x1_sg U69269 ( .A(n46644), .B(n44835), .X(n39951) );
  nand_x1_sg U69270 ( .A(n46650), .B(n45851), .X(n39965) );
  nand_x1_sg U69271 ( .A(n46646), .B(n45897), .X(n39967) );
  nand_x1_sg U69272 ( .A(n46654), .B(n45849), .X(n39969) );
  nand_x1_sg U69273 ( .A(n46644), .B(n45847), .X(n39971) );
  nand_x1_sg U69274 ( .A(n46655), .B(n45845), .X(n39973) );
  nand_x1_sg U69275 ( .A(n46653), .B(n45885), .X(n39975) );
  nand_x1_sg U69276 ( .A(n46654), .B(n45843), .X(n39977) );
  nand_x1_sg U69277 ( .A(n46645), .B(n45841), .X(n39979) );
  nand_x1_sg U69278 ( .A(n46657), .B(n45839), .X(n39981) );
  nand_x1_sg U69279 ( .A(n46641), .B(n45837), .X(n39983) );
  nand_x1_sg U69280 ( .A(n45629), .B(n46654), .X(n39987) );
  nand_x1_sg U69281 ( .A(n46648), .B(n44857), .X(n39991) );
  nand_x1_sg U69282 ( .A(n46647), .B(n44795), .X(n40001) );
  nand_x1_sg U69283 ( .A(n46651), .B(n45835), .X(n40005) );
  nand_x1_sg U69284 ( .A(n46654), .B(n45911), .X(n40007) );
  nand_x1_sg U69285 ( .A(n46657), .B(n45833), .X(n40009) );
  nand_x1_sg U69286 ( .A(n46646), .B(n45831), .X(n40011) );
  nand_x1_sg U69287 ( .A(n46644), .B(n45829), .X(n40013) );
  nand_x1_sg U69288 ( .A(n46643), .B(n45891), .X(n40015) );
  nand_x1_sg U69289 ( .A(n46651), .B(n45827), .X(n40017) );
  nand_x1_sg U69290 ( .A(n46647), .B(n45825), .X(n40019) );
  nand_x1_sg U69291 ( .A(n46650), .B(n45823), .X(n40021) );
  nand_x1_sg U69292 ( .A(n46653), .B(n45821), .X(n40023) );
  nand_x1_sg U69293 ( .A(n45627), .B(n46642), .X(n40027) );
  nand_x1_sg U69294 ( .A(n46641), .B(n44845), .X(n40031) );
  nand_x1_sg U69295 ( .A(n46653), .B(n45819), .X(n40045) );
  nand_x1_sg U69296 ( .A(n46655), .B(n45907), .X(n40047) );
  nand_x1_sg U69297 ( .A(n46650), .B(n45817), .X(n40049) );
  nand_x1_sg U69298 ( .A(n46657), .B(n45881), .X(n40051) );
  nand_x1_sg U69299 ( .A(n46657), .B(n45815), .X(n40053) );
  nand_x1_sg U69300 ( .A(n46648), .B(n45917), .X(n40055) );
  nand_x1_sg U69301 ( .A(n46657), .B(n45813), .X(n40057) );
  nand_x1_sg U69302 ( .A(n46647), .B(n45811), .X(n40059) );
  nand_x1_sg U69303 ( .A(n46646), .B(n45809), .X(n40061) );
  nand_x1_sg U69304 ( .A(n46657), .B(n45807), .X(n40063) );
  nand_x1_sg U69305 ( .A(n45625), .B(n46641), .X(n40067) );
  nand_x1_sg U69306 ( .A(n46648), .B(n44855), .X(n40071) );
  nand_x1_sg U69307 ( .A(n46654), .B(n44839), .X(n40081) );
  nand_x1_sg U69308 ( .A(n46657), .B(n45805), .X(n40085) );
  nand_x1_sg U69309 ( .A(n46657), .B(n45909), .X(n40087) );
  nand_x1_sg U69310 ( .A(n46648), .B(n45803), .X(n40089) );
  nand_x1_sg U69311 ( .A(n46655), .B(n45875), .X(n40091) );
  nand_x1_sg U69312 ( .A(n46650), .B(n45801), .X(n40093) );
  nand_x1_sg U69313 ( .A(n46657), .B(n45901), .X(n40095) );
  nand_x1_sg U69314 ( .A(n46647), .B(n45799), .X(n40097) );
  nand_x1_sg U69315 ( .A(n46657), .B(n45797), .X(n40099) );
  nand_x1_sg U69316 ( .A(n46651), .B(n45795), .X(n40101) );
  nand_x1_sg U69317 ( .A(n46659), .B(n45793), .X(n40103) );
  nand_x1_sg U69318 ( .A(n45623), .B(n46648), .X(n40107) );
  nand_x1_sg U69319 ( .A(n46655), .B(n44867), .X(n40111) );
  nand_x1_sg U69320 ( .A(n46648), .B(n44817), .X(n40121) );
  nand_x1_sg U69321 ( .A(n46645), .B(n45791), .X(n40125) );
  nand_x1_sg U69322 ( .A(n46643), .B(n45937), .X(n40127) );
  nand_x1_sg U69323 ( .A(n46648), .B(n45789), .X(n40129) );
  nand_x1_sg U69324 ( .A(n46646), .B(n45787), .X(n40131) );
  nand_x1_sg U69325 ( .A(n46655), .B(n45923), .X(n40133) );
  nand_x1_sg U69326 ( .A(n46644), .B(n45785), .X(n40135) );
  nand_x1_sg U69327 ( .A(n46643), .B(n45867), .X(n40137) );
  nand_x1_sg U69328 ( .A(n46644), .B(n45783), .X(n40139) );
  nand_x1_sg U69329 ( .A(n46655), .B(n45781), .X(n40141) );
  nand_x1_sg U69330 ( .A(n46643), .B(n45779), .X(n40143) );
  nand_x1_sg U69331 ( .A(n45621), .B(n46651), .X(n40147) );
  nand_x1_sg U69332 ( .A(n46655), .B(n44843), .X(n40151) );
  nand_x1_sg U69333 ( .A(n46652), .B(n45777), .X(n40165) );
  nand_x1_sg U69334 ( .A(n46650), .B(n45905), .X(n40167) );
  nand_x1_sg U69335 ( .A(n46653), .B(n45775), .X(n40169) );
  nand_x1_sg U69336 ( .A(n46657), .B(n45879), .X(n40171) );
  nand_x1_sg U69337 ( .A(n46650), .B(n45773), .X(n40173) );
  nand_x1_sg U69338 ( .A(n46642), .B(n45915), .X(n40175) );
  nand_x1_sg U69339 ( .A(n46657), .B(n45771), .X(n40177) );
  nand_x1_sg U69340 ( .A(n46642), .B(n45769), .X(n40179) );
  nand_x1_sg U69341 ( .A(n46655), .B(n45767), .X(n40181) );
  nand_x1_sg U69342 ( .A(n46653), .B(n45765), .X(n40183) );
  nand_x1_sg U69343 ( .A(n45619), .B(n46657), .X(n40187) );
  nand_x1_sg U69344 ( .A(n46653), .B(n44847), .X(n40191) );
  nand_x1_sg U69345 ( .A(n46653), .B(n44791), .X(n40201) );
  nand_x1_sg U69346 ( .A(n46657), .B(n45763), .X(n40205) );
  nand_x1_sg U69347 ( .A(n46659), .B(n45919), .X(n40207) );
  nand_x1_sg U69348 ( .A(n46652), .B(n45761), .X(n40209) );
  nand_x1_sg U69349 ( .A(n46654), .B(n45759), .X(n40211) );
  nand_x1_sg U69350 ( .A(n46650), .B(n45757), .X(n40213) );
  nand_x1_sg U69351 ( .A(n46655), .B(n45899), .X(n40215) );
  nand_x1_sg U69352 ( .A(n46647), .B(n45755), .X(n40217) );
  nand_x1_sg U69353 ( .A(n46650), .B(n45753), .X(n40219) );
  nand_x1_sg U69354 ( .A(n46653), .B(n45751), .X(n40221) );
  nand_x1_sg U69355 ( .A(n46653), .B(n45749), .X(n40223) );
  nand_x1_sg U69356 ( .A(n45617), .B(n46647), .X(n40227) );
  nand_x1_sg U69357 ( .A(n46654), .B(n44841), .X(n40231) );
  nand_x1_sg U69358 ( .A(n46653), .B(n45747), .X(n40245) );
  nand_x1_sg U69359 ( .A(n46648), .B(n45903), .X(n40247) );
  nand_x1_sg U69360 ( .A(n46648), .B(n45745), .X(n40249) );
  nand_x1_sg U69361 ( .A(n46646), .B(n45877), .X(n40251) );
  nand_x1_sg U69362 ( .A(n46654), .B(n45743), .X(n40253) );
  nand_x1_sg U69363 ( .A(n46651), .B(n45913), .X(n40255) );
  nand_x1_sg U69364 ( .A(n46650), .B(n45741), .X(n40257) );
  nand_x1_sg U69365 ( .A(n46653), .B(n45739), .X(n40259) );
  nand_x1_sg U69366 ( .A(n46645), .B(n45737), .X(n40261) );
  nand_x1_sg U69367 ( .A(n46648), .B(n45735), .X(n40263) );
  nand_x1_sg U69368 ( .A(n45615), .B(n46655), .X(n40267) );
  nand_x1_sg U69369 ( .A(n46642), .B(n44831), .X(n40271) );
  nand_x1_sg U69370 ( .A(n46643), .B(n45733), .X(n40285) );
  nand_x1_sg U69371 ( .A(n46657), .B(n45935), .X(n40287) );
  nand_x1_sg U69372 ( .A(n46641), .B(n45731), .X(n40289) );
  nand_x1_sg U69373 ( .A(n46657), .B(n45729), .X(n40291) );
  nand_x1_sg U69374 ( .A(n46651), .B(n45929), .X(n40293) );
  nand_x1_sg U69375 ( .A(n46652), .B(n45727), .X(n40295) );
  nand_x1_sg U69376 ( .A(n46652), .B(n45873), .X(n40297) );
  nand_x1_sg U69377 ( .A(n46648), .B(n45725), .X(n40299) );
  nand_x1_sg U69378 ( .A(n46655), .B(n45723), .X(n40301) );
  nand_x1_sg U69379 ( .A(n46651), .B(n45721), .X(n40303) );
  nand_x1_sg U69380 ( .A(n45613), .B(n46651), .X(n40307) );
  nand_x1_sg U69381 ( .A(n46646), .B(n44815), .X(n40311) );
  nand_x1_sg U69382 ( .A(n46642), .B(n44837), .X(n40313) );
  nand_x1_sg U69383 ( .A(n46653), .B(n45579), .X(n39909) );
  nand_x1_sg U69384 ( .A(n46655), .B(n45565), .X(n40229) );
  nand_x1_sg U69385 ( .A(n46642), .B(n45563), .X(n40269) );
  nand_x1_sg U69386 ( .A(n46642), .B(n45553), .X(n40309) );
  nand_x1_sg U69387 ( .A(n46645), .B(n45571), .X(n39949) );
  nand_x1_sg U69388 ( .A(n46648), .B(n45555), .X(n39989) );
  nand_x1_sg U69389 ( .A(n46646), .B(n45569), .X(n40029) );
  nand_x1_sg U69390 ( .A(n46650), .B(n45573), .X(n40109) );
  nand_x1_sg U69391 ( .A(n46657), .B(n45567), .X(n40149) );
  nand_x1_sg U69392 ( .A(n46654), .B(n45557), .X(n40189) );
  nand_x1_sg U69393 ( .A(n46652), .B(n46191), .X(n39713) );
  nand_x1_sg U69394 ( .A(n46652), .B(n46193), .X(n39715) );
  nand_x1_sg U69395 ( .A(n46655), .B(n46065), .X(n40355) );
  nand_x1_sg U69396 ( .A(n46641), .B(n46057), .X(n40357) );
  nand_x1_sg U69397 ( .A(n46641), .B(n46039), .X(n40361) );
  nand_x1_sg U69398 ( .A(n46652), .B(n46079), .X(n40395) );
  nand_x1_sg U69399 ( .A(n46652), .B(n45231), .X(n40403) );
  nand_x1_sg U69400 ( .A(n46657), .B(n46069), .X(n40435) );
  nand_x1_sg U69401 ( .A(n46652), .B(n46061), .X(n40437) );
  nand_x1_sg U69402 ( .A(n46657), .B(n46037), .X(n40441) );
  nand_x1_sg U69403 ( .A(n46646), .B(n45247), .X(n40345) );
  nand_x1_sg U69404 ( .A(n46645), .B(n45297), .X(n40353) );
  nand_x1_sg U69405 ( .A(n46655), .B(n45253), .X(n40385) );
  nand_x1_sg U69406 ( .A(n46657), .B(n45311), .X(n40393) );
  nand_x1_sg U69407 ( .A(n46653), .B(n45289), .X(n40397) );
  nand_x1_sg U69408 ( .A(n46641), .B(n45279), .X(n40399) );
  nand_x1_sg U69409 ( .A(n46652), .B(n45245), .X(n40425) );
  nand_x1_sg U69410 ( .A(n46651), .B(n45295), .X(n40433) );
  nand_x1_sg U69411 ( .A(n46641), .B(n45991), .X(n40359) );
  nand_x1_sg U69412 ( .A(n46641), .B(n45979), .X(n40363) );
  nand_x1_sg U69413 ( .A(n46651), .B(n45989), .X(n40439) );
  nand_x1_sg U69414 ( .A(n46652), .B(n45977), .X(n40443) );
  nand_x1_sg U69415 ( .A(n46647), .B(n46133), .X(n39317) );
  nand_x1_sg U69416 ( .A(n46647), .B(n46187), .X(n39319) );
  nand_x1_sg U69417 ( .A(n46647), .B(n46131), .X(n39323) );
  nand_x1_sg U69418 ( .A(n46645), .B(n46087), .X(n39345) );
  nand_x1_sg U69419 ( .A(n46647), .B(n46165), .X(n39353) );
  nand_x1_sg U69420 ( .A(n46646), .B(n46105), .X(n39385) );
  nand_x1_sg U69421 ( .A(n46646), .B(n46185), .X(n39393) );
  nand_x1_sg U69422 ( .A(n46652), .B(n46139), .X(n39397) );
  nand_x1_sg U69423 ( .A(n46653), .B(n46153), .X(n39399) );
  nand_x1_sg U69424 ( .A(n46642), .B(n46127), .X(n39403) );
  nand_x1_sg U69425 ( .A(n46645), .B(n46109), .X(n39425) );
  nand_x1_sg U69426 ( .A(n46645), .B(n46183), .X(n39433) );
  nand_x1_sg U69427 ( .A(n46645), .B(n46115), .X(n39465) );
  nand_x1_sg U69428 ( .A(n46645), .B(n46177), .X(n39473) );
  nand_x1_sg U69429 ( .A(n46644), .B(n46151), .X(n39477) );
  nand_x1_sg U69430 ( .A(n46644), .B(n46129), .X(n39479) );
  nand_x1_sg U69431 ( .A(n46644), .B(n46119), .X(n39483) );
  nand_x1_sg U69432 ( .A(n46644), .B(n46107), .X(n39505) );
  nand_x1_sg U69433 ( .A(n46643), .B(n46173), .X(n39513) );
  nand_x1_sg U69434 ( .A(n46643), .B(n46169), .X(n39517) );
  nand_x1_sg U69435 ( .A(n46643), .B(n46141), .X(n39519) );
  nand_x1_sg U69436 ( .A(n46643), .B(n46149), .X(n39521) );
  nand_x1_sg U69437 ( .A(n46651), .B(n46095), .X(n39545) );
  nand_x1_sg U69438 ( .A(n46653), .B(n46181), .X(n39553) );
  nand_x1_sg U69439 ( .A(n46642), .B(n46113), .X(n39585) );
  nand_x1_sg U69440 ( .A(n46642), .B(n46167), .X(n39593) );
  nand_x1_sg U69441 ( .A(n46650), .B(n46143), .X(n39597) );
  nand_x1_sg U69442 ( .A(n46641), .B(n46161), .X(n39599) );
  nand_x1_sg U69443 ( .A(n46647), .B(n46125), .X(n39603) );
  nand_x1_sg U69444 ( .A(n46655), .B(n46103), .X(n39625) );
  nand_x1_sg U69445 ( .A(n46651), .B(n46179), .X(n39633) );
  nand_x1_sg U69446 ( .A(n46653), .B(n46111), .X(n39665) );
  nand_x1_sg U69447 ( .A(n46653), .B(n46159), .X(n39673) );
  nand_x1_sg U69448 ( .A(n46652), .B(n46101), .X(n39705) );
  nand_x1_sg U69449 ( .A(n46653), .B(n46117), .X(n39717) );
  nand_x1_sg U69450 ( .A(n46645), .B(n46093), .X(n39745) );
  nand_x1_sg U69451 ( .A(n46651), .B(n46157), .X(n39753) );
  nand_x1_sg U69452 ( .A(n46643), .B(n46099), .X(n39785) );
  nand_x1_sg U69453 ( .A(n46642), .B(n46171), .X(n39793) );
  nand_x1_sg U69454 ( .A(n46651), .B(n46147), .X(n39797) );
  nand_x1_sg U69455 ( .A(n46651), .B(n46137), .X(n39799) );
  nand_x1_sg U69456 ( .A(n46651), .B(n46123), .X(n39803) );
  nand_x1_sg U69457 ( .A(n46653), .B(n46019), .X(n39351) );
  nand_x1_sg U69458 ( .A(n46646), .B(n46017), .X(n39391) );
  nand_x1_sg U69459 ( .A(n46655), .B(n46011), .X(n39431) );
  nand_x1_sg U69460 ( .A(n46645), .B(n46015), .X(n39471) );
  nand_x1_sg U69461 ( .A(n46643), .B(n46023), .X(n39511) );
  nand_x1_sg U69462 ( .A(n46652), .B(n46009), .X(n39551) );
  nand_x1_sg U69463 ( .A(n46648), .B(n46013), .X(n39591) );
  nand_x1_sg U69464 ( .A(n46647), .B(n46007), .X(n39631) );
  nand_x1_sg U69465 ( .A(n46642), .B(n46005), .X(n39671) );
  nand_x1_sg U69466 ( .A(n46648), .B(n45985), .X(n39711) );
  nand_x1_sg U69467 ( .A(n46646), .B(n45987), .X(n39719) );
  nand_x1_sg U69468 ( .A(n46645), .B(n45983), .X(n39723) );
  nand_x1_sg U69469 ( .A(n46644), .B(n46003), .X(n39751) );
  nand_x1_sg U69470 ( .A(n46648), .B(n46021), .X(n39791) );
  nand_x1_sg U69471 ( .A(n46646), .B(n45967), .X(n39349) );
  nand_x1_sg U69472 ( .A(n46646), .B(n45951), .X(n39389) );
  nand_x1_sg U69473 ( .A(n46644), .B(n45965), .X(n39429) );
  nand_x1_sg U69474 ( .A(n46643), .B(n45971), .X(n39509) );
  nand_x1_sg U69475 ( .A(n46647), .B(n45963), .X(n39549) );
  nand_x1_sg U69476 ( .A(n46654), .B(n45959), .X(n39589) );
  nand_x1_sg U69477 ( .A(n46641), .B(n45961), .X(n39629) );
  nand_x1_sg U69478 ( .A(n46650), .B(n45957), .X(n39669) );
  nand_x1_sg U69479 ( .A(n46652), .B(n45949), .X(n39709) );
  nand_x1_sg U69480 ( .A(n46651), .B(n45955), .X(n39749) );
  nand_x1_sg U69481 ( .A(n46653), .B(n45969), .X(n39789) );
  nand_x1_sg U69482 ( .A(n46650), .B(n45719), .X(n40325) );
  nand_x1_sg U69483 ( .A(n46641), .B(n45939), .X(n40327) );
  nand_x1_sg U69484 ( .A(n46650), .B(n45717), .X(n40329) );
  nand_x1_sg U69485 ( .A(n46650), .B(n45715), .X(n40331) );
  nand_x1_sg U69486 ( .A(n46641), .B(n45713), .X(n40333) );
  nand_x1_sg U69487 ( .A(n46641), .B(n45711), .X(n40335) );
  nand_x1_sg U69488 ( .A(n46650), .B(n45709), .X(n40337) );
  nand_x1_sg U69489 ( .A(n46641), .B(n45707), .X(n40339) );
  nand_x1_sg U69490 ( .A(n46643), .B(n45705), .X(n40341) );
  nand_x1_sg U69491 ( .A(n46641), .B(n45703), .X(n40343) );
  nand_x1_sg U69492 ( .A(n45611), .B(n46653), .X(n40347) );
  nand_x1_sg U69493 ( .A(n46646), .B(n44829), .X(n40351) );
  nand_x1_sg U69494 ( .A(n46641), .B(n45701), .X(n40365) );
  nand_x1_sg U69495 ( .A(n46641), .B(n45933), .X(n40367) );
  nand_x1_sg U69496 ( .A(n46641), .B(n45699), .X(n40369) );
  nand_x1_sg U69497 ( .A(n46641), .B(n45697), .X(n40371) );
  nand_x1_sg U69498 ( .A(n46641), .B(n45927), .X(n40373) );
  nand_x1_sg U69499 ( .A(n46650), .B(n45695), .X(n40375) );
  nand_x1_sg U69500 ( .A(n46647), .B(n45871), .X(n40377) );
  nand_x1_sg U69501 ( .A(n46641), .B(n45693), .X(n40379) );
  nand_x1_sg U69502 ( .A(n46641), .B(n45691), .X(n40381) );
  nand_x1_sg U69503 ( .A(n46648), .B(n45689), .X(n40383) );
  nand_x1_sg U69504 ( .A(n45609), .B(n46641), .X(n40387) );
  nand_x1_sg U69505 ( .A(n46650), .B(n44863), .X(n40391) );
  nand_x1_sg U69506 ( .A(n46654), .B(n44861), .X(n40401) );
  nand_x1_sg U69507 ( .A(n46655), .B(n45687), .X(n40405) );
  nand_x1_sg U69508 ( .A(n46648), .B(n45943), .X(n40407) );
  nand_x1_sg U69509 ( .A(n46651), .B(n45685), .X(n40409) );
  nand_x1_sg U69510 ( .A(n46648), .B(n45683), .X(n40411) );
  nand_x1_sg U69511 ( .A(n46648), .B(n45681), .X(n40413) );
  nand_x1_sg U69512 ( .A(n46648), .B(n45889), .X(n40415) );
  nand_x1_sg U69513 ( .A(n46650), .B(n45895), .X(n40417) );
  nand_x1_sg U69514 ( .A(n46641), .B(n45679), .X(n40419) );
  nand_x1_sg U69515 ( .A(n46646), .B(n45677), .X(n40421) );
  nand_x1_sg U69516 ( .A(n46652), .B(n45675), .X(n40423) );
  nand_x1_sg U69517 ( .A(n45607), .B(n46657), .X(n40427) );
  nand_x1_sg U69518 ( .A(n46657), .B(n44827), .X(n40431) );
  nand_x1_sg U69519 ( .A(n46657), .B(n45673), .X(n40445) );
  nand_x1_sg U69520 ( .A(n46651), .B(n45931), .X(n40447) );
  nand_x1_sg U69521 ( .A(n46652), .B(n45671), .X(n40449) );
  nand_x1_sg U69522 ( .A(n46651), .B(n45669), .X(n40451) );
  nand_x1_sg U69523 ( .A(n46651), .B(n45561), .X(n40349) );
  nand_x1_sg U69524 ( .A(n46655), .B(n45575), .X(n40389) );
  nand_x1_sg U69525 ( .A(n46654), .B(n45559), .X(n40429) );
  nand_x1_sg U69526 ( .A(n46647), .B(n45635), .X(n39321) );
  nand_x1_sg U69527 ( .A(n46647), .B(n45125), .X(n39325) );
  nand_x1_sg U69528 ( .A(n46647), .B(n45207), .X(n39327) );
  nand_x1_sg U69529 ( .A(n46647), .B(n45123), .X(n39329) );
  nand_x1_sg U69530 ( .A(n46647), .B(n45121), .X(n39331) );
  nand_x1_sg U69531 ( .A(n46647), .B(n45119), .X(n39333) );
  nand_x1_sg U69532 ( .A(n46646), .B(n45183), .X(n39335) );
  nand_x1_sg U69533 ( .A(n46647), .B(n45117), .X(n39337) );
  nand_x1_sg U69534 ( .A(n46645), .B(n45115), .X(n39339) );
  nand_x1_sg U69535 ( .A(n46642), .B(n45145), .X(n39341) );
  nand_x1_sg U69536 ( .A(n46643), .B(n45127), .X(n39343) );
  nand_x1_sg U69537 ( .A(n44787), .B(n46645), .X(n39347) );
  nand_x1_sg U69538 ( .A(n46654), .B(n44897), .X(n39355) );
  nand_x1_sg U69539 ( .A(n46655), .B(n44905), .X(n39357) );
  nand_x1_sg U69540 ( .A(n46654), .B(n44819), .X(n39359) );
  nand_x1_sg U69541 ( .A(n46648), .B(n44793), .X(n39361) );
  nand_x1_sg U69542 ( .A(n46647), .B(n44907), .X(n39363) );
  nand_x1_sg U69543 ( .A(n46648), .B(n45113), .X(n39365) );
  nand_x1_sg U69544 ( .A(n46647), .B(n45159), .X(n39367) );
  nand_x1_sg U69545 ( .A(n46654), .B(n45111), .X(n39369) );
  nand_x1_sg U69546 ( .A(n46655), .B(n45109), .X(n39371) );
  nand_x1_sg U69547 ( .A(n46654), .B(n45107), .X(n39373) );
  nand_x1_sg U69548 ( .A(n46654), .B(n45147), .X(n39375) );
  nand_x1_sg U69549 ( .A(n46651), .B(n45105), .X(n39377) );
  nand_x1_sg U69550 ( .A(n46654), .B(n45103), .X(n39379) );
  nand_x1_sg U69551 ( .A(n46646), .B(n45101), .X(n39381) );
  nand_x1_sg U69552 ( .A(n46646), .B(n45099), .X(n39383) );
  nand_x1_sg U69553 ( .A(n44785), .B(n46646), .X(n39387) );
  nand_x1_sg U69554 ( .A(n46646), .B(n44885), .X(n39395) );
  nand_x1_sg U69555 ( .A(n46654), .B(n45639), .X(n39401) );
  nand_x1_sg U69556 ( .A(n46655), .B(n45097), .X(n39405) );
  nand_x1_sg U69557 ( .A(n46641), .B(n45173), .X(n39407) );
  nand_x1_sg U69558 ( .A(n46648), .B(n45095), .X(n39409) );
  nand_x1_sg U69559 ( .A(n46651), .B(n45093), .X(n39411) );
  nand_x1_sg U69560 ( .A(n46643), .B(n45091), .X(n39413) );
  nand_x1_sg U69561 ( .A(n46644), .B(n45153), .X(n39415) );
  nand_x1_sg U69562 ( .A(n46644), .B(n45089), .X(n39417) );
  nand_x1_sg U69563 ( .A(n46643), .B(n45087), .X(n39419) );
  nand_x1_sg U69564 ( .A(n46644), .B(n45085), .X(n39421) );
  nand_x1_sg U69565 ( .A(n46643), .B(n45083), .X(n39423) );
  nand_x1_sg U69566 ( .A(n44783), .B(n46644), .X(n39427) );
  nand_x1_sg U69567 ( .A(n46645), .B(n44873), .X(n39435) );
  nand_x1_sg U69568 ( .A(n46644), .B(n44853), .X(n39437) );
  nand_x1_sg U69569 ( .A(n46645), .B(n44825), .X(n39439) );
  nand_x1_sg U69570 ( .A(n46644), .B(n44313), .X(n39441) );
  nand_x1_sg U69571 ( .A(n46644), .B(n44319), .X(n39443) );
  nand_x1_sg U69572 ( .A(n46645), .B(n45081), .X(n39445) );
  nand_x1_sg U69573 ( .A(n46644), .B(n45169), .X(n39447) );
  nand_x1_sg U69574 ( .A(n46645), .B(n45079), .X(n39449) );
  nand_x1_sg U69575 ( .A(n46644), .B(n45143), .X(n39451) );
  nand_x1_sg U69576 ( .A(n46645), .B(n45077), .X(n39453) );
  nand_x1_sg U69577 ( .A(n46655), .B(n45179), .X(n39455) );
  nand_x1_sg U69578 ( .A(n46655), .B(n45075), .X(n39457) );
  nand_x1_sg U69579 ( .A(n46645), .B(n45073), .X(n39459) );
  nand_x1_sg U69580 ( .A(n46645), .B(n45071), .X(n39461) );
  nand_x1_sg U69581 ( .A(n46645), .B(n45069), .X(n39463) );
  nand_x1_sg U69582 ( .A(n44781), .B(n46645), .X(n39467) );
  nand_x1_sg U69583 ( .A(n46645), .B(n44877), .X(n39475) );
  nand_x1_sg U69584 ( .A(n46644), .B(n45641), .X(n39481) );
  nand_x1_sg U69585 ( .A(n46644), .B(n45067), .X(n39485) );
  nand_x1_sg U69586 ( .A(n46644), .B(n45171), .X(n39487) );
  nand_x1_sg U69587 ( .A(n46644), .B(n45065), .X(n39489) );
  nand_x1_sg U69588 ( .A(n46644), .B(n45137), .X(n39491) );
  nand_x1_sg U69589 ( .A(n46645), .B(n45063), .X(n39493) );
  nand_x1_sg U69590 ( .A(n46645), .B(n45163), .X(n39495) );
  nand_x1_sg U69591 ( .A(n46644), .B(n45061), .X(n39497) );
  nand_x1_sg U69592 ( .A(n46655), .B(n45059), .X(n39499) );
  nand_x1_sg U69593 ( .A(n46645), .B(n45057), .X(n39501) );
  nand_x1_sg U69594 ( .A(n46644), .B(n45055), .X(n39503) );
  nand_x1_sg U69595 ( .A(n44779), .B(n46644), .X(n39507) );
  nand_x1_sg U69596 ( .A(n46643), .B(n44901), .X(n39515) );
  nand_x1_sg U69597 ( .A(n46643), .B(n45633), .X(n39523) );
  nand_x1_sg U69598 ( .A(n46644), .B(n45053), .X(n39525) );
  nand_x1_sg U69599 ( .A(n46651), .B(n45199), .X(n39527) );
  nand_x1_sg U69600 ( .A(n46653), .B(n45051), .X(n39529) );
  nand_x1_sg U69601 ( .A(n46652), .B(n45049), .X(n39531) );
  nand_x1_sg U69602 ( .A(n46641), .B(n45185), .X(n39533) );
  nand_x1_sg U69603 ( .A(n46648), .B(n45047), .X(n39535) );
  nand_x1_sg U69604 ( .A(n46654), .B(n45129), .X(n39537) );
  nand_x1_sg U69605 ( .A(n46647), .B(n45045), .X(n39539) );
  nand_x1_sg U69606 ( .A(n46642), .B(n45043), .X(n39541) );
  nand_x1_sg U69607 ( .A(n46650), .B(n45041), .X(n39543) );
  nand_x1_sg U69608 ( .A(n44777), .B(n46646), .X(n39547) );
  nand_x1_sg U69609 ( .A(n46650), .B(n44871), .X(n39555) );
  nand_x1_sg U69610 ( .A(n46642), .B(n44851), .X(n39557) );
  nand_x1_sg U69611 ( .A(n46641), .B(n44823), .X(n39559) );
  nand_x1_sg U69612 ( .A(n46647), .B(n44311), .X(n39561) );
  nand_x1_sg U69613 ( .A(n46648), .B(n44317), .X(n39563) );
  nand_x1_sg U69614 ( .A(n46654), .B(n45039), .X(n39565) );
  nand_x1_sg U69615 ( .A(n46642), .B(n45167), .X(n39567) );
  nand_x1_sg U69616 ( .A(n46646), .B(n45037), .X(n39569) );
  nand_x1_sg U69617 ( .A(n46643), .B(n45141), .X(n39571) );
  nand_x1_sg U69618 ( .A(n46642), .B(n45035), .X(n39573) );
  nand_x1_sg U69619 ( .A(n46642), .B(n45177), .X(n39575) );
  nand_x1_sg U69620 ( .A(n46642), .B(n45033), .X(n39577) );
  nand_x1_sg U69621 ( .A(n46642), .B(n45031), .X(n39579) );
  nand_x1_sg U69622 ( .A(n46650), .B(n45029), .X(n39581) );
  nand_x1_sg U69623 ( .A(n46641), .B(n45027), .X(n39583) );
  nand_x1_sg U69624 ( .A(n44775), .B(n46647), .X(n39587) );
  nand_x1_sg U69625 ( .A(n46642), .B(n44887), .X(n39595) );
  nand_x1_sg U69626 ( .A(n46652), .B(n45637), .X(n39601) );
  nand_x1_sg U69627 ( .A(n46646), .B(n45025), .X(n39605) );
  nand_x1_sg U69628 ( .A(n46644), .B(n45181), .X(n39607) );
  nand_x1_sg U69629 ( .A(n46650), .B(n45023), .X(n39609) );
  nand_x1_sg U69630 ( .A(n46644), .B(n45021), .X(n39611) );
  nand_x1_sg U69631 ( .A(n46654), .B(n45019), .X(n39613) );
  nand_x1_sg U69632 ( .A(n46651), .B(n45161), .X(n39615) );
  nand_x1_sg U69633 ( .A(n46651), .B(n45017), .X(n39617) );
  nand_x1_sg U69634 ( .A(n46653), .B(n45015), .X(n39619) );
  nand_x1_sg U69635 ( .A(n46643), .B(n45013), .X(n39621) );
  nand_x1_sg U69636 ( .A(n46651), .B(n45011), .X(n39623) );
  nand_x1_sg U69637 ( .A(n44773), .B(n46652), .X(n39627) );
  nand_x1_sg U69638 ( .A(n46648), .B(n44869), .X(n39635) );
  nand_x1_sg U69639 ( .A(n46642), .B(n44849), .X(n39637) );
  nand_x1_sg U69640 ( .A(n46642), .B(n44821), .X(n39639) );
  nand_x1_sg U69641 ( .A(n46642), .B(n44309), .X(n39641) );
  nand_x1_sg U69642 ( .A(n46642), .B(n44315), .X(n39643) );
  nand_x1_sg U69643 ( .A(n46642), .B(n45009), .X(n39645) );
  nand_x1_sg U69644 ( .A(n46642), .B(n45165), .X(n39647) );
  nand_x1_sg U69645 ( .A(n46642), .B(n45007), .X(n39649) );
  nand_x1_sg U69646 ( .A(n46642), .B(n45139), .X(n39651) );
  nand_x1_sg U69647 ( .A(n46653), .B(n45005), .X(n39653) );
  nand_x1_sg U69648 ( .A(n46642), .B(n45175), .X(n39655) );
  nand_x1_sg U69649 ( .A(n46645), .B(n45003), .X(n39657) );
  nand_x1_sg U69650 ( .A(n46642), .B(n45001), .X(n39659) );
  nand_x1_sg U69651 ( .A(n46646), .B(n44999), .X(n39661) );
  nand_x1_sg U69652 ( .A(n46642), .B(n44997), .X(n39663) );
  nand_x1_sg U69653 ( .A(n44771), .B(n46643), .X(n39667) );
  nand_x1_sg U69654 ( .A(n46653), .B(n44891), .X(n39675) );
  nand_x1_sg U69655 ( .A(n46642), .B(n44881), .X(n39677) );
  nand_x1_sg U69656 ( .A(n46653), .B(n44807), .X(n39679) );
  nand_x1_sg U69657 ( .A(n46642), .B(n44813), .X(n39681) );
  nand_x1_sg U69658 ( .A(n46654), .B(n44801), .X(n39683) );
  nand_x1_sg U69659 ( .A(n46652), .B(n44995), .X(n39685) );
  nand_x1_sg U69660 ( .A(n46643), .B(n45197), .X(n39687) );
  nand_x1_sg U69661 ( .A(n46655), .B(n44993), .X(n39689) );
  nand_x1_sg U69662 ( .A(n46642), .B(n44991), .X(n39691) );
  nand_x1_sg U69663 ( .A(n46646), .B(n45191), .X(n39693) );
  nand_x1_sg U69664 ( .A(n46644), .B(n44989), .X(n39695) );
  nand_x1_sg U69665 ( .A(n46644), .B(n45135), .X(n39697) );
  nand_x1_sg U69666 ( .A(n46644), .B(n44987), .X(n39699) );
  nand_x1_sg U69667 ( .A(n46650), .B(n44985), .X(n39701) );
  nand_x1_sg U69668 ( .A(n46641), .B(n44983), .X(n39703) );
  nand_x1_sg U69669 ( .A(n44769), .B(n46647), .X(n39707) );
  nand_x1_sg U69670 ( .A(n46643), .B(n44833), .X(n39721) );
  nand_x1_sg U69671 ( .A(n46644), .B(n44981), .X(n39725) );
  nand_x1_sg U69672 ( .A(n46650), .B(n45201), .X(n39727) );
  nand_x1_sg U69673 ( .A(n46643), .B(n44979), .X(n39729) );
  nand_x1_sg U69674 ( .A(n46645), .B(n44977), .X(n39731) );
  nand_x1_sg U69675 ( .A(n46644), .B(n44975), .X(n39733) );
  nand_x1_sg U69676 ( .A(n46645), .B(n44973), .X(n39735) );
  nand_x1_sg U69677 ( .A(n46652), .B(n44971), .X(n39737) );
  nand_x1_sg U69678 ( .A(n46646), .B(n44969), .X(n39739) );
  nand_x1_sg U69679 ( .A(n46654), .B(n44967), .X(n39741) );
  nand_x1_sg U69680 ( .A(n46643), .B(n44965), .X(n39743) );
  nand_x1_sg U69681 ( .A(n44767), .B(n46650), .X(n39747) );
  nand_x1_sg U69682 ( .A(n46653), .B(n44889), .X(n39755) );
  nand_x1_sg U69683 ( .A(n46650), .B(n44879), .X(n39757) );
  nand_x1_sg U69684 ( .A(n46641), .B(n44805), .X(n39759) );
  nand_x1_sg U69685 ( .A(n46647), .B(n44811), .X(n39761) );
  nand_x1_sg U69686 ( .A(n46648), .B(n44799), .X(n39763) );
  nand_x1_sg U69687 ( .A(n46654), .B(n44963), .X(n39765) );
  nand_x1_sg U69688 ( .A(n46646), .B(n45195), .X(n39767) );
  nand_x1_sg U69689 ( .A(n46645), .B(n44961), .X(n39769) );
  nand_x1_sg U69690 ( .A(n46643), .B(n44959), .X(n39771) );
  nand_x1_sg U69691 ( .A(n46651), .B(n45189), .X(n39773) );
  nand_x1_sg U69692 ( .A(n46645), .B(n44957), .X(n39775) );
  nand_x1_sg U69693 ( .A(n46651), .B(n45133), .X(n39777) );
  nand_x1_sg U69694 ( .A(n46653), .B(n44955), .X(n39779) );
  nand_x1_sg U69695 ( .A(n46650), .B(n44953), .X(n39781) );
  nand_x1_sg U69696 ( .A(n46641), .B(n44951), .X(n39783) );
  nand_x1_sg U69697 ( .A(n44765), .B(n46647), .X(n39787) );
  nand_x1_sg U69698 ( .A(n46654), .B(n44895), .X(n39795) );
  nand_x1_sg U69699 ( .A(n46655), .B(n45645), .X(n39801) );
  nand_x1_sg U69700 ( .A(n46646), .B(n44949), .X(n39805) );
  nand_x1_sg U69701 ( .A(n46647), .B(n45205), .X(n39807) );
  nand_x1_sg U69702 ( .A(n46645), .B(n44947), .X(n39809) );
  nand_x1_sg U69703 ( .A(n46647), .B(n44945), .X(n39811) );
  nand_x1_sg U69704 ( .A(n46645), .B(n45581), .X(n39469) );
  nand_x1_sg U69705 ( .A(n46657), .B(n46200), .X(n40511) );
  nand_x1_sg U69706 ( .A(n46650), .B(n46195), .X(n40513) );
  nand_x1_sg U69707 ( .A(n46641), .B(n46081), .X(n40475) );
  nand_x1_sg U69708 ( .A(n46651), .B(n45229), .X(n40483) );
  nand_x1_sg U69709 ( .A(n46643), .B(n45251), .X(n40465) );
  nand_x1_sg U69710 ( .A(n46652), .B(n45315), .X(n40473) );
  nand_x1_sg U69711 ( .A(n46644), .B(n45287), .X(n40477) );
  nand_x1_sg U69712 ( .A(n46654), .B(n45277), .X(n40479) );
  nand_x1_sg U69713 ( .A(n46651), .B(n45243), .X(n40505) );
  nand_x1_sg U69714 ( .A(n46650), .B(n45925), .X(n40453) );
  nand_x1_sg U69715 ( .A(n46641), .B(n45667), .X(n40455) );
  nand_x1_sg U69716 ( .A(n46641), .B(n45869), .X(n40457) );
  nand_x1_sg U69717 ( .A(n46654), .B(n45665), .X(n40459) );
  nand_x1_sg U69718 ( .A(n46641), .B(n45663), .X(n40461) );
  nand_x1_sg U69719 ( .A(n46641), .B(n45661), .X(n40463) );
  nand_x1_sg U69720 ( .A(n45605), .B(n46641), .X(n40467) );
  nand_x1_sg U69721 ( .A(n46655), .B(n44875), .X(n40471) );
  nand_x1_sg U69722 ( .A(n46643), .B(n44859), .X(n40481) );
  nand_x1_sg U69723 ( .A(n46644), .B(n45659), .X(n40485) );
  nand_x1_sg U69724 ( .A(n46651), .B(n45941), .X(n40487) );
  nand_x1_sg U69725 ( .A(n46643), .B(n45657), .X(n40489) );
  nand_x1_sg U69726 ( .A(n46653), .B(n45655), .X(n40491) );
  nand_x1_sg U69727 ( .A(n46646), .B(n45653), .X(n40493) );
  nand_x1_sg U69728 ( .A(n46641), .B(n45887), .X(n40495) );
  nand_x1_sg U69729 ( .A(n46645), .B(n45893), .X(n40497) );
  nand_x1_sg U69730 ( .A(n46653), .B(n45651), .X(n40499) );
  nand_x1_sg U69731 ( .A(n46652), .B(n45649), .X(n40501) );
  nand_x1_sg U69732 ( .A(n46643), .B(n45647), .X(n40503) );
  nand_x1_sg U69733 ( .A(n45603), .B(n46653), .X(n40507) );
  nand_x1_sg U69734 ( .A(n46651), .B(n45577), .X(n40469) );
  nand_x1_sg U69735 ( .A(n46648), .B(n46163), .X(n39313) );
  nand_x1_sg U69736 ( .A(n46648), .B(n46027), .X(n39311) );
  nand_x1_sg U69737 ( .A(n46648), .B(n45975), .X(n39309) );
  nand_x1_sg U69738 ( .A(n46648), .B(n44903), .X(n39315) );
  nand_x4_sg U69739 ( .A(n40516), .B(input_ready), .X(n39303) );
  nor_x1_sg U69740 ( .A(state[0]), .B(state[1]), .X(n40516) );
  nand_x1_sg U69741 ( .A(n39297), .B(state[0]), .X(n39293) );
  nor_x1_sg U69742 ( .A(n39296), .B(n39297), .X(n39295) );
  nand_x1_sg U69743 ( .A(n39297), .B(state[1]), .X(n39298) );
  nand_x1_sg U69744 ( .A(n39296), .B(n46576), .X(n39299) );
  nor_x1_sg U69745 ( .A(n40721), .B(n24417), .X(n24459) );
  nor_x1_sg U69746 ( .A(n40722), .B(n32083), .X(n32125) );
  nor_x1_sg U69747 ( .A(n52681), .B(n27043), .X(n27042) );
  nand_x1_sg U69748 ( .A(n46191), .B(n28394), .X(n28453) );
  nand_x1_sg U69749 ( .A(n28389), .B(n46193), .X(n28450) );
  nand_x2_sg U69750 ( .A(n8345), .B(n30515), .X(n30514) );
  nand_x2_sg U69751 ( .A(n8645), .B(n22849), .X(n22848) );
  nand_x2_sg U69752 ( .A(n8765), .B(n22809), .X(n22810) );
  nand_x2_sg U69753 ( .A(n8465), .B(n30475), .X(n30476) );
  nand_x2_sg U69754 ( .A(n8349), .B(n31391), .X(n31390) );
  nand_x2_sg U69755 ( .A(n8649), .B(n23725), .X(n23724) );
  nand_x2_sg U69756 ( .A(n8347), .B(n30996), .X(n30995) );
  nand_x2_sg U69757 ( .A(n8647), .B(n23330), .X(n23329) );
  nand_x2_sg U69758 ( .A(n8767), .B(n23290), .X(n23291) );
  nand_x2_sg U69759 ( .A(n8769), .B(n23685), .X(n23686) );
  nand_x2_sg U69760 ( .A(n8771), .B(n24009), .X(n24010) );
  nand_x2_sg U69761 ( .A(n8467), .B(n30956), .X(n30957) );
  nand_x2_sg U69762 ( .A(n8469), .B(n31351), .X(n31352) );
  nand_x2_sg U69763 ( .A(n8471), .B(n31675), .X(n31676) );
  nand_x2_sg U69764 ( .A(n8773), .B(n24269), .X(n24270) );
  nand_x2_sg U69765 ( .A(n8473), .B(n31935), .X(n31936) );
  nor_x1_sg U69766 ( .A(n51159), .B(n45209), .X(n28390) );
  nand_x1_sg U69767 ( .A(n26130), .B(n46127), .X(n26203) );
  nand_x1_sg U69768 ( .A(n26687), .B(n46119), .X(n26760) );
  nand_x1_sg U69769 ( .A(n46125), .B(n27525), .X(n27598) );
  nand_x1_sg U69770 ( .A(n46131), .B(n25569), .X(n25644) );
  nand_x1_sg U69771 ( .A(n28921), .B(n46123), .X(n28994) );
  nand_x1_sg U69772 ( .A(n29482), .B(n46121), .X(n29555) );
  nand_x1_sg U69773 ( .A(n28383), .B(n46117), .X(n28447) );
  nand_x4_sg U69774 ( .A(n45947), .B(n51043), .X(n26725) );
  nor_x1_sg U69775 ( .A(n51069), .B(n46033), .X(n26968) );
  nand_x1_sg U69776 ( .A(n46033), .B(n51069), .X(n26969) );
  nor_x1_sg U69777 ( .A(n50973), .B(n45237), .X(n25571) );
  nand_x1_sg U69778 ( .A(n45237), .B(n50973), .X(n25572) );
  nor_x1_sg U69779 ( .A(n51011), .B(n45235), .X(n26132) );
  nand_x1_sg U69780 ( .A(n45235), .B(n51011), .X(n26133) );
  nor_x1_sg U69781 ( .A(n51107), .B(n45233), .X(n27527) );
  nand_x1_sg U69782 ( .A(n45233), .B(n51107), .X(n27528) );
  nor_x1_sg U69783 ( .A(n51201), .B(n45231), .X(n28923) );
  nand_x1_sg U69784 ( .A(n45231), .B(n51201), .X(n28924) );
  nor_x1_sg U69785 ( .A(n51239), .B(n45229), .X(n29484) );
  nand_x1_sg U69786 ( .A(n45229), .B(n51239), .X(n29485) );
  nor_x1_sg U69787 ( .A(n51050), .B(n45227), .X(n26689) );
  nand_x1_sg U69788 ( .A(n45227), .B(n51050), .X(n26690) );
  nor_x1_sg U69789 ( .A(n40853), .B(n23637), .X(n23636) );
  nor_x1_sg U69790 ( .A(n40854), .B(n31303), .X(n31302) );
  nor_x1_sg U69791 ( .A(n40855), .B(n31285), .X(n31284) );
  nor_x1_sg U69792 ( .A(n40856), .B(n23619), .X(n23618) );
  nor_x1_sg U69793 ( .A(n41151), .B(n8350), .X(n31319) );
  nor_x1_sg U69794 ( .A(n41203), .B(n8650), .X(n23653) );
  nor_x1_sg U69795 ( .A(n41886), .B(n8344), .X(n30511) );
  nor_x1_sg U69796 ( .A(n41888), .B(n8644), .X(n22845) );
  nor_x1_sg U69797 ( .A(n40857), .B(n49401), .X(n31272) );
  nor_x1_sg U69798 ( .A(n40858), .B(n50260), .X(n23606) );
  nor_x1_sg U69799 ( .A(n40859), .B(n41195), .X(n24376) );
  nor_x1_sg U69800 ( .A(n40860), .B(n41205), .X(n32042) );
  nor_x1_sg U69801 ( .A(n40861), .B(n41201), .X(n23500) );
  nor_x1_sg U69802 ( .A(n40862), .B(n41199), .X(n23861) );
  nor_x1_sg U69803 ( .A(n40863), .B(n41197), .X(n24158) );
  nor_x1_sg U69804 ( .A(n40864), .B(n41153), .X(n24361) );
  nor_x1_sg U69805 ( .A(n40865), .B(n41160), .X(n32027) );
  nor_x1_sg U69806 ( .A(n40866), .B(n41211), .X(n31166) );
  nor_x1_sg U69807 ( .A(n40867), .B(n41209), .X(n31527) );
  nor_x1_sg U69808 ( .A(n40868), .B(n41207), .X(n31824) );
  nand_x1_sg U69809 ( .A(n43759), .B(n51162), .X(n28373) );
  nand_x4_sg U69810 ( .A(n45835), .B(n51012), .X(n26127) );
  nand_x4_sg U69811 ( .A(n45805), .B(n51051), .X(n26684) );
  nand_x4_sg U69812 ( .A(n45763), .B(n51108), .X(n27522) );
  nand_x4_sg U69813 ( .A(n45863), .B(n50974), .X(n25566) );
  nand_x4_sg U69814 ( .A(n45859), .B(n50977), .X(n25550) );
  nand_x4_sg U69815 ( .A(n45857), .B(n50978), .X(n25544) );
  nand_x4_sg U69816 ( .A(n45719), .B(n51164), .X(n28361) );
  nand_x4_sg U69817 ( .A(n45687), .B(n51202), .X(n28918) );
  nand_x4_sg U69818 ( .A(n45659), .B(n51240), .X(n29479) );
  nand_x4_sg U69819 ( .A(n45861), .B(n50976), .X(n25554) );
  nand_x4_sg U69820 ( .A(n45717), .B(n51166), .X(n28349) );
  nand_x4_sg U69821 ( .A(n45685), .B(n51204), .X(n28906) );
  nand_x4_sg U69822 ( .A(n45657), .B(n51242), .X(n29467) );
  nand_x4_sg U69823 ( .A(n45945), .B(n50975), .X(n25560) );
  nand_x4_sg U69824 ( .A(n45939), .B(n51165), .X(n28355) );
  nand_x4_sg U69825 ( .A(n45943), .B(n51203), .X(n28912) );
  nand_x4_sg U69826 ( .A(n45941), .B(n51241), .X(n29473) );
  nand_x4_sg U69827 ( .A(n45897), .B(n50994), .X(n25841) );
  nand_x4_sg U69828 ( .A(n45907), .B(n51032), .X(n26400) );
  nand_x4_sg U69829 ( .A(n45937), .B(n51071), .X(n26957) );
  nand_x4_sg U69830 ( .A(n45905), .B(n51090), .X(n27237) );
  nand_x4_sg U69831 ( .A(n45903), .B(n51128), .X(n27795) );
  nand_x4_sg U69832 ( .A(n45935), .B(n51147), .X(n28076) );
  nand_x4_sg U69833 ( .A(n45933), .B(n51184), .X(n28634) );
  nand_x4_sg U69834 ( .A(n45931), .B(n51222), .X(n29195) );
  nand_x4_sg U69835 ( .A(n45851), .B(n50993), .X(n25847) );
  nand_x4_sg U69836 ( .A(n45819), .B(n51031), .X(n26406) );
  nand_x4_sg U69837 ( .A(n45791), .B(n51070), .X(n26963) );
  nand_x4_sg U69838 ( .A(n45777), .B(n51089), .X(n27243) );
  nand_x4_sg U69839 ( .A(n45747), .B(n51127), .X(n27801) );
  nand_x4_sg U69840 ( .A(n45733), .B(n51146), .X(n28082) );
  nand_x4_sg U69841 ( .A(n45701), .B(n51183), .X(n28640) );
  nand_x4_sg U69842 ( .A(n45673), .B(n51221), .X(n29201) );
  nand_x4_sg U69843 ( .A(n45865), .B(n50983), .X(n25613) );
  nand_x4_sg U69844 ( .A(n45749), .B(n51117), .X(n27569) );
  nand_x4_sg U69845 ( .A(n45883), .B(n50982), .X(n25619) );
  nand_x4_sg U69846 ( .A(n45837), .B(n51002), .X(n25894) );
  nand_x4_sg U69847 ( .A(n45821), .B(n51021), .X(n26174) );
  nand_x4_sg U69848 ( .A(n45825), .B(n51019), .X(n26085) );
  nand_x4_sg U69849 ( .A(n45807), .B(n51040), .X(n26453) );
  nand_x4_sg U69850 ( .A(n45811), .B(n51038), .X(n26364) );
  nand_x4_sg U69851 ( .A(n45793), .B(n51060), .X(n26731) );
  nand_x4_sg U69852 ( .A(n45797), .B(n51058), .X(n26642) );
  nand_x4_sg U69853 ( .A(n45779), .B(n51079), .X(n27010) );
  nand_x4_sg U69854 ( .A(n45765), .B(n51098), .X(n27290) );
  nand_x4_sg U69855 ( .A(n45769), .B(n51096), .X(n27201) );
  nand_x4_sg U69856 ( .A(n45751), .B(n51116), .X(n27575) );
  nand_x4_sg U69857 ( .A(n45735), .B(n51136), .X(n27848) );
  nand_x4_sg U69858 ( .A(n45739), .B(n51134), .X(n27759) );
  nand_x4_sg U69859 ( .A(n45721), .B(n51155), .X(n28129) );
  nand_x4_sg U69860 ( .A(n45703), .B(n51173), .X(n28408) );
  nand_x4_sg U69861 ( .A(n45689), .B(n51192), .X(n28687) );
  nand_x4_sg U69862 ( .A(n45675), .B(n51211), .X(n28965) );
  nand_x4_sg U69863 ( .A(n45661), .B(n51230), .X(n29248) );
  nand_x4_sg U69864 ( .A(n45647), .B(n51249), .X(n29526) );
  nand_x4_sg U69865 ( .A(n45839), .B(n51001), .X(n25900) );
  nand_x4_sg U69866 ( .A(n45823), .B(n51020), .X(n26180) );
  nand_x4_sg U69867 ( .A(n45827), .B(n51018), .X(n26091) );
  nand_x4_sg U69868 ( .A(n45809), .B(n51039), .X(n26459) );
  nand_x4_sg U69869 ( .A(n45813), .B(n51037), .X(n26370) );
  nand_x4_sg U69870 ( .A(n45795), .B(n51059), .X(n26737) );
  nand_x4_sg U69871 ( .A(n45799), .B(n51057), .X(n26648) );
  nand_x4_sg U69872 ( .A(n45781), .B(n51078), .X(n27016) );
  nand_x4_sg U69873 ( .A(n45767), .B(n51097), .X(n27296) );
  nand_x4_sg U69874 ( .A(n45771), .B(n51095), .X(n27207) );
  nand_x4_sg U69875 ( .A(n45737), .B(n51135), .X(n27854) );
  nand_x4_sg U69876 ( .A(n45741), .B(n51133), .X(n27765) );
  nand_x4_sg U69877 ( .A(n45723), .B(n51154), .X(n28135) );
  nand_x4_sg U69878 ( .A(n45705), .B(n51172), .X(n28414) );
  nand_x4_sg U69879 ( .A(n45691), .B(n51191), .X(n28693) );
  nand_x4_sg U69880 ( .A(n45677), .B(n51210), .X(n28971) );
  nand_x4_sg U69881 ( .A(n45663), .B(n51229), .X(n29254) );
  nand_x4_sg U69882 ( .A(n45649), .B(n51248), .X(n29532) );
  nand_x4_sg U69883 ( .A(n45921), .B(n50979), .X(n25538) );
  nand_x4_sg U69884 ( .A(n45855), .B(n50980), .X(n25532) );
  nand_x4_sg U69885 ( .A(n45849), .B(n50995), .X(n25835) );
  nand_x4_sg U69886 ( .A(n45847), .B(n50996), .X(n25829) );
  nand_x4_sg U69887 ( .A(n45845), .B(n50997), .X(n25823) );
  nand_x4_sg U69888 ( .A(n45885), .B(n50998), .X(n25817) );
  nand_x4_sg U69889 ( .A(n45843), .B(n50999), .X(n25811) );
  nand_x4_sg U69890 ( .A(n45911), .B(n51013), .X(n26121) );
  nand_x4_sg U69891 ( .A(n45833), .B(n51014), .X(n26115) );
  nand_x4_sg U69892 ( .A(n45831), .B(n51015), .X(n26109) );
  nand_x4_sg U69893 ( .A(n45829), .B(n51016), .X(n26103) );
  nand_x4_sg U69894 ( .A(n45891), .B(n51017), .X(n26097) );
  nand_x4_sg U69895 ( .A(n45817), .B(n51033), .X(n26394) );
  nand_x4_sg U69896 ( .A(n45881), .B(n51034), .X(n26388) );
  nand_x4_sg U69897 ( .A(n45815), .B(n51035), .X(n26382) );
  nand_x4_sg U69898 ( .A(n45917), .B(n51036), .X(n26376) );
  nand_x4_sg U69899 ( .A(n45909), .B(n51052), .X(n26678) );
  nand_x4_sg U69900 ( .A(n45803), .B(n51053), .X(n26672) );
  nand_x4_sg U69901 ( .A(n45875), .B(n51054), .X(n26666) );
  nand_x4_sg U69902 ( .A(n45801), .B(n51055), .X(n26660) );
  nand_x4_sg U69903 ( .A(n45901), .B(n51056), .X(n26654) );
  nand_x4_sg U69904 ( .A(n45789), .B(n51072), .X(n26951) );
  nand_x4_sg U69905 ( .A(n45787), .B(n51073), .X(n26945) );
  nand_x4_sg U69906 ( .A(n45923), .B(n51074), .X(n26939) );
  nand_x4_sg U69907 ( .A(n45785), .B(n51075), .X(n26933) );
  nand_x4_sg U69908 ( .A(n45867), .B(n51076), .X(n26927) );
  nand_x4_sg U69909 ( .A(n45775), .B(n51091), .X(n27231) );
  nand_x4_sg U69910 ( .A(n45879), .B(n51092), .X(n27225) );
  nand_x4_sg U69911 ( .A(n45773), .B(n51093), .X(n27219) );
  nand_x4_sg U69912 ( .A(n45915), .B(n51094), .X(n27213) );
  nand_x4_sg U69913 ( .A(n45919), .B(n51109), .X(n27516) );
  nand_x4_sg U69914 ( .A(n45761), .B(n51110), .X(n27510) );
  nand_x4_sg U69915 ( .A(n45759), .B(n51111), .X(n27504) );
  nand_x4_sg U69916 ( .A(n45757), .B(n51112), .X(n27498) );
  nand_x4_sg U69917 ( .A(n45899), .B(n51113), .X(n27492) );
  nand_x4_sg U69918 ( .A(n45755), .B(n51114), .X(n27486) );
  nand_x4_sg U69919 ( .A(n45745), .B(n51129), .X(n27789) );
  nand_x4_sg U69920 ( .A(n45877), .B(n51130), .X(n27783) );
  nand_x4_sg U69921 ( .A(n45743), .B(n51131), .X(n27777) );
  nand_x4_sg U69922 ( .A(n45913), .B(n51132), .X(n27771) );
  nand_x4_sg U69923 ( .A(n45731), .B(n51148), .X(n28070) );
  nand_x4_sg U69924 ( .A(n45729), .B(n51149), .X(n28064) );
  nand_x4_sg U69925 ( .A(n45929), .B(n51150), .X(n28058) );
  nand_x4_sg U69926 ( .A(n45727), .B(n51151), .X(n28052) );
  nand_x4_sg U69927 ( .A(n45873), .B(n51152), .X(n28046) );
  nand_x4_sg U69928 ( .A(n45715), .B(n51167), .X(n28345) );
  nand_x4_sg U69929 ( .A(n45713), .B(n51168), .X(n28339) );
  nand_x4_sg U69930 ( .A(n45711), .B(n51169), .X(n28333) );
  nand_x4_sg U69931 ( .A(n45709), .B(n51170), .X(n28327) );
  nand_x4_sg U69932 ( .A(n45699), .B(n51185), .X(n28628) );
  nand_x4_sg U69933 ( .A(n45697), .B(n51186), .X(n28622) );
  nand_x4_sg U69934 ( .A(n45927), .B(n51187), .X(n28616) );
  nand_x4_sg U69935 ( .A(n45695), .B(n51188), .X(n28610) );
  nand_x4_sg U69936 ( .A(n45871), .B(n51189), .X(n28604) );
  nand_x4_sg U69937 ( .A(n45683), .B(n51205), .X(n28902) );
  nand_x4_sg U69938 ( .A(n45681), .B(n51206), .X(n28896) );
  nand_x4_sg U69939 ( .A(n45889), .B(n51207), .X(n28890) );
  nand_x4_sg U69940 ( .A(n45895), .B(n51208), .X(n28884) );
  nand_x4_sg U69941 ( .A(n45671), .B(n51223), .X(n29189) );
  nand_x4_sg U69942 ( .A(n45669), .B(n51224), .X(n29183) );
  nand_x4_sg U69943 ( .A(n45925), .B(n51225), .X(n29177) );
  nand_x4_sg U69944 ( .A(n45667), .B(n51226), .X(n29171) );
  nand_x4_sg U69945 ( .A(n45869), .B(n51227), .X(n29165) );
  nand_x4_sg U69946 ( .A(n45655), .B(n51243), .X(n29463) );
  nand_x4_sg U69947 ( .A(n45653), .B(n51244), .X(n29457) );
  nand_x4_sg U69948 ( .A(n45887), .B(n51245), .X(n29451) );
  nand_x4_sg U69949 ( .A(n45893), .B(n51246), .X(n29445) );
  nand_x4_sg U69950 ( .A(n45651), .B(n51247), .X(n29439) );
  nand_x4_sg U69951 ( .A(n45853), .B(n50981), .X(n25526) );
  nand_x4_sg U69952 ( .A(n45841), .B(n51000), .X(n25805) );
  nand_x4_sg U69953 ( .A(n45783), .B(n51077), .X(n26921) );
  nand_x4_sg U69954 ( .A(n45753), .B(n51115), .X(n27480) );
  nand_x4_sg U69955 ( .A(n45725), .B(n51153), .X(n28040) );
  nand_x4_sg U69956 ( .A(n45707), .B(n51171), .X(n28321) );
  nand_x4_sg U69957 ( .A(n45693), .B(n51190), .X(n28598) );
  nand_x4_sg U69958 ( .A(n45679), .B(n51209), .X(n28878) );
  nand_x4_sg U69959 ( .A(n45665), .B(n51228), .X(n29159) );
  nand_x2_sg U69960 ( .A(n8622), .B(n10252), .X(n23169) );
  nand_x2_sg U69961 ( .A(n8582), .B(n10260), .X(n22670) );
  nand_x2_sg U69962 ( .A(n8322), .B(n25360), .X(n30835) );
  nand_x2_sg U69963 ( .A(n8282), .B(n25367), .X(n30336) );
  nand_x2_sg U69964 ( .A(n8562), .B(n10257), .X(n22401) );
  nand_x2_sg U69965 ( .A(n8262), .B(n25364), .X(n30066) );
  nand_x2_sg U69966 ( .A(n8402), .B(n25349), .X(n31590) );
  nand_x2_sg U69967 ( .A(n8542), .B(n10279), .X(n22244) );
  nand_x2_sg U69968 ( .A(n8242), .B(n25385), .X(n29909) );
  nand_x2_sg U69969 ( .A(n8522), .B(n10280), .X(n22053) );
  nand_x2_sg U69970 ( .A(n8702), .B(n10241), .X(n23924) );
  nand_x2_sg U69971 ( .A(n8222), .B(n25386), .X(n29718) );
  nand_x2_sg U69972 ( .A(n8602), .B(n10255), .X(n22921) );
  nand_x2_sg U69973 ( .A(n8642), .B(n10240), .X(n23384) );
  nand_x2_sg U69974 ( .A(n8302), .B(n25363), .X(n30587) );
  nand_x2_sg U69975 ( .A(n8342), .B(n25353), .X(n31050) );
  nand_x2_sg U69976 ( .A(n8762), .B(n10273), .X(n24309) );
  nand_x2_sg U69977 ( .A(n8362), .B(n25382), .X(n31248) );
  nand_x2_sg U69978 ( .A(n8722), .B(n10272), .X(n24068) );
  nand_x2_sg U69979 ( .A(n8462), .B(n25379), .X(n31975) );
  nand_x2_sg U69980 ( .A(n8662), .B(n10276), .X(n23582) );
  nand_x2_sg U69981 ( .A(n8422), .B(n25378), .X(n31734) );
  nand_x1_sg U69982 ( .A(n44321), .B(n45633), .X(n27040) );
  nand_x1_sg U69983 ( .A(n45969), .B(n54605), .X(n28955) );
  nand_x1_sg U69984 ( .A(n45973), .B(n55173), .X(n29516) );
  nand_x1_sg U69985 ( .A(n45951), .B(n51810), .X(n26164) );
  nand_x1_sg U69986 ( .A(n45959), .B(n53198), .X(n27559) );
  nand_x1_sg U69987 ( .A(n45967), .B(n51528), .X(n25884) );
  nand_x1_sg U69988 ( .A(n45965), .B(n52086), .X(n26443) );
  nand_x1_sg U69989 ( .A(n45963), .B(n52920), .X(n27280) );
  nand_x1_sg U69990 ( .A(n45961), .B(n53478), .X(n27838) );
  nand_x2_sg U69991 ( .A(n8565), .B(n50907), .X(n22871) );
  nand_x2_sg U69992 ( .A(n8265), .B(n50048), .X(n30537) );
  nand_x2_sg U69993 ( .A(n8566), .B(n50859), .X(n22874) );
  nand_x2_sg U69994 ( .A(n8567), .B(n50815), .X(n22877) );
  nand_x2_sg U69995 ( .A(n8266), .B(n50000), .X(n30540) );
  nand_x2_sg U69996 ( .A(n8267), .B(n49956), .X(n30543) );
  nand_x2_sg U69997 ( .A(n8738), .B(n50313), .X(n24298) );
  nand_x2_sg U69998 ( .A(n8739), .B(n50268), .X(n24301) );
  nand_x2_sg U69999 ( .A(n8438), .B(n49454), .X(n31964) );
  nand_x2_sg U70000 ( .A(n8439), .B(n49409), .X(n31967) );
  nand_x2_sg U70001 ( .A(n8736), .B(n50407), .X(n24292) );
  nand_x2_sg U70002 ( .A(n8436), .B(n49548), .X(n31958) );
  nand_x2_sg U70003 ( .A(n8580), .B(n50206), .X(n22916) );
  nand_x2_sg U70004 ( .A(n8280), .B(n49347), .X(n30582) );
  nand_x2_sg U70005 ( .A(n8571), .B(n50625), .X(n22889) );
  nand_x2_sg U70006 ( .A(n8693), .B(n50542), .X(n24042) );
  nand_x2_sg U70007 ( .A(n8577), .B(n50342), .X(n22907) );
  nand_x2_sg U70008 ( .A(n8579), .B(n50250), .X(n22913) );
  nand_x2_sg U70009 ( .A(n8700), .B(n50218), .X(n24063) );
  nand_x2_sg U70010 ( .A(n8271), .B(n49766), .X(n30555) );
  nand_x2_sg U70011 ( .A(n8277), .B(n49483), .X(n30573) );
  nand_x2_sg U70012 ( .A(n8279), .B(n49391), .X(n30579) );
  nand_x2_sg U70013 ( .A(n8486), .B(n50851), .X(n22006) );
  nand_x2_sg U70014 ( .A(n8487), .B(n50806), .X(n22009) );
  nand_x2_sg U70015 ( .A(n8568), .B(n50767), .X(n22880) );
  nand_x2_sg U70016 ( .A(n8488), .B(n50758), .X(n22012) );
  nand_x2_sg U70017 ( .A(n8569), .B(n50720), .X(n22883) );
  nand_x2_sg U70018 ( .A(n8489), .B(n50711), .X(n22015) );
  nand_x2_sg U70019 ( .A(n8570), .B(n50672), .X(n22886) );
  nand_x2_sg U70020 ( .A(n8490), .B(n50663), .X(n22018) );
  nand_x2_sg U70021 ( .A(n8491), .B(n50616), .X(n22021) );
  nand_x2_sg U70022 ( .A(n8572), .B(n50576), .X(n22892) );
  nand_x2_sg U70023 ( .A(n8492), .B(n50567), .X(n22024) );
  nand_x2_sg U70024 ( .A(n8573), .B(n50529), .X(n22895) );
  nand_x2_sg U70025 ( .A(n8493), .B(n50520), .X(n22027) );
  nand_x2_sg U70026 ( .A(n8574), .B(n50482), .X(n22898) );
  nand_x2_sg U70027 ( .A(n8494), .B(n50473), .X(n22030) );
  nand_x2_sg U70028 ( .A(n8575), .B(n50436), .X(n22901) );
  nand_x2_sg U70029 ( .A(n8495), .B(n50427), .X(n22033) );
  nand_x2_sg U70030 ( .A(n8697), .B(n50354), .X(n24054) );
  nand_x2_sg U70031 ( .A(n8576), .B(n50389), .X(n22904) );
  nand_x2_sg U70032 ( .A(n8496), .B(n50380), .X(n22036) );
  nand_x2_sg U70033 ( .A(n8497), .B(n50333), .X(n22039) );
  nand_x2_sg U70034 ( .A(n8699), .B(n50263), .X(n24060) );
  nand_x2_sg U70035 ( .A(n8578), .B(n50296), .X(n22910) );
  nand_x2_sg U70036 ( .A(n8498), .B(n50287), .X(n22042) );
  nand_x2_sg U70037 ( .A(n8499), .B(n50241), .X(n22045) );
  nand_x2_sg U70038 ( .A(n8500), .B(n50197), .X(n22048) );
  nand_x2_sg U70039 ( .A(n8186), .B(n49992), .X(n29671) );
  nand_x2_sg U70040 ( .A(n8187), .B(n49947), .X(n29674) );
  nand_x2_sg U70041 ( .A(n8268), .B(n49908), .X(n30546) );
  nand_x2_sg U70042 ( .A(n8188), .B(n49899), .X(n29677) );
  nand_x2_sg U70043 ( .A(n8269), .B(n49861), .X(n30549) );
  nand_x2_sg U70044 ( .A(n8189), .B(n49852), .X(n29680) );
  nand_x2_sg U70045 ( .A(n8270), .B(n49813), .X(n30552) );
  nand_x2_sg U70046 ( .A(n8190), .B(n49804), .X(n29683) );
  nand_x2_sg U70047 ( .A(n8191), .B(n49757), .X(n29686) );
  nand_x2_sg U70048 ( .A(n8272), .B(n49717), .X(n30558) );
  nand_x2_sg U70049 ( .A(n8192), .B(n49708), .X(n29689) );
  nand_x2_sg U70050 ( .A(n8273), .B(n49670), .X(n30561) );
  nand_x2_sg U70051 ( .A(n8193), .B(n49661), .X(n29692) );
  nand_x2_sg U70052 ( .A(n8274), .B(n49623), .X(n30564) );
  nand_x2_sg U70053 ( .A(n8194), .B(n49614), .X(n29695) );
  nand_x2_sg U70054 ( .A(n8275), .B(n49577), .X(n30567) );
  nand_x2_sg U70055 ( .A(n8195), .B(n49568), .X(n29698) );
  nand_x2_sg U70056 ( .A(n8276), .B(n49530), .X(n30570) );
  nand_x2_sg U70057 ( .A(n8196), .B(n49521), .X(n29701) );
  nand_x2_sg U70058 ( .A(n8197), .B(n49474), .X(n29704) );
  nand_x2_sg U70059 ( .A(n8278), .B(n49437), .X(n30576) );
  nand_x2_sg U70060 ( .A(n8198), .B(n49428), .X(n29707) );
  nand_x2_sg U70061 ( .A(n8199), .B(n49382), .X(n29710) );
  nand_x2_sg U70062 ( .A(n8200), .B(n49338), .X(n29713) );
  nand_x2_sg U70063 ( .A(n8694), .B(n50494), .X(n24045) );
  nand_x2_sg U70064 ( .A(n8695), .B(n50448), .X(n24048) );
  nand_x2_sg U70065 ( .A(n8696), .B(n50402), .X(n24051) );
  nand_x2_sg U70066 ( .A(n8698), .B(n50308), .X(n24057) );
  nand_x2_sg U70067 ( .A(n8393), .B(n49683), .X(n31708) );
  nand_x2_sg U70068 ( .A(n8394), .B(n49635), .X(n31711) );
  nand_x2_sg U70069 ( .A(n8395), .B(n49589), .X(n31714) );
  nand_x2_sg U70070 ( .A(n8396), .B(n49543), .X(n31717) );
  nand_x2_sg U70071 ( .A(n8397), .B(n49495), .X(n31720) );
  nand_x2_sg U70072 ( .A(n8398), .B(n49449), .X(n31723) );
  nand_x2_sg U70073 ( .A(n8399), .B(n49404), .X(n31726) );
  nand_x2_sg U70074 ( .A(n8400), .B(n49359), .X(n31729) );
  nand_x2_sg U70075 ( .A(n8737), .B(n50359), .X(n24295) );
  nand_x2_sg U70076 ( .A(n8437), .B(n49500), .X(n31961) );
  nand_x2_sg U70077 ( .A(n8740), .B(n50223), .X(n24304) );
  nand_x2_sg U70078 ( .A(n8735), .B(n50453), .X(n24289) );
  nand_x2_sg U70079 ( .A(n8435), .B(n49594), .X(n31955) );
  nand_x2_sg U70080 ( .A(n8440), .B(n49364), .X(n31970) );
  nand_x2_sg U70081 ( .A(n8734), .B(n50499), .X(n24286) );
  nand_x2_sg U70082 ( .A(n8729), .B(n50689), .X(n23699) );
  nand_x2_sg U70083 ( .A(n8731), .B(n50598), .X(n24023) );
  nand_x2_sg U70084 ( .A(n8733), .B(n50546), .X(n24283) );
  nand_x2_sg U70085 ( .A(n8727), .B(n50781), .X(n23304) );
  nand_x2_sg U70086 ( .A(n8728), .B(n50735), .X(n23509) );
  nand_x2_sg U70087 ( .A(n8730), .B(n50644), .X(n23870) );
  nand_x2_sg U70088 ( .A(n8732), .B(n50552), .X(n24167) );
  nand_x2_sg U70089 ( .A(n8434), .B(n49640), .X(n31952) );
  nand_x2_sg U70090 ( .A(n8726), .B(n50825), .X(n23078) );
  nand_x2_sg U70091 ( .A(n8433), .B(n49687), .X(n31949) );
  nand_x2_sg U70092 ( .A(n8725), .B(n50869), .X(n22823) );
  nand_x2_sg U70093 ( .A(n8425), .B(n50010), .X(n30489) );
  nand_x2_sg U70094 ( .A(n8426), .B(n49966), .X(n30744) );
  nand_x2_sg U70095 ( .A(n8427), .B(n49922), .X(n30970) );
  nand_x2_sg U70096 ( .A(n8428), .B(n49876), .X(n31175) );
  nand_x2_sg U70097 ( .A(n8429), .B(n49830), .X(n31365) );
  nand_x2_sg U70098 ( .A(n8430), .B(n49785), .X(n31536) );
  nand_x2_sg U70099 ( .A(n8431), .B(n49739), .X(n31689) );
  nand_x2_sg U70100 ( .A(n8432), .B(n49693), .X(n31833) );
  nand_x2_sg U70101 ( .A(n8618), .B(n50301), .X(n23373) );
  nand_x2_sg U70102 ( .A(n8620), .B(n50211), .X(n23379) );
  nand_x2_sg U70103 ( .A(n8318), .B(n49442), .X(n31039) );
  nand_x2_sg U70104 ( .A(n8320), .B(n49352), .X(n31045) );
  nand_x2_sg U70105 ( .A(n8529), .B(n50716), .X(n22363) );
  nand_x2_sg U70106 ( .A(n8530), .B(n50668), .X(n22366) );
  nand_x2_sg U70107 ( .A(n8531), .B(n50621), .X(n22369) );
  nand_x2_sg U70108 ( .A(n8532), .B(n50572), .X(n22372) );
  nand_x2_sg U70109 ( .A(n8613), .B(n50534), .X(n23358) );
  nand_x2_sg U70110 ( .A(n8533), .B(n50525), .X(n22375) );
  nand_x2_sg U70111 ( .A(n8614), .B(n50487), .X(n23361) );
  nand_x2_sg U70112 ( .A(n8534), .B(n50478), .X(n22378) );
  nand_x2_sg U70113 ( .A(n8615), .B(n50441), .X(n23364) );
  nand_x2_sg U70114 ( .A(n8535), .B(n50432), .X(n22381) );
  nand_x2_sg U70115 ( .A(n8616), .B(n50394), .X(n23367) );
  nand_x2_sg U70116 ( .A(n8536), .B(n50385), .X(n22384) );
  nand_x2_sg U70117 ( .A(n8617), .B(n50347), .X(n23370) );
  nand_x2_sg U70118 ( .A(n8537), .B(n50338), .X(n22387) );
  nand_x2_sg U70119 ( .A(n8538), .B(n50292), .X(n22390) );
  nand_x2_sg U70120 ( .A(n8619), .B(n50255), .X(n23376) );
  nand_x2_sg U70121 ( .A(n8539), .B(n50246), .X(n22393) );
  nand_x2_sg U70122 ( .A(n8540), .B(n50202), .X(n22396) );
  nand_x2_sg U70123 ( .A(n8229), .B(n49857), .X(n30028) );
  nand_x2_sg U70124 ( .A(n8230), .B(n49809), .X(n30031) );
  nand_x2_sg U70125 ( .A(n8231), .B(n49762), .X(n30034) );
  nand_x2_sg U70126 ( .A(n8232), .B(n49713), .X(n30037) );
  nand_x2_sg U70127 ( .A(n8313), .B(n49675), .X(n31024) );
  nand_x2_sg U70128 ( .A(n8233), .B(n49666), .X(n30040) );
  nand_x2_sg U70129 ( .A(n8314), .B(n49628), .X(n31027) );
  nand_x2_sg U70130 ( .A(n8234), .B(n49619), .X(n30043) );
  nand_x2_sg U70131 ( .A(n8315), .B(n49582), .X(n31030) );
  nand_x2_sg U70132 ( .A(n8235), .B(n49573), .X(n30046) );
  nand_x2_sg U70133 ( .A(n8316), .B(n49535), .X(n31033) );
  nand_x2_sg U70134 ( .A(n8236), .B(n49526), .X(n30049) );
  nand_x2_sg U70135 ( .A(n8317), .B(n49488), .X(n31036) );
  nand_x2_sg U70136 ( .A(n8237), .B(n49479), .X(n30052) );
  nand_x2_sg U70137 ( .A(n8238), .B(n49433), .X(n30055) );
  nand_x2_sg U70138 ( .A(n8319), .B(n49396), .X(n31042) );
  nand_x2_sg U70139 ( .A(n8239), .B(n49387), .X(n30058) );
  nand_x2_sg U70140 ( .A(n8240), .B(n49343), .X(n30061) );
  nand_x2_sg U70141 ( .A(n8528), .B(n50763), .X(n22360) );
  nand_x2_sg U70142 ( .A(n8612), .B(n50581), .X(n23355) );
  nand_x2_sg U70143 ( .A(n8228), .B(n49904), .X(n30025) );
  nand_x2_sg U70144 ( .A(n8312), .B(n49722), .X(n31021) );
  nand_x2_sg U70145 ( .A(n8527), .B(n50811), .X(n22357) );
  nand_x2_sg U70146 ( .A(n8611), .B(n50630), .X(n23352) );
  nand_x2_sg U70147 ( .A(n8227), .B(n49952), .X(n30022) );
  nand_x2_sg U70148 ( .A(n8311), .B(n49771), .X(n31018) );
  nand_x2_sg U70149 ( .A(n8526), .B(n50855), .X(n22354) );
  nand_x2_sg U70150 ( .A(n8610), .B(n50677), .X(n23349) );
  nand_x2_sg U70151 ( .A(n8226), .B(n49996), .X(n30019) );
  nand_x2_sg U70152 ( .A(n8310), .B(n49818), .X(n31015) );
  nand_x2_sg U70153 ( .A(n8525), .B(n50895), .X(n22188) );
  nand_x2_sg U70154 ( .A(n8605), .B(n50888), .X(n22859) );
  nand_x2_sg U70155 ( .A(n8609), .B(n50725), .X(n23346) );
  nand_x2_sg U70156 ( .A(n8225), .B(n50036), .X(n29853) );
  nand_x2_sg U70157 ( .A(n8305), .B(n50029), .X(n30525) );
  nand_x2_sg U70158 ( .A(n8309), .B(n49866), .X(n31012) );
  nand_x2_sg U70159 ( .A(n8606), .B(n50843), .X(n23116) );
  nand_x2_sg U70160 ( .A(n8607), .B(n50819), .X(n23340) );
  nand_x2_sg U70161 ( .A(n8608), .B(n50771), .X(n23343) );
  nand_x2_sg U70162 ( .A(n8306), .B(n49984), .X(n30782) );
  nand_x2_sg U70163 ( .A(n8307), .B(n49960), .X(n31006) );
  nand_x2_sg U70164 ( .A(n8308), .B(n49912), .X(n31009) );
  nand_x2_sg U70165 ( .A(n8687), .B(n50788), .X(n23317) );
  nand_x2_sg U70166 ( .A(n8689), .B(n50696), .X(n23712) );
  nand_x2_sg U70167 ( .A(n8691), .B(n50638), .X(n24036) );
  nand_x2_sg U70168 ( .A(n8686), .B(n50832), .X(n23091) );
  nand_x2_sg U70169 ( .A(n8688), .B(n50742), .X(n23522) );
  nand_x2_sg U70170 ( .A(n8690), .B(n50651), .X(n23883) );
  nand_x2_sg U70171 ( .A(n8692), .B(n50588), .X(n24039) );
  nand_x2_sg U70172 ( .A(n8685), .B(n50876), .X(n22836) );
  nand_x2_sg U70173 ( .A(n8485), .B(n50900), .X(n22003) );
  nand_x2_sg U70174 ( .A(n8185), .B(n50041), .X(n29668) );
  nand_x2_sg U70175 ( .A(n8385), .B(n50017), .X(n30502) );
  nand_x2_sg U70176 ( .A(n8386), .B(n49973), .X(n30757) );
  nand_x2_sg U70177 ( .A(n8387), .B(n49929), .X(n30983) );
  nand_x2_sg U70178 ( .A(n8388), .B(n49883), .X(n31188) );
  nand_x2_sg U70179 ( .A(n8389), .B(n49837), .X(n31378) );
  nand_x2_sg U70180 ( .A(n8390), .B(n49792), .X(n31549) );
  nand_x2_sg U70181 ( .A(n8391), .B(n49779), .X(n31702) );
  nand_x2_sg U70182 ( .A(n8392), .B(n49729), .X(n31705) );
  nand_x2_sg U70183 ( .A(n25869), .B(n50989), .X(n25931) );
  nand_x1_sg U70184 ( .A(n51540), .B(n44905), .X(n25933) );
  nand_x2_sg U70185 ( .A(n26428), .B(n51027), .X(n26490) );
  nand_x1_sg U70186 ( .A(n52097), .B(n44853), .X(n26492) );
  nand_x2_sg U70187 ( .A(n27265), .B(n51085), .X(n27327) );
  nand_x1_sg U70188 ( .A(n52931), .B(n44851), .X(n27329) );
  nand_x2_sg U70189 ( .A(n27823), .B(n51123), .X(n27885) );
  nand_x1_sg U70190 ( .A(n53489), .B(n44849), .X(n27887) );
  nand_x2_sg U70191 ( .A(n25857), .B(n50991), .X(n25925) );
  nand_x1_sg U70192 ( .A(n44793), .B(n51557), .X(n25927) );
  nand_x2_sg U70193 ( .A(n26416), .B(n51029), .X(n26484) );
  nand_x1_sg U70194 ( .A(n44313), .B(n52114), .X(n26486) );
  nand_x2_sg U70195 ( .A(n27253), .B(n51087), .X(n27321) );
  nand_x1_sg U70196 ( .A(n44311), .B(n52948), .X(n27323) );
  nand_x2_sg U70197 ( .A(n27811), .B(n51125), .X(n27879) );
  nand_x1_sg U70198 ( .A(n44309), .B(n53506), .X(n27881) );
  nand_x2_sg U70199 ( .A(n28104), .B(n51142), .X(n28166) );
  nand_x1_sg U70200 ( .A(n53769), .B(n44881), .X(n28168) );
  nand_x2_sg U70201 ( .A(n28662), .B(n51179), .X(n28724) );
  nand_x1_sg U70202 ( .A(n54334), .B(n44879), .X(n28726) );
  nand_x2_sg U70203 ( .A(n29223), .B(n51217), .X(n29285) );
  nand_x1_sg U70204 ( .A(n54902), .B(n44883), .X(n29287) );
  nand_x2_sg U70205 ( .A(n28092), .B(n51144), .X(n28160) );
  nand_x1_sg U70206 ( .A(n44813), .B(n53785), .X(n28162) );
  nand_x2_sg U70207 ( .A(n28650), .B(n51181), .X(n28718) );
  nand_x1_sg U70208 ( .A(n44811), .B(n54350), .X(n28720) );
  nand_x2_sg U70209 ( .A(n29211), .B(n51219), .X(n29279) );
  nand_x1_sg U70210 ( .A(n44809), .B(n54918), .X(n29281) );
  nand_x2_sg U70211 ( .A(n28934), .B(n51199), .X(n28999) );
  nand_x1_sg U70212 ( .A(n46137), .B(n54625), .X(n29001) );
  nand_x2_sg U70213 ( .A(n29495), .B(n51237), .X(n29560) );
  nand_x1_sg U70214 ( .A(n46135), .B(n55193), .X(n29562) );
  nand_x2_sg U70215 ( .A(n26700), .B(n51048), .X(n26765) );
  nand_x1_sg U70216 ( .A(n52383), .B(n46129), .X(n26767) );
  nand_x2_sg U70217 ( .A(n25582), .B(n50971), .X(n25649) );
  nand_x1_sg U70218 ( .A(n46187), .B(n51271), .X(n25651) );
  nand_x2_sg U70219 ( .A(n27538), .B(n51105), .X(n27603) );
  nand_x1_sg U70220 ( .A(n46161), .B(n53219), .X(n27605) );
  nand_x2_sg U70221 ( .A(n26143), .B(n51009), .X(n26208) );
  nand_x1_sg U70222 ( .A(n46153), .B(n51831), .X(n26210) );
  nand_x2_sg U70223 ( .A(n28456), .B(n54042), .X(n28455) );
  nand_x1_sg U70224 ( .A(n28401), .B(n51158), .X(n28456) );
  nand_x2_sg U70225 ( .A(n26979), .B(n51067), .X(n27044) );
  nand_x1_sg U70226 ( .A(n52660), .B(n46141), .X(n27046) );
  nand_x2_sg U70227 ( .A(n28371), .B(n51162), .X(n28439) );
  nand_x1_sg U70228 ( .A(n54067), .B(n44833), .X(n28441) );
  nand_x2_sg U70229 ( .A(n25862), .B(n50990), .X(n25928) );
  nand_x2_sg U70230 ( .A(n26421), .B(n51028), .X(n26487) );
  nand_x2_sg U70231 ( .A(n27258), .B(n51086), .X(n27324) );
  nand_x2_sg U70232 ( .A(n27816), .B(n51124), .X(n27882) );
  nand_x2_sg U70233 ( .A(n28097), .B(n51143), .X(n28163) );
  nand_x2_sg U70234 ( .A(n28655), .B(n51180), .X(n28721) );
  nand_x2_sg U70235 ( .A(n29216), .B(n51218), .X(n29282) );
  nand_x2_sg U70236 ( .A(n8621), .B(n23383), .X(n23382) );
  nand_x1_sg U70237 ( .A(n23176), .B(n23172), .X(n23383) );
  nand_x2_sg U70238 ( .A(n8321), .B(n31049), .X(n31048) );
  nand_x1_sg U70239 ( .A(n30842), .B(n30838), .X(n31049) );
  nand_x2_sg U70240 ( .A(n8741), .B(n24308), .X(n24307) );
  nand_x1_sg U70241 ( .A(n24209), .B(n24205), .X(n24308) );
  nand_x2_sg U70242 ( .A(n8561), .B(n22669), .X(n22668) );
  nand_x2_sg U70243 ( .A(n10213), .B(n50122), .X(n22667) );
  nand_x1_sg U70244 ( .A(n22407), .B(n50151), .X(n22669) );
  nand_x2_sg U70245 ( .A(n8261), .B(n30335), .X(n30334) );
  nand_x2_sg U70246 ( .A(n25321), .B(n49263), .X(n30333) );
  nand_x1_sg U70247 ( .A(n30072), .B(n49292), .X(n30335) );
  nand_x2_sg U70248 ( .A(n8541), .B(n22400), .X(n22399) );
  nand_x1_sg U70249 ( .A(n22251), .B(n22247), .X(n22400) );
  nand_x2_sg U70250 ( .A(n8241), .B(n30065), .X(n30064) );
  nand_x1_sg U70251 ( .A(n29916), .B(n29912), .X(n30065) );
  nand_x2_sg U70252 ( .A(n8441), .B(n31974), .X(n31973) );
  nand_x1_sg U70253 ( .A(n31875), .B(n31871), .X(n31974) );
  nand_x2_sg U70254 ( .A(n8681), .B(n23923), .X(n23922) );
  nand_x2_sg U70255 ( .A(n10200), .B(n50115), .X(n23921) );
  nand_x1_sg U70256 ( .A(n23769), .B(n50145), .X(n23923) );
  nand_x2_sg U70257 ( .A(n8581), .B(n22920), .X(n22919) );
  nand_x1_sg U70258 ( .A(n22677), .B(n22673), .X(n22920) );
  nand_x2_sg U70259 ( .A(n8401), .B(n31733), .X(n31732) );
  nand_x1_sg U70260 ( .A(n31597), .B(n31593), .X(n31733) );
  nand_x2_sg U70261 ( .A(n8281), .B(n30586), .X(n30585) );
  nand_x1_sg U70262 ( .A(n30343), .B(n30339), .X(n30586) );
  nand_x2_sg U70263 ( .A(n8641), .B(n23581), .X(n23580) );
  nand_x2_sg U70264 ( .A(n10197), .B(n50118), .X(n23579) );
  nand_x1_sg U70265 ( .A(n23390), .B(n50147), .X(n23581) );
  nand_x2_sg U70266 ( .A(n8381), .B(n31589), .X(n31588) );
  nand_x2_sg U70267 ( .A(n25307), .B(n49256), .X(n31587) );
  nand_x1_sg U70268 ( .A(n31435), .B(n49286), .X(n31589) );
  nand_x2_sg U70269 ( .A(n8341), .B(n31247), .X(n31246) );
  nand_x2_sg U70270 ( .A(n25308), .B(n49259), .X(n31245) );
  nand_x1_sg U70271 ( .A(n31056), .B(n49288), .X(n31247) );
  nand_x2_sg U70272 ( .A(n8701), .B(n24067), .X(n24066) );
  nand_x1_sg U70273 ( .A(n23931), .B(n23927), .X(n24067) );
  nand_x2_sg U70274 ( .A(n8585), .B(n22866), .X(n22865) );
  nand_x2_sg U70275 ( .A(n50890), .B(n22867), .X(n22864) );
  nand_x1_sg U70276 ( .A(n50861), .B(n9443), .X(n22866) );
  nand_x2_sg U70277 ( .A(n8285), .B(n30532), .X(n30531) );
  nand_x2_sg U70278 ( .A(n50031), .B(n30533), .X(n30530) );
  nand_x1_sg U70279 ( .A(n50002), .B(n24551), .X(n30532) );
  nand_x2_sg U70280 ( .A(n8501), .B(n22052), .X(n22051) );
  nand_x2_sg U70281 ( .A(n50154), .B(n50125), .X(n22050) );
  nand_x1_sg U70282 ( .A(n10230), .B(n10226), .X(n22052) );
  nand_x2_sg U70283 ( .A(n8201), .B(n29717), .X(n29716) );
  nand_x2_sg U70284 ( .A(n49295), .B(n49266), .X(n29715) );
  nand_x1_sg U70285 ( .A(n25338), .B(n25334), .X(n29717) );
  nand_x2_sg U70286 ( .A(n24449), .B(n40791), .X(n24448) );
  nand_x2_sg U70287 ( .A(n8775), .B(n50364), .X(n24447) );
  nand_x1_sg U70288 ( .A(n24441), .B(n40797), .X(n24449) );
  nand_x2_sg U70289 ( .A(n32115), .B(n40792), .X(n32114) );
  nand_x2_sg U70290 ( .A(n8475), .B(n49505), .X(n32113) );
  nand_x1_sg U70291 ( .A(n32107), .B(n40798), .X(n32115) );
  nand_x2_sg U70292 ( .A(n23064), .B(n40727), .X(n23063) );
  nand_x2_sg U70293 ( .A(n8766), .B(n50776), .X(n23062) );
  nand_x1_sg U70294 ( .A(n23065), .B(n40743), .X(n23064) );
  nand_x2_sg U70295 ( .A(n23495), .B(n40728), .X(n23494) );
  nand_x2_sg U70296 ( .A(n8768), .B(n50684), .X(n23493) );
  nand_x1_sg U70297 ( .A(n23496), .B(n40744), .X(n23495) );
  nand_x2_sg U70298 ( .A(n23856), .B(n40729), .X(n23855) );
  nand_x2_sg U70299 ( .A(n8770), .B(n50593), .X(n23854) );
  nand_x1_sg U70300 ( .A(n23857), .B(n40745), .X(n23856) );
  nand_x2_sg U70301 ( .A(n24153), .B(n40730), .X(n24152) );
  nand_x2_sg U70302 ( .A(n8772), .B(n50502), .X(n24151) );
  nand_x1_sg U70303 ( .A(n24154), .B(n40746), .X(n24153) );
  nand_x2_sg U70304 ( .A(n30730), .B(n40733), .X(n30729) );
  nand_x2_sg U70305 ( .A(n8466), .B(n49917), .X(n30728) );
  nand_x1_sg U70306 ( .A(n30731), .B(n40749), .X(n30730) );
  nand_x2_sg U70307 ( .A(n31161), .B(n40734), .X(n31160) );
  nand_x2_sg U70308 ( .A(n8468), .B(n49825), .X(n31159) );
  nand_x1_sg U70309 ( .A(n31162), .B(n40750), .X(n31161) );
  nand_x2_sg U70310 ( .A(n31522), .B(n40735), .X(n31521) );
  nand_x2_sg U70311 ( .A(n8470), .B(n49734), .X(n31520) );
  nand_x1_sg U70312 ( .A(n31523), .B(n40751), .X(n31522) );
  nand_x2_sg U70313 ( .A(n31819), .B(n40731), .X(n31818) );
  nand_x2_sg U70314 ( .A(n8472), .B(n49643), .X(n31817) );
  nand_x1_sg U70315 ( .A(n31820), .B(n40747), .X(n31819) );
  nand_x2_sg U70316 ( .A(n8774), .B(n24372), .X(n24369) );
  nor_x1_sg U70317 ( .A(n24371), .B(out_L2[8]), .X(n24370) );
  nand_x2_sg U70318 ( .A(n8474), .B(n32038), .X(n32035) );
  nor_x1_sg U70319 ( .A(n32037), .B(out_L1[8]), .X(n32036) );
  nand_x2_sg U70320 ( .A(n8601), .B(n23168), .X(n23167) );
  nand_x2_sg U70321 ( .A(n22924), .B(n50120), .X(n23166) );
  nand_x1_sg U70322 ( .A(n22928), .B(n50149), .X(n23168) );
  nand_x2_sg U70323 ( .A(n8521), .B(n22243), .X(n22242) );
  nand_x2_sg U70324 ( .A(n22056), .B(n50124), .X(n22241) );
  nand_x1_sg U70325 ( .A(n22060), .B(n50153), .X(n22243) );
  nand_x2_sg U70326 ( .A(n8301), .B(n30834), .X(n30833) );
  nand_x2_sg U70327 ( .A(n30590), .B(n49261), .X(n30832) );
  nand_x1_sg U70328 ( .A(n30594), .B(n49290), .X(n30834) );
  nand_x2_sg U70329 ( .A(n8221), .B(n29908), .X(n29907) );
  nand_x2_sg U70330 ( .A(n29721), .B(n49265), .X(n29906) );
  nand_x1_sg U70331 ( .A(n29725), .B(n49294), .X(n29908) );
  nand_x2_sg U70332 ( .A(n8761), .B(n24400), .X(n24399) );
  nand_x2_sg U70333 ( .A(n24312), .B(n50110), .X(n24398) );
  nand_x1_sg U70334 ( .A(n24316), .B(n50141), .X(n24400) );
  nand_x2_sg U70335 ( .A(n8461), .B(n32066), .X(n32065) );
  nand_x2_sg U70336 ( .A(n31978), .B(n49251), .X(n32064) );
  nand_x1_sg U70337 ( .A(n31982), .B(n49282), .X(n32066) );
  nand_x2_sg U70338 ( .A(n8421), .B(n31867), .X(n31866) );
  nand_x2_sg U70339 ( .A(n31737), .B(n49254), .X(n31865) );
  nand_x1_sg U70340 ( .A(n31741), .B(n49284), .X(n31867) );
  nand_x2_sg U70341 ( .A(n8661), .B(n23762), .X(n23761) );
  nand_x1_sg U70342 ( .A(n23588), .B(n10220), .X(n23762) );
  nand_x2_sg U70343 ( .A(n8721), .B(n24201), .X(n24200) );
  nand_x2_sg U70344 ( .A(n24071), .B(n50113), .X(n24199) );
  nand_x1_sg U70345 ( .A(n24075), .B(n50143), .X(n24201) );
  nand_x2_sg U70346 ( .A(n8361), .B(n31428), .X(n31427) );
  nand_x1_sg U70347 ( .A(n31254), .B(n25328), .X(n31428) );
  nand_x2_sg U70348 ( .A(n8547), .B(n50813), .X(n22626) );
  nand_x2_sg U70349 ( .A(n9544), .B(n22491), .X(n22625) );
  nand_x2_sg U70350 ( .A(n8247), .B(n49954), .X(n30292) );
  nand_x2_sg U70351 ( .A(n24652), .B(n30156), .X(n30291) );
  nand_x2_sg U70352 ( .A(n8546), .B(n50857), .X(n22623) );
  nand_x2_sg U70353 ( .A(n9495), .B(n22497), .X(n22622) );
  nand_x2_sg U70354 ( .A(n8246), .B(n49998), .X(n30289) );
  nand_x2_sg U70355 ( .A(n24603), .B(n30162), .X(n30288) );
  nand_x2_sg U70356 ( .A(n8545), .B(n50905), .X(n22620) );
  nand_x2_sg U70357 ( .A(n9446), .B(n22350), .X(n22619) );
  nand_x2_sg U70358 ( .A(n8245), .B(n50046), .X(n30286) );
  nand_x2_sg U70359 ( .A(n24554), .B(n30015), .X(n30285) );
  nand_x2_sg U70360 ( .A(n8550), .B(n50670), .X(n22635) );
  nand_x2_sg U70361 ( .A(n9688), .B(n22473), .X(n22634) );
  nand_x2_sg U70362 ( .A(n8551), .B(n50623), .X(n22638) );
  nand_x2_sg U70363 ( .A(n9735), .B(n22467), .X(n22637) );
  nand_x2_sg U70364 ( .A(n8552), .B(n50574), .X(n22641) );
  nand_x2_sg U70365 ( .A(n9783), .B(n22461), .X(n22640) );
  nand_x2_sg U70366 ( .A(n8553), .B(n50527), .X(n22644) );
  nand_x2_sg U70367 ( .A(n9831), .B(n22455), .X(n22643) );
  nand_x2_sg U70368 ( .A(n8554), .B(n50480), .X(n22647) );
  nand_x2_sg U70369 ( .A(n9879), .B(n22449), .X(n22646) );
  nand_x2_sg U70370 ( .A(n8555), .B(n50434), .X(n22650) );
  nand_x2_sg U70371 ( .A(n9927), .B(n22443), .X(n22649) );
  nand_x2_sg U70372 ( .A(n8556), .B(n50387), .X(n22653) );
  nand_x2_sg U70373 ( .A(n9975), .B(n22437), .X(n22652) );
  nand_x2_sg U70374 ( .A(n8557), .B(n50340), .X(n22656) );
  nand_x2_sg U70375 ( .A(n10024), .B(n22431), .X(n22655) );
  nand_x2_sg U70376 ( .A(n8558), .B(n50294), .X(n22659) );
  nand_x2_sg U70377 ( .A(n10072), .B(n22425), .X(n22658) );
  nand_x2_sg U70378 ( .A(n8559), .B(n50248), .X(n22662) );
  nand_x2_sg U70379 ( .A(n10121), .B(n22419), .X(n22661) );
  nand_x2_sg U70380 ( .A(n8560), .B(n50204), .X(n22665) );
  nand_x2_sg U70381 ( .A(n10170), .B(n22413), .X(n22664) );
  nand_x2_sg U70382 ( .A(n8250), .B(n49811), .X(n30301) );
  nand_x2_sg U70383 ( .A(n24796), .B(n30138), .X(n30300) );
  nand_x2_sg U70384 ( .A(n8251), .B(n49764), .X(n30304) );
  nand_x2_sg U70385 ( .A(n24843), .B(n30132), .X(n30303) );
  nand_x2_sg U70386 ( .A(n8252), .B(n49715), .X(n30307) );
  nand_x2_sg U70387 ( .A(n24891), .B(n30126), .X(n30306) );
  nand_x2_sg U70388 ( .A(n8253), .B(n49668), .X(n30310) );
  nand_x2_sg U70389 ( .A(n24939), .B(n30120), .X(n30309) );
  nand_x2_sg U70390 ( .A(n8254), .B(n49621), .X(n30313) );
  nand_x2_sg U70391 ( .A(n24987), .B(n30114), .X(n30312) );
  nand_x2_sg U70392 ( .A(n8255), .B(n49575), .X(n30316) );
  nand_x2_sg U70393 ( .A(n25035), .B(n30108), .X(n30315) );
  nand_x2_sg U70394 ( .A(n8256), .B(n49528), .X(n30319) );
  nand_x2_sg U70395 ( .A(n25083), .B(n30102), .X(n30318) );
  nand_x2_sg U70396 ( .A(n8257), .B(n49481), .X(n30322) );
  nand_x2_sg U70397 ( .A(n25132), .B(n30096), .X(n30321) );
  nand_x2_sg U70398 ( .A(n8258), .B(n49435), .X(n30325) );
  nand_x2_sg U70399 ( .A(n25180), .B(n30090), .X(n30324) );
  nand_x2_sg U70400 ( .A(n8259), .B(n49389), .X(n30328) );
  nand_x2_sg U70401 ( .A(n25229), .B(n30084), .X(n30327) );
  nand_x2_sg U70402 ( .A(n8260), .B(n49345), .X(n30331) );
  nand_x2_sg U70403 ( .A(n25278), .B(n30078), .X(n30330) );
  nand_x2_sg U70404 ( .A(n8549), .B(n50718), .X(n22632) );
  nand_x2_sg U70405 ( .A(n9640), .B(n22479), .X(n22631) );
  nand_x2_sg U70406 ( .A(n8249), .B(n49859), .X(n30298) );
  nand_x2_sg U70407 ( .A(n24748), .B(n30144), .X(n30297) );
  nand_x2_sg U70408 ( .A(n8548), .B(n50765), .X(n22629) );
  nand_x2_sg U70409 ( .A(n9592), .B(n22485), .X(n22628) );
  nand_x2_sg U70410 ( .A(n8248), .B(n49906), .X(n30295) );
  nand_x2_sg U70411 ( .A(n24700), .B(n30150), .X(n30294) );
  nand_x2_sg U70412 ( .A(n8675), .B(n50446), .X(n23904) );
  nand_x2_sg U70413 ( .A(n9911), .B(n23805), .X(n23903) );
  nand_x2_sg U70414 ( .A(n8676), .B(n50400), .X(n23907) );
  nand_x2_sg U70415 ( .A(n9959), .B(n23799), .X(n23906) );
  nand_x2_sg U70416 ( .A(n8373), .B(n49681), .X(n31564) );
  nand_x2_sg U70417 ( .A(n24923), .B(n31483), .X(n31563) );
  nand_x2_sg U70418 ( .A(n8374), .B(n49633), .X(n31567) );
  nand_x2_sg U70419 ( .A(n24971), .B(n31477), .X(n31566) );
  nand_x2_sg U70420 ( .A(n8375), .B(n49587), .X(n31570) );
  nand_x2_sg U70421 ( .A(n25019), .B(n31471), .X(n31569) );
  nand_x2_sg U70422 ( .A(n8376), .B(n49541), .X(n31573) );
  nand_x2_sg U70423 ( .A(n25067), .B(n31465), .X(n31572) );
  nand_x2_sg U70424 ( .A(n8377), .B(n49493), .X(n31576) );
  nand_x2_sg U70425 ( .A(n25116), .B(n31459), .X(n31575) );
  nand_x2_sg U70426 ( .A(n8378), .B(n49447), .X(n31579) );
  nand_x2_sg U70427 ( .A(n25164), .B(n31453), .X(n31578) );
  nand_x2_sg U70428 ( .A(n8379), .B(n49402), .X(n31582) );
  nand_x2_sg U70429 ( .A(n25213), .B(n31447), .X(n31581) );
  nand_x2_sg U70430 ( .A(n8380), .B(n49357), .X(n31585) );
  nand_x2_sg U70431 ( .A(n25262), .B(n31441), .X(n31584) );
  nand_x2_sg U70432 ( .A(n8674), .B(n50492), .X(n23901) );
  nand_x2_sg U70433 ( .A(n9863), .B(n23811), .X(n23900) );
  nand_x2_sg U70434 ( .A(n8678), .B(n50306), .X(n23913) );
  nand_x2_sg U70435 ( .A(n10056), .B(n23787), .X(n23912) );
  nand_x2_sg U70436 ( .A(n8673), .B(n50540), .X(n23898) );
  nand_x2_sg U70437 ( .A(n9815), .B(n23817), .X(n23897) );
  nand_x2_sg U70438 ( .A(n8677), .B(n50352), .X(n23910) );
  nand_x2_sg U70439 ( .A(n10008), .B(n23793), .X(n23909) );
  nand_x2_sg U70440 ( .A(n8679), .B(n50261), .X(n23916) );
  nand_x2_sg U70441 ( .A(n10105), .B(n23781), .X(n23915) );
  nand_x2_sg U70442 ( .A(n8680), .B(n50216), .X(n23919) );
  nand_x2_sg U70443 ( .A(n10154), .B(n23775), .X(n23918) );
  nand_x2_sg U70444 ( .A(n8665), .B(n50879), .X(n22842) );
  nand_x2_sg U70445 ( .A(n9429), .B(n22844), .X(n22841) );
  nand_x2_sg U70446 ( .A(n8365), .B(n50020), .X(n30508) );
  nand_x2_sg U70447 ( .A(n24537), .B(n30510), .X(n30507) );
  nand_x2_sg U70448 ( .A(n8367), .B(n49932), .X(n30989) );
  nand_x2_sg U70449 ( .A(n24635), .B(n30991), .X(n30988) );
  nand_x2_sg U70450 ( .A(n8369), .B(n49840), .X(n31384) );
  nand_x2_sg U70451 ( .A(n24732), .B(n31386), .X(n31383) );
  nand_x2_sg U70452 ( .A(n8371), .B(n49777), .X(n31558) );
  nand_x2_sg U70453 ( .A(n24827), .B(n31495), .X(n31557) );
  nand_x2_sg U70454 ( .A(n8366), .B(n49976), .X(n30763) );
  nand_x2_sg U70455 ( .A(n24586), .B(n30765), .X(n30762) );
  nand_x2_sg U70456 ( .A(n8368), .B(n49886), .X(n31194) );
  nand_x2_sg U70457 ( .A(n24684), .B(n31196), .X(n31193) );
  nand_x2_sg U70458 ( .A(n8370), .B(n49823), .X(n31555) );
  nand_x2_sg U70459 ( .A(n24780), .B(n31501), .X(n31554) );
  nand_x2_sg U70460 ( .A(n8372), .B(n49727), .X(n31561) );
  nand_x2_sg U70461 ( .A(n24875), .B(n31489), .X(n31560) );
  nand_x2_sg U70462 ( .A(n8667), .B(n50791), .X(n23323) );
  nand_x2_sg U70463 ( .A(n9527), .B(n23325), .X(n23322) );
  nand_x2_sg U70464 ( .A(n8669), .B(n50699), .X(n23718) );
  nand_x2_sg U70465 ( .A(n9624), .B(n23720), .X(n23717) );
  nand_x2_sg U70466 ( .A(n8671), .B(n50636), .X(n23892) );
  nand_x2_sg U70467 ( .A(n9719), .B(n23829), .X(n23891) );
  nand_x2_sg U70468 ( .A(n8666), .B(n50835), .X(n23097) );
  nand_x2_sg U70469 ( .A(n9478), .B(n23099), .X(n23096) );
  nand_x2_sg U70470 ( .A(n8668), .B(n50745), .X(n23528) );
  nand_x2_sg U70471 ( .A(n9576), .B(n23530), .X(n23527) );
  nand_x2_sg U70472 ( .A(n8670), .B(n50682), .X(n23889) );
  nand_x2_sg U70473 ( .A(n9672), .B(n23835), .X(n23888) );
  nand_x2_sg U70474 ( .A(n8672), .B(n50586), .X(n23895) );
  nand_x2_sg U70475 ( .A(n9767), .B(n23823), .X(n23894) );
  nand_x4_sg U70476 ( .A(n28396), .B(n54048), .X(n28393) );
  nand_x1_sg U70477 ( .A(n46191), .B(n54047), .X(n28396) );
  nor_x1_sg U70478 ( .A(n54047), .B(n46191), .X(n28397) );
  nand_x2_sg U70479 ( .A(n8630), .B(n50679), .X(n23547) );
  nand_x2_sg U70480 ( .A(n9668), .B(n23456), .X(n23546) );
  nand_x2_sg U70481 ( .A(n8330), .B(n49820), .X(n31213) );
  nand_x2_sg U70482 ( .A(n24781), .B(n31122), .X(n31212) );
  nand_x2_sg U70483 ( .A(n8640), .B(n50213), .X(n23577) );
  nand_x2_sg U70484 ( .A(n10150), .B(n23396), .X(n23576) );
  nand_x2_sg U70485 ( .A(n8340), .B(n49354), .X(n31243) );
  nand_x2_sg U70486 ( .A(n25263), .B(n31062), .X(n31242) );
  nand_x2_sg U70487 ( .A(n8626), .B(n50840), .X(n23110) );
  nand_x2_sg U70488 ( .A(n9474), .B(n23112), .X(n23109) );
  nand_x2_sg U70489 ( .A(n8628), .B(n50773), .X(n23541) );
  nand_x2_sg U70490 ( .A(n9572), .B(n23468), .X(n23540) );
  nand_x2_sg U70491 ( .A(n8326), .B(n49981), .X(n30776) );
  nand_x2_sg U70492 ( .A(n24587), .B(n30778), .X(n30775) );
  nand_x2_sg U70493 ( .A(n8328), .B(n49914), .X(n31207) );
  nand_x2_sg U70494 ( .A(n24685), .B(n31134), .X(n31206) );
  nand_x2_sg U70495 ( .A(n8625), .B(n50885), .X(n22853) );
  nand_x2_sg U70496 ( .A(n9425), .B(n22855), .X(n22852) );
  nand_x2_sg U70497 ( .A(n8627), .B(n50797), .X(n23334) );
  nand_x2_sg U70498 ( .A(n9523), .B(n23336), .X(n23333) );
  nand_x2_sg U70499 ( .A(n8629), .B(n50727), .X(n23544) );
  nand_x2_sg U70500 ( .A(n9620), .B(n23462), .X(n23543) );
  nand_x2_sg U70501 ( .A(n8631), .B(n50632), .X(n23550) );
  nand_x2_sg U70502 ( .A(n9715), .B(n23450), .X(n23549) );
  nand_x2_sg U70503 ( .A(n8632), .B(n50583), .X(n23553) );
  nand_x2_sg U70504 ( .A(n9763), .B(n23444), .X(n23552) );
  nand_x2_sg U70505 ( .A(n8633), .B(n50536), .X(n23556) );
  nand_x2_sg U70506 ( .A(n9811), .B(n23438), .X(n23555) );
  nand_x2_sg U70507 ( .A(n8634), .B(n50489), .X(n23559) );
  nand_x2_sg U70508 ( .A(n9859), .B(n23432), .X(n23558) );
  nand_x2_sg U70509 ( .A(n8635), .B(n50443), .X(n23562) );
  nand_x2_sg U70510 ( .A(n9907), .B(n23426), .X(n23561) );
  nand_x2_sg U70511 ( .A(n8636), .B(n50396), .X(n23565) );
  nand_x2_sg U70512 ( .A(n9955), .B(n23420), .X(n23564) );
  nand_x2_sg U70513 ( .A(n8637), .B(n50349), .X(n23568) );
  nand_x2_sg U70514 ( .A(n10004), .B(n23414), .X(n23567) );
  nand_x2_sg U70515 ( .A(n8638), .B(n50303), .X(n23571) );
  nand_x2_sg U70516 ( .A(n10052), .B(n23408), .X(n23570) );
  nand_x2_sg U70517 ( .A(n8639), .B(n50257), .X(n23574) );
  nand_x2_sg U70518 ( .A(n10101), .B(n23402), .X(n23573) );
  nand_x2_sg U70519 ( .A(n8325), .B(n50026), .X(n30519) );
  nand_x2_sg U70520 ( .A(n24538), .B(n30521), .X(n30518) );
  nand_x2_sg U70521 ( .A(n8327), .B(n49938), .X(n31000) );
  nand_x2_sg U70522 ( .A(n24636), .B(n31002), .X(n30999) );
  nand_x2_sg U70523 ( .A(n8329), .B(n49868), .X(n31210) );
  nand_x2_sg U70524 ( .A(n24733), .B(n31128), .X(n31209) );
  nand_x2_sg U70525 ( .A(n8331), .B(n49773), .X(n31216) );
  nand_x2_sg U70526 ( .A(n24828), .B(n31116), .X(n31215) );
  nand_x2_sg U70527 ( .A(n8332), .B(n49724), .X(n31219) );
  nand_x2_sg U70528 ( .A(n24876), .B(n31110), .X(n31218) );
  nand_x2_sg U70529 ( .A(n8333), .B(n49677), .X(n31222) );
  nand_x2_sg U70530 ( .A(n24924), .B(n31104), .X(n31221) );
  nand_x2_sg U70531 ( .A(n8334), .B(n49630), .X(n31225) );
  nand_x2_sg U70532 ( .A(n24972), .B(n31098), .X(n31224) );
  nand_x2_sg U70533 ( .A(n8335), .B(n49584), .X(n31228) );
  nand_x2_sg U70534 ( .A(n25020), .B(n31092), .X(n31227) );
  nand_x2_sg U70535 ( .A(n8336), .B(n49537), .X(n31231) );
  nand_x2_sg U70536 ( .A(n25068), .B(n31086), .X(n31230) );
  nand_x2_sg U70537 ( .A(n8337), .B(n49490), .X(n31234) );
  nand_x2_sg U70538 ( .A(n25117), .B(n31080), .X(n31233) );
  nand_x2_sg U70539 ( .A(n8338), .B(n49444), .X(n31237) );
  nand_x2_sg U70540 ( .A(n25165), .B(n31074), .X(n31236) );
  nand_x2_sg U70541 ( .A(n8339), .B(n49398), .X(n31240) );
  nand_x2_sg U70542 ( .A(n25214), .B(n31068), .X(n31239) );
  nand_x2_sg U70543 ( .A(n8707), .B(n50785), .X(n23310) );
  nand_x2_sg U70544 ( .A(n23313), .B(n23312), .X(n23309) );
  nand_x2_sg U70545 ( .A(n8709), .B(n50693), .X(n23705) );
  nand_x2_sg U70546 ( .A(n23708), .B(n23707), .X(n23704) );
  nand_x2_sg U70547 ( .A(n8711), .B(n50602), .X(n24029) );
  nand_x2_sg U70548 ( .A(n24032), .B(n24031), .X(n24028) );
  nand_x2_sg U70549 ( .A(n8706), .B(n50829), .X(n23084) );
  nand_x2_sg U70550 ( .A(n23087), .B(n23086), .X(n23083) );
  nand_x2_sg U70551 ( .A(n8708), .B(n50739), .X(n23515) );
  nand_x2_sg U70552 ( .A(n23518), .B(n23517), .X(n23514) );
  nand_x2_sg U70553 ( .A(n8710), .B(n50648), .X(n23876) );
  nand_x2_sg U70554 ( .A(n23879), .B(n23878), .X(n23875) );
  nand_x2_sg U70555 ( .A(n8712), .B(n50590), .X(n24173) );
  nand_x2_sg U70556 ( .A(n24135), .B(n24138), .X(n24172) );
  nand_x2_sg U70557 ( .A(n8705), .B(n50873), .X(n22829) );
  nand_x2_sg U70558 ( .A(n22832), .B(n22831), .X(n22828) );
  nand_x2_sg U70559 ( .A(n8505), .B(n50902), .X(n22194) );
  nand_x2_sg U70560 ( .A(n22169), .B(n22172), .X(n22193) );
  nand_x2_sg U70561 ( .A(n8205), .B(n50043), .X(n29859) );
  nand_x2_sg U70562 ( .A(n29834), .B(n29837), .X(n29858) );
  nand_x2_sg U70563 ( .A(n8405), .B(n50014), .X(n30495) );
  nand_x2_sg U70564 ( .A(n30498), .B(n30497), .X(n30494) );
  nand_x2_sg U70565 ( .A(n8406), .B(n49970), .X(n30750) );
  nand_x2_sg U70566 ( .A(n30753), .B(n30752), .X(n30749) );
  nand_x2_sg U70567 ( .A(n8407), .B(n49926), .X(n30976) );
  nand_x2_sg U70568 ( .A(n30979), .B(n30978), .X(n30975) );
  nand_x2_sg U70569 ( .A(n8408), .B(n49880), .X(n31181) );
  nand_x2_sg U70570 ( .A(n31184), .B(n31183), .X(n31180) );
  nand_x2_sg U70571 ( .A(n8409), .B(n49834), .X(n31371) );
  nand_x2_sg U70572 ( .A(n31374), .B(n31373), .X(n31370) );
  nand_x2_sg U70573 ( .A(n8410), .B(n49789), .X(n31542) );
  nand_x2_sg U70574 ( .A(n31545), .B(n31544), .X(n31541) );
  nand_x2_sg U70575 ( .A(n8411), .B(n49743), .X(n31695) );
  nand_x2_sg U70576 ( .A(n31698), .B(n31697), .X(n31694) );
  nand_x2_sg U70577 ( .A(n8412), .B(n49731), .X(n31839) );
  nand_x2_sg U70578 ( .A(n31801), .B(n31804), .X(n31838) );
  nand_x2_sg U70579 ( .A(n8713), .B(n24177), .X(n24176) );
  nand_x2_sg U70580 ( .A(n24128), .B(n24131), .X(n24175) );
  nand_x1_sg U70581 ( .A(n50496), .B(n50508), .X(n24177) );
  nand_x2_sg U70582 ( .A(n8506), .B(n22198), .X(n22197) );
  nand_x2_sg U70583 ( .A(n22162), .B(n22165), .X(n22196) );
  nand_x1_sg U70584 ( .A(n50808), .B(n50849), .X(n22198) );
  nand_x2_sg U70585 ( .A(n8206), .B(n29863), .X(n29862) );
  nand_x2_sg U70586 ( .A(n29827), .B(n29830), .X(n29861) );
  nand_x1_sg U70587 ( .A(n49949), .B(n49990), .X(n29863) );
  nand_x2_sg U70588 ( .A(n8413), .B(n31843), .X(n31842) );
  nand_x2_sg U70589 ( .A(n31794), .B(n31797), .X(n31841) );
  nand_x1_sg U70590 ( .A(n49637), .B(n49649), .X(n31843) );
  nand_x2_sg U70591 ( .A(n8745), .B(n22817), .X(n22816) );
  nand_x2_sg U70592 ( .A(n22818), .B(n22819), .X(n22815) );
  nand_x1_sg U70593 ( .A(n50824), .B(n50866), .X(n22817) );
  nand_x2_sg U70594 ( .A(n8445), .B(n30483), .X(n30482) );
  nand_x2_sg U70595 ( .A(n30484), .B(n30485), .X(n30481) );
  nand_x1_sg U70596 ( .A(n49965), .B(n50007), .X(n30483) );
  nand_x2_sg U70597 ( .A(n8586), .B(n23123), .X(n23122) );
  nand_x2_sg U70598 ( .A(n50845), .B(n23031), .X(n23121) );
  nand_x1_sg U70599 ( .A(n50817), .B(n9492), .X(n23123) );
  nand_x2_sg U70600 ( .A(n8587), .B(n23126), .X(n23125) );
  nand_x2_sg U70601 ( .A(n50800), .B(n23025), .X(n23124) );
  nand_x1_sg U70602 ( .A(n50769), .B(n9541), .X(n23126) );
  nand_x2_sg U70603 ( .A(n8286), .B(n30789), .X(n30788) );
  nand_x2_sg U70604 ( .A(n49986), .B(n30697), .X(n30787) );
  nand_x1_sg U70605 ( .A(n49958), .B(n24600), .X(n30789) );
  nand_x2_sg U70606 ( .A(n8287), .B(n30792), .X(n30791) );
  nand_x2_sg U70607 ( .A(n49941), .B(n30691), .X(n30790) );
  nand_x1_sg U70608 ( .A(n49910), .B(n24649), .X(n30792) );
  nand_x2_sg U70609 ( .A(n8759), .B(n24394), .X(n24393) );
  nand_x2_sg U70610 ( .A(n40648), .B(n24329), .X(n24392) );
  nand_x1_sg U70611 ( .A(n50225), .B(n10127), .X(n24394) );
  nand_x2_sg U70612 ( .A(n8459), .B(n32060), .X(n32059) );
  nand_x2_sg U70613 ( .A(n40698), .B(n31995), .X(n32058) );
  nand_x1_sg U70614 ( .A(n49366), .B(n25235), .X(n32060) );
  nand_x2_sg U70615 ( .A(n8758), .B(n24391), .X(n24390) );
  nand_x2_sg U70616 ( .A(n50273), .B(n24335), .X(n24389) );
  nand_x1_sg U70617 ( .A(n50270), .B(n10078), .X(n24391) );
  nand_x2_sg U70618 ( .A(n8458), .B(n32057), .X(n32056) );
  nand_x2_sg U70619 ( .A(n49414), .B(n32001), .X(n32055) );
  nand_x1_sg U70620 ( .A(n49411), .B(n25186), .X(n32057) );
  nand_x2_sg U70621 ( .A(n8756), .B(n24385), .X(n24384) );
  nand_x2_sg U70622 ( .A(n50366), .B(n24348), .X(n24383) );
  nand_x1_sg U70623 ( .A(n50361), .B(n9981), .X(n24385) );
  nand_x2_sg U70624 ( .A(n8456), .B(n32051), .X(n32050) );
  nand_x2_sg U70625 ( .A(n49507), .B(n32014), .X(n32049) );
  nand_x1_sg U70626 ( .A(n49502), .B(n25089), .X(n32051) );
  nand_x1_sg U70627 ( .A(n45235), .B(n26203), .X(n26202) );
  nor_x1_sg U70628 ( .A(n26130), .B(n46127), .X(n26204) );
  nand_x1_sg U70629 ( .A(n45227), .B(n26760), .X(n26759) );
  nor_x1_sg U70630 ( .A(n26687), .B(n46119), .X(n26761) );
  nand_x1_sg U70631 ( .A(n45233), .B(n27598), .X(n27597) );
  nor_x1_sg U70632 ( .A(n27525), .B(n46125), .X(n27599) );
  nand_x1_sg U70633 ( .A(n45237), .B(n25644), .X(n25643) );
  nor_x1_sg U70634 ( .A(n25569), .B(n46131), .X(n25645) );
  nand_x4_sg U70635 ( .A(n26771), .B(n26772), .X(n26706) );
  nand_x1_sg U70636 ( .A(n26712), .B(n51046), .X(n26771) );
  nand_x1_sg U70637 ( .A(n46071), .B(n26773), .X(n26772) );
  nand_x1_sg U70638 ( .A(n52370), .B(n44877), .X(n26773) );
  nand_x1_sg U70639 ( .A(n45231), .B(n28994), .X(n28993) );
  nor_x1_sg U70640 ( .A(n28921), .B(n46123), .X(n28995) );
  nand_x1_sg U70641 ( .A(n45229), .B(n29555), .X(n29554) );
  nor_x1_sg U70642 ( .A(n29482), .B(n46121), .X(n29556) );
  nand_x1_sg U70643 ( .A(n46063), .B(n25936), .X(n25935) );
  nand_x1_sg U70644 ( .A(n51535), .B(n44897), .X(n25936) );
  nand_x1_sg U70645 ( .A(n46055), .B(n26495), .X(n26494) );
  nand_x1_sg U70646 ( .A(n52093), .B(n44873), .X(n26495) );
  nand_x1_sg U70647 ( .A(n46053), .B(n27332), .X(n27331) );
  nand_x1_sg U70648 ( .A(n52927), .B(n44871), .X(n27332) );
  nand_x1_sg U70649 ( .A(n46051), .B(n27890), .X(n27889) );
  nand_x1_sg U70650 ( .A(n53485), .B(n44869), .X(n27890) );
  nand_x4_sg U70651 ( .A(n29005), .B(n29006), .X(n28940) );
  nand_x1_sg U70652 ( .A(n28946), .B(n51197), .X(n29005) );
  nand_x1_sg U70653 ( .A(n46079), .B(n29007), .X(n29006) );
  nand_x1_sg U70654 ( .A(n44895), .B(n54612), .X(n29007) );
  nand_x4_sg U70655 ( .A(n29566), .B(n29567), .X(n29501) );
  nand_x1_sg U70656 ( .A(n29507), .B(n51235), .X(n29566) );
  nand_x1_sg U70657 ( .A(n46081), .B(n29568), .X(n29567) );
  nand_x1_sg U70658 ( .A(n44899), .B(n55180), .X(n29568) );
  nand_x4_sg U70659 ( .A(n25655), .B(n25656), .X(n25588) );
  nand_x1_sg U70660 ( .A(n25594), .B(n50969), .X(n25655) );
  nand_x1_sg U70661 ( .A(n46085), .B(n25657), .X(n25656) );
  nand_x1_sg U70662 ( .A(n44903), .B(n51259), .X(n25657) );
  nand_x4_sg U70663 ( .A(n27609), .B(n27610), .X(n27544) );
  nand_x1_sg U70664 ( .A(n27550), .B(n51103), .X(n27609) );
  nand_x1_sg U70665 ( .A(n46075), .B(n27611), .X(n27610) );
  nand_x1_sg U70666 ( .A(n44887), .B(n53205), .X(n27611) );
  nand_x4_sg U70667 ( .A(n26214), .B(n26215), .X(n26149) );
  nand_x1_sg U70668 ( .A(n26155), .B(n51007), .X(n26214) );
  nand_x1_sg U70669 ( .A(n46073), .B(n26216), .X(n26215) );
  nand_x1_sg U70670 ( .A(n44885), .B(n51817), .X(n26216) );
  nand_x1_sg U70671 ( .A(n46067), .B(n28171), .X(n28170) );
  nand_x1_sg U70672 ( .A(n53763), .B(n44891), .X(n28171) );
  nand_x1_sg U70673 ( .A(n46065), .B(n28729), .X(n28728) );
  nand_x1_sg U70674 ( .A(n54328), .B(n44889), .X(n28729) );
  nand_x1_sg U70675 ( .A(n46069), .B(n29290), .X(n29289) );
  nand_x1_sg U70676 ( .A(n54896), .B(n44893), .X(n29290) );
  nand_x4_sg U70677 ( .A(n27050), .B(n27051), .X(n26985) );
  nand_x1_sg U70678 ( .A(n26991), .B(n51065), .X(n27050) );
  nand_x1_sg U70679 ( .A(n46083), .B(n27052), .X(n27051) );
  nand_x1_sg U70680 ( .A(n52646), .B(n44901), .X(n27052) );
  nand_x1_sg U70681 ( .A(n46033), .B(n27040), .X(n27039) );
  nand_x1_sg U70682 ( .A(n45971), .B(n52639), .X(n27000) );
  nand_x1_sg U70683 ( .A(n45957), .B(n53756), .X(n28119) );
  nand_x1_sg U70684 ( .A(n45955), .B(n54321), .X(n28677) );
  nand_x1_sg U70685 ( .A(n45953), .B(n54889), .X(n29238) );
  nand_x1_sg U70686 ( .A(n45975), .B(n51252), .X(n25603) );
  nand_x1_sg U70687 ( .A(n45949), .B(n54040), .X(n28398) );
  nand_x4_sg U70688 ( .A(n25940), .B(n25941), .X(n25880) );
  nand_x1_sg U70689 ( .A(n46019), .B(n51529), .X(n25940) );
  nand_x1_sg U70690 ( .A(n25887), .B(n50986), .X(n25942) );
  nand_x4_sg U70691 ( .A(n27615), .B(n27616), .X(n27555) );
  nand_x1_sg U70692 ( .A(n46013), .B(n53199), .X(n27615) );
  nand_x1_sg U70693 ( .A(n27562), .B(n51101), .X(n27617) );
  nand_x4_sg U70694 ( .A(n25661), .B(n25662), .X(n25599) );
  nand_x1_sg U70695 ( .A(n46027), .B(n51253), .X(n25661) );
  nand_x1_sg U70696 ( .A(n25606), .B(n50967), .X(n25663) );
  nand_x4_sg U70697 ( .A(n26777), .B(n26778), .X(n26717) );
  nand_x1_sg U70698 ( .A(n46015), .B(n26725), .X(n26777) );
  nand_x1_sg U70699 ( .A(n52364), .B(n51044), .X(n26779) );
  nand_x4_sg U70700 ( .A(n29011), .B(n29012), .X(n28951) );
  nand_x1_sg U70701 ( .A(n46021), .B(n54606), .X(n29011) );
  nand_x1_sg U70702 ( .A(n28958), .B(n51195), .X(n29013) );
  nand_x4_sg U70703 ( .A(n29572), .B(n29573), .X(n29512) );
  nand_x1_sg U70704 ( .A(n46025), .B(n55174), .X(n29572) );
  nand_x1_sg U70705 ( .A(n29519), .B(n51233), .X(n29574) );
  nand_x4_sg U70706 ( .A(n28175), .B(n28176), .X(n28115) );
  nand_x1_sg U70707 ( .A(n46005), .B(n53757), .X(n28175) );
  nand_x1_sg U70708 ( .A(n28122), .B(n51139), .X(n28177) );
  nand_x4_sg U70709 ( .A(n28733), .B(n28734), .X(n28673) );
  nand_x1_sg U70710 ( .A(n46003), .B(n54322), .X(n28733) );
  nand_x1_sg U70711 ( .A(n28680), .B(n51176), .X(n28735) );
  nand_x4_sg U70712 ( .A(n29294), .B(n29295), .X(n29234) );
  nand_x1_sg U70713 ( .A(n46001), .B(n54890), .X(n29294) );
  nand_x1_sg U70714 ( .A(n29241), .B(n51214), .X(n29296) );
  nand_x4_sg U70715 ( .A(n27056), .B(n27057), .X(n26996) );
  nand_x1_sg U70716 ( .A(n46023), .B(n52640), .X(n27056) );
  nand_x1_sg U70717 ( .A(n27003), .B(n51063), .X(n27058) );
  nand_x4_sg U70718 ( .A(n26220), .B(n26221), .X(n26160) );
  nand_x1_sg U70719 ( .A(n46017), .B(n51811), .X(n26220) );
  nand_x1_sg U70720 ( .A(n26167), .B(n51005), .X(n26222) );
  nand_x4_sg U70721 ( .A(n26499), .B(n26500), .X(n26439) );
  nand_x1_sg U70722 ( .A(n46011), .B(n52087), .X(n26499) );
  nand_x1_sg U70723 ( .A(n26446), .B(n51024), .X(n26501) );
  nand_x4_sg U70724 ( .A(n27336), .B(n27337), .X(n27276) );
  nand_x1_sg U70725 ( .A(n46009), .B(n52921), .X(n27336) );
  nand_x1_sg U70726 ( .A(n27283), .B(n51082), .X(n27338) );
  nand_x4_sg U70727 ( .A(n27894), .B(n27895), .X(n27834) );
  nand_x1_sg U70728 ( .A(n46007), .B(n53479), .X(n27894) );
  nand_x1_sg U70729 ( .A(n27841), .B(n51120), .X(n27896) );
  nand_x1_sg U70730 ( .A(n42805), .B(n51045), .X(n26774) );
  nand_x1_sg U70731 ( .A(n45317), .B(n26776), .X(n26775) );
  nand_x1_sg U70732 ( .A(n46177), .B(n26717), .X(n26776) );
  nand_x1_sg U70733 ( .A(n52375), .B(n46151), .X(n26770) );
  nand_x1_sg U70734 ( .A(n42833), .B(n51196), .X(n29008) );
  nand_x1_sg U70735 ( .A(n45311), .B(n29010), .X(n29009) );
  nand_x1_sg U70736 ( .A(n46171), .B(n28951), .X(n29010) );
  nand_x1_sg U70737 ( .A(n42831), .B(n51234), .X(n29569) );
  nand_x1_sg U70738 ( .A(n45315), .B(n29571), .X(n29570) );
  nand_x1_sg U70739 ( .A(n46175), .B(n29512), .X(n29571) );
  nand_x1_sg U70740 ( .A(n42829), .B(n50968), .X(n25658) );
  nand_x1_sg U70741 ( .A(n45303), .B(n25660), .X(n25659) );
  nand_x1_sg U70742 ( .A(n46163), .B(n25599), .X(n25660) );
  nand_x1_sg U70743 ( .A(n42823), .B(n50987), .X(n25937) );
  nand_x1_sg U70744 ( .A(n45305), .B(n25939), .X(n25938) );
  nand_x1_sg U70745 ( .A(n46165), .B(n25880), .X(n25939) );
  nand_x1_sg U70746 ( .A(n42821), .B(n51025), .X(n26496) );
  nand_x1_sg U70747 ( .A(n45323), .B(n26498), .X(n26497) );
  nand_x1_sg U70748 ( .A(n46183), .B(n26439), .X(n26498) );
  nand_x1_sg U70749 ( .A(n42819), .B(n51083), .X(n27333) );
  nand_x1_sg U70750 ( .A(n45321), .B(n27335), .X(n27334) );
  nand_x1_sg U70751 ( .A(n46181), .B(n27276), .X(n27335) );
  nand_x1_sg U70752 ( .A(n42817), .B(n51121), .X(n27891) );
  nand_x1_sg U70753 ( .A(n45319), .B(n27893), .X(n27892) );
  nand_x1_sg U70754 ( .A(n46179), .B(n27834), .X(n27893) );
  nand_x1_sg U70755 ( .A(n42825), .B(n51006), .X(n26217) );
  nand_x1_sg U70756 ( .A(n45325), .B(n26219), .X(n26218) );
  nand_x1_sg U70757 ( .A(n46185), .B(n26160), .X(n26219) );
  nand_x1_sg U70758 ( .A(n42827), .B(n51102), .X(n27612) );
  nand_x1_sg U70759 ( .A(n45307), .B(n27614), .X(n27613) );
  nand_x1_sg U70760 ( .A(n46167), .B(n27555), .X(n27614) );
  nand_x1_sg U70761 ( .A(n42841), .B(n51140), .X(n28172) );
  nand_x1_sg U70762 ( .A(n45299), .B(n28174), .X(n28173) );
  nand_x1_sg U70763 ( .A(n46159), .B(n28115), .X(n28174) );
  nand_x1_sg U70764 ( .A(n42839), .B(n51177), .X(n28730) );
  nand_x1_sg U70765 ( .A(n45297), .B(n28732), .X(n28731) );
  nand_x1_sg U70766 ( .A(n46157), .B(n28673), .X(n28732) );
  nand_x1_sg U70767 ( .A(n42837), .B(n51215), .X(n29291) );
  nand_x1_sg U70768 ( .A(n45295), .B(n29293), .X(n29292) );
  nand_x1_sg U70769 ( .A(n46155), .B(n29234), .X(n29293) );
  nand_x1_sg U70770 ( .A(n42835), .B(n51064), .X(n27053) );
  nand_x1_sg U70771 ( .A(n45313), .B(n27055), .X(n27054) );
  nand_x1_sg U70772 ( .A(n46173), .B(n26996), .X(n27055) );
  nand_x4_sg U70773 ( .A(n28445), .B(n28446), .X(n28377) );
  nand_x1_sg U70774 ( .A(n54057), .B(n51160), .X(n28445) );
  nand_x1_sg U70775 ( .A(n45271), .B(n28447), .X(n28446) );
  nand_x1_sg U70776 ( .A(n46147), .B(n54618), .X(n29004) );
  nand_x1_sg U70777 ( .A(n46145), .B(n55186), .X(n29565) );
  nand_x1_sg U70778 ( .A(n46133), .B(n51264), .X(n25654) );
  nand_x1_sg U70779 ( .A(n46143), .B(n53211), .X(n27608) );
  nand_x1_sg U70780 ( .A(n46139), .B(n51823), .X(n26213) );
  nand_x1_sg U70781 ( .A(n52652), .B(n46169), .X(n27049) );
  nand_x2_sg U70782 ( .A(n8760), .B(n24397), .X(n24396) );
  nand_x2_sg U70783 ( .A(n24320), .B(n24323), .X(n24395) );
  nand_x1_sg U70784 ( .A(n50176), .B(n50183), .X(n24397) );
  nand_x2_sg U70785 ( .A(n8460), .B(n32063), .X(n32062) );
  nand_x2_sg U70786 ( .A(n31986), .B(n31989), .X(n32061) );
  nand_x1_sg U70787 ( .A(n49317), .B(n49324), .X(n32063) );
  nand_x2_sg U70788 ( .A(n8600), .B(n23165), .X(n23164) );
  nand_x2_sg U70789 ( .A(n22932), .B(n22935), .X(n23163) );
  nand_x1_sg U70790 ( .A(n50162), .B(n50191), .X(n23165) );
  nand_x2_sg U70791 ( .A(n8300), .B(n30831), .X(n30830) );
  nand_x2_sg U70792 ( .A(n30598), .B(n30601), .X(n30829) );
  nand_x1_sg U70793 ( .A(n49303), .B(n49332), .X(n30831) );
  nand_x2_sg U70794 ( .A(n8720), .B(n24198), .X(n24197) );
  nand_x2_sg U70795 ( .A(n24079), .B(n24082), .X(n24196) );
  nand_x1_sg U70796 ( .A(n50172), .B(n50185), .X(n24198) );
  nand_x2_sg U70797 ( .A(n8520), .B(n22240), .X(n22239) );
  nand_x2_sg U70798 ( .A(n22064), .B(n22067), .X(n22238) );
  nand_x1_sg U70799 ( .A(n50156), .B(n50195), .X(n22240) );
  nand_x2_sg U70800 ( .A(n8220), .B(n29905), .X(n29904) );
  nand_x2_sg U70801 ( .A(n29729), .B(n29732), .X(n29903) );
  nand_x1_sg U70802 ( .A(n49297), .B(n49336), .X(n29905) );
  nand_x2_sg U70803 ( .A(n8420), .B(n31864), .X(n31863) );
  nand_x2_sg U70804 ( .A(n31745), .B(n31748), .X(n31862) );
  nand_x1_sg U70805 ( .A(n49313), .B(n49326), .X(n31864) );
  nand_x2_sg U70806 ( .A(n8757), .B(n24388), .X(n24387) );
  nand_x2_sg U70807 ( .A(n24339), .B(n24342), .X(n24386) );
  nand_x1_sg U70808 ( .A(n50315), .B(n50319), .X(n24388) );
  nand_x2_sg U70809 ( .A(n8457), .B(n32054), .X(n32053) );
  nand_x2_sg U70810 ( .A(n32005), .B(n32008), .X(n32052) );
  nand_x1_sg U70811 ( .A(n49456), .B(n49460), .X(n32054) );
  nand_x2_sg U70812 ( .A(n8719), .B(n24195), .X(n24194) );
  nand_x2_sg U70813 ( .A(n24086), .B(n24089), .X(n24193) );
  nand_x1_sg U70814 ( .A(n50220), .B(n50229), .X(n24195) );
  nand_x2_sg U70815 ( .A(n8716), .B(n24186), .X(n24185) );
  nand_x2_sg U70816 ( .A(n24107), .B(n24110), .X(n24184) );
  nand_x1_sg U70817 ( .A(n50356), .B(n50368), .X(n24186) );
  nand_x2_sg U70818 ( .A(n8718), .B(n24192), .X(n24191) );
  nand_x2_sg U70819 ( .A(n24093), .B(n24096), .X(n24190) );
  nand_x1_sg U70820 ( .A(n50265), .B(n50275), .X(n24192) );
  nand_x2_sg U70821 ( .A(n8416), .B(n31852), .X(n31851) );
  nand_x2_sg U70822 ( .A(n31773), .B(n31776), .X(n31850) );
  nand_x1_sg U70823 ( .A(n49497), .B(n49509), .X(n31852) );
  nand_x2_sg U70824 ( .A(n8418), .B(n31858), .X(n31857) );
  nand_x2_sg U70825 ( .A(n31759), .B(n31762), .X(n31856) );
  nand_x1_sg U70826 ( .A(n49406), .B(n49416), .X(n31858) );
  nand_x2_sg U70827 ( .A(n8419), .B(n31861), .X(n31860) );
  nand_x2_sg U70828 ( .A(n31752), .B(n31755), .X(n31859) );
  nand_x1_sg U70829 ( .A(n49361), .B(n49370), .X(n31861) );
  nand_x2_sg U70830 ( .A(n8717), .B(n24189), .X(n24188) );
  nand_x2_sg U70831 ( .A(n24100), .B(n24103), .X(n24187) );
  nand_x1_sg U70832 ( .A(n50310), .B(n50321), .X(n24189) );
  nand_x2_sg U70833 ( .A(n8417), .B(n31855), .X(n31854) );
  nand_x2_sg U70834 ( .A(n31766), .B(n31769), .X(n31853) );
  nand_x1_sg U70835 ( .A(n49451), .B(n49462), .X(n31855) );
  nand_x2_sg U70836 ( .A(n8591), .B(n23138), .X(n23137) );
  nand_x2_sg U70837 ( .A(n22995), .B(n22998), .X(n23136) );
  nand_x1_sg U70838 ( .A(n50578), .B(n50610), .X(n23138) );
  nand_x2_sg U70839 ( .A(n8597), .B(n23156), .X(n23155) );
  nand_x2_sg U70840 ( .A(n22953), .B(n22956), .X(n23154) );
  nand_x1_sg U70841 ( .A(n50298), .B(n50327), .X(n23156) );
  nand_x2_sg U70842 ( .A(n8599), .B(n23162), .X(n23161) );
  nand_x2_sg U70843 ( .A(n22939), .B(n22942), .X(n23160) );
  nand_x1_sg U70844 ( .A(n50208), .B(n50235), .X(n23162) );
  nand_x2_sg U70845 ( .A(n8291), .B(n30804), .X(n30803) );
  nand_x2_sg U70846 ( .A(n30661), .B(n30664), .X(n30802) );
  nand_x1_sg U70847 ( .A(n49719), .B(n49751), .X(n30804) );
  nand_x2_sg U70848 ( .A(n8297), .B(n30822), .X(n30821) );
  nand_x2_sg U70849 ( .A(n30619), .B(n30622), .X(n30820) );
  nand_x1_sg U70850 ( .A(n49439), .B(n49468), .X(n30822) );
  nand_x2_sg U70851 ( .A(n8299), .B(n30828), .X(n30827) );
  nand_x2_sg U70852 ( .A(n30605), .B(n30608), .X(n30826) );
  nand_x1_sg U70853 ( .A(n49349), .B(n49376), .X(n30828) );
  nand_x2_sg U70854 ( .A(n8507), .B(n22201), .X(n22200) );
  nand_x2_sg U70855 ( .A(n22155), .B(n22158), .X(n22199) );
  nand_x1_sg U70856 ( .A(n50760), .B(n50804), .X(n22201) );
  nand_x2_sg U70857 ( .A(n8588), .B(n23129), .X(n23128) );
  nand_x2_sg U70858 ( .A(n23016), .B(n23019), .X(n23127) );
  nand_x1_sg U70859 ( .A(n50722), .B(n50752), .X(n23129) );
  nand_x2_sg U70860 ( .A(n8508), .B(n22204), .X(n22203) );
  nand_x2_sg U70861 ( .A(n22148), .B(n22151), .X(n22202) );
  nand_x1_sg U70862 ( .A(n50713), .B(n50756), .X(n22204) );
  nand_x2_sg U70863 ( .A(n8589), .B(n23132), .X(n23131) );
  nand_x2_sg U70864 ( .A(n23009), .B(n23012), .X(n23130) );
  nand_x1_sg U70865 ( .A(n50674), .B(n50705), .X(n23132) );
  nand_x2_sg U70866 ( .A(n8509), .B(n22207), .X(n22206) );
  nand_x2_sg U70867 ( .A(n22141), .B(n22144), .X(n22205) );
  nand_x1_sg U70868 ( .A(n50665), .B(n50709), .X(n22207) );
  nand_x2_sg U70869 ( .A(n8590), .B(n23135), .X(n23134) );
  nand_x2_sg U70870 ( .A(n23002), .B(n23005), .X(n23133) );
  nand_x1_sg U70871 ( .A(n50627), .B(n50658), .X(n23135) );
  nand_x2_sg U70872 ( .A(n8510), .B(n22210), .X(n22209) );
  nand_x2_sg U70873 ( .A(n22134), .B(n22137), .X(n22208) );
  nand_x1_sg U70874 ( .A(n50618), .B(n50661), .X(n22210) );
  nand_x2_sg U70875 ( .A(n8511), .B(n22213), .X(n22212) );
  nand_x2_sg U70876 ( .A(n22127), .B(n22130), .X(n22211) );
  nand_x1_sg U70877 ( .A(n50569), .B(n50614), .X(n22213) );
  nand_x2_sg U70878 ( .A(n8592), .B(n23141), .X(n23140) );
  nand_x2_sg U70879 ( .A(n22988), .B(n22991), .X(n23139) );
  nand_x1_sg U70880 ( .A(n50531), .B(n50561), .X(n23141) );
  nand_x2_sg U70881 ( .A(n8512), .B(n22216), .X(n22215) );
  nand_x2_sg U70882 ( .A(n22120), .B(n22123), .X(n22214) );
  nand_x1_sg U70883 ( .A(n50522), .B(n50565), .X(n22216) );
  nand_x2_sg U70884 ( .A(n8593), .B(n23144), .X(n23143) );
  nand_x2_sg U70885 ( .A(n22981), .B(n22984), .X(n23142) );
  nand_x1_sg U70886 ( .A(n50484), .B(n50514), .X(n23144) );
  nand_x2_sg U70887 ( .A(n8513), .B(n22219), .X(n22218) );
  nand_x2_sg U70888 ( .A(n22113), .B(n22116), .X(n22217) );
  nand_x1_sg U70889 ( .A(n50475), .B(n50518), .X(n22219) );
  nand_x2_sg U70890 ( .A(n8594), .B(n23147), .X(n23146) );
  nand_x2_sg U70891 ( .A(n22974), .B(n22977), .X(n23145) );
  nand_x1_sg U70892 ( .A(n50438), .B(n50467), .X(n23147) );
  nand_x2_sg U70893 ( .A(n8514), .B(n22222), .X(n22221) );
  nand_x2_sg U70894 ( .A(n22106), .B(n22109), .X(n22220) );
  nand_x1_sg U70895 ( .A(n50429), .B(n50471), .X(n22222) );
  nand_x2_sg U70896 ( .A(n8595), .B(n23150), .X(n23149) );
  nand_x2_sg U70897 ( .A(n22967), .B(n22970), .X(n23148) );
  nand_x1_sg U70898 ( .A(n50391), .B(n50421), .X(n23150) );
  nand_x2_sg U70899 ( .A(n8515), .B(n22225), .X(n22224) );
  nand_x2_sg U70900 ( .A(n22099), .B(n22102), .X(n22223) );
  nand_x1_sg U70901 ( .A(n50382), .B(n50425), .X(n22225) );
  nand_x2_sg U70902 ( .A(n8596), .B(n23153), .X(n23152) );
  nand_x2_sg U70903 ( .A(n22960), .B(n22963), .X(n23151) );
  nand_x1_sg U70904 ( .A(n50344), .B(n50374), .X(n23153) );
  nand_x2_sg U70905 ( .A(n8516), .B(n22228), .X(n22227) );
  nand_x2_sg U70906 ( .A(n22092), .B(n22095), .X(n22226) );
  nand_x1_sg U70907 ( .A(n50335), .B(n50378), .X(n22228) );
  nand_x2_sg U70908 ( .A(n8517), .B(n22231), .X(n22230) );
  nand_x2_sg U70909 ( .A(n22085), .B(n22088), .X(n22229) );
  nand_x1_sg U70910 ( .A(n50289), .B(n50331), .X(n22231) );
  nand_x2_sg U70911 ( .A(n8598), .B(n23159), .X(n23158) );
  nand_x2_sg U70912 ( .A(n22946), .B(n22949), .X(n23157) );
  nand_x1_sg U70913 ( .A(n50252), .B(n50281), .X(n23159) );
  nand_x2_sg U70914 ( .A(n8518), .B(n22234), .X(n22233) );
  nand_x2_sg U70915 ( .A(n22078), .B(n22081), .X(n22232) );
  nand_x1_sg U70916 ( .A(n50243), .B(n50285), .X(n22234) );
  nand_x2_sg U70917 ( .A(n8519), .B(n22237), .X(n22236) );
  nand_x2_sg U70918 ( .A(n22071), .B(n22074), .X(n22235) );
  nand_x1_sg U70919 ( .A(n50199), .B(n50239), .X(n22237) );
  nand_x2_sg U70920 ( .A(n8207), .B(n29866), .X(n29865) );
  nand_x2_sg U70921 ( .A(n29820), .B(n29823), .X(n29864) );
  nand_x1_sg U70922 ( .A(n49901), .B(n49945), .X(n29866) );
  nand_x2_sg U70923 ( .A(n8288), .B(n30795), .X(n30794) );
  nand_x2_sg U70924 ( .A(n30682), .B(n30685), .X(n30793) );
  nand_x1_sg U70925 ( .A(n49863), .B(n49893), .X(n30795) );
  nand_x2_sg U70926 ( .A(n8208), .B(n29869), .X(n29868) );
  nand_x2_sg U70927 ( .A(n29813), .B(n29816), .X(n29867) );
  nand_x1_sg U70928 ( .A(n49854), .B(n49897), .X(n29869) );
  nand_x2_sg U70929 ( .A(n8289), .B(n30798), .X(n30797) );
  nand_x2_sg U70930 ( .A(n30675), .B(n30678), .X(n30796) );
  nand_x1_sg U70931 ( .A(n49815), .B(n49846), .X(n30798) );
  nand_x2_sg U70932 ( .A(n8209), .B(n29872), .X(n29871) );
  nand_x2_sg U70933 ( .A(n29806), .B(n29809), .X(n29870) );
  nand_x1_sg U70934 ( .A(n49806), .B(n49850), .X(n29872) );
  nand_x2_sg U70935 ( .A(n8290), .B(n30801), .X(n30800) );
  nand_x2_sg U70936 ( .A(n30668), .B(n30671), .X(n30799) );
  nand_x1_sg U70937 ( .A(n49768), .B(n49799), .X(n30801) );
  nand_x2_sg U70938 ( .A(n8210), .B(n29875), .X(n29874) );
  nand_x2_sg U70939 ( .A(n29799), .B(n29802), .X(n29873) );
  nand_x1_sg U70940 ( .A(n49759), .B(n49802), .X(n29875) );
  nand_x2_sg U70941 ( .A(n8211), .B(n29878), .X(n29877) );
  nand_x2_sg U70942 ( .A(n29792), .B(n29795), .X(n29876) );
  nand_x1_sg U70943 ( .A(n49710), .B(n49755), .X(n29878) );
  nand_x2_sg U70944 ( .A(n8292), .B(n30807), .X(n30806) );
  nand_x2_sg U70945 ( .A(n30654), .B(n30657), .X(n30805) );
  nand_x1_sg U70946 ( .A(n49672), .B(n49702), .X(n30807) );
  nand_x2_sg U70947 ( .A(n8212), .B(n29881), .X(n29880) );
  nand_x2_sg U70948 ( .A(n29785), .B(n29788), .X(n29879) );
  nand_x1_sg U70949 ( .A(n49663), .B(n49706), .X(n29881) );
  nand_x2_sg U70950 ( .A(n8293), .B(n30810), .X(n30809) );
  nand_x2_sg U70951 ( .A(n30647), .B(n30650), .X(n30808) );
  nand_x1_sg U70952 ( .A(n49625), .B(n49655), .X(n30810) );
  nand_x2_sg U70953 ( .A(n8213), .B(n29884), .X(n29883) );
  nand_x2_sg U70954 ( .A(n29778), .B(n29781), .X(n29882) );
  nand_x1_sg U70955 ( .A(n49616), .B(n49659), .X(n29884) );
  nand_x2_sg U70956 ( .A(n8294), .B(n30813), .X(n30812) );
  nand_x2_sg U70957 ( .A(n30640), .B(n30643), .X(n30811) );
  nand_x1_sg U70958 ( .A(n49579), .B(n49608), .X(n30813) );
  nand_x2_sg U70959 ( .A(n8214), .B(n29887), .X(n29886) );
  nand_x2_sg U70960 ( .A(n29771), .B(n29774), .X(n29885) );
  nand_x1_sg U70961 ( .A(n49570), .B(n49612), .X(n29887) );
  nand_x2_sg U70962 ( .A(n8295), .B(n30816), .X(n30815) );
  nand_x2_sg U70963 ( .A(n30633), .B(n30636), .X(n30814) );
  nand_x1_sg U70964 ( .A(n49532), .B(n49562), .X(n30816) );
  nand_x2_sg U70965 ( .A(n8215), .B(n29890), .X(n29889) );
  nand_x2_sg U70966 ( .A(n29764), .B(n29767), .X(n29888) );
  nand_x1_sg U70967 ( .A(n49523), .B(n49566), .X(n29890) );
  nand_x2_sg U70968 ( .A(n8296), .B(n30819), .X(n30818) );
  nand_x2_sg U70969 ( .A(n30626), .B(n30629), .X(n30817) );
  nand_x1_sg U70970 ( .A(n49485), .B(n49515), .X(n30819) );
  nand_x2_sg U70971 ( .A(n8216), .B(n29893), .X(n29892) );
  nand_x2_sg U70972 ( .A(n29757), .B(n29760), .X(n29891) );
  nand_x1_sg U70973 ( .A(n49476), .B(n49519), .X(n29893) );
  nand_x2_sg U70974 ( .A(n8217), .B(n29896), .X(n29895) );
  nand_x2_sg U70975 ( .A(n29750), .B(n29753), .X(n29894) );
  nand_x1_sg U70976 ( .A(n49430), .B(n49472), .X(n29896) );
  nand_x2_sg U70977 ( .A(n8298), .B(n30825), .X(n30824) );
  nand_x2_sg U70978 ( .A(n30612), .B(n30615), .X(n30823) );
  nand_x1_sg U70979 ( .A(n49393), .B(n49422), .X(n30825) );
  nand_x2_sg U70980 ( .A(n8218), .B(n29899), .X(n29898) );
  nand_x2_sg U70981 ( .A(n29743), .B(n29746), .X(n29897) );
  nand_x1_sg U70982 ( .A(n49384), .B(n49426), .X(n29899) );
  nand_x2_sg U70983 ( .A(n8219), .B(n29902), .X(n29901) );
  nand_x2_sg U70984 ( .A(n29736), .B(n29739), .X(n29900) );
  nand_x1_sg U70985 ( .A(n49340), .B(n49380), .X(n29902) );
  nand_x2_sg U70986 ( .A(n8714), .B(n24180), .X(n24179) );
  nand_x2_sg U70987 ( .A(n24121), .B(n24124), .X(n24178) );
  nand_x1_sg U70988 ( .A(n50450), .B(n50461), .X(n24180) );
  nand_x2_sg U70989 ( .A(n8715), .B(n24183), .X(n24182) );
  nand_x2_sg U70990 ( .A(n24114), .B(n24117), .X(n24181) );
  nand_x1_sg U70991 ( .A(n50404), .B(n50415), .X(n24183) );
  nand_x2_sg U70992 ( .A(n8414), .B(n31846), .X(n31845) );
  nand_x2_sg U70993 ( .A(n31787), .B(n31790), .X(n31844) );
  nand_x1_sg U70994 ( .A(n49591), .B(n49602), .X(n31846) );
  nand_x2_sg U70995 ( .A(n8415), .B(n31849), .X(n31848) );
  nand_x2_sg U70996 ( .A(n31780), .B(n31783), .X(n31847) );
  nand_x1_sg U70997 ( .A(n49545), .B(n49556), .X(n31849) );
  nand_x1_sg U70998 ( .A(n54081), .B(n45983), .X(n28438) );
  nand_x1_sg U70999 ( .A(n54058), .B(n45987), .X(n28444) );
  nand_x4_sg U71000 ( .A(n51574), .B(n25858), .X(n25856) );
  nand_x1_sg U71001 ( .A(n43757), .B(n50991), .X(n25858) );
  nor_x1_sg U71002 ( .A(n50991), .B(n46035), .X(n25859) );
  nand_x4_sg U71003 ( .A(n52131), .B(n26417), .X(n26415) );
  nand_x1_sg U71004 ( .A(n43753), .B(n51029), .X(n26417) );
  nor_x1_sg U71005 ( .A(n51029), .B(n45225), .X(n26418) );
  nand_x4_sg U71006 ( .A(n52965), .B(n27254), .X(n27252) );
  nand_x1_sg U71007 ( .A(n43751), .B(n51087), .X(n27254) );
  nor_x1_sg U71008 ( .A(n51087), .B(n45223), .X(n27255) );
  nand_x4_sg U71009 ( .A(n53523), .B(n27812), .X(n27810) );
  nand_x1_sg U71010 ( .A(n43749), .B(n51125), .X(n27812) );
  nor_x1_sg U71011 ( .A(n51125), .B(n45221), .X(n27813) );
  nand_x4_sg U71012 ( .A(n53800), .B(n28093), .X(n28091) );
  nand_x1_sg U71013 ( .A(n43779), .B(n51144), .X(n28093) );
  nor_x1_sg U71014 ( .A(n51144), .B(n46041), .X(n28094) );
  nand_x4_sg U71015 ( .A(n54365), .B(n28651), .X(n28649) );
  nand_x1_sg U71016 ( .A(n43777), .B(n51181), .X(n28651) );
  nor_x1_sg U71017 ( .A(n51181), .B(n46039), .X(n28652) );
  nand_x4_sg U71018 ( .A(n54933), .B(n29212), .X(n29210) );
  nand_x1_sg U71019 ( .A(n43775), .B(n51219), .X(n29212) );
  nor_x1_sg U71020 ( .A(n51219), .B(n46037), .X(n29213) );
  nand_x4_sg U71021 ( .A(n26974), .B(n26975), .X(n26972) );
  nand_x1_sg U71022 ( .A(n44817), .B(n51068), .X(n26975) );
  nand_x1_sg U71023 ( .A(n46149), .B(n52681), .X(n26974) );
  nand_x4_sg U71024 ( .A(n25624), .B(n25625), .X(n25621) );
  nand_x1_sg U71025 ( .A(n25627), .B(n50984), .X(n25624) );
  nand_x1_sg U71026 ( .A(n45241), .B(n25626), .X(n25625) );
  nand_x1_sg U71027 ( .A(n51515), .B(n46087), .X(n25626) );
  nand_x4_sg U71028 ( .A(n25905), .B(n25906), .X(n25902) );
  nand_x1_sg U71029 ( .A(n11693), .B(n51003), .X(n25905) );
  nand_x1_sg U71030 ( .A(n45259), .B(n25907), .X(n25906) );
  nand_x1_sg U71031 ( .A(n51795), .B(n46105), .X(n25907) );
  nand_x4_sg U71032 ( .A(n26185), .B(n26186), .X(n26182) );
  nand_x1_sg U71033 ( .A(n12472), .B(n51022), .X(n26185) );
  nand_x1_sg U71034 ( .A(n45263), .B(n26187), .X(n26186) );
  nand_x1_sg U71035 ( .A(n52071), .B(n46109), .X(n26187) );
  nand_x4_sg U71036 ( .A(n26464), .B(n26465), .X(n26461) );
  nand_x1_sg U71037 ( .A(n13253), .B(n51041), .X(n26464) );
  nand_x1_sg U71038 ( .A(n45269), .B(n26466), .X(n26465) );
  nand_x1_sg U71039 ( .A(n52349), .B(n46115), .X(n26466) );
  nand_x4_sg U71040 ( .A(n26742), .B(n26743), .X(n26739) );
  nand_x1_sg U71041 ( .A(n14033), .B(n51061), .X(n26742) );
  nand_x1_sg U71042 ( .A(n45261), .B(n26744), .X(n26743) );
  nand_x1_sg U71043 ( .A(n52624), .B(n46107), .X(n26744) );
  nand_x4_sg U71044 ( .A(n27021), .B(n27022), .X(n27018) );
  nand_x1_sg U71045 ( .A(n14805), .B(n51080), .X(n27021) );
  nand_x1_sg U71046 ( .A(n45249), .B(n27023), .X(n27022) );
  nand_x1_sg U71047 ( .A(n52905), .B(n46095), .X(n27023) );
  nand_x4_sg U71048 ( .A(n27301), .B(n27302), .X(n27298) );
  nand_x1_sg U71049 ( .A(n15586), .B(n51099), .X(n27301) );
  nand_x1_sg U71050 ( .A(n45267), .B(n27303), .X(n27302) );
  nand_x1_sg U71051 ( .A(n53183), .B(n46113), .X(n27303) );
  nand_x4_sg U71052 ( .A(n27580), .B(n27581), .X(n27577) );
  nand_x1_sg U71053 ( .A(n16367), .B(n51118), .X(n27580) );
  nand_x1_sg U71054 ( .A(n45257), .B(n27582), .X(n27581) );
  nand_x1_sg U71055 ( .A(n53463), .B(n46103), .X(n27582) );
  nand_x4_sg U71056 ( .A(n27859), .B(n27860), .X(n27856) );
  nand_x1_sg U71057 ( .A(n17152), .B(n51137), .X(n27859) );
  nand_x1_sg U71058 ( .A(n45265), .B(n27861), .X(n27860) );
  nand_x1_sg U71059 ( .A(n53741), .B(n46111), .X(n27861) );
  nand_x4_sg U71060 ( .A(n28140), .B(n28141), .X(n28137) );
  nand_x1_sg U71061 ( .A(n17926), .B(n51156), .X(n28140) );
  nand_x1_sg U71062 ( .A(n45255), .B(n28142), .X(n28141) );
  nand_x1_sg U71063 ( .A(n54025), .B(n46101), .X(n28142) );
  nand_x4_sg U71064 ( .A(n28419), .B(n28420), .X(n28416) );
  nand_x1_sg U71065 ( .A(n18695), .B(n51174), .X(n28419) );
  nand_x1_sg U71066 ( .A(n45247), .B(n28421), .X(n28420) );
  nand_x1_sg U71067 ( .A(n54306), .B(n46093), .X(n28421) );
  nand_x4_sg U71068 ( .A(n28698), .B(n28699), .X(n28695) );
  nand_x1_sg U71069 ( .A(n19471), .B(n51193), .X(n28698) );
  nand_x1_sg U71070 ( .A(n45253), .B(n28700), .X(n28699) );
  nand_x1_sg U71071 ( .A(n54590), .B(n46099), .X(n28700) );
  nand_x4_sg U71072 ( .A(n28976), .B(n28977), .X(n28973) );
  nand_x1_sg U71073 ( .A(n20241), .B(n51212), .X(n28976) );
  nand_x1_sg U71074 ( .A(n45245), .B(n28978), .X(n28977) );
  nand_x1_sg U71075 ( .A(n54874), .B(n46091), .X(n28978) );
  nand_x4_sg U71076 ( .A(n29259), .B(n29260), .X(n29256) );
  nand_x1_sg U71077 ( .A(n21015), .B(n51231), .X(n29259) );
  nand_x1_sg U71078 ( .A(n45251), .B(n29261), .X(n29260) );
  nand_x1_sg U71079 ( .A(n55158), .B(n46097), .X(n29261) );
  nand_x4_sg U71080 ( .A(n29537), .B(n29538), .X(n29534) );
  nand_x1_sg U71081 ( .A(n21786), .B(n51250), .X(n29537) );
  nand_x1_sg U71082 ( .A(n45243), .B(n29539), .X(n29538) );
  nand_x1_sg U71083 ( .A(n55442), .B(n46089), .X(n29539) );
  nand_x4_sg U71084 ( .A(n22609), .B(n22610), .X(n22607) );
  nand_x1_sg U71085 ( .A(n9393), .B(n22612), .X(n22609) );
  nand_x4_sg U71086 ( .A(n21999), .B(n22000), .X(n21997) );
  nand_x1_sg U71087 ( .A(n9383), .B(n9412), .X(n21999) );
  nand_x4_sg U71088 ( .A(n30275), .B(n30276), .X(n30273) );
  nand_x1_sg U71089 ( .A(n24506), .B(n30278), .X(n30275) );
  nand_x4_sg U71090 ( .A(n29664), .B(n29665), .X(n29662) );
  nand_x1_sg U71091 ( .A(n24498), .B(n24521), .X(n29664) );
  nand_x4_sg U71092 ( .A(n22551), .B(n22552), .X(n22549) );
  nand_x1_sg U71093 ( .A(n9372), .B(n22554), .X(n22551) );
  nand_x4_sg U71094 ( .A(n30217), .B(n30218), .X(n30215) );
  nand_x1_sg U71095 ( .A(n24483), .B(n30220), .X(n30217) );
  nand_x2_sg U71096 ( .A(n24467), .B(n40732), .X(n24466) );
  nand_x2_sg U71097 ( .A(n8781), .B(n50108), .X(n24465) );
  nand_x1_sg U71098 ( .A(n24404), .B(n40748), .X(n24467) );
  nand_x2_sg U71099 ( .A(n32133), .B(n40736), .X(n32132) );
  nand_x2_sg U71100 ( .A(n8481), .B(n49249), .X(n32131) );
  nand_x1_sg U71101 ( .A(n32070), .B(n40752), .X(n32133) );
  nand_x4_sg U71102 ( .A(n21985), .B(n21986), .X(n21983) );
  nand_x1_sg U71103 ( .A(n9414), .B(n21988), .X(n21985) );
  nand_x4_sg U71104 ( .A(n22595), .B(n22596), .X(n22593) );
  nand_x1_sg U71105 ( .A(n9384), .B(n22598), .X(n22595) );
  nand_x4_sg U71106 ( .A(n29650), .B(n29651), .X(n29648) );
  nand_x1_sg U71107 ( .A(n24523), .B(n29653), .X(n29650) );
  nand_x4_sg U71108 ( .A(n30261), .B(n30262), .X(n30259) );
  nand_x1_sg U71109 ( .A(n24499), .B(n30264), .X(n30261) );
  nand_x4_sg U71110 ( .A(n22566), .B(n22567), .X(n22564) );
  nand_x1_sg U71111 ( .A(n9366), .B(n22569), .X(n22566) );
  nand_x4_sg U71112 ( .A(n30232), .B(n30233), .X(n30230) );
  nand_x1_sg U71113 ( .A(n24484), .B(n30235), .X(n30232) );
  nand_x4_sg U71114 ( .A(n28099), .B(n28100), .X(n28096) );
  nand_x1_sg U71115 ( .A(n44807), .B(n53786), .X(n28099) );
  nand_x1_sg U71116 ( .A(n45993), .B(n51143), .X(n28100) );
  nand_x4_sg U71117 ( .A(n28657), .B(n28658), .X(n28654) );
  nand_x1_sg U71118 ( .A(n44805), .B(n54351), .X(n28657) );
  nand_x1_sg U71119 ( .A(n45991), .B(n51180), .X(n28658) );
  nand_x4_sg U71120 ( .A(n29218), .B(n29219), .X(n29215) );
  nand_x1_sg U71121 ( .A(n44803), .B(n54919), .X(n29218) );
  nand_x1_sg U71122 ( .A(n45989), .B(n51218), .X(n29219) );
  nand_x4_sg U71123 ( .A(n25864), .B(n25865), .X(n25861) );
  nand_x1_sg U71124 ( .A(n44819), .B(n51558), .X(n25864) );
  nand_x1_sg U71125 ( .A(n46031), .B(n50990), .X(n25865) );
  nand_x4_sg U71126 ( .A(n26423), .B(n26424), .X(n26420) );
  nand_x1_sg U71127 ( .A(n44825), .B(n52115), .X(n26423) );
  nand_x1_sg U71128 ( .A(n45999), .B(n51028), .X(n26424) );
  nand_x4_sg U71129 ( .A(n27260), .B(n27261), .X(n27257) );
  nand_x1_sg U71130 ( .A(n44823), .B(n52949), .X(n27260) );
  nand_x1_sg U71131 ( .A(n45997), .B(n51086), .X(n27261) );
  nand_x4_sg U71132 ( .A(n27818), .B(n27819), .X(n27815) );
  nand_x1_sg U71133 ( .A(n44821), .B(n53507), .X(n27818) );
  nand_x1_sg U71134 ( .A(n45995), .B(n51124), .X(n27819) );
  nand_x4_sg U71135 ( .A(n28366), .B(n28367), .X(n28363) );
  nand_x1_sg U71136 ( .A(n45983), .B(n54095), .X(n28366) );
  nand_x1_sg U71137 ( .A(n45211), .B(n51163), .X(n28367) );
  nand_x4_sg U71138 ( .A(n28087), .B(n28088), .X(n28084) );
  nand_x1_sg U71139 ( .A(n44801), .B(n53812), .X(n28087) );
  nand_x1_sg U71140 ( .A(n45981), .B(n51145), .X(n28088) );
  nand_x4_sg U71141 ( .A(n28645), .B(n28646), .X(n28642) );
  nand_x1_sg U71142 ( .A(n44799), .B(n54377), .X(n28645) );
  nand_x1_sg U71143 ( .A(n45979), .B(n51182), .X(n28646) );
  nand_x4_sg U71144 ( .A(n29206), .B(n29207), .X(n29203) );
  nand_x1_sg U71145 ( .A(n44797), .B(n54945), .X(n29206) );
  nand_x1_sg U71146 ( .A(n45977), .B(n51220), .X(n29207) );
  nand_x4_sg U71147 ( .A(n25852), .B(n25853), .X(n25849) );
  nand_x1_sg U71148 ( .A(n44907), .B(n51586), .X(n25852) );
  nand_x1_sg U71149 ( .A(n46029), .B(n50992), .X(n25853) );
  nand_x4_sg U71150 ( .A(n26411), .B(n26412), .X(n26408) );
  nand_x1_sg U71151 ( .A(n44319), .B(n52144), .X(n26411) );
  nand_x1_sg U71152 ( .A(n45217), .B(n51030), .X(n26412) );
  nand_x4_sg U71153 ( .A(n27248), .B(n27249), .X(n27245) );
  nand_x1_sg U71154 ( .A(n44317), .B(n52978), .X(n27248) );
  nand_x1_sg U71155 ( .A(n45215), .B(n51088), .X(n27249) );
  nand_x4_sg U71156 ( .A(n27806), .B(n27807), .X(n27803) );
  nand_x1_sg U71157 ( .A(n44315), .B(n53536), .X(n27806) );
  nand_x1_sg U71158 ( .A(n45213), .B(n51126), .X(n27807) );
  nand_x1_sg U71159 ( .A(n42847), .B(n51142), .X(n28105) );
  nor_x1_sg U71160 ( .A(n51142), .B(n46059), .X(n28106) );
  nand_x1_sg U71161 ( .A(n42845), .B(n51179), .X(n28663) );
  nor_x1_sg U71162 ( .A(n51179), .B(n46057), .X(n28664) );
  nand_x1_sg U71163 ( .A(n42843), .B(n51217), .X(n29224) );
  nor_x1_sg U71164 ( .A(n51217), .B(n46061), .X(n29225) );
  nand_x1_sg U71165 ( .A(n46073), .B(n51007), .X(n26156) );
  nor_x1_sg U71166 ( .A(n51007), .B(n46073), .X(n26157) );
  nand_x1_sg U71167 ( .A(n46071), .B(n51046), .X(n26713) );
  nor_x1_sg U71168 ( .A(n51046), .B(n46071), .X(n26714) );
  nand_x1_sg U71169 ( .A(n46067), .B(n51141), .X(n28111) );
  nor_x1_sg U71170 ( .A(n51141), .B(n46067), .X(n28112) );
  nand_x1_sg U71171 ( .A(n46065), .B(n51178), .X(n28669) );
  nor_x1_sg U71172 ( .A(n51178), .B(n46065), .X(n28670) );
  nand_x1_sg U71173 ( .A(n46079), .B(n51197), .X(n28947) );
  nor_x1_sg U71174 ( .A(n51197), .B(n46079), .X(n28948) );
  nand_x1_sg U71175 ( .A(n46069), .B(n51216), .X(n29230) );
  nor_x1_sg U71176 ( .A(n51216), .B(n46069), .X(n29231) );
  nand_x1_sg U71177 ( .A(n46081), .B(n51235), .X(n29508) );
  nor_x1_sg U71178 ( .A(n51235), .B(n46081), .X(n29509) );
  nand_x1_sg U71179 ( .A(n46085), .B(n50969), .X(n25595) );
  nor_x1_sg U71180 ( .A(n50969), .B(n46085), .X(n25596) );
  nand_x1_sg U71181 ( .A(n43781), .B(n50989), .X(n25870) );
  nor_x1_sg U71182 ( .A(n50989), .B(n46077), .X(n25871) );
  nand_x1_sg U71183 ( .A(n46063), .B(n50988), .X(n25876) );
  nor_x1_sg U71184 ( .A(n50988), .B(n46063), .X(n25877) );
  nand_x1_sg U71185 ( .A(n43765), .B(n51027), .X(n26429) );
  nor_x1_sg U71186 ( .A(n51027), .B(n46049), .X(n26430) );
  nand_x1_sg U71187 ( .A(n46055), .B(n51026), .X(n26435) );
  nor_x1_sg U71188 ( .A(n51026), .B(n46055), .X(n26436) );
  nand_x1_sg U71189 ( .A(n43763), .B(n51085), .X(n27266) );
  nor_x1_sg U71190 ( .A(n51085), .B(n46047), .X(n27267) );
  nand_x1_sg U71191 ( .A(n46053), .B(n51084), .X(n27272) );
  nor_x1_sg U71192 ( .A(n51084), .B(n46053), .X(n27273) );
  nand_x1_sg U71193 ( .A(n43761), .B(n51123), .X(n27824) );
  nor_x1_sg U71194 ( .A(n51123), .B(n46045), .X(n27825) );
  nand_x1_sg U71195 ( .A(n46051), .B(n51122), .X(n27830) );
  nor_x1_sg U71196 ( .A(n51122), .B(n46051), .X(n27831) );
  nand_x1_sg U71197 ( .A(n46083), .B(n51065), .X(n26992) );
  nor_x1_sg U71198 ( .A(n51065), .B(n46083), .X(n26993) );
  nand_x1_sg U71199 ( .A(n46075), .B(n51103), .X(n27551) );
  nor_x1_sg U71200 ( .A(n51103), .B(n46075), .X(n27552) );
  nand_x2_sg U71201 ( .A(n8777), .B(n40564), .X(n24453) );
  nand_x2_sg U71202 ( .A(n24455), .B(n40793), .X(n24454) );
  nand_x2_sg U71203 ( .A(n8477), .B(n40576), .X(n32119) );
  nand_x2_sg U71204 ( .A(n32121), .B(n40794), .X(n32120) );
  nand_x1_sg U71205 ( .A(n44863), .B(n51195), .X(n28961) );
  nand_x1_sg U71206 ( .A(n46021), .B(n54607), .X(n28960) );
  nand_x1_sg U71207 ( .A(n44875), .B(n51233), .X(n29522) );
  nand_x1_sg U71208 ( .A(n46025), .B(n55175), .X(n29521) );
  nand_x1_sg U71209 ( .A(n44867), .B(n51063), .X(n27006) );
  nand_x1_sg U71210 ( .A(n46023), .B(n52641), .X(n27005) );
  nand_x1_sg U71211 ( .A(n44831), .B(n51139), .X(n28125) );
  nand_x1_sg U71212 ( .A(n46005), .B(n53758), .X(n28124) );
  nand_x1_sg U71213 ( .A(n44815), .B(n51158), .X(n28404) );
  nand_x1_sg U71214 ( .A(n45985), .B(n54042), .X(n28403) );
  nand_x1_sg U71215 ( .A(n44829), .B(n51176), .X(n28683) );
  nand_x1_sg U71216 ( .A(n46003), .B(n54323), .X(n28682) );
  nand_x1_sg U71217 ( .A(n44827), .B(n51214), .X(n29244) );
  nand_x1_sg U71218 ( .A(n46001), .B(n54891), .X(n29243) );
  nand_x1_sg U71219 ( .A(n44845), .B(n51024), .X(n26449) );
  nand_x1_sg U71220 ( .A(n46011), .B(n52088), .X(n26448) );
  nand_x1_sg U71221 ( .A(n44843), .B(n51082), .X(n27286) );
  nand_x1_sg U71222 ( .A(n46009), .B(n52922), .X(n27285) );
  nand_x1_sg U71223 ( .A(n44841), .B(n51120), .X(n27844) );
  nand_x1_sg U71224 ( .A(n46007), .B(n53480), .X(n27843) );
  nand_x1_sg U71225 ( .A(n44857), .B(n51005), .X(n26170) );
  nand_x1_sg U71226 ( .A(n46017), .B(n51812), .X(n26169) );
  nand_x1_sg U71227 ( .A(n44855), .B(n51044), .X(n26727) );
  nand_x1_sg U71228 ( .A(n46015), .B(n52365), .X(n26726) );
  nand_x1_sg U71229 ( .A(n44835), .B(n50986), .X(n25890) );
  nand_x1_sg U71230 ( .A(n46019), .B(n51530), .X(n25889) );
  nand_x1_sg U71231 ( .A(n44847), .B(n51101), .X(n27565) );
  nand_x1_sg U71232 ( .A(n46013), .B(n53200), .X(n27564) );
  nand_x1_sg U71233 ( .A(n45987), .B(n54068), .X(n28378) );
  nand_x1_sg U71234 ( .A(n45219), .B(n51161), .X(n28379) );
  nand_x1_sg U71235 ( .A(n44865), .B(n50967), .X(n25609) );
  nand_x1_sg U71236 ( .A(n46027), .B(n51254), .X(n25608) );
  nand_x4_sg U71237 ( .A(n28929), .B(n28930), .X(n28927) );
  nand_x1_sg U71238 ( .A(n45645), .B(n54645), .X(n28929) );
  nand_x1_sg U71239 ( .A(n44861), .B(n51200), .X(n28930) );
  nand_x4_sg U71240 ( .A(n29490), .B(n29491), .X(n29488) );
  nand_x1_sg U71241 ( .A(n45643), .B(n55213), .X(n29490) );
  nand_x1_sg U71242 ( .A(n44859), .B(n51238), .X(n29491) );
  nand_x4_sg U71243 ( .A(n26695), .B(n26696), .X(n26693) );
  nand_x1_sg U71244 ( .A(n45641), .B(n52404), .X(n26695) );
  nand_x1_sg U71245 ( .A(n44839), .B(n51049), .X(n26696) );
  nand_x4_sg U71246 ( .A(n25577), .B(n25578), .X(n25575) );
  nand_x1_sg U71247 ( .A(n45635), .B(n51291), .X(n25577) );
  nand_x1_sg U71248 ( .A(n44789), .B(n50972), .X(n25578) );
  nand_x4_sg U71249 ( .A(n27533), .B(n27534), .X(n27531) );
  nand_x1_sg U71250 ( .A(n45637), .B(n53238), .X(n27533) );
  nand_x1_sg U71251 ( .A(n44791), .B(n51106), .X(n27534) );
  nand_x4_sg U71252 ( .A(n26138), .B(n26139), .X(n26136) );
  nand_x1_sg U71253 ( .A(n45639), .B(n51852), .X(n26138) );
  nand_x1_sg U71254 ( .A(n44795), .B(n51010), .X(n26139) );
  nand_x4_sg U71255 ( .A(n24380), .B(n24381), .X(n24362) );
  nand_x1_sg U71256 ( .A(n50409), .B(n50413), .X(n24382) );
  nand_x4_sg U71257 ( .A(n32046), .B(n32047), .X(n32028) );
  nand_x1_sg U71258 ( .A(n49550), .B(n49554), .X(n32048) );
  nand_x4_sg U71259 ( .A(n23501), .B(n23502), .X(n23300) );
  nand_x1_sg U71260 ( .A(n50688), .B(n50733), .X(n23503) );
  nand_x4_sg U71261 ( .A(n23862), .B(n23863), .X(n23695) );
  nand_x1_sg U71262 ( .A(n50597), .B(n50642), .X(n23864) );
  nand_x4_sg U71263 ( .A(n24159), .B(n24160), .X(n24019) );
  nand_x1_sg U71264 ( .A(n50506), .B(n50550), .X(n24161) );
  nand_x2_sg U71265 ( .A(n8746), .B(n23072), .X(n23071) );
  nand_x2_sg U71266 ( .A(n23073), .B(n23074), .X(n23070) );
  nand_x1_sg U71267 ( .A(n50780), .B(n50823), .X(n23072) );
  nand_x2_sg U71268 ( .A(n8446), .B(n30738), .X(n30737) );
  nand_x2_sg U71269 ( .A(n30739), .B(n30740), .X(n30736) );
  nand_x1_sg U71270 ( .A(n49921), .B(n49964), .X(n30738) );
  nand_x4_sg U71271 ( .A(n31167), .B(n31168), .X(n30966) );
  nand_x1_sg U71272 ( .A(n49829), .B(n49874), .X(n31169) );
  nand_x4_sg U71273 ( .A(n31528), .B(n31529), .X(n31361) );
  nand_x1_sg U71274 ( .A(n49738), .B(n49783), .X(n31530) );
  nand_x4_sg U71275 ( .A(n31825), .B(n31826), .X(n31685) );
  nand_x1_sg U71276 ( .A(n49647), .B(n49691), .X(n31827) );
  nand_x4_sg U71277 ( .A(n24377), .B(n24378), .X(n24279) );
  nand_x1_sg U71278 ( .A(n41153), .B(n50459), .X(n24379) );
  nand_x2_sg U71279 ( .A(n8749), .B(n23693), .X(n23692) );
  nand_x2_sg U71280 ( .A(n23694), .B(n23695), .X(n23691) );
  nand_x1_sg U71281 ( .A(n41199), .B(n50687), .X(n23693) );
  nand_x2_sg U71282 ( .A(n8751), .B(n24017), .X(n24016) );
  nand_x2_sg U71283 ( .A(n24018), .B(n24019), .X(n24015) );
  nand_x1_sg U71284 ( .A(n41197), .B(n50596), .X(n24017) );
  nand_x2_sg U71285 ( .A(n8747), .B(n23298), .X(n23297) );
  nand_x2_sg U71286 ( .A(n23299), .B(n23300), .X(n23296) );
  nand_x1_sg U71287 ( .A(n41201), .B(n50779), .X(n23298) );
  nand_x4_sg U71288 ( .A(n32043), .B(n32044), .X(n31945) );
  nand_x1_sg U71289 ( .A(n41160), .B(n49600), .X(n32045) );
  nand_x2_sg U71290 ( .A(n8447), .B(n30964), .X(n30963) );
  nand_x2_sg U71291 ( .A(n30965), .B(n30966), .X(n30962) );
  nand_x1_sg U71292 ( .A(n41211), .B(n49920), .X(n30964) );
  nand_x2_sg U71293 ( .A(n8449), .B(n31359), .X(n31358) );
  nand_x2_sg U71294 ( .A(n31360), .B(n31361), .X(n31357) );
  nand_x1_sg U71295 ( .A(n41209), .B(n49828), .X(n31359) );
  nand_x2_sg U71296 ( .A(n8451), .B(n31683), .X(n31682) );
  nand_x2_sg U71297 ( .A(n31684), .B(n31685), .X(n31681) );
  nand_x1_sg U71298 ( .A(n41207), .B(n49737), .X(n31683) );
  nand_x2_sg U71299 ( .A(n8753), .B(n24277), .X(n24276) );
  nand_x2_sg U71300 ( .A(n24278), .B(n24279), .X(n24275) );
  nand_x1_sg U71301 ( .A(n41195), .B(n50505), .X(n24277) );
  nand_x2_sg U71302 ( .A(n8453), .B(n31943), .X(n31942) );
  nand_x2_sg U71303 ( .A(n31944), .B(n31945), .X(n31941) );
  nand_x1_sg U71304 ( .A(n41205), .B(n49646), .X(n31943) );
  nand_x4_sg U71305 ( .A(n22602), .B(n22603), .X(n22600) );
  nand_x1_sg U71306 ( .A(n50933), .B(n22605), .X(n22602) );
  nand_x4_sg U71307 ( .A(n21992), .B(n21993), .X(n21990) );
  nand_x1_sg U71308 ( .A(n50943), .B(n21995), .X(n21992) );
  nand_x4_sg U71309 ( .A(n30268), .B(n30269), .X(n30266) );
  nand_x1_sg U71310 ( .A(n50074), .B(n30271), .X(n30268) );
  nand_x4_sg U71311 ( .A(n29657), .B(n29658), .X(n29655) );
  nand_x1_sg U71312 ( .A(n50084), .B(n29660), .X(n29657) );
  nand_x4_sg U71313 ( .A(n22544), .B(n22545), .X(n22542) );
  nand_x1_sg U71314 ( .A(n50910), .B(n22547), .X(n22544) );
  nand_x4_sg U71315 ( .A(n30210), .B(n30211), .X(n30208) );
  nand_x1_sg U71316 ( .A(n50051), .B(n30213), .X(n30210) );
  nand_x4_sg U71317 ( .A(n25628), .B(n25629), .X(n25622) );
  nand_x1_sg U71318 ( .A(n44787), .B(n51523), .X(n25628) );
  nand_x1_sg U71319 ( .A(n45631), .B(n50985), .X(n25629) );
  nand_x4_sg U71320 ( .A(n25908), .B(n25909), .X(n25903) );
  nand_x1_sg U71321 ( .A(n44785), .B(n51805), .X(n25908) );
  nand_x1_sg U71322 ( .A(n45629), .B(n51004), .X(n25909) );
  nand_x4_sg U71323 ( .A(n26188), .B(n26189), .X(n26183) );
  nand_x1_sg U71324 ( .A(n44783), .B(n52081), .X(n26188) );
  nand_x1_sg U71325 ( .A(n45627), .B(n51023), .X(n26189) );
  nand_x4_sg U71326 ( .A(n26467), .B(n26468), .X(n26462) );
  nand_x1_sg U71327 ( .A(n44781), .B(n52359), .X(n26467) );
  nand_x1_sg U71328 ( .A(n45625), .B(n51042), .X(n26468) );
  nand_x4_sg U71329 ( .A(n26745), .B(n26746), .X(n26740) );
  nand_x1_sg U71330 ( .A(n44779), .B(n52634), .X(n26745) );
  nand_x1_sg U71331 ( .A(n45623), .B(n51062), .X(n26746) );
  nand_x4_sg U71332 ( .A(n27024), .B(n27025), .X(n27019) );
  nand_x1_sg U71333 ( .A(n44777), .B(n52915), .X(n27024) );
  nand_x1_sg U71334 ( .A(n45621), .B(n51081), .X(n27025) );
  nand_x4_sg U71335 ( .A(n27304), .B(n27305), .X(n27299) );
  nand_x1_sg U71336 ( .A(n44775), .B(n53193), .X(n27304) );
  nand_x1_sg U71337 ( .A(n45619), .B(n51100), .X(n27305) );
  nand_x4_sg U71338 ( .A(n27583), .B(n27584), .X(n27578) );
  nand_x1_sg U71339 ( .A(n44773), .B(n53473), .X(n27583) );
  nand_x1_sg U71340 ( .A(n45617), .B(n51119), .X(n27584) );
  nand_x4_sg U71341 ( .A(n27862), .B(n27863), .X(n27857) );
  nand_x1_sg U71342 ( .A(n44771), .B(n53751), .X(n27862) );
  nand_x1_sg U71343 ( .A(n45615), .B(n51138), .X(n27863) );
  nand_x4_sg U71344 ( .A(n28143), .B(n28144), .X(n28138) );
  nand_x1_sg U71345 ( .A(n44769), .B(n54035), .X(n28143) );
  nand_x1_sg U71346 ( .A(n45613), .B(n51157), .X(n28144) );
  nand_x4_sg U71347 ( .A(n28422), .B(n28423), .X(n28417) );
  nand_x1_sg U71348 ( .A(n44767), .B(n54316), .X(n28422) );
  nand_x1_sg U71349 ( .A(n45611), .B(n51175), .X(n28423) );
  nand_x4_sg U71350 ( .A(n28701), .B(n28702), .X(n28696) );
  nand_x1_sg U71351 ( .A(n44765), .B(n54600), .X(n28701) );
  nand_x1_sg U71352 ( .A(n45609), .B(n51194), .X(n28702) );
  nand_x4_sg U71353 ( .A(n28979), .B(n28980), .X(n28974) );
  nand_x1_sg U71354 ( .A(n44763), .B(n54884), .X(n28979) );
  nand_x1_sg U71355 ( .A(n45607), .B(n51213), .X(n28980) );
  nand_x4_sg U71356 ( .A(n29262), .B(n29263), .X(n29257) );
  nand_x1_sg U71357 ( .A(n44761), .B(n55168), .X(n29262) );
  nand_x1_sg U71358 ( .A(n45605), .B(n51232), .X(n29263) );
  nand_x4_sg U71359 ( .A(n29540), .B(n29541), .X(n29535) );
  nand_x1_sg U71360 ( .A(n44759), .B(n55452), .X(n29540) );
  nand_x1_sg U71361 ( .A(n45603), .B(n51251), .X(n29541) );
  nand_x4_sg U71362 ( .A(n31387), .B(n31388), .X(n31330) );
  nand_x1_sg U71363 ( .A(n31203), .B(n40809), .X(n31387) );
  nand_x4_sg U71364 ( .A(n23721), .B(n23722), .X(n23664) );
  nand_x1_sg U71365 ( .A(n23537), .B(n40810), .X(n23721) );
  nand_x4_sg U71366 ( .A(n30992), .B(n30993), .X(n30935) );
  nand_x1_sg U71367 ( .A(n30772), .B(n40811), .X(n30992) );
  nand_x4_sg U71368 ( .A(n23326), .B(n23327), .X(n23269) );
  nand_x1_sg U71369 ( .A(n23106), .B(n40812), .X(n23326) );
  nand_x4_sg U71370 ( .A(n22580), .B(n22581), .X(n22579) );
  nand_x1_sg U71371 ( .A(n43187), .B(n41888), .X(n22580) );
  nand_x1_sg U71372 ( .A(n22583), .B(n50925), .X(n22582) );
  nand_x4_sg U71373 ( .A(n30246), .B(n30247), .X(n30245) );
  nand_x1_sg U71374 ( .A(n43183), .B(n41886), .X(n30246) );
  nand_x1_sg U71375 ( .A(n30249), .B(n50066), .X(n30248) );
  nand_x4_sg U71376 ( .A(n22535), .B(n22536), .X(n22532) );
  nand_x1_sg U71377 ( .A(n8764), .B(n41213), .X(n22535) );
  nand_x1_sg U71378 ( .A(n22538), .B(n40740), .X(n22537) );
  nand_x4_sg U71379 ( .A(n30201), .B(n30202), .X(n30198) );
  nand_x1_sg U71380 ( .A(n8464), .B(n41212), .X(n30201) );
  nand_x1_sg U71381 ( .A(n30204), .B(n40742), .X(n30203) );
  nand_x1_sg U71382 ( .A(n23390), .B(n40813), .X(n23388) );
  nand_x1_sg U71383 ( .A(n8641), .B(n50118), .X(n23389) );
  nand_x1_sg U71384 ( .A(n31056), .B(n40814), .X(n31054) );
  nand_x1_sg U71385 ( .A(n8341), .B(n49259), .X(n31055) );
  nand_x1_sg U71386 ( .A(n23176), .B(n40815), .X(n23174) );
  nand_x1_sg U71387 ( .A(n8621), .B(n50119), .X(n23175) );
  nand_x1_sg U71388 ( .A(n30842), .B(n40816), .X(n30840) );
  nand_x1_sg U71389 ( .A(n8321), .B(n49260), .X(n30841) );
  nand_x1_sg U71390 ( .A(n22928), .B(n40817), .X(n22926) );
  nand_x1_sg U71391 ( .A(n8601), .B(n50120), .X(n22927) );
  nand_x1_sg U71392 ( .A(n22677), .B(n40818), .X(n22675) );
  nand_x1_sg U71393 ( .A(n8581), .B(n50121), .X(n22676) );
  nand_x1_sg U71394 ( .A(n30594), .B(n40819), .X(n30592) );
  nand_x1_sg U71395 ( .A(n8301), .B(n49261), .X(n30593) );
  nand_x1_sg U71396 ( .A(n30343), .B(n40820), .X(n30341) );
  nand_x1_sg U71397 ( .A(n8281), .B(n49262), .X(n30342) );
  nand_x1_sg U71398 ( .A(n22407), .B(n40821), .X(n22405) );
  nand_x1_sg U71399 ( .A(n8561), .B(n50122), .X(n22406) );
  nand_x1_sg U71400 ( .A(n24209), .B(n40822), .X(n24207) );
  nand_x1_sg U71401 ( .A(n8741), .B(n50111), .X(n24208) );
  nand_x1_sg U71402 ( .A(n30072), .B(n40823), .X(n30070) );
  nand_x1_sg U71403 ( .A(n8261), .B(n49263), .X(n30071) );
  nand_x1_sg U71404 ( .A(n31435), .B(n40824), .X(n31433) );
  nand_x1_sg U71405 ( .A(n8381), .B(n49256), .X(n31434) );
  nand_x1_sg U71406 ( .A(n22251), .B(n40825), .X(n22249) );
  nand_x1_sg U71407 ( .A(n8541), .B(n50123), .X(n22250) );
  nand_x1_sg U71408 ( .A(n29916), .B(n40826), .X(n29914) );
  nand_x1_sg U71409 ( .A(n8241), .B(n49264), .X(n29915) );
  nand_x1_sg U71410 ( .A(n22060), .B(n40827), .X(n22058) );
  nand_x1_sg U71411 ( .A(n8521), .B(n50124), .X(n22059) );
  nand_x1_sg U71412 ( .A(n23931), .B(n40828), .X(n23929) );
  nand_x1_sg U71413 ( .A(n8701), .B(n50114), .X(n23930) );
  nand_x1_sg U71414 ( .A(n29725), .B(n40829), .X(n29723) );
  nand_x1_sg U71415 ( .A(n8221), .B(n49265), .X(n29724) );
  nand_x1_sg U71416 ( .A(n31875), .B(n40830), .X(n31873) );
  nand_x1_sg U71417 ( .A(n8441), .B(n49252), .X(n31874) );
  nand_x1_sg U71418 ( .A(n23769), .B(n40831), .X(n23767) );
  nand_x1_sg U71419 ( .A(n8681), .B(n50115), .X(n23768) );
  nand_x1_sg U71420 ( .A(n31597), .B(n40832), .X(n31595) );
  nand_x1_sg U71421 ( .A(n8401), .B(n49255), .X(n31596) );
  nand_x1_sg U71422 ( .A(n24316), .B(n40833), .X(n24314) );
  nand_x1_sg U71423 ( .A(n8761), .B(n50110), .X(n24315) );
  nand_x1_sg U71424 ( .A(n31254), .B(n40834), .X(n31252) );
  nand_x1_sg U71425 ( .A(n8361), .B(n49258), .X(n31253) );
  nand_x1_sg U71426 ( .A(n24075), .B(n40835), .X(n24073) );
  nand_x1_sg U71427 ( .A(n8721), .B(n50113), .X(n24074) );
  nand_x1_sg U71428 ( .A(n31982), .B(n40836), .X(n31980) );
  nand_x1_sg U71429 ( .A(n8461), .B(n49251), .X(n31981) );
  nand_x1_sg U71430 ( .A(n31741), .B(n40837), .X(n31739) );
  nand_x1_sg U71431 ( .A(n8421), .B(n49254), .X(n31740) );
  nand_x1_sg U71432 ( .A(n23588), .B(n40838), .X(n23586) );
  nand_x1_sg U71433 ( .A(n8661), .B(n50117), .X(n23587) );
  nand_x4_sg U71434 ( .A(n24373), .B(n50503), .X(n24368) );
  nand_x1_sg U71435 ( .A(n8773), .B(n40841), .X(n24373) );
  nor_x1_sg U71436 ( .A(n40841), .B(n8773), .X(n24374) );
  nand_x4_sg U71437 ( .A(n23066), .B(n50864), .X(n23061) );
  nand_x1_sg U71438 ( .A(n8765), .B(n40842), .X(n23066) );
  nor_x1_sg U71439 ( .A(n40842), .B(n8765), .X(n23067) );
  nand_x4_sg U71440 ( .A(n23497), .B(n50777), .X(n23492) );
  nand_x1_sg U71441 ( .A(n8767), .B(n40843), .X(n23497) );
  nor_x1_sg U71442 ( .A(n40843), .B(n8767), .X(n23498) );
  nand_x4_sg U71443 ( .A(n23858), .B(n50685), .X(n23853) );
  nand_x1_sg U71444 ( .A(n8769), .B(n40844), .X(n23858) );
  nor_x1_sg U71445 ( .A(n40844), .B(n8769), .X(n23859) );
  nand_x4_sg U71446 ( .A(n24155), .B(n50594), .X(n24150) );
  nand_x1_sg U71447 ( .A(n8771), .B(n40845), .X(n24155) );
  nor_x1_sg U71448 ( .A(n40845), .B(n8771), .X(n24156) );
  nand_x4_sg U71449 ( .A(n32039), .B(n49644), .X(n32034) );
  nand_x1_sg U71450 ( .A(n8473), .B(n40846), .X(n32039) );
  nor_x1_sg U71451 ( .A(n40846), .B(n8473), .X(n32040) );
  nand_x4_sg U71452 ( .A(n30732), .B(n50005), .X(n30727) );
  nand_x1_sg U71453 ( .A(n8465), .B(n40847), .X(n30732) );
  nor_x1_sg U71454 ( .A(n40847), .B(n8465), .X(n30733) );
  nand_x4_sg U71455 ( .A(n31163), .B(n49918), .X(n31158) );
  nand_x1_sg U71456 ( .A(n8467), .B(n40848), .X(n31163) );
  nor_x1_sg U71457 ( .A(n40848), .B(n8467), .X(n31164) );
  nand_x4_sg U71458 ( .A(n31524), .B(n49826), .X(n31519) );
  nand_x1_sg U71459 ( .A(n8469), .B(n40849), .X(n31524) );
  nor_x1_sg U71460 ( .A(n40849), .B(n8469), .X(n31525) );
  nand_x4_sg U71461 ( .A(n31821), .B(n49735), .X(n31816) );
  nand_x1_sg U71462 ( .A(n8471), .B(n40850), .X(n31821) );
  nor_x1_sg U71463 ( .A(n40850), .B(n8471), .X(n31822) );
  nand_x1_sg U71464 ( .A(out_L2[2]), .B(n40723), .X(n24412) );
  nor_x1_sg U71465 ( .A(n40723), .B(out_L2[2]), .X(n24413) );
  nand_x1_sg U71466 ( .A(out_L1[2]), .B(n40724), .X(n32078) );
  nor_x1_sg U71467 ( .A(n40724), .B(out_L1[2]), .X(n32079) );
  nand_x4_sg U71468 ( .A(n31423), .B(n31424), .X(n31267) );
  nand_x1_sg U71469 ( .A(n31258), .B(n31261), .X(n31423) );
  nand_x1_sg U71470 ( .A(n49308), .B(n49329), .X(n31425) );
  nand_x4_sg U71471 ( .A(n23757), .B(n23758), .X(n23601) );
  nand_x1_sg U71472 ( .A(n23592), .B(n23595), .X(n23757) );
  nand_x1_sg U71473 ( .A(n50167), .B(n50188), .X(n23759) );
  nand_x4_sg U71474 ( .A(n50816), .B(n22765), .X(n22764) );
  nor_x1_sg U71475 ( .A(n22766), .B(n8566), .X(n22767) );
  nand_x4_sg U71476 ( .A(n50001), .B(n30437), .X(n30436) );
  nor_x1_sg U71477 ( .A(n30438), .B(n8265), .X(n30439) );
  nand_x4_sg U71478 ( .A(n50626), .B(n22741), .X(n22740) );
  nor_x1_sg U71479 ( .A(n22742), .B(n8570), .X(n22743) );
  nand_x4_sg U71480 ( .A(n50251), .B(n22693), .X(n22692) );
  nor_x1_sg U71481 ( .A(n22694), .B(n8578), .X(n22695) );
  nand_x4_sg U71482 ( .A(n50207), .B(n22687), .X(n22686) );
  nor_x1_sg U71483 ( .A(n22688), .B(n8579), .X(n22689) );
  nand_x4_sg U71484 ( .A(n49767), .B(n30407), .X(n30406) );
  nor_x1_sg U71485 ( .A(n30408), .B(n8270), .X(n30409) );
  nand_x4_sg U71486 ( .A(n49484), .B(n30371), .X(n30370) );
  nor_x1_sg U71487 ( .A(n30372), .B(n8276), .X(n30373) );
  nand_x4_sg U71488 ( .A(n49392), .B(n30359), .X(n30358) );
  nor_x1_sg U71489 ( .A(n30360), .B(n8278), .X(n30361) );
  nand_x4_sg U71490 ( .A(n49348), .B(n30353), .X(n30352) );
  nor_x1_sg U71491 ( .A(n30354), .B(n8279), .X(n30355) );
  nand_x4_sg U71492 ( .A(n50314), .B(n24231), .X(n24230) );
  nor_x1_sg U71493 ( .A(n24232), .B(n8737), .X(n24233) );
  nand_x4_sg U71494 ( .A(n50224), .B(n24219), .X(n24218) );
  nor_x1_sg U71495 ( .A(n24220), .B(n8739), .X(n24221) );
  nand_x4_sg U71496 ( .A(n50408), .B(n24243), .X(n24242) );
  nor_x1_sg U71497 ( .A(n24244), .B(n8735), .X(n24245) );
  nand_x4_sg U71498 ( .A(n50908), .B(n22868), .X(n22776) );
  nor_x1_sg U71499 ( .A(n22612), .B(n8564), .X(n22869) );
  nand_x4_sg U71500 ( .A(n50049), .B(n30534), .X(n30442) );
  nor_x1_sg U71501 ( .A(n30278), .B(n8264), .X(n30535) );
  nand_x4_sg U71502 ( .A(n50860), .B(n22771), .X(n22770) );
  nor_x1_sg U71503 ( .A(n22772), .B(n8565), .X(n22773) );
  nand_x4_sg U71504 ( .A(n49957), .B(n30431), .X(n30430) );
  nor_x1_sg U71505 ( .A(n30432), .B(n8266), .X(n30433) );
  nand_x4_sg U71506 ( .A(n50343), .B(n22705), .X(n22704) );
  nor_x1_sg U71507 ( .A(n22706), .B(n8576), .X(n22707) );
  nand_x4_sg U71508 ( .A(n50360), .B(n24237), .X(n24236) );
  nor_x1_sg U71509 ( .A(n24238), .B(n8736), .X(n24239) );
  nand_x4_sg U71510 ( .A(n50269), .B(n24225), .X(n24224) );
  nor_x1_sg U71511 ( .A(n24226), .B(n8738), .X(n24227) );
  nand_x4_sg U71512 ( .A(n49501), .B(n31903), .X(n31902) );
  nor_x1_sg U71513 ( .A(n31904), .B(n8436), .X(n31905) );
  nand_x4_sg U71514 ( .A(n49455), .B(n31897), .X(n31896) );
  nor_x1_sg U71515 ( .A(n31898), .B(n8437), .X(n31899) );
  nand_x4_sg U71516 ( .A(n49410), .B(n31891), .X(n31890) );
  nor_x1_sg U71517 ( .A(n31892), .B(n8438), .X(n31893) );
  nand_x4_sg U71518 ( .A(n50543), .B(n23983), .X(n23982) );
  nor_x1_sg U71519 ( .A(n23984), .B(n8692), .X(n23985) );
  nand_x4_sg U71520 ( .A(n50355), .B(n23959), .X(n23958) );
  nor_x1_sg U71521 ( .A(n23960), .B(n8696), .X(n23961) );
  nand_x4_sg U71522 ( .A(n50264), .B(n23947), .X(n23946) );
  nor_x1_sg U71523 ( .A(n23948), .B(n8698), .X(n23949) );
  nand_x4_sg U71524 ( .A(n50219), .B(n23941), .X(n23940) );
  nor_x1_sg U71525 ( .A(n23942), .B(n8699), .X(n23943) );
  nand_x4_sg U71526 ( .A(n50852), .B(n9461), .X(n9460) );
  nor_x1_sg U71527 ( .A(n9462), .B(n8485), .X(n9463) );
  nand_x4_sg U71528 ( .A(n50807), .B(n9510), .X(n9509) );
  nor_x1_sg U71529 ( .A(n9511), .B(n8486), .X(n9512) );
  nand_x4_sg U71530 ( .A(n50768), .B(n22759), .X(n22758) );
  nor_x1_sg U71531 ( .A(n22760), .B(n8567), .X(n22761) );
  nand_x4_sg U71532 ( .A(n50759), .B(n9559), .X(n9558) );
  nor_x1_sg U71533 ( .A(n9560), .B(n8487), .X(n9561) );
  nand_x4_sg U71534 ( .A(n50721), .B(n22753), .X(n22752) );
  nor_x1_sg U71535 ( .A(n22754), .B(n8568), .X(n22755) );
  nand_x4_sg U71536 ( .A(n50712), .B(n9607), .X(n9606) );
  nor_x1_sg U71537 ( .A(n9608), .B(n8488), .X(n9609) );
  nand_x4_sg U71538 ( .A(n50673), .B(n22747), .X(n22746) );
  nor_x1_sg U71539 ( .A(n22748), .B(n8569), .X(n22749) );
  nand_x4_sg U71540 ( .A(n50664), .B(n9655), .X(n9654) );
  nor_x1_sg U71541 ( .A(n9656), .B(n8489), .X(n9657) );
  nand_x4_sg U71542 ( .A(n50617), .B(n9702), .X(n9701) );
  nor_x1_sg U71543 ( .A(n9703), .B(n8490), .X(n9704) );
  nand_x4_sg U71544 ( .A(n50577), .B(n22735), .X(n22734) );
  nor_x1_sg U71545 ( .A(n22736), .B(n8571), .X(n22737) );
  nand_x4_sg U71546 ( .A(n50568), .B(n9750), .X(n9749) );
  nor_x1_sg U71547 ( .A(n9751), .B(n8491), .X(n9752) );
  nand_x4_sg U71548 ( .A(n50530), .B(n22729), .X(n22728) );
  nor_x1_sg U71549 ( .A(n22730), .B(n8572), .X(n22731) );
  nand_x4_sg U71550 ( .A(n50521), .B(n9798), .X(n9797) );
  nor_x1_sg U71551 ( .A(n9799), .B(n8492), .X(n9800) );
  nand_x4_sg U71552 ( .A(n50483), .B(n22723), .X(n22722) );
  nor_x1_sg U71553 ( .A(n22724), .B(n8573), .X(n22725) );
  nand_x4_sg U71554 ( .A(n50474), .B(n9846), .X(n9845) );
  nor_x1_sg U71555 ( .A(n9847), .B(n8493), .X(n9848) );
  nand_x4_sg U71556 ( .A(n50437), .B(n22717), .X(n22716) );
  nor_x1_sg U71557 ( .A(n22718), .B(n8574), .X(n22719) );
  nand_x4_sg U71558 ( .A(n50428), .B(n9894), .X(n9893) );
  nor_x1_sg U71559 ( .A(n9895), .B(n8494), .X(n9896) );
  nand_x4_sg U71560 ( .A(n50390), .B(n22711), .X(n22710) );
  nor_x1_sg U71561 ( .A(n22712), .B(n8575), .X(n22713) );
  nand_x4_sg U71562 ( .A(n50381), .B(n9942), .X(n9941) );
  nor_x1_sg U71563 ( .A(n9943), .B(n8495), .X(n9944) );
  nand_x4_sg U71564 ( .A(n50334), .B(n9991), .X(n9990) );
  nor_x1_sg U71565 ( .A(n9992), .B(n8496), .X(n9993) );
  nand_x4_sg U71566 ( .A(n50297), .B(n22699), .X(n22698) );
  nor_x1_sg U71567 ( .A(n22700), .B(n8577), .X(n22701) );
  nand_x4_sg U71568 ( .A(n50288), .B(n10039), .X(n10038) );
  nor_x1_sg U71569 ( .A(n10040), .B(n8497), .X(n10041) );
  nand_x4_sg U71570 ( .A(n50242), .B(n10088), .X(n10087) );
  nor_x1_sg U71571 ( .A(n10089), .B(n8498), .X(n10090) );
  nand_x4_sg U71572 ( .A(n50198), .B(n10137), .X(n10136) );
  nor_x1_sg U71573 ( .A(n10138), .B(n8499), .X(n10139) );
  nand_x4_sg U71574 ( .A(n49993), .B(n24569), .X(n24568) );
  nor_x1_sg U71575 ( .A(n24570), .B(n8185), .X(n24571) );
  nand_x4_sg U71576 ( .A(n49948), .B(n24618), .X(n24617) );
  nor_x1_sg U71577 ( .A(n24619), .B(n8186), .X(n24620) );
  nand_x4_sg U71578 ( .A(n49909), .B(n30425), .X(n30424) );
  nor_x1_sg U71579 ( .A(n30426), .B(n8267), .X(n30427) );
  nand_x4_sg U71580 ( .A(n49900), .B(n24667), .X(n24666) );
  nor_x1_sg U71581 ( .A(n24668), .B(n8187), .X(n24669) );
  nand_x4_sg U71582 ( .A(n49862), .B(n30419), .X(n30418) );
  nor_x1_sg U71583 ( .A(n30420), .B(n8268), .X(n30421) );
  nand_x4_sg U71584 ( .A(n49853), .B(n24715), .X(n24714) );
  nor_x1_sg U71585 ( .A(n24716), .B(n8188), .X(n24717) );
  nand_x4_sg U71586 ( .A(n49814), .B(n30413), .X(n30412) );
  nor_x1_sg U71587 ( .A(n30414), .B(n8269), .X(n30415) );
  nand_x4_sg U71588 ( .A(n49805), .B(n24763), .X(n24762) );
  nor_x1_sg U71589 ( .A(n24764), .B(n8189), .X(n24765) );
  nand_x4_sg U71590 ( .A(n49758), .B(n24810), .X(n24809) );
  nor_x1_sg U71591 ( .A(n24811), .B(n8190), .X(n24812) );
  nand_x4_sg U71592 ( .A(n49718), .B(n30401), .X(n30400) );
  nor_x1_sg U71593 ( .A(n30402), .B(n8271), .X(n30403) );
  nand_x4_sg U71594 ( .A(n49709), .B(n24858), .X(n24857) );
  nor_x1_sg U71595 ( .A(n24859), .B(n8191), .X(n24860) );
  nand_x4_sg U71596 ( .A(n49671), .B(n30395), .X(n30394) );
  nor_x1_sg U71597 ( .A(n30396), .B(n8272), .X(n30397) );
  nand_x4_sg U71598 ( .A(n49662), .B(n24906), .X(n24905) );
  nor_x1_sg U71599 ( .A(n24907), .B(n8192), .X(n24908) );
  nand_x4_sg U71600 ( .A(n49624), .B(n30389), .X(n30388) );
  nor_x1_sg U71601 ( .A(n30390), .B(n8273), .X(n30391) );
  nand_x4_sg U71602 ( .A(n49615), .B(n24954), .X(n24953) );
  nor_x1_sg U71603 ( .A(n24955), .B(n8193), .X(n24956) );
  nand_x4_sg U71604 ( .A(n49578), .B(n30383), .X(n30382) );
  nor_x1_sg U71605 ( .A(n30384), .B(n8274), .X(n30385) );
  nand_x4_sg U71606 ( .A(n49569), .B(n25002), .X(n25001) );
  nor_x1_sg U71607 ( .A(n25003), .B(n8194), .X(n25004) );
  nand_x4_sg U71608 ( .A(n49531), .B(n30377), .X(n30376) );
  nor_x1_sg U71609 ( .A(n30378), .B(n8275), .X(n30379) );
  nand_x4_sg U71610 ( .A(n49522), .B(n25050), .X(n25049) );
  nor_x1_sg U71611 ( .A(n25051), .B(n8195), .X(n25052) );
  nand_x4_sg U71612 ( .A(n49475), .B(n25099), .X(n25098) );
  nor_x1_sg U71613 ( .A(n25100), .B(n8196), .X(n25101) );
  nand_x4_sg U71614 ( .A(n49438), .B(n30365), .X(n30364) );
  nor_x1_sg U71615 ( .A(n30366), .B(n8277), .X(n30367) );
  nand_x4_sg U71616 ( .A(n49429), .B(n25147), .X(n25146) );
  nor_x1_sg U71617 ( .A(n25148), .B(n8197), .X(n25149) );
  nand_x4_sg U71618 ( .A(n49383), .B(n25196), .X(n25195) );
  nor_x1_sg U71619 ( .A(n25197), .B(n8198), .X(n25198) );
  nand_x4_sg U71620 ( .A(n49339), .B(n25245), .X(n25244) );
  nor_x1_sg U71621 ( .A(n25246), .B(n8199), .X(n25247) );
  nand_x4_sg U71622 ( .A(n50495), .B(n23977), .X(n23976) );
  nor_x1_sg U71623 ( .A(n23978), .B(n8693), .X(n23979) );
  nand_x4_sg U71624 ( .A(n50449), .B(n23971), .X(n23970) );
  nor_x1_sg U71625 ( .A(n23972), .B(n8694), .X(n23973) );
  nand_x4_sg U71626 ( .A(n50403), .B(n23965), .X(n23964) );
  nor_x1_sg U71627 ( .A(n23966), .B(n8695), .X(n23967) );
  nand_x4_sg U71628 ( .A(n50309), .B(n23953), .X(n23952) );
  nor_x1_sg U71629 ( .A(n23954), .B(n8697), .X(n23955) );
  nand_x4_sg U71630 ( .A(n49684), .B(n31649), .X(n31648) );
  nor_x1_sg U71631 ( .A(n31650), .B(n8392), .X(n31651) );
  nand_x4_sg U71632 ( .A(n49636), .B(n31643), .X(n31642) );
  nor_x1_sg U71633 ( .A(n31644), .B(n8393), .X(n31645) );
  nand_x4_sg U71634 ( .A(n49590), .B(n31637), .X(n31636) );
  nor_x1_sg U71635 ( .A(n31638), .B(n8394), .X(n31639) );
  nand_x4_sg U71636 ( .A(n49544), .B(n31631), .X(n31630) );
  nor_x1_sg U71637 ( .A(n31632), .B(n8395), .X(n31633) );
  nand_x4_sg U71638 ( .A(n49496), .B(n31625), .X(n31624) );
  nor_x1_sg U71639 ( .A(n31626), .B(n8396), .X(n31627) );
  nand_x4_sg U71640 ( .A(n49450), .B(n31619), .X(n31618) );
  nor_x1_sg U71641 ( .A(n31620), .B(n8397), .X(n31621) );
  nand_x4_sg U71642 ( .A(n49405), .B(n31613), .X(n31612) );
  nor_x1_sg U71643 ( .A(n31614), .B(n8398), .X(n31615) );
  nand_x4_sg U71644 ( .A(n49360), .B(n31607), .X(n31606) );
  nor_x1_sg U71645 ( .A(n31608), .B(n8399), .X(n31609) );
  nand_x4_sg U71646 ( .A(n50782), .B(n23301), .X(n23281) );
  nor_x1_sg U71647 ( .A(n23080), .B(n8726), .X(n23302) );
  nand_x4_sg U71648 ( .A(n50690), .B(n23696), .X(n23676) );
  nor_x1_sg U71649 ( .A(n23511), .B(n8728), .X(n23697) );
  nand_x4_sg U71650 ( .A(n50599), .B(n24020), .X(n24000) );
  nor_x1_sg U71651 ( .A(n23872), .B(n8730), .X(n24021) );
  nand_x4_sg U71652 ( .A(n50582), .B(n23234), .X(n23233) );
  nor_x1_sg U71653 ( .A(n23235), .B(n8611), .X(n23236) );
  nand_x4_sg U71654 ( .A(n50547), .B(n24280), .X(n24260) );
  nor_x1_sg U71655 ( .A(n24169), .B(n8732), .X(n24281) );
  nand_x4_sg U71656 ( .A(n50500), .B(n24255), .X(n24254) );
  nor_x1_sg U71657 ( .A(n24256), .B(n8733), .X(n24257) );
  nand_x4_sg U71658 ( .A(n50302), .B(n23198), .X(n23197) );
  nor_x1_sg U71659 ( .A(n23199), .B(n8617), .X(n23200) );
  nand_x4_sg U71660 ( .A(n50212), .B(n23186), .X(n23185) );
  nor_x1_sg U71661 ( .A(n23187), .B(n8619), .X(n23188) );
  nand_x4_sg U71662 ( .A(n49723), .B(n30900), .X(n30899) );
  nor_x1_sg U71663 ( .A(n30901), .B(n8311), .X(n30902) );
  nand_x4_sg U71664 ( .A(n49443), .B(n30864), .X(n30863) );
  nor_x1_sg U71665 ( .A(n30865), .B(n8317), .X(n30866) );
  nand_x4_sg U71666 ( .A(n49353), .B(n30852), .X(n30851) );
  nor_x1_sg U71667 ( .A(n30853), .B(n8319), .X(n30854) );
  nand_x4_sg U71668 ( .A(n50877), .B(n22833), .X(n22794) );
  nor_x1_sg U71669 ( .A(n22569), .B(n8684), .X(n22834) );
  nand_x4_sg U71670 ( .A(n50889), .B(n22856), .X(n22781) );
  nor_x1_sg U71671 ( .A(n22598), .B(n8604), .X(n22857) );
  nand_x4_sg U71672 ( .A(n50812), .B(n22339), .X(n22338) );
  nor_x1_sg U71673 ( .A(n22340), .B(n8526), .X(n22341) );
  nand_x4_sg U71674 ( .A(n50764), .B(n22333), .X(n22332) );
  nor_x1_sg U71675 ( .A(n22334), .B(n8527), .X(n22335) );
  nand_x4_sg U71676 ( .A(n50726), .B(n23252), .X(n23251) );
  nor_x1_sg U71677 ( .A(n23253), .B(n8608), .X(n23254) );
  nand_x4_sg U71678 ( .A(n50717), .B(n22327), .X(n22326) );
  nor_x1_sg U71679 ( .A(n22328), .B(n8528), .X(n22329) );
  nand_x4_sg U71680 ( .A(n50678), .B(n23246), .X(n23245) );
  nor_x1_sg U71681 ( .A(n23247), .B(n8609), .X(n23248) );
  nand_x4_sg U71682 ( .A(n50669), .B(n22321), .X(n22320) );
  nor_x1_sg U71683 ( .A(n22322), .B(n8529), .X(n22323) );
  nand_x4_sg U71684 ( .A(n50631), .B(n23240), .X(n23239) );
  nor_x1_sg U71685 ( .A(n23241), .B(n8610), .X(n23242) );
  nand_x4_sg U71686 ( .A(n50622), .B(n22315), .X(n22314) );
  nor_x1_sg U71687 ( .A(n22316), .B(n8530), .X(n22317) );
  nand_x4_sg U71688 ( .A(n50573), .B(n22309), .X(n22308) );
  nor_x1_sg U71689 ( .A(n22310), .B(n8531), .X(n22311) );
  nand_x4_sg U71690 ( .A(n50535), .B(n23228), .X(n23227) );
  nor_x1_sg U71691 ( .A(n23229), .B(n8612), .X(n23230) );
  nand_x4_sg U71692 ( .A(n50526), .B(n22303), .X(n22302) );
  nor_x1_sg U71693 ( .A(n22304), .B(n8532), .X(n22305) );
  nand_x4_sg U71694 ( .A(n50488), .B(n23222), .X(n23221) );
  nor_x1_sg U71695 ( .A(n23223), .B(n8613), .X(n23224) );
  nand_x4_sg U71696 ( .A(n50479), .B(n22297), .X(n22296) );
  nor_x1_sg U71697 ( .A(n22298), .B(n8533), .X(n22299) );
  nand_x4_sg U71698 ( .A(n50442), .B(n23216), .X(n23215) );
  nor_x1_sg U71699 ( .A(n23217), .B(n8614), .X(n23218) );
  nand_x4_sg U71700 ( .A(n50433), .B(n22291), .X(n22290) );
  nor_x1_sg U71701 ( .A(n22292), .B(n8534), .X(n22293) );
  nand_x4_sg U71702 ( .A(n50395), .B(n23210), .X(n23209) );
  nor_x1_sg U71703 ( .A(n23211), .B(n8615), .X(n23212) );
  nand_x4_sg U71704 ( .A(n50386), .B(n22285), .X(n22284) );
  nor_x1_sg U71705 ( .A(n22286), .B(n8535), .X(n22287) );
  nand_x4_sg U71706 ( .A(n50348), .B(n23204), .X(n23203) );
  nor_x1_sg U71707 ( .A(n23205), .B(n8616), .X(n23206) );
  nand_x4_sg U71708 ( .A(n50339), .B(n22279), .X(n22278) );
  nor_x1_sg U71709 ( .A(n22280), .B(n8536), .X(n22281) );
  nand_x4_sg U71710 ( .A(n50293), .B(n22273), .X(n22272) );
  nor_x1_sg U71711 ( .A(n22274), .B(n8537), .X(n22275) );
  nand_x4_sg U71712 ( .A(n50256), .B(n23192), .X(n23191) );
  nor_x1_sg U71713 ( .A(n23193), .B(n8618), .X(n23194) );
  nand_x4_sg U71714 ( .A(n50247), .B(n22267), .X(n22266) );
  nor_x1_sg U71715 ( .A(n22268), .B(n8538), .X(n22269) );
  nand_x4_sg U71716 ( .A(n50203), .B(n22261), .X(n22260) );
  nor_x1_sg U71717 ( .A(n22262), .B(n8539), .X(n22263) );
  nand_x4_sg U71718 ( .A(n50030), .B(n30522), .X(n30447) );
  nor_x1_sg U71719 ( .A(n30264), .B(n8304), .X(n30523) );
  nand_x4_sg U71720 ( .A(n49953), .B(n30004), .X(n30003) );
  nor_x1_sg U71721 ( .A(n30005), .B(n8226), .X(n30006) );
  nand_x4_sg U71722 ( .A(n49905), .B(n29998), .X(n29997) );
  nor_x1_sg U71723 ( .A(n29999), .B(n8227), .X(n30000) );
  nand_x4_sg U71724 ( .A(n49867), .B(n30918), .X(n30917) );
  nor_x1_sg U71725 ( .A(n30919), .B(n8308), .X(n30920) );
  nand_x4_sg U71726 ( .A(n49858), .B(n29992), .X(n29991) );
  nor_x1_sg U71727 ( .A(n29993), .B(n8228), .X(n29994) );
  nand_x4_sg U71728 ( .A(n49819), .B(n30912), .X(n30911) );
  nor_x1_sg U71729 ( .A(n30913), .B(n8309), .X(n30914) );
  nand_x4_sg U71730 ( .A(n49810), .B(n29986), .X(n29985) );
  nor_x1_sg U71731 ( .A(n29987), .B(n8229), .X(n29988) );
  nand_x4_sg U71732 ( .A(n49772), .B(n30906), .X(n30905) );
  nor_x1_sg U71733 ( .A(n30907), .B(n8310), .X(n30908) );
  nand_x4_sg U71734 ( .A(n49763), .B(n29980), .X(n29979) );
  nor_x1_sg U71735 ( .A(n29981), .B(n8230), .X(n29982) );
  nand_x4_sg U71736 ( .A(n49714), .B(n29974), .X(n29973) );
  nor_x1_sg U71737 ( .A(n29975), .B(n8231), .X(n29976) );
  nand_x4_sg U71738 ( .A(n49676), .B(n30894), .X(n30893) );
  nor_x1_sg U71739 ( .A(n30895), .B(n8312), .X(n30896) );
  nand_x4_sg U71740 ( .A(n49667), .B(n29968), .X(n29967) );
  nor_x1_sg U71741 ( .A(n29969), .B(n8232), .X(n29970) );
  nand_x4_sg U71742 ( .A(n49629), .B(n30888), .X(n30887) );
  nor_x1_sg U71743 ( .A(n30889), .B(n8313), .X(n30890) );
  nand_x4_sg U71744 ( .A(n49620), .B(n29962), .X(n29961) );
  nor_x1_sg U71745 ( .A(n29963), .B(n8233), .X(n29964) );
  nand_x4_sg U71746 ( .A(n49583), .B(n30882), .X(n30881) );
  nor_x1_sg U71747 ( .A(n30883), .B(n8314), .X(n30884) );
  nand_x4_sg U71748 ( .A(n49574), .B(n29956), .X(n29955) );
  nor_x1_sg U71749 ( .A(n29957), .B(n8234), .X(n29958) );
  nand_x4_sg U71750 ( .A(n49536), .B(n30876), .X(n30875) );
  nor_x1_sg U71751 ( .A(n30877), .B(n8315), .X(n30878) );
  nand_x4_sg U71752 ( .A(n49527), .B(n29950), .X(n29949) );
  nor_x1_sg U71753 ( .A(n29951), .B(n8235), .X(n29952) );
  nand_x4_sg U71754 ( .A(n49489), .B(n30870), .X(n30869) );
  nor_x1_sg U71755 ( .A(n30871), .B(n8316), .X(n30872) );
  nand_x4_sg U71756 ( .A(n49480), .B(n29944), .X(n29943) );
  nor_x1_sg U71757 ( .A(n29945), .B(n8236), .X(n29946) );
  nand_x4_sg U71758 ( .A(n49434), .B(n29938), .X(n29937) );
  nor_x1_sg U71759 ( .A(n29939), .B(n8237), .X(n29940) );
  nand_x4_sg U71760 ( .A(n49397), .B(n30858), .X(n30857) );
  nor_x1_sg U71761 ( .A(n30859), .B(n8318), .X(n30860) );
  nand_x4_sg U71762 ( .A(n49388), .B(n29932), .X(n29931) );
  nor_x1_sg U71763 ( .A(n29933), .B(n8238), .X(n29934) );
  nand_x4_sg U71764 ( .A(n49344), .B(n29926), .X(n29925) );
  nor_x1_sg U71765 ( .A(n29927), .B(n8239), .X(n29928) );
  nand_x4_sg U71766 ( .A(n50856), .B(n22351), .X(n22344) );
  nor_x1_sg U71767 ( .A(n22190), .B(n8525), .X(n22352) );
  nand_x4_sg U71768 ( .A(n49997), .B(n30016), .X(n30009) );
  nor_x1_sg U71769 ( .A(n29855), .B(n8225), .X(n30017) );
  nand_x4_sg U71770 ( .A(n50870), .B(n22820), .X(n22800) );
  nor_x1_sg U71771 ( .A(n22554), .B(n8724), .X(n22821) );
  nand_x4_sg U71772 ( .A(n50826), .B(n23075), .X(n23055) );
  nor_x1_sg U71773 ( .A(n22825), .B(n8725), .X(n23076) );
  nand_x4_sg U71774 ( .A(n50736), .B(n23506), .X(n23486) );
  nor_x1_sg U71775 ( .A(n23306), .B(n8727), .X(n23507) );
  nand_x4_sg U71776 ( .A(n50645), .B(n23867), .X(n23847) );
  nor_x1_sg U71777 ( .A(n23701), .B(n8729), .X(n23868) );
  nand_x4_sg U71778 ( .A(n50553), .B(n24164), .X(n24144) );
  nor_x1_sg U71779 ( .A(n24025), .B(n8731), .X(n24165) );
  nand_x4_sg U71780 ( .A(n50454), .B(n24249), .X(n24248) );
  nor_x1_sg U71781 ( .A(n24250), .B(n8734), .X(n24251) );
  nand_x4_sg U71782 ( .A(n49688), .B(n31946), .X(n31926) );
  nor_x1_sg U71783 ( .A(n31835), .B(n8432), .X(n31947) );
  nand_x4_sg U71784 ( .A(n49641), .B(n31921), .X(n31920) );
  nor_x1_sg U71785 ( .A(n31922), .B(n8433), .X(n31923) );
  nand_x4_sg U71786 ( .A(n49595), .B(n31915), .X(n31914) );
  nor_x1_sg U71787 ( .A(n31916), .B(n8434), .X(n31917) );
  nand_x4_sg U71788 ( .A(n49549), .B(n31909), .X(n31908) );
  nor_x1_sg U71789 ( .A(n31910), .B(n8435), .X(n31911) );
  nand_x4_sg U71790 ( .A(n49365), .B(n31885), .X(n31884) );
  nor_x1_sg U71791 ( .A(n31886), .B(n8439), .X(n31887) );
  nand_x4_sg U71792 ( .A(n50789), .B(n23314), .X(n23275) );
  nor_x1_sg U71793 ( .A(n23093), .B(n8686), .X(n23315) );
  nand_x4_sg U71794 ( .A(n50697), .B(n23709), .X(n23670) );
  nor_x1_sg U71795 ( .A(n23524), .B(n8688), .X(n23710) );
  nand_x4_sg U71796 ( .A(n50639), .B(n24033), .X(n23994) );
  nor_x1_sg U71797 ( .A(n23885), .B(n8690), .X(n24034) );
  nand_x4_sg U71798 ( .A(n50896), .B(n22185), .X(n22177) );
  nor_x1_sg U71799 ( .A(n21988), .B(n8524), .X(n22186) );
  nand_x4_sg U71800 ( .A(n50037), .B(n29850), .X(n29842) );
  nor_x1_sg U71801 ( .A(n29653), .B(n8224), .X(n29851) );
  nand_x4_sg U71802 ( .A(n50011), .B(n30486), .X(n30466) );
  nor_x1_sg U71803 ( .A(n30220), .B(n8424), .X(n30487) );
  nand_x4_sg U71804 ( .A(n49967), .B(n30741), .X(n30721) );
  nor_x1_sg U71805 ( .A(n30491), .B(n8425), .X(n30742) );
  nand_x4_sg U71806 ( .A(n49923), .B(n30967), .X(n30947) );
  nor_x1_sg U71807 ( .A(n30746), .B(n8426), .X(n30968) );
  nand_x4_sg U71808 ( .A(n49877), .B(n31172), .X(n31152) );
  nor_x1_sg U71809 ( .A(n30972), .B(n8427), .X(n31173) );
  nand_x4_sg U71810 ( .A(n49831), .B(n31362), .X(n31342) );
  nor_x1_sg U71811 ( .A(n31177), .B(n8428), .X(n31363) );
  nand_x4_sg U71812 ( .A(n49786), .B(n31533), .X(n31513) );
  nor_x1_sg U71813 ( .A(n31367), .B(n8429), .X(n31534) );
  nand_x4_sg U71814 ( .A(n49740), .B(n31686), .X(n31666) );
  nor_x1_sg U71815 ( .A(n31538), .B(n8430), .X(n31687) );
  nand_x4_sg U71816 ( .A(n49694), .B(n31830), .X(n31810) );
  nor_x1_sg U71817 ( .A(n31691), .B(n8431), .X(n31831) );
  nand_x4_sg U71818 ( .A(n50833), .B(n23088), .X(n23049) );
  nor_x1_sg U71819 ( .A(n22838), .B(n8685), .X(n23089) );
  nand_x4_sg U71820 ( .A(n50743), .B(n23519), .X(n23480) );
  nor_x1_sg U71821 ( .A(n23319), .B(n8687), .X(n23520) );
  nand_x4_sg U71822 ( .A(n50652), .B(n23880), .X(n23841) );
  nor_x1_sg U71823 ( .A(n23714), .B(n8689), .X(n23881) );
  nand_x4_sg U71824 ( .A(n50589), .B(n23989), .X(n23988) );
  nor_x1_sg U71825 ( .A(n23990), .B(n8691), .X(n23991) );
  nand_x4_sg U71826 ( .A(n50901), .B(n9411), .X(n9410) );
  nor_x1_sg U71827 ( .A(n9412), .B(n8484), .X(n9413) );
  nand_x4_sg U71828 ( .A(n50042), .B(n24520), .X(n24519) );
  nor_x1_sg U71829 ( .A(n24521), .B(n8184), .X(n24522) );
  nand_x4_sg U71830 ( .A(n50844), .B(n23113), .X(n23036) );
  nor_x1_sg U71831 ( .A(n22861), .B(n8605), .X(n23114) );
  nand_x4_sg U71832 ( .A(n50820), .B(n23337), .X(n23262) );
  nor_x1_sg U71833 ( .A(n23118), .B(n8606), .X(n23338) );
  nand_x4_sg U71834 ( .A(n50772), .B(n23258), .X(n23256) );
  nor_x1_sg U71835 ( .A(n23259), .B(n8607), .X(n23260) );
  nand_x4_sg U71836 ( .A(n49985), .B(n30779), .X(n30702) );
  nor_x1_sg U71837 ( .A(n30527), .B(n8305), .X(n30780) );
  nand_x4_sg U71838 ( .A(n49961), .B(n31003), .X(n30928) );
  nor_x1_sg U71839 ( .A(n30784), .B(n8306), .X(n31004) );
  nand_x4_sg U71840 ( .A(n49913), .B(n30924), .X(n30922) );
  nor_x1_sg U71841 ( .A(n30925), .B(n8307), .X(n30926) );
  nand_x4_sg U71842 ( .A(n50018), .B(n30499), .X(n30460) );
  nor_x1_sg U71843 ( .A(n30235), .B(n8384), .X(n30500) );
  nand_x4_sg U71844 ( .A(n49974), .B(n30754), .X(n30715) );
  nor_x1_sg U71845 ( .A(n30504), .B(n8385), .X(n30755) );
  nand_x4_sg U71846 ( .A(n49930), .B(n30980), .X(n30941) );
  nor_x1_sg U71847 ( .A(n30759), .B(n8386), .X(n30981) );
  nand_x4_sg U71848 ( .A(n49884), .B(n31185), .X(n31146) );
  nor_x1_sg U71849 ( .A(n30985), .B(n8387), .X(n31186) );
  nand_x4_sg U71850 ( .A(n49838), .B(n31375), .X(n31336) );
  nor_x1_sg U71851 ( .A(n31190), .B(n8388), .X(n31376) );
  nand_x4_sg U71852 ( .A(n49793), .B(n31546), .X(n31507) );
  nor_x1_sg U71853 ( .A(n31380), .B(n8389), .X(n31547) );
  nand_x4_sg U71854 ( .A(n49780), .B(n31699), .X(n31660) );
  nor_x1_sg U71855 ( .A(n31551), .B(n8390), .X(n31700) );
  nand_x4_sg U71856 ( .A(n49730), .B(n31655), .X(n31654) );
  nor_x1_sg U71857 ( .A(n31656), .B(n8391), .X(n31657) );
  nand_x4_sg U71858 ( .A(n50165), .B(n23180), .X(n23179) );
  nor_x1_sg U71859 ( .A(n23181), .B(n8620), .X(n23182) );
  nand_x4_sg U71860 ( .A(n49306), .B(n30846), .X(n30845) );
  nor_x1_sg U71861 ( .A(n30847), .B(n8320), .X(n30848) );
  nand_x4_sg U71862 ( .A(n50175), .B(n24213), .X(n24212) );
  nor_x1_sg U71863 ( .A(n24214), .B(n8740), .X(n24215) );
  nand_x4_sg U71864 ( .A(n50159), .B(n22255), .X(n22254) );
  nor_x1_sg U71865 ( .A(n22256), .B(n8540), .X(n22257) );
  nand_x4_sg U71866 ( .A(n49300), .B(n29920), .X(n29919) );
  nor_x1_sg U71867 ( .A(n29921), .B(n8240), .X(n29922) );
  nand_x4_sg U71868 ( .A(n49316), .B(n31879), .X(n31878) );
  nor_x1_sg U71869 ( .A(n31880), .B(n8440), .X(n31881) );
  nand_x4_sg U71870 ( .A(n49312), .B(n31601), .X(n31600) );
  nor_x1_sg U71871 ( .A(n31602), .B(n8400), .X(n31603) );
  nand_x4_sg U71872 ( .A(n50161), .B(n22681), .X(n22680) );
  nor_x1_sg U71873 ( .A(n22682), .B(n8580), .X(n22683) );
  nand_x4_sg U71874 ( .A(n49302), .B(n30347), .X(n30346) );
  nor_x1_sg U71875 ( .A(n30348), .B(n8280), .X(n30349) );
  nand_x4_sg U71876 ( .A(n50171), .B(n23935), .X(n23934) );
  nor_x1_sg U71877 ( .A(n23936), .B(n8700), .X(n23937) );
  nand_x4_sg U71878 ( .A(n50155), .B(n10184), .X(n10183) );
  nor_x1_sg U71879 ( .A(n10185), .B(n8500), .X(n10186) );
  nand_x4_sg U71880 ( .A(n49296), .B(n25292), .X(n25291) );
  nor_x1_sg U71881 ( .A(n25293), .B(n8200), .X(n25294) );
  nand_x4_sg U71882 ( .A(n50914), .B(n22548), .X(n22526) );
  nor_x1_sg U71883 ( .A(n22549), .B(n8723), .X(n22550) );
  nand_x4_sg U71884 ( .A(n50055), .B(n30214), .X(n30192) );
  nor_x1_sg U71885 ( .A(n30215), .B(n8423), .X(n30216) );
  nand_x4_sg U71886 ( .A(n50937), .B(n22606), .X(n22503) );
  nor_x1_sg U71887 ( .A(n22607), .B(n8563), .X(n22608) );
  nand_x4_sg U71888 ( .A(n50948), .B(n21996), .X(n21974) );
  nor_x1_sg U71889 ( .A(n21997), .B(n8483), .X(n21998) );
  nand_x4_sg U71890 ( .A(n50078), .B(n30272), .X(n30169) );
  nor_x1_sg U71891 ( .A(n30273), .B(n8263), .X(n30274) );
  nand_x4_sg U71892 ( .A(n50089), .B(n29661), .X(n29639) );
  nor_x1_sg U71893 ( .A(n29662), .B(n8183), .X(n29663) );
  nand_x4_sg U71894 ( .A(n50941), .B(n21982), .X(n21980) );
  nor_x1_sg U71895 ( .A(n21983), .B(n8523), .X(n21984) );
  nand_x4_sg U71896 ( .A(n50931), .B(n22592), .X(n22508) );
  nor_x1_sg U71897 ( .A(n22593), .B(n8603), .X(n22594) );
  nand_x4_sg U71898 ( .A(n50082), .B(n29647), .X(n29645) );
  nor_x1_sg U71899 ( .A(n29648), .B(n8223), .X(n29649) );
  nand_x4_sg U71900 ( .A(n50072), .B(n30258), .X(n30174) );
  nor_x1_sg U71901 ( .A(n30259), .B(n8303), .X(n30260) );
  nand_x4_sg U71902 ( .A(n50920), .B(n22563), .X(n22521) );
  nor_x1_sg U71903 ( .A(n22564), .B(n8683), .X(n22565) );
  nand_x4_sg U71904 ( .A(n50061), .B(n30229), .X(n30187) );
  nor_x1_sg U71905 ( .A(n30230), .B(n8383), .X(n30231) );
  nand_x4_sg U71906 ( .A(n50935), .B(n22599), .X(n22505) );
  nor_x1_sg U71907 ( .A(n22600), .B(n8583), .X(n22601) );
  nand_x4_sg U71908 ( .A(n50945), .B(n21989), .X(n21976) );
  nor_x1_sg U71909 ( .A(n21990), .B(n8503), .X(n21991) );
  nand_x4_sg U71910 ( .A(n50076), .B(n30265), .X(n30171) );
  nor_x1_sg U71911 ( .A(n30266), .B(n8283), .X(n30267) );
  nand_x4_sg U71912 ( .A(n50086), .B(n29654), .X(n29641) );
  nor_x1_sg U71913 ( .A(n29655), .B(n8203), .X(n29656) );
  nand_x4_sg U71914 ( .A(n50912), .B(n22541), .X(n22529) );
  nor_x1_sg U71915 ( .A(n22542), .B(n8743), .X(n22543) );
  nand_x4_sg U71916 ( .A(n50053), .B(n30207), .X(n30195) );
  nor_x1_sg U71917 ( .A(n30208), .B(n8443), .X(n30209) );
  nand_x4_sg U71918 ( .A(n49400), .B(n31420), .X(n31273) );
  nand_x1_sg U71919 ( .A(n49356), .B(n25238), .X(n31421) );
  nand_x4_sg U71920 ( .A(n50259), .B(n23754), .X(n23607) );
  nand_x1_sg U71921 ( .A(n50215), .B(n10130), .X(n23755) );
  nand_x4_sg U71922 ( .A(n50918), .B(n22555), .X(n22523) );
  nor_x1_sg U71923 ( .A(n22556), .B(n8703), .X(n22557) );
  nand_x4_sg U71924 ( .A(n50059), .B(n30221), .X(n30189) );
  nor_x1_sg U71925 ( .A(n30222), .B(n8403), .X(n30223) );
  nand_x4_sg U71926 ( .A(n31392), .B(n31393), .X(n31327) );
  nand_x1_sg U71927 ( .A(n43179), .B(n41151), .X(n31392) );
  nand_x1_sg U71928 ( .A(n31321), .B(n49796), .X(n31394) );
  nand_x4_sg U71929 ( .A(n23726), .B(n23727), .X(n23661) );
  nand_x1_sg U71930 ( .A(n43191), .B(n41203), .X(n23726) );
  nand_x1_sg U71931 ( .A(n23655), .B(n50655), .X(n23728) );
  nand_x4_sg U71932 ( .A(n30769), .B(n30770), .X(n30768) );
  nand_x1_sg U71933 ( .A(n49979), .B(n49936), .X(n30769) );
  nand_x1_sg U71934 ( .A(n30772), .B(n24611), .X(n30771) );
  nand_x4_sg U71935 ( .A(n31200), .B(n31201), .X(n31199) );
  nand_x1_sg U71936 ( .A(n49889), .B(n49871), .X(n31200) );
  nand_x1_sg U71937 ( .A(n31203), .B(n24708), .X(n31202) );
  nand_x4_sg U71938 ( .A(n23103), .B(n23104), .X(n23102) );
  nand_x1_sg U71939 ( .A(n50838), .B(n50795), .X(n23103) );
  nand_x1_sg U71940 ( .A(n23106), .B(n9503), .X(n23105) );
  nand_x4_sg U71941 ( .A(n23534), .B(n23535), .X(n23533) );
  nand_x1_sg U71942 ( .A(n50748), .B(n50730), .X(n23534) );
  nand_x1_sg U71943 ( .A(n23537), .B(n9600), .X(n23536) );
  nand_x4_sg U71944 ( .A(n22616), .B(n22617), .X(n22615) );
  nand_x4_sg U71945 ( .A(n30282), .B(n30283), .X(n30281) );
  nand_x4_sg U71946 ( .A(n22573), .B(n22574), .X(n22572) );
  nand_x4_sg U71947 ( .A(n30239), .B(n30240), .X(n30238) );
  nand_x1_sg U71948 ( .A(n8501), .B(n50125), .X(n10229) );
  nand_x1_sg U71949 ( .A(n10230), .B(n40839), .X(n10228) );
  nand_x1_sg U71950 ( .A(n8201), .B(n49266), .X(n25337) );
  nand_x1_sg U71951 ( .A(n25338), .B(n40840), .X(n25336) );
  nand_x4_sg U71952 ( .A(n22588), .B(n22589), .X(n22587) );
  nand_x4_sg U71953 ( .A(n30254), .B(n30255), .X(n30253) );
  nand_x4_sg U71954 ( .A(n22558), .B(n22559), .X(n22556) );
  nand_x4_sg U71955 ( .A(n30224), .B(n30225), .X(n30222) );
  nand_x4_sg U71956 ( .A(n24436), .B(n24437), .X(n24434) );
  nand_x1_sg U71957 ( .A(out_L2[6]), .B(n40851), .X(n24437) );
  nand_x4_sg U71958 ( .A(n32102), .B(n32103), .X(n32100) );
  nand_x1_sg U71959 ( .A(out_L1[6]), .B(n40852), .X(n32103) );
  nand_x4_sg U71960 ( .A(n22811), .B(n22812), .X(n22806) );
  nand_x1_sg U71961 ( .A(n8764), .B(n40739), .X(n22811) );
  nand_x1_sg U71962 ( .A(out_L2[18]), .B(n40740), .X(n22812) );
  nand_x4_sg U71963 ( .A(n30477), .B(n30478), .X(n30472) );
  nand_x1_sg U71964 ( .A(n8464), .B(n40741), .X(n30477) );
  nand_x1_sg U71965 ( .A(out_L1[18]), .B(n40742), .X(n30478) );
  nand_x4_sg U71966 ( .A(n24468), .B(n24469), .X(n24446) );
  nand_x4_sg U71967 ( .A(n32134), .B(n32135), .X(n32112) );
  nand_x4_sg U71968 ( .A(n22539), .B(n22540), .X(n22533) );
  nand_x4_sg U71969 ( .A(n30205), .B(n30206), .X(n30199) );
  nand_x1_sg U71970 ( .A(n8766), .B(n40727), .X(n23292) );
  nand_x1_sg U71971 ( .A(out_L2[16]), .B(n40743), .X(n23293) );
  nand_x1_sg U71972 ( .A(n8768), .B(n40728), .X(n23687) );
  nand_x1_sg U71973 ( .A(out_L2[14]), .B(n40744), .X(n23688) );
  nand_x1_sg U71974 ( .A(n8770), .B(n40729), .X(n24011) );
  nand_x1_sg U71975 ( .A(out_L2[12]), .B(n40745), .X(n24012) );
  nand_x1_sg U71976 ( .A(n8772), .B(n40730), .X(n24271) );
  nand_x1_sg U71977 ( .A(out_L2[10]), .B(n40746), .X(n24272) );
  nand_x1_sg U71978 ( .A(n8472), .B(n40731), .X(n31937) );
  nand_x1_sg U71979 ( .A(out_L1[10]), .B(n40747), .X(n31938) );
  nand_x1_sg U71980 ( .A(n8781), .B(n40732), .X(n24406) );
  nand_x1_sg U71981 ( .A(out_L2[1]), .B(n40748), .X(n24407) );
  nand_x1_sg U71982 ( .A(n8466), .B(n40733), .X(n30958) );
  nand_x1_sg U71983 ( .A(out_L1[16]), .B(n40749), .X(n30959) );
  nand_x1_sg U71984 ( .A(n8468), .B(n40734), .X(n31353) );
  nand_x1_sg U71985 ( .A(out_L1[14]), .B(n40750), .X(n31354) );
  nand_x1_sg U71986 ( .A(n8470), .B(n40735), .X(n31677) );
  nand_x1_sg U71987 ( .A(out_L1[12]), .B(n40751), .X(n31678) );
  nand_x1_sg U71988 ( .A(n8481), .B(n40736), .X(n32072) );
  nand_x1_sg U71989 ( .A(out_L1[1]), .B(n40752), .X(n32073) );
  inv_x8_sg U71990 ( .A(n44160), .X(n46203) );
  inv_x8_sg U71991 ( .A(n46203), .X(n46204) );
  inv_x8_sg U71992 ( .A(n43788), .X(n46205) );
  inv_x8_sg U71993 ( .A(n46205), .X(n46206) );
  inv_x8_sg U71994 ( .A(n43852), .X(n46207) );
  inv_x8_sg U71995 ( .A(n46207), .X(n46208) );
  inv_x8_sg U71996 ( .A(n44162), .X(n46209) );
  inv_x8_sg U71997 ( .A(n46209), .X(n46210) );
  inv_x8_sg U71998 ( .A(n43807), .X(n46211) );
  inv_x8_sg U71999 ( .A(n46211), .X(n46212) );
  inv_x8_sg U72000 ( .A(n43767), .X(n46213) );
  inv_x8_sg U72001 ( .A(n46213), .X(n46214) );
  inv_x8_sg U72002 ( .A(n43854), .X(n46215) );
  inv_x8_sg U72003 ( .A(n46215), .X(n46216) );
  inv_x8_sg U72004 ( .A(n44164), .X(n46217) );
  inv_x8_sg U72005 ( .A(n46217), .X(n46218) );
  inv_x8_sg U72006 ( .A(n43790), .X(n46219) );
  inv_x8_sg U72007 ( .A(n46219), .X(n46220) );
  inv_x8_sg U72008 ( .A(n43786), .X(n46221) );
  inv_x8_sg U72009 ( .A(n46221), .X(n46222) );
  inv_x8_sg U72010 ( .A(n43809), .X(n46223) );
  inv_x8_sg U72011 ( .A(n46223), .X(n46224) );
  inv_x8_sg U72012 ( .A(n43792), .X(n46225) );
  inv_x8_sg U72013 ( .A(n46225), .X(n46226) );
  inv_x8_sg U72014 ( .A(n44168), .X(n46227) );
  inv_x8_sg U72015 ( .A(n46227), .X(n46228) );
  inv_x8_sg U72016 ( .A(n44166), .X(n46229) );
  inv_x8_sg U72017 ( .A(n46229), .X(n46230) );
  inv_x8_sg U72018 ( .A(n44158), .X(n46231) );
  inv_x8_sg U72019 ( .A(n46231), .X(n46232) );
  nand_x8_sg U72020 ( .A(n46235), .B(n25388), .X(n46233) );
  nand_x8_sg U72021 ( .A(n46235), .B(n25388), .X(n46234) );
  inv_x8_sg U72022 ( .A(n25394), .X(n46235) );
  inv_x8_sg U72023 ( .A(n46235), .X(n46236) );
  nand_x8_sg U72024 ( .A(n25388), .B(n46236), .X(n46237) );
  nand_x8_sg U72025 ( .A(n25388), .B(n46236), .X(n46238) );
  inv_x8_sg U72026 ( .A(n46239), .X(n46240) );
  inv_x8_sg U72027 ( .A(n21527), .X(n55256) );
  inv_x8_sg U72028 ( .A(n21391), .X(n46241) );
  inv_x8_sg U72029 ( .A(n46241), .X(n46242) );
  inv_x8_sg U72030 ( .A(n46243), .X(n46244) );
  inv_x8_sg U72031 ( .A(n46244), .X(n55228) );
  inv_x8_sg U72032 ( .A(n46245), .X(n46246) );
  inv_x8_sg U72033 ( .A(n46246), .X(n55215) );
  inv_x8_sg U72034 ( .A(n46247), .X(n46248) );
  inv_x8_sg U72035 ( .A(n46248), .X(n55202) );
  inv_x8_sg U72036 ( .A(n21280), .X(n46249) );
  inv_x8_sg U72037 ( .A(n46249), .X(n46250) );
  inv_x8_sg U72038 ( .A(n21269), .X(n46251) );
  inv_x8_sg U72039 ( .A(n46251), .X(n46252) );
  inv_x8_sg U72040 ( .A(n46253), .X(n46254) );
  inv_x8_sg U72041 ( .A(n46254), .X(n55182) );
  inv_x8_sg U72042 ( .A(n21155), .X(n46255) );
  inv_x8_sg U72043 ( .A(n46255), .X(n46256) );
  inv_x8_sg U72044 ( .A(n46257), .X(n46258) );
  inv_x8_sg U72045 ( .A(n46259), .X(n46260) );
  inv_x8_sg U72046 ( .A(n46260), .X(n46261) );
  inv_x8_sg U72047 ( .A(n46262), .X(n46263) );
  inv_x8_sg U72048 ( .A(n20757), .X(n46264) );
  inv_x8_sg U72049 ( .A(n46266), .X(n54947) );
  inv_x8_sg U72050 ( .A(n20613), .X(n54960) );
  inv_x8_sg U72051 ( .A(n46265), .X(n46266) );
  inv_x8_sg U72052 ( .A(n46268), .X(n54921) );
  inv_x8_sg U72053 ( .A(n20685), .X(n54935) );
  inv_x8_sg U72054 ( .A(n46267), .X(n46268) );
  inv_x8_sg U72055 ( .A(n20506), .X(n46269) );
  inv_x8_sg U72056 ( .A(n46269), .X(n46270) );
  inv_x8_sg U72057 ( .A(n46274), .X(n54898) );
  inv_x8_sg U72058 ( .A(n20497), .X(n46271) );
  inv_x8_sg U72059 ( .A(n46271), .X(n46272) );
  inv_x8_sg U72060 ( .A(n46273), .X(n46274) );
  inv_x8_sg U72061 ( .A(n20382), .X(n46275) );
  inv_x8_sg U72062 ( .A(n46275), .X(n46276) );
  inv_x8_sg U72063 ( .A(n46277), .X(n46278) );
  inv_x8_sg U72064 ( .A(n46279), .X(n46280) );
  inv_x8_sg U72065 ( .A(n46280), .X(n46281) );
  inv_x8_sg U72066 ( .A(n46282), .X(n46283) );
  inv_x8_sg U72067 ( .A(n46284), .X(n46285) );
  inv_x8_sg U72068 ( .A(n19982), .X(n54688) );
  inv_x8_sg U72069 ( .A(n19846), .X(n46286) );
  inv_x8_sg U72070 ( .A(n46286), .X(n46287) );
  inv_x8_sg U72071 ( .A(n46288), .X(n46289) );
  inv_x8_sg U72072 ( .A(n46289), .X(n54660) );
  inv_x8_sg U72073 ( .A(n46290), .X(n46291) );
  inv_x8_sg U72074 ( .A(n46291), .X(n54647) );
  inv_x8_sg U72075 ( .A(n46292), .X(n46293) );
  inv_x8_sg U72076 ( .A(n46293), .X(n54634) );
  inv_x8_sg U72077 ( .A(n19735), .X(n46294) );
  inv_x8_sg U72078 ( .A(n46294), .X(n46295) );
  inv_x8_sg U72079 ( .A(n19724), .X(n46296) );
  inv_x8_sg U72080 ( .A(n46296), .X(n46297) );
  inv_x8_sg U72081 ( .A(n46298), .X(n46299) );
  inv_x8_sg U72082 ( .A(n46299), .X(n54614) );
  inv_x8_sg U72083 ( .A(n19610), .X(n46300) );
  inv_x8_sg U72084 ( .A(n46300), .X(n46301) );
  inv_x8_sg U72085 ( .A(n46302), .X(n46303) );
  inv_x8_sg U72086 ( .A(n46304), .X(n46305) );
  inv_x8_sg U72087 ( .A(n46305), .X(n46306) );
  inv_x8_sg U72088 ( .A(n46307), .X(n46308) );
  inv_x8_sg U72089 ( .A(n19213), .X(n46309) );
  inv_x8_sg U72090 ( .A(n46311), .X(n54379) );
  inv_x8_sg U72091 ( .A(n19069), .X(n54392) );
  inv_x8_sg U72092 ( .A(n46310), .X(n46311) );
  inv_x8_sg U72093 ( .A(n46313), .X(n54353) );
  inv_x8_sg U72094 ( .A(n19141), .X(n54367) );
  inv_x8_sg U72095 ( .A(n46312), .X(n46313) );
  inv_x8_sg U72096 ( .A(n18962), .X(n46314) );
  inv_x8_sg U72097 ( .A(n46314), .X(n46315) );
  inv_x8_sg U72098 ( .A(n46319), .X(n54330) );
  inv_x8_sg U72099 ( .A(n18953), .X(n46316) );
  inv_x8_sg U72100 ( .A(n46316), .X(n46317) );
  inv_x8_sg U72101 ( .A(n46318), .X(n46319) );
  inv_x8_sg U72102 ( .A(n18838), .X(n46320) );
  inv_x8_sg U72103 ( .A(n46320), .X(n46321) );
  inv_x8_sg U72104 ( .A(n46322), .X(n46323) );
  inv_x8_sg U72105 ( .A(n46324), .X(n46325) );
  inv_x8_sg U72106 ( .A(n46325), .X(n46326) );
  inv_x8_sg U72107 ( .A(n19608), .X(n46327) );
  inv_x8_sg U72108 ( .A(n46328), .X(n46329) );
  inv_x8_sg U72109 ( .A(n18437), .X(n54124) );
  inv_x8_sg U72110 ( .A(n46331), .X(n54109) );
  inv_x8_sg U72111 ( .A(n46330), .X(n46331) );
  inv_x8_sg U72112 ( .A(n46333), .X(n54097) );
  inv_x8_sg U72113 ( .A(n46332), .X(n46333) );
  inv_x8_sg U72114 ( .A(n46334), .X(n46335) );
  inv_x8_sg U72115 ( .A(n46335), .X(n54084) );
  inv_x8_sg U72116 ( .A(n46336), .X(n46337) );
  inv_x8_sg U72117 ( .A(n46337), .X(n54070) );
  inv_x8_sg U72118 ( .A(n46338), .X(n46339) );
  inv_x8_sg U72119 ( .A(n46339), .X(n46340) );
  inv_x8_sg U72120 ( .A(n46348), .X(n46341) );
  inv_x8_sg U72121 ( .A(n46342), .X(n46343) );
  inv_x8_sg U72122 ( .A(n46343), .X(n46344) );
  inv_x8_sg U72123 ( .A(n43858), .X(n46345) );
  inv_x8_sg U72124 ( .A(n46345), .X(n46346) );
  inv_x8_sg U72125 ( .A(n46347), .X(n46348) );
  inv_x8_sg U72126 ( .A(n46349), .X(n46350) );
  inv_x8_sg U72127 ( .A(n46351), .X(n46352) );
  inv_x8_sg U72128 ( .A(n46352), .X(n46353) );
  inv_x8_sg U72129 ( .A(n46354), .X(n46355) );
  inv_x8_sg U72130 ( .A(n17668), .X(n46356) );
  inv_x8_sg U72131 ( .A(n46358), .X(n53814) );
  inv_x8_sg U72132 ( .A(n17524), .X(n53827) );
  inv_x8_sg U72133 ( .A(n46357), .X(n46358) );
  inv_x8_sg U72134 ( .A(n46360), .X(n53788) );
  inv_x8_sg U72135 ( .A(n17596), .X(n53802) );
  inv_x8_sg U72136 ( .A(n46359), .X(n46360) );
  inv_x8_sg U72137 ( .A(n17417), .X(n46361) );
  inv_x8_sg U72138 ( .A(n46361), .X(n46362) );
  inv_x8_sg U72139 ( .A(n46366), .X(n53765) );
  inv_x8_sg U72140 ( .A(n17408), .X(n46363) );
  inv_x8_sg U72141 ( .A(n46363), .X(n46364) );
  inv_x8_sg U72142 ( .A(n46365), .X(n46366) );
  inv_x8_sg U72143 ( .A(n17293), .X(n46367) );
  inv_x8_sg U72144 ( .A(n46367), .X(n46368) );
  inv_x8_sg U72145 ( .A(n46369), .X(n46370) );
  inv_x8_sg U72146 ( .A(n46371), .X(n46372) );
  inv_x8_sg U72147 ( .A(n46372), .X(n46373) );
  inv_x8_sg U72148 ( .A(n46374), .X(n46375) );
  inv_x8_sg U72149 ( .A(n16854), .X(n53579) );
  inv_x8_sg U72150 ( .A(n16894), .X(n46376) );
  inv_x8_sg U72151 ( .A(n16725), .X(n46377) );
  inv_x8_sg U72152 ( .A(n46378), .X(n46379) );
  inv_x8_sg U72153 ( .A(n46379), .X(n53548) );
  inv_x8_sg U72154 ( .A(n46383), .X(n53509) );
  inv_x8_sg U72155 ( .A(n46380), .X(n46381) );
  inv_x8_sg U72156 ( .A(n46381), .X(n53525) );
  inv_x8_sg U72157 ( .A(n46382), .X(n46383) );
  inv_x8_sg U72158 ( .A(n46387), .X(n53492) );
  inv_x8_sg U72159 ( .A(n16633), .X(n46384) );
  inv_x8_sg U72160 ( .A(n46384), .X(n46385) );
  inv_x8_sg U72161 ( .A(n46386), .X(n46387) );
  inv_x8_sg U72162 ( .A(n43888), .X(n46388) );
  inv_x8_sg U72163 ( .A(n46388), .X(n46389) );
  inv_x8_sg U72164 ( .A(n16510), .X(n46390) );
  inv_x8_sg U72165 ( .A(n46390), .X(n46391) );
  inv_x8_sg U72166 ( .A(n46392), .X(n46393) );
  inv_x8_sg U72167 ( .A(n46394), .X(n46395) );
  inv_x8_sg U72168 ( .A(n46395), .X(n46396) );
  inv_x8_sg U72169 ( .A(n46397), .X(n46398) );
  inv_x8_sg U72170 ( .A(n16109), .X(n53282) );
  inv_x8_sg U72171 ( .A(n46399), .X(n46400) );
  inv_x8_sg U72172 ( .A(n46400), .X(n53266) );
  inv_x8_sg U72173 ( .A(n46401), .X(n46402) );
  inv_x8_sg U72174 ( .A(n46402), .X(n53253) );
  inv_x8_sg U72175 ( .A(n15925), .X(n53240) );
  inv_x8_sg U72176 ( .A(n46403), .X(n46404) );
  inv_x8_sg U72177 ( .A(n46404), .X(n53227) );
  inv_x8_sg U72178 ( .A(n15852), .X(n46405) );
  inv_x8_sg U72179 ( .A(n46405), .X(n46406) );
  inv_x8_sg U72180 ( .A(n46409), .X(n53214) );
  inv_x8_sg U72181 ( .A(n46413), .X(n46407) );
  inv_x8_sg U72182 ( .A(n46408), .X(n46409) );
  inv_x8_sg U72183 ( .A(n46410), .X(n46411) );
  inv_x8_sg U72184 ( .A(n46411), .X(n53207) );
  inv_x8_sg U72185 ( .A(n46412), .X(n46413) );
  inv_x8_sg U72186 ( .A(n46414), .X(n46415) );
  inv_x8_sg U72187 ( .A(n15847), .X(n46416) );
  inv_x8_sg U72188 ( .A(n46416), .X(n46417) );
  inv_x8_sg U72189 ( .A(n46418), .X(n46419) );
  inv_x8_sg U72190 ( .A(n15288), .X(n53021) );
  inv_x8_sg U72191 ( .A(n15328), .X(n46420) );
  inv_x8_sg U72192 ( .A(n15159), .X(n46421) );
  inv_x8_sg U72193 ( .A(n46422), .X(n46423) );
  inv_x8_sg U72194 ( .A(n46423), .X(n52990) );
  inv_x8_sg U72195 ( .A(n46427), .X(n52951) );
  inv_x8_sg U72196 ( .A(n46424), .X(n46425) );
  inv_x8_sg U72197 ( .A(n46425), .X(n52967) );
  inv_x8_sg U72198 ( .A(n46426), .X(n46427) );
  inv_x8_sg U72199 ( .A(n46431), .X(n52934) );
  inv_x8_sg U72200 ( .A(n15067), .X(n46428) );
  inv_x8_sg U72201 ( .A(n46428), .X(n46429) );
  inv_x8_sg U72202 ( .A(n46430), .X(n46431) );
  inv_x8_sg U72203 ( .A(n43892), .X(n46432) );
  inv_x8_sg U72204 ( .A(n46432), .X(n46433) );
  inv_x8_sg U72205 ( .A(n14944), .X(n46434) );
  inv_x8_sg U72206 ( .A(n46434), .X(n46435) );
  inv_x8_sg U72207 ( .A(n46436), .X(n46437) );
  inv_x8_sg U72208 ( .A(n46438), .X(n46439) );
  inv_x8_sg U72209 ( .A(n46439), .X(n46440) );
  inv_x8_sg U72210 ( .A(n46441), .X(n46442) );
  inv_x8_sg U72211 ( .A(n14547), .X(n46443) );
  inv_x8_sg U72212 ( .A(n14411), .X(n52707) );
  inv_x8_sg U72213 ( .A(n46444), .X(n46445) );
  inv_x8_sg U72214 ( .A(n46445), .X(n52695) );
  inv_x8_sg U72215 ( .A(n46446), .X(n46447) );
  inv_x8_sg U72216 ( .A(n46447), .X(n52683) );
  inv_x8_sg U72217 ( .A(n46448), .X(n46449) );
  inv_x8_sg U72218 ( .A(n46449), .X(n52670) );
  inv_x8_sg U72219 ( .A(n46454), .X(n52655) );
  inv_x8_sg U72220 ( .A(n14300), .X(n46450) );
  inv_x8_sg U72221 ( .A(n46450), .X(n46451) );
  inv_x8_sg U72222 ( .A(n46458), .X(n46452) );
  inv_x8_sg U72223 ( .A(n46453), .X(n46454) );
  inv_x8_sg U72224 ( .A(n46455), .X(n46456) );
  inv_x8_sg U72225 ( .A(n46456), .X(n52648) );
  inv_x8_sg U72226 ( .A(n46457), .X(n46458) );
  inv_x8_sg U72227 ( .A(n46459), .X(n46460) );
  inv_x8_sg U72228 ( .A(n46461), .X(n46462) );
  inv_x8_sg U72229 ( .A(n46462), .X(n46463) );
  inv_x8_sg U72230 ( .A(n46464), .X(n46465) );
  inv_x8_sg U72231 ( .A(n13735), .X(n52463) );
  inv_x8_sg U72232 ( .A(n13775), .X(n52447) );
  inv_x8_sg U72233 ( .A(n46466), .X(n46467) );
  inv_x8_sg U72234 ( .A(n46467), .X(n52430) );
  inv_x8_sg U72235 ( .A(n13604), .X(n46468) );
  inv_x8_sg U72236 ( .A(n46468), .X(n46469) );
  inv_x8_sg U72237 ( .A(n46470), .X(n46471) );
  inv_x8_sg U72238 ( .A(n46471), .X(n52406) );
  inv_x8_sg U72239 ( .A(n46472), .X(n46473) );
  inv_x8_sg U72240 ( .A(n46473), .X(n52391) );
  inv_x8_sg U72241 ( .A(n13518), .X(n46474) );
  inv_x8_sg U72242 ( .A(n46474), .X(n46475) );
  inv_x8_sg U72243 ( .A(n46477), .X(n52378) );
  inv_x8_sg U72244 ( .A(n46476), .X(n46477) );
  inv_x8_sg U72245 ( .A(n43884), .X(n46478) );
  inv_x8_sg U72246 ( .A(n46478), .X(n46479) );
  inv_x8_sg U72247 ( .A(n13395), .X(n46480) );
  inv_x8_sg U72248 ( .A(n46480), .X(n46481) );
  inv_x8_sg U72249 ( .A(n46482), .X(n46483) );
  inv_x8_sg U72250 ( .A(n44285), .X(n46484) );
  inv_x8_sg U72251 ( .A(n46484), .X(n46485) );
  inv_x8_sg U72252 ( .A(n46486), .X(n46487) );
  inv_x8_sg U72253 ( .A(n12955), .X(n52187) );
  inv_x8_sg U72254 ( .A(n12995), .X(n46488) );
  inv_x8_sg U72255 ( .A(n12826), .X(n46489) );
  inv_x8_sg U72256 ( .A(n46490), .X(n46491) );
  inv_x8_sg U72257 ( .A(n46491), .X(n52156) );
  inv_x8_sg U72258 ( .A(n46495), .X(n52117) );
  inv_x8_sg U72259 ( .A(n46492), .X(n46493) );
  inv_x8_sg U72260 ( .A(n46493), .X(n52133) );
  inv_x8_sg U72261 ( .A(n46494), .X(n46495) );
  inv_x8_sg U72262 ( .A(n46499), .X(n52100) );
  inv_x8_sg U72263 ( .A(n12734), .X(n46496) );
  inv_x8_sg U72264 ( .A(n46496), .X(n46497) );
  inv_x8_sg U72265 ( .A(n46498), .X(n46499) );
  inv_x8_sg U72266 ( .A(n43896), .X(n46500) );
  inv_x8_sg U72267 ( .A(n46500), .X(n46501) );
  inv_x8_sg U72268 ( .A(n12611), .X(n46502) );
  inv_x8_sg U72269 ( .A(n46502), .X(n46503) );
  inv_x8_sg U72270 ( .A(n46504), .X(n46505) );
  inv_x8_sg U72271 ( .A(n46506), .X(n46507) );
  inv_x8_sg U72272 ( .A(n46507), .X(n46508) );
  inv_x8_sg U72273 ( .A(n46509), .X(n46510) );
  inv_x8_sg U72274 ( .A(n12174), .X(n51911) );
  inv_x8_sg U72275 ( .A(n12214), .X(n51896) );
  inv_x8_sg U72276 ( .A(n46511), .X(n46512) );
  inv_x8_sg U72277 ( .A(n46512), .X(n51879) );
  inv_x8_sg U72278 ( .A(n12043), .X(n46513) );
  inv_x8_sg U72279 ( .A(n46513), .X(n46514) );
  inv_x8_sg U72280 ( .A(n12030), .X(n51854) );
  inv_x8_sg U72281 ( .A(n46515), .X(n46516) );
  inv_x8_sg U72282 ( .A(n46516), .X(n51839) );
  inv_x8_sg U72283 ( .A(n11957), .X(n46517) );
  inv_x8_sg U72284 ( .A(n46517), .X(n46518) );
  inv_x8_sg U72285 ( .A(n46521), .X(n51826) );
  inv_x8_sg U72286 ( .A(n46525), .X(n46519) );
  inv_x8_sg U72287 ( .A(n46520), .X(n46521) );
  inv_x8_sg U72288 ( .A(n46522), .X(n46523) );
  inv_x8_sg U72289 ( .A(n46523), .X(n51819) );
  inv_x8_sg U72290 ( .A(n46524), .X(n46525) );
  inv_x8_sg U72291 ( .A(n46526), .X(n46527) );
  inv_x8_sg U72292 ( .A(n11952), .X(n46528) );
  inv_x8_sg U72293 ( .A(n46528), .X(n46529) );
  inv_x8_sg U72294 ( .A(n46530), .X(n46531) );
  inv_x8_sg U72295 ( .A(n11394), .X(n51630) );
  inv_x8_sg U72296 ( .A(n11434), .X(n46532) );
  inv_x8_sg U72297 ( .A(n11265), .X(n46533) );
  inv_x8_sg U72298 ( .A(n46534), .X(n46535) );
  inv_x8_sg U72299 ( .A(n46535), .X(n51598) );
  inv_x8_sg U72300 ( .A(n46539), .X(n51560) );
  inv_x8_sg U72301 ( .A(n11240), .X(n46536) );
  inv_x8_sg U72302 ( .A(n46536), .X(n46537) );
  inv_x8_sg U72303 ( .A(n46538), .X(n46539) );
  inv_x8_sg U72304 ( .A(n46543), .X(n51543) );
  inv_x8_sg U72305 ( .A(n11173), .X(n46540) );
  inv_x8_sg U72306 ( .A(n46540), .X(n46541) );
  inv_x8_sg U72307 ( .A(n46542), .X(n46543) );
  inv_x8_sg U72308 ( .A(n46544), .X(n46545) );
  inv_x8_sg U72309 ( .A(n46545), .X(n51537) );
  inv_x8_sg U72310 ( .A(n11050), .X(n46546) );
  inv_x8_sg U72311 ( .A(n46546), .X(n46547) );
  inv_x8_sg U72312 ( .A(n46548), .X(n46549) );
  inv_x8_sg U72313 ( .A(n46550), .X(n46551) );
  inv_x8_sg U72314 ( .A(n46551), .X(n46552) );
  inv_x8_sg U72315 ( .A(n11831), .X(n46553) );
  inv_x8_sg U72316 ( .A(n46554), .X(n46555) );
  inv_x8_sg U72317 ( .A(n46556), .X(n46557) );
  inv_x8_sg U72318 ( .A(n10655), .X(n51334) );
  inv_x8_sg U72319 ( .A(n10519), .X(n46558) );
  inv_x8_sg U72320 ( .A(n46558), .X(n46559) );
  inv_x8_sg U72321 ( .A(n46560), .X(n46561) );
  inv_x8_sg U72322 ( .A(n46561), .X(n51306) );
  inv_x8_sg U72323 ( .A(n10518), .X(n51293) );
  inv_x8_sg U72324 ( .A(n46562), .X(n46563) );
  inv_x8_sg U72325 ( .A(n46563), .X(n51280) );
  inv_x8_sg U72326 ( .A(n10408), .X(n46564) );
  inv_x8_sg U72327 ( .A(n46564), .X(n46565) );
  inv_x8_sg U72328 ( .A(n46572), .X(n46566) );
  inv_x8_sg U72329 ( .A(n10397), .X(n46567) );
  inv_x8_sg U72330 ( .A(n46567), .X(n46568) );
  inv_x8_sg U72331 ( .A(n43872), .X(n46569) );
  inv_x8_sg U72332 ( .A(n46569), .X(n46570) );
  inv_x8_sg U72333 ( .A(n46571), .X(n46572) );
  inv_x8_sg U72334 ( .A(n10403), .X(n46573) );
  inv_x8_sg U72335 ( .A(n46573), .X(n46574) );
  inv_x8_sg U72336 ( .A(n46578), .X(n46575) );
  inv_x8_sg U72337 ( .A(n39300), .X(n46576) );
  nand_x8_sg U72338 ( .A(n11831), .B(n24470), .X(n46577) );
  nand_x8_sg U72339 ( .A(n11831), .B(n24470), .X(n46578) );
  inv_x8_sg U72340 ( .A(n11830), .X(n46579) );
  inv_x8_sg U72341 ( .A(n46579), .X(n46580) );
  inv_x8_sg U72342 ( .A(n46581), .X(n46582) );
  inv_x8_sg U72343 ( .A(n44717), .X(n46583) );
  inv_x8_sg U72344 ( .A(n46583), .X(n46584) );
  inv_x8_sg U72345 ( .A(n46586), .X(n46585) );
  inv_x8_sg U72346 ( .A(n46588), .X(n46587) );
  inv_x8_sg U72347 ( .A(n46590), .X(n46589) );
  inv_x8_sg U72348 ( .A(n46592), .X(n46591) );
  inv_x8_sg U72349 ( .A(n27901), .X(n46592) );
  inv_x8_sg U72350 ( .A(n46594), .X(n46593) );
  inv_x8_sg U72351 ( .A(n46597), .X(n46596) );
  inv_x8_sg U72352 ( .A(n46599), .X(n46598) );
  inv_x8_sg U72353 ( .A(n46601), .X(n46600) );
  inv_x8_sg U72354 ( .A(n10281), .X(n46602) );
  inv_x8_sg U72355 ( .A(n46604), .X(n46603) );
  inv_x8_sg U72356 ( .A(n10256), .X(n46607) );
  inv_x8_sg U72357 ( .A(n46609), .X(n46608) );
  inv_x8_sg U72358 ( .A(n25667), .X(n46611) );
  inv_x8_sg U72359 ( .A(n46613), .X(n46612) );
  inv_x8_sg U72360 ( .A(n25388), .X(n46615) );
  inv_x8_sg U72361 ( .A(n46617), .X(n46616) );
  inv_x8_sg U72362 ( .A(n46620), .X(n46619) );
  inv_x8_sg U72363 ( .A(n46622), .X(n46621) );
  inv_x8_sg U72364 ( .A(n46624), .X(n46623) );
  inv_x8_sg U72365 ( .A(n26783), .X(n46625) );
  inv_x8_sg U72366 ( .A(n46637), .X(n46626) );
  inv_x8_sg U72367 ( .A(n46633), .X(n46627) );
  inv_x8_sg U72368 ( .A(n46633), .X(n46628) );
  inv_x8_sg U72369 ( .A(n46633), .X(n46629) );
  inv_x8_sg U72370 ( .A(n46637), .X(n46631) );
  inv_x8_sg U72371 ( .A(n46637), .X(n46632) );
  inv_x8_sg U72372 ( .A(n46635), .X(n46633) );
  inv_x8_sg U72373 ( .A(n46637), .X(n46634) );
  inv_x8_sg U72374 ( .A(n46637), .X(n46635) );
  inv_x8_sg U72375 ( .A(n46638), .X(n46637) );
  inv_x8_sg U72376 ( .A(n46639), .X(n46638) );
  inv_x8_sg U72377 ( .A(n46656), .X(n46641) );
  inv_x8_sg U72378 ( .A(n46649), .X(n46642) );
  inv_x8_sg U72379 ( .A(n46649), .X(n46643) );
  inv_x8_sg U72380 ( .A(n46649), .X(n46644) );
  inv_x8_sg U72381 ( .A(n46656), .X(n46645) );
  inv_x8_sg U72382 ( .A(n46649), .X(n46646) );
  inv_x8_sg U72383 ( .A(n46649), .X(n46647) );
  inv_x8_sg U72384 ( .A(n46656), .X(n46648) );
  inv_x8_sg U72385 ( .A(n46657), .X(n46649) );
  inv_x8_sg U72386 ( .A(n46649), .X(n46650) );
  inv_x8_sg U72387 ( .A(n46656), .X(n46651) );
  inv_x8_sg U72388 ( .A(n46656), .X(n46652) );
  inv_x8_sg U72389 ( .A(n46656), .X(n46653) );
  inv_x8_sg U72390 ( .A(n46656), .X(n46654) );
  inv_x8_sg U72391 ( .A(n46656), .X(n46655) );
  inv_x8_sg U72392 ( .A(n46657), .X(n46656) );
  inv_x8_sg U72393 ( .A(n46658), .X(n46657) );
  inv_x8_sg U72394 ( .A(n46673), .X(n46672) );
  inv_x4_sg U72395 ( .A(n40909), .X(n46673) );
  inv_x2_sg U74971 ( .A(n29426), .X(n55454) );
  inv_x2_sg U74972 ( .A(n29422), .X(n55629) );
  inv_x2_sg U74973 ( .A(n29413), .X(n55628) );
  inv_x2_sg U74974 ( .A(n29412), .X(n55456) );
  inv_x2_sg U74975 ( .A(n29408), .X(n55627) );
  inv_x2_sg U74976 ( .A(n29401), .X(n55779) );
  inv_x2_sg U74977 ( .A(n43815), .X(n55626) );
  inv_x2_sg U74978 ( .A(n29387), .X(n55778) );
  inv_x2_sg U74979 ( .A(n43900), .X(n55625) );
  inv_x2_sg U74980 ( .A(n29373), .X(n55777) );
  inv_x2_sg U74981 ( .A(n44040), .X(n55624) );
  inv_x2_sg U74982 ( .A(n29358), .X(n55776) );
  inv_x2_sg U74983 ( .A(n44217), .X(n55623) );
  inv_x2_sg U74984 ( .A(n29347), .X(n55238) );
  inv_x2_sg U74985 ( .A(n44479), .X(n55622) );
  inv_x2_sg U74986 ( .A(n29337), .X(n55775) );
  inv_x2_sg U74987 ( .A(n29335), .X(n55212) );
  inv_x2_sg U74988 ( .A(n29329), .X(n55774) );
  inv_x2_sg U74989 ( .A(n29322), .X(n55773) );
  inv_x2_sg U74990 ( .A(n29315), .X(n55772) );
  inv_x2_sg U74991 ( .A(n29308), .X(n55771) );
  inv_x2_sg U74992 ( .A(n29536), .X(n55453) );
  inv_x2_sg U74993 ( .A(n29302), .X(n55770) );
  inv_x2_sg U74994 ( .A(n29144), .X(n55170) );
  inv_x2_sg U74995 ( .A(n29140), .X(n55621) );
  inv_x2_sg U74996 ( .A(n29131), .X(n55620) );
  inv_x2_sg U74997 ( .A(n29130), .X(n55172) );
  inv_x2_sg U74998 ( .A(n29126), .X(n55619) );
  inv_x2_sg U74999 ( .A(n29119), .X(n55769) );
  inv_x2_sg U75000 ( .A(n43817), .X(n55618) );
  inv_x2_sg U75001 ( .A(n29105), .X(n55768) );
  inv_x2_sg U75002 ( .A(n43902), .X(n55617) );
  inv_x2_sg U75003 ( .A(n29091), .X(n55767) );
  inv_x2_sg U75004 ( .A(n43904), .X(n55616) );
  inv_x2_sg U75005 ( .A(n29077), .X(n55766) );
  inv_x2_sg U75006 ( .A(n44219), .X(n55615) );
  inv_x2_sg U75007 ( .A(n29066), .X(n54949) );
  inv_x2_sg U75008 ( .A(n44042), .X(n55614) );
  inv_x2_sg U75009 ( .A(n29056), .X(n55765) );
  inv_x2_sg U75010 ( .A(n29054), .X(n54922) );
  inv_x2_sg U75011 ( .A(n29048), .X(n55764) );
  inv_x2_sg U75012 ( .A(n29041), .X(n55763) );
  inv_x2_sg U75013 ( .A(n29034), .X(n55762) );
  inv_x2_sg U75014 ( .A(n29027), .X(n55761) );
  inv_x2_sg U75015 ( .A(n29258), .X(n55169) );
  inv_x2_sg U75016 ( .A(n29021), .X(n55760) );
  inv_x2_sg U75017 ( .A(n29149), .X(n55783) );
  inv_x2_sg U75018 ( .A(n28865), .X(n54886) );
  inv_x2_sg U75019 ( .A(n28861), .X(n55613) );
  inv_x2_sg U75020 ( .A(n28852), .X(n55612) );
  inv_x2_sg U75021 ( .A(n28851), .X(n54888) );
  inv_x2_sg U75022 ( .A(n28847), .X(n55611) );
  inv_x2_sg U75023 ( .A(n28840), .X(n55759) );
  inv_x2_sg U75024 ( .A(n44044), .X(n55610) );
  inv_x2_sg U75025 ( .A(n28826), .X(n55758) );
  inv_x2_sg U75026 ( .A(n44221), .X(n55609) );
  inv_x2_sg U75027 ( .A(n28812), .X(n55757) );
  inv_x2_sg U75028 ( .A(n44223), .X(n55608) );
  inv_x2_sg U75029 ( .A(n28797), .X(n55756) );
  inv_x2_sg U75030 ( .A(n44225), .X(n55607) );
  inv_x2_sg U75031 ( .A(n28786), .X(n54670) );
  inv_x2_sg U75032 ( .A(n44481), .X(n55606) );
  inv_x2_sg U75033 ( .A(n28776), .X(n55755) );
  inv_x2_sg U75034 ( .A(n28774), .X(n54644) );
  inv_x2_sg U75035 ( .A(n28768), .X(n55754) );
  inv_x2_sg U75036 ( .A(n28761), .X(n55753) );
  inv_x2_sg U75037 ( .A(n28754), .X(n55752) );
  inv_x2_sg U75038 ( .A(n28747), .X(n55751) );
  inv_x2_sg U75039 ( .A(n28975), .X(n54885) );
  inv_x2_sg U75040 ( .A(n28741), .X(n55750) );
  inv_x2_sg U75041 ( .A(n26358), .X(n55780) );
  inv_x2_sg U75042 ( .A(n28585), .X(n54602) );
  inv_x2_sg U75043 ( .A(n28581), .X(n55605) );
  inv_x2_sg U75044 ( .A(n28572), .X(n55604) );
  inv_x2_sg U75045 ( .A(n28571), .X(n54604) );
  inv_x2_sg U75046 ( .A(n28567), .X(n55603) );
  inv_x2_sg U75047 ( .A(n28560), .X(n55749) );
  inv_x2_sg U75048 ( .A(n43906), .X(n55602) );
  inv_x2_sg U75049 ( .A(n28546), .X(n55748) );
  inv_x2_sg U75050 ( .A(n43819), .X(n55601) );
  inv_x2_sg U75051 ( .A(n28532), .X(n55747) );
  inv_x2_sg U75052 ( .A(n43821), .X(n55600) );
  inv_x2_sg U75053 ( .A(n28518), .X(n55746) );
  inv_x2_sg U75054 ( .A(n43908), .X(n55599) );
  inv_x2_sg U75055 ( .A(n28507), .X(n54381) );
  inv_x2_sg U75056 ( .A(n44046), .X(n55598) );
  inv_x2_sg U75057 ( .A(n28497), .X(n55745) );
  inv_x2_sg U75058 ( .A(n28495), .X(n54354) );
  inv_x2_sg U75059 ( .A(n28489), .X(n55744) );
  inv_x2_sg U75060 ( .A(n28482), .X(n55743) );
  inv_x2_sg U75061 ( .A(n28475), .X(n55742) );
  inv_x2_sg U75062 ( .A(n28468), .X(n55741) );
  inv_x2_sg U75063 ( .A(n28697), .X(n54601) );
  inv_x2_sg U75064 ( .A(n28462), .X(n55740) );
  inv_x2_sg U75065 ( .A(n28307), .X(n54318) );
  inv_x2_sg U75066 ( .A(n28303), .X(n55597) );
  inv_x2_sg U75067 ( .A(n28294), .X(n55596) );
  inv_x2_sg U75068 ( .A(n28293), .X(n54320) );
  inv_x2_sg U75069 ( .A(n28289), .X(n55595) );
  inv_x2_sg U75070 ( .A(n28282), .X(n55739) );
  inv_x2_sg U75071 ( .A(n44227), .X(n55594) );
  inv_x2_sg U75072 ( .A(n28268), .X(n55738) );
  inv_x2_sg U75073 ( .A(n43910), .X(n55593) );
  inv_x2_sg U75074 ( .A(n28254), .X(n55737) );
  inv_x2_sg U75075 ( .A(n44483), .X(n55592) );
  inv_x2_sg U75076 ( .A(n28239), .X(n55736) );
  inv_x2_sg U75077 ( .A(n44485), .X(n55591) );
  inv_x2_sg U75078 ( .A(n28228), .X(n54098) );
  inv_x2_sg U75079 ( .A(n43912), .X(n55590) );
  inv_x2_sg U75080 ( .A(n28218), .X(n55735) );
  inv_x2_sg U75081 ( .A(n28216), .X(n54080) );
  inv_x2_sg U75082 ( .A(n28210), .X(n55734) );
  inv_x2_sg U75083 ( .A(n28203), .X(n55733) );
  inv_x2_sg U75084 ( .A(n28196), .X(n55732) );
  inv_x2_sg U75085 ( .A(n28189), .X(n55731) );
  inv_x2_sg U75086 ( .A(n28418), .X(n54317) );
  inv_x2_sg U75087 ( .A(n28183), .X(n55730) );
  inv_x2_sg U75088 ( .A(n28027), .X(n54037) );
  inv_x2_sg U75089 ( .A(n28023), .X(n55589) );
  inv_x2_sg U75090 ( .A(n28014), .X(n55588) );
  inv_x2_sg U75091 ( .A(n28013), .X(n54039) );
  inv_x2_sg U75092 ( .A(n28009), .X(n55587) );
  inv_x2_sg U75093 ( .A(n28002), .X(n55729) );
  inv_x2_sg U75094 ( .A(n43794), .X(n55586) );
  inv_x2_sg U75095 ( .A(n27988), .X(n55728) );
  inv_x2_sg U75096 ( .A(n43823), .X(n55585) );
  inv_x2_sg U75097 ( .A(n27974), .X(n55727) );
  inv_x2_sg U75098 ( .A(n43914), .X(n55584) );
  inv_x2_sg U75099 ( .A(n27960), .X(n55726) );
  inv_x2_sg U75100 ( .A(n44229), .X(n55583) );
  inv_x2_sg U75101 ( .A(n27949), .X(n53816) );
  inv_x2_sg U75102 ( .A(n44048), .X(n55582) );
  inv_x2_sg U75103 ( .A(n27939), .X(n55725) );
  inv_x2_sg U75104 ( .A(n27937), .X(n53789) );
  inv_x2_sg U75105 ( .A(n27931), .X(n55724) );
  inv_x2_sg U75106 ( .A(n27924), .X(n55723) );
  inv_x2_sg U75107 ( .A(n27917), .X(n55722) );
  inv_x2_sg U75108 ( .A(n27910), .X(n55721) );
  inv_x2_sg U75109 ( .A(n28139), .X(n54036) );
  inv_x2_sg U75110 ( .A(n27904), .X(n55720) );
  inv_x2_sg U75111 ( .A(n27748), .X(n53753) );
  inv_x2_sg U75112 ( .A(n27744), .X(n55581) );
  inv_x2_sg U75113 ( .A(n27735), .X(n55580) );
  inv_x2_sg U75114 ( .A(n27734), .X(n53755) );
  inv_x2_sg U75115 ( .A(n27730), .X(n55579) );
  inv_x2_sg U75116 ( .A(n27722), .X(n55719) );
  inv_x2_sg U75117 ( .A(n43769), .X(n55578) );
  inv_x2_sg U75118 ( .A(n27708), .X(n55718) );
  inv_x2_sg U75119 ( .A(n43796), .X(n55577) );
  inv_x2_sg U75120 ( .A(n27694), .X(n55717) );
  inv_x2_sg U75121 ( .A(n44231), .X(n55576) );
  inv_x2_sg U75122 ( .A(n27680), .X(n55716) );
  inv_x2_sg U75123 ( .A(n44487), .X(n55575) );
  inv_x2_sg U75124 ( .A(n27669), .X(n53538) );
  inv_x2_sg U75125 ( .A(n44050), .X(n55574) );
  inv_x2_sg U75126 ( .A(n27659), .X(n55715) );
  inv_x2_sg U75127 ( .A(n27657), .X(n53510) );
  inv_x2_sg U75128 ( .A(n27651), .X(n55714) );
  inv_x2_sg U75129 ( .A(n27644), .X(n55713) );
  inv_x2_sg U75130 ( .A(n27637), .X(n55712) );
  inv_x2_sg U75131 ( .A(n27630), .X(n55711) );
  inv_x2_sg U75132 ( .A(n27858), .X(n53752) );
  inv_x2_sg U75133 ( .A(n27624), .X(n55710) );
  inv_x2_sg U75134 ( .A(n27467), .X(n53475) );
  inv_x2_sg U75135 ( .A(n27463), .X(n55573) );
  inv_x2_sg U75136 ( .A(n27454), .X(n55572) );
  inv_x2_sg U75137 ( .A(n27453), .X(n53477) );
  inv_x2_sg U75138 ( .A(n27449), .X(n55571) );
  inv_x2_sg U75139 ( .A(n27442), .X(n55709) );
  inv_x2_sg U75140 ( .A(n27428), .X(n55708) );
  inv_x2_sg U75141 ( .A(n43825), .X(n55570) );
  inv_x2_sg U75142 ( .A(n27414), .X(n55707) );
  inv_x2_sg U75143 ( .A(n43916), .X(n55569) );
  inv_x2_sg U75144 ( .A(n27400), .X(n55706) );
  inv_x2_sg U75145 ( .A(n45487), .X(n55568) );
  inv_x2_sg U75146 ( .A(n27389), .X(n53263) );
  inv_x2_sg U75147 ( .A(n44489), .X(n55567) );
  inv_x2_sg U75148 ( .A(n27379), .X(n55705) );
  inv_x2_sg U75149 ( .A(n27377), .X(n53237) );
  inv_x2_sg U75150 ( .A(n27371), .X(n55704) );
  inv_x2_sg U75151 ( .A(n27364), .X(n55703) );
  inv_x2_sg U75152 ( .A(n27357), .X(n55702) );
  inv_x2_sg U75153 ( .A(n27350), .X(n55701) );
  inv_x2_sg U75154 ( .A(n27579), .X(n53474) );
  inv_x2_sg U75155 ( .A(n27344), .X(n55700) );
  inv_x2_sg U75156 ( .A(n27188), .X(n53195) );
  inv_x2_sg U75157 ( .A(n27184), .X(n55566) );
  inv_x2_sg U75158 ( .A(n27175), .X(n55565) );
  inv_x2_sg U75159 ( .A(n27174), .X(n53197) );
  inv_x2_sg U75160 ( .A(n27170), .X(n55564) );
  inv_x2_sg U75161 ( .A(n27162), .X(n55699) );
  inv_x2_sg U75162 ( .A(n43918), .X(n55563) );
  inv_x2_sg U75163 ( .A(n27148), .X(n55698) );
  inv_x2_sg U75164 ( .A(n43827), .X(n55562) );
  inv_x2_sg U75165 ( .A(n27134), .X(n55697) );
  inv_x2_sg U75166 ( .A(n44233), .X(n55561) );
  inv_x2_sg U75167 ( .A(n27120), .X(n55696) );
  inv_x2_sg U75168 ( .A(n44491), .X(n55560) );
  inv_x2_sg U75169 ( .A(n27109), .X(n52980) );
  inv_x2_sg U75170 ( .A(n44052), .X(n55559) );
  inv_x2_sg U75171 ( .A(n27099), .X(n55695) );
  inv_x2_sg U75172 ( .A(n27097), .X(n52952) );
  inv_x2_sg U75173 ( .A(n27091), .X(n55694) );
  inv_x2_sg U75174 ( .A(n27084), .X(n55693) );
  inv_x2_sg U75175 ( .A(n27077), .X(n55692) );
  inv_x2_sg U75176 ( .A(n27070), .X(n55691) );
  inv_x2_sg U75177 ( .A(n27300), .X(n53194) );
  inv_x2_sg U75178 ( .A(n27064), .X(n55690) );
  inv_x2_sg U75179 ( .A(n26908), .X(n52917) );
  inv_x2_sg U75180 ( .A(n26904), .X(n55558) );
  inv_x2_sg U75181 ( .A(n26895), .X(n55557) );
  inv_x2_sg U75182 ( .A(n26894), .X(n52919) );
  inv_x2_sg U75183 ( .A(n26890), .X(n55556) );
  inv_x2_sg U75184 ( .A(n26883), .X(n55689) );
  inv_x2_sg U75185 ( .A(n43829), .X(n55555) );
  inv_x2_sg U75186 ( .A(n26869), .X(n55688) );
  inv_x2_sg U75187 ( .A(n43920), .X(n55554) );
  inv_x2_sg U75188 ( .A(n26855), .X(n55687) );
  inv_x2_sg U75189 ( .A(n44054), .X(n55553) );
  inv_x2_sg U75190 ( .A(n26841), .X(n55686) );
  inv_x2_sg U75191 ( .A(n44235), .X(n55552) );
  inv_x2_sg U75192 ( .A(n26830), .X(n52704) );
  inv_x2_sg U75193 ( .A(n43922), .X(n55551) );
  inv_x2_sg U75194 ( .A(n26820), .X(n55685) );
  inv_x2_sg U75195 ( .A(n26818), .X(n52680) );
  inv_x2_sg U75196 ( .A(n26812), .X(n55684) );
  inv_x2_sg U75197 ( .A(n26805), .X(n55683) );
  inv_x2_sg U75198 ( .A(n26798), .X(n55682) );
  inv_x2_sg U75199 ( .A(n26791), .X(n55681) );
  inv_x2_sg U75200 ( .A(n27020), .X(n52916) );
  inv_x2_sg U75201 ( .A(n26785), .X(n55680) );
  inv_x2_sg U75202 ( .A(n26631), .X(n52636) );
  inv_x2_sg U75203 ( .A(n26627), .X(n55550) );
  inv_x2_sg U75204 ( .A(n26618), .X(n55549) );
  inv_x2_sg U75205 ( .A(n26617), .X(n52638) );
  inv_x2_sg U75206 ( .A(n26613), .X(n55548) );
  inv_x2_sg U75207 ( .A(n26605), .X(n55679) );
  inv_x2_sg U75208 ( .A(n44237), .X(n55547) );
  inv_x2_sg U75209 ( .A(n26591), .X(n55678) );
  inv_x2_sg U75210 ( .A(n43924), .X(n55546) );
  inv_x2_sg U75211 ( .A(n26577), .X(n55677) );
  inv_x2_sg U75212 ( .A(n43926), .X(n55545) );
  inv_x2_sg U75213 ( .A(n26563), .X(n55676) );
  inv_x2_sg U75214 ( .A(n44493), .X(n55544) );
  inv_x2_sg U75215 ( .A(n26552), .X(n52427) );
  inv_x2_sg U75216 ( .A(n44056), .X(n55543) );
  inv_x2_sg U75217 ( .A(n26542), .X(n55675) );
  inv_x2_sg U75218 ( .A(n26540), .X(n52403) );
  inv_x2_sg U75219 ( .A(n26534), .X(n55674) );
  inv_x2_sg U75220 ( .A(n26527), .X(n55673) );
  inv_x2_sg U75221 ( .A(n26520), .X(n55672) );
  inv_x2_sg U75222 ( .A(n26513), .X(n55671) );
  inv_x2_sg U75223 ( .A(n26741), .X(n52635) );
  inv_x2_sg U75224 ( .A(n26507), .X(n55670) );
  inv_x2_sg U75225 ( .A(n26352), .X(n52361) );
  inv_x2_sg U75226 ( .A(n26348), .X(n55542) );
  inv_x2_sg U75227 ( .A(n26339), .X(n55541) );
  inv_x2_sg U75228 ( .A(n26338), .X(n52363) );
  inv_x2_sg U75229 ( .A(n26334), .X(n55540) );
  inv_x2_sg U75230 ( .A(n26326), .X(n55669) );
  inv_x2_sg U75231 ( .A(n43928), .X(n55539) );
  inv_x2_sg U75232 ( .A(n26312), .X(n55668) );
  inv_x2_sg U75233 ( .A(n43831), .X(n55538) );
  inv_x2_sg U75234 ( .A(n26298), .X(n55667) );
  inv_x2_sg U75235 ( .A(n44239), .X(n55537) );
  inv_x2_sg U75236 ( .A(n26284), .X(n55666) );
  inv_x2_sg U75237 ( .A(n44495), .X(n55536) );
  inv_x2_sg U75238 ( .A(n26273), .X(n52146) );
  inv_x2_sg U75239 ( .A(n44058), .X(n55535) );
  inv_x2_sg U75240 ( .A(n26263), .X(n55665) );
  inv_x2_sg U75241 ( .A(n26261), .X(n52118) );
  inv_x2_sg U75242 ( .A(n26255), .X(n55664) );
  inv_x2_sg U75243 ( .A(n26248), .X(n55663) );
  inv_x2_sg U75244 ( .A(n26241), .X(n55662) );
  inv_x2_sg U75245 ( .A(n26234), .X(n55661) );
  inv_x2_sg U75246 ( .A(n26463), .X(n52360) );
  inv_x2_sg U75247 ( .A(n26228), .X(n55660) );
  inv_x2_sg U75248 ( .A(n26071), .X(n52083) );
  inv_x2_sg U75249 ( .A(n26067), .X(n55534) );
  inv_x2_sg U75250 ( .A(n26058), .X(n55533) );
  inv_x2_sg U75251 ( .A(n26057), .X(n52085) );
  inv_x2_sg U75252 ( .A(n26053), .X(n55532) );
  inv_x2_sg U75253 ( .A(n26045), .X(n55659) );
  inv_x2_sg U75254 ( .A(n26031), .X(n55658) );
  inv_x2_sg U75255 ( .A(n43833), .X(n55531) );
  inv_x2_sg U75256 ( .A(n26017), .X(n55657) );
  inv_x2_sg U75257 ( .A(n43930), .X(n55530) );
  inv_x2_sg U75258 ( .A(n26003), .X(n55656) );
  inv_x2_sg U75259 ( .A(n44241), .X(n55529) );
  inv_x2_sg U75260 ( .A(n25992), .X(n51876) );
  inv_x2_sg U75261 ( .A(n44497), .X(n55528) );
  inv_x2_sg U75262 ( .A(n25982), .X(n55655) );
  inv_x2_sg U75263 ( .A(n25980), .X(n51851) );
  inv_x2_sg U75264 ( .A(n25974), .X(n55654) );
  inv_x2_sg U75265 ( .A(n25967), .X(n55653) );
  inv_x2_sg U75266 ( .A(n25960), .X(n55652) );
  inv_x2_sg U75267 ( .A(n25953), .X(n55651) );
  inv_x2_sg U75268 ( .A(n26184), .X(n52082) );
  inv_x2_sg U75269 ( .A(n25947), .X(n55650) );
  inv_x2_sg U75270 ( .A(n26076), .X(n55781) );
  inv_x2_sg U75271 ( .A(n25792), .X(n51807) );
  inv_x2_sg U75272 ( .A(n25788), .X(n55527) );
  inv_x2_sg U75273 ( .A(n25779), .X(n55526) );
  inv_x2_sg U75274 ( .A(n25778), .X(n51809) );
  inv_x2_sg U75275 ( .A(n25774), .X(n55525) );
  inv_x2_sg U75276 ( .A(n25767), .X(n55649) );
  inv_x2_sg U75277 ( .A(n25753), .X(n55648) );
  inv_x2_sg U75278 ( .A(n44060), .X(n55524) );
  inv_x2_sg U75279 ( .A(n25739), .X(n55647) );
  inv_x2_sg U75280 ( .A(n43932), .X(n55523) );
  inv_x2_sg U75281 ( .A(n25725), .X(n55646) );
  inv_x2_sg U75282 ( .A(n44499), .X(n55522) );
  inv_x2_sg U75283 ( .A(n25714), .X(n51588) );
  inv_x2_sg U75284 ( .A(n44062), .X(n55521) );
  inv_x2_sg U75285 ( .A(n25704), .X(n55645) );
  inv_x2_sg U75286 ( .A(n25702), .X(n51561) );
  inv_x2_sg U75287 ( .A(n25696), .X(n55644) );
  inv_x2_sg U75288 ( .A(n25689), .X(n55643) );
  inv_x2_sg U75289 ( .A(n25682), .X(n55642) );
  inv_x2_sg U75290 ( .A(n25675), .X(n55641) );
  inv_x2_sg U75291 ( .A(n25904), .X(n51806) );
  inv_x2_sg U75292 ( .A(n25669), .X(n55640) );
  inv_x2_sg U75293 ( .A(n25516), .X(n55782) );
  inv_x2_sg U75294 ( .A(n25514), .X(n51525) );
  inv_x2_sg U75295 ( .A(n25510), .X(n55520) );
  inv_x2_sg U75296 ( .A(n25501), .X(n55519) );
  inv_x2_sg U75297 ( .A(n25500), .X(n51527) );
  inv_x2_sg U75298 ( .A(n25496), .X(n55518) );
  inv_x2_sg U75299 ( .A(n25489), .X(n55639) );
  inv_x2_sg U75300 ( .A(n43835), .X(n55517) );
  inv_x2_sg U75301 ( .A(n25475), .X(n55638) );
  inv_x2_sg U75302 ( .A(n43934), .X(n55516) );
  inv_x2_sg U75303 ( .A(n25461), .X(n55637) );
  inv_x2_sg U75304 ( .A(n44064), .X(n55515) );
  inv_x2_sg U75305 ( .A(n25446), .X(n55636) );
  inv_x2_sg U75306 ( .A(n44243), .X(n55514) );
  inv_x2_sg U75307 ( .A(n25435), .X(n51316) );
  inv_x2_sg U75308 ( .A(n44501), .X(n55513) );
  inv_x2_sg U75309 ( .A(n25425), .X(n55635) );
  inv_x2_sg U75310 ( .A(n25423), .X(n51290) );
  inv_x2_sg U75311 ( .A(n25417), .X(n55634) );
  inv_x2_sg U75312 ( .A(n25410), .X(n55633) );
  inv_x2_sg U75313 ( .A(n25403), .X(n55632) );
  inv_x2_sg U75314 ( .A(n25396), .X(n55631) );
  inv_x2_sg U75315 ( .A(n25623), .X(n51524) );
  inv_x2_sg U75316 ( .A(n25389), .X(n55630) );
  inv_x2_sg U75317 ( .A(n25338), .X(n49266) );
  inv_x2_sg U75318 ( .A(n44066), .X(n49299) );
  inv_x2_sg U75319 ( .A(n29731), .X(n49298) );
  inv_x2_sg U75320 ( .A(n44531), .X(n49342) );
  inv_x2_sg U75321 ( .A(n29738), .X(n49341) );
  inv_x2_sg U75322 ( .A(n44533), .X(n49386) );
  inv_x2_sg U75323 ( .A(n29745), .X(n49385) );
  inv_x2_sg U75324 ( .A(n44535), .X(n49432) );
  inv_x2_sg U75325 ( .A(n29752), .X(n49431) );
  inv_x2_sg U75326 ( .A(n44539), .X(n49478) );
  inv_x2_sg U75327 ( .A(n29759), .X(n49477) );
  inv_x2_sg U75328 ( .A(n44541), .X(n49525) );
  inv_x2_sg U75329 ( .A(n29766), .X(n49524) );
  inv_x2_sg U75330 ( .A(n44545), .X(n49572) );
  inv_x2_sg U75331 ( .A(n29773), .X(n49571) );
  inv_x2_sg U75332 ( .A(n44549), .X(n49618) );
  inv_x2_sg U75333 ( .A(n29780), .X(n49617) );
  inv_x2_sg U75334 ( .A(n44553), .X(n49665) );
  inv_x2_sg U75335 ( .A(n29787), .X(n49664) );
  inv_x2_sg U75336 ( .A(n44557), .X(n49712) );
  inv_x2_sg U75337 ( .A(n29794), .X(n49711) );
  inv_x2_sg U75338 ( .A(n44561), .X(n49761) );
  inv_x2_sg U75339 ( .A(n29801), .X(n49760) );
  inv_x2_sg U75340 ( .A(n44563), .X(n49808) );
  inv_x2_sg U75341 ( .A(n29808), .X(n49807) );
  inv_x2_sg U75342 ( .A(n44567), .X(n49856) );
  inv_x2_sg U75343 ( .A(n29815), .X(n49855) );
  inv_x2_sg U75344 ( .A(n44571), .X(n49903) );
  inv_x2_sg U75345 ( .A(n29822), .X(n49902) );
  inv_x2_sg U75346 ( .A(n44573), .X(n49951) );
  inv_x2_sg U75347 ( .A(n29829), .X(n49950) );
  inv_x2_sg U75348 ( .A(n44575), .X(n49995) );
  inv_x2_sg U75349 ( .A(n29836), .X(n49994) );
  inv_x2_sg U75350 ( .A(n44529), .X(n50045) );
  inv_x2_sg U75351 ( .A(n29848), .X(n50047) );
  inv_x2_sg U75352 ( .A(n29857), .X(n50044) );
  inv_x2_sg U75353 ( .A(n30008), .X(n50038) );
  inv_x2_sg U75354 ( .A(n30014), .X(n49999) );
  inv_x2_sg U75355 ( .A(n30077), .X(n49301) );
  inv_x2_sg U75356 ( .A(n30083), .X(n49346) );
  inv_x2_sg U75357 ( .A(n30089), .X(n49390) );
  inv_x2_sg U75358 ( .A(n30095), .X(n49436) );
  inv_x2_sg U75359 ( .A(n30101), .X(n49482) );
  inv_x2_sg U75360 ( .A(n30107), .X(n49529) );
  inv_x2_sg U75361 ( .A(n30113), .X(n49576) );
  inv_x2_sg U75362 ( .A(n30119), .X(n49622) );
  inv_x2_sg U75363 ( .A(n30125), .X(n49669) );
  inv_x2_sg U75364 ( .A(n30131), .X(n49716) );
  inv_x2_sg U75365 ( .A(n30137), .X(n49765) );
  inv_x2_sg U75366 ( .A(n30143), .X(n49812) );
  inv_x2_sg U75367 ( .A(n30149), .X(n49860) );
  inv_x2_sg U75368 ( .A(n30155), .X(n49907) );
  inv_x2_sg U75369 ( .A(n30161), .X(n49955) );
  inv_x2_sg U75370 ( .A(n30237), .X(n50064) );
  inv_x2_sg U75371 ( .A(n30244), .X(n50092) );
  inv_x2_sg U75372 ( .A(n30252), .X(n50069) );
  inv_x2_sg U75373 ( .A(n30280), .X(n50091) );
  inv_x2_sg U75374 ( .A(n25321), .X(n49292) );
  inv_x2_sg U75375 ( .A(n30345), .X(n49333) );
  inv_x2_sg U75376 ( .A(n30351), .X(n49377) );
  inv_x2_sg U75377 ( .A(n30357), .X(n49423) );
  inv_x2_sg U75378 ( .A(n30363), .X(n49469) );
  inv_x2_sg U75379 ( .A(n30369), .X(n49516) );
  inv_x2_sg U75380 ( .A(n30375), .X(n49563) );
  inv_x2_sg U75381 ( .A(n30381), .X(n49609) );
  inv_x2_sg U75382 ( .A(n30387), .X(n49656) );
  inv_x2_sg U75383 ( .A(n30393), .X(n49703) );
  inv_x2_sg U75384 ( .A(n30399), .X(n49752) );
  inv_x2_sg U75385 ( .A(n30405), .X(n49800) );
  inv_x2_sg U75386 ( .A(n30411), .X(n49847) );
  inv_x2_sg U75387 ( .A(n30417), .X(n49894) );
  inv_x2_sg U75388 ( .A(n30423), .X(n49942) );
  inv_x2_sg U75389 ( .A(n30429), .X(n49987) );
  inv_x2_sg U75390 ( .A(n30435), .X(n50034) );
  inv_x2_sg U75391 ( .A(n30441), .X(n50079) );
  inv_x2_sg U75392 ( .A(n44631), .X(n50033) );
  inv_x2_sg U75393 ( .A(n30456), .X(n50065) );
  inv_x2_sg U75394 ( .A(n30459), .X(n50062) );
  inv_x2_sg U75395 ( .A(n45527), .X(n50016) );
  inv_x2_sg U75396 ( .A(n30465), .X(n50056) );
  inv_x2_sg U75397 ( .A(n44623), .X(n50009) );
  inv_x2_sg U75398 ( .A(n30472), .X(n50050) );
  inv_x2_sg U75399 ( .A(n30480), .X(n50008) );
  inv_x2_sg U75400 ( .A(n30484), .X(n50007) );
  inv_x2_sg U75401 ( .A(n30493), .X(n50015) );
  inv_x2_sg U75402 ( .A(n30506), .X(n50021) );
  inv_x2_sg U75403 ( .A(n30454), .X(n50067) );
  inv_x2_sg U75404 ( .A(n30517), .X(n50027) );
  inv_x2_sg U75405 ( .A(n30529), .X(n50032) );
  inv_x2_sg U75406 ( .A(n44068), .X(n49305) );
  inv_x2_sg U75407 ( .A(n30600), .X(n49304) );
  inv_x2_sg U75408 ( .A(n44649), .X(n49351) );
  inv_x2_sg U75409 ( .A(n30607), .X(n49350) );
  inv_x2_sg U75410 ( .A(n44635), .X(n49395) );
  inv_x2_sg U75411 ( .A(n30614), .X(n49394) );
  inv_x2_sg U75412 ( .A(n44537), .X(n49441) );
  inv_x2_sg U75413 ( .A(n30621), .X(n49440) );
  inv_x2_sg U75414 ( .A(n44637), .X(n49487) );
  inv_x2_sg U75415 ( .A(n30628), .X(n49486) );
  inv_x2_sg U75416 ( .A(n44543), .X(n49534) );
  inv_x2_sg U75417 ( .A(n30635), .X(n49533) );
  inv_x2_sg U75418 ( .A(n44547), .X(n49581) );
  inv_x2_sg U75419 ( .A(n30642), .X(n49580) );
  inv_x2_sg U75420 ( .A(n44551), .X(n49627) );
  inv_x2_sg U75421 ( .A(n30649), .X(n49626) );
  inv_x2_sg U75422 ( .A(n44555), .X(n49674) );
  inv_x2_sg U75423 ( .A(n30656), .X(n49673) );
  inv_x2_sg U75424 ( .A(n44559), .X(n49721) );
  inv_x2_sg U75425 ( .A(n30663), .X(n49720) );
  inv_x2_sg U75426 ( .A(n44639), .X(n49770) );
  inv_x2_sg U75427 ( .A(n30670), .X(n49769) );
  inv_x2_sg U75428 ( .A(n44565), .X(n49817) );
  inv_x2_sg U75429 ( .A(n30677), .X(n49816) );
  inv_x2_sg U75430 ( .A(n44569), .X(n49865) );
  inv_x2_sg U75431 ( .A(n30684), .X(n49864) );
  inv_x2_sg U75432 ( .A(n30690), .X(n49911) );
  inv_x2_sg U75433 ( .A(n30696), .X(n49959) );
  inv_x2_sg U75434 ( .A(n30714), .X(n50019) );
  inv_x2_sg U75435 ( .A(n45517), .X(n49972) );
  inv_x2_sg U75436 ( .A(n30720), .X(n50012) );
  inv_x2_sg U75437 ( .A(n30726), .X(n50006) );
  inv_x2_sg U75438 ( .A(n30739), .X(n49964) );
  inv_x2_sg U75439 ( .A(n30748), .X(n49971) );
  inv_x2_sg U75440 ( .A(n30761), .X(n49977) );
  inv_x2_sg U75441 ( .A(n30712), .X(n50022) );
  inv_x2_sg U75442 ( .A(n30709), .X(n50025) );
  inv_x2_sg U75443 ( .A(n30774), .X(n49982) );
  inv_x2_sg U75444 ( .A(n30786), .X(n50003) );
  inv_x2_sg U75445 ( .A(n30934), .X(n49980) );
  inv_x2_sg U75446 ( .A(n30940), .X(n49975) );
  inv_x2_sg U75447 ( .A(n45511), .X(n49928) );
  inv_x2_sg U75448 ( .A(n30946), .X(n49968) );
  inv_x2_sg U75449 ( .A(n30731), .X(n49917) );
  inv_x2_sg U75450 ( .A(n30965), .X(n49920) );
  inv_x2_sg U75451 ( .A(n30974), .X(n49927) );
  inv_x2_sg U75452 ( .A(n30987), .X(n49933) );
  inv_x2_sg U75453 ( .A(n30772), .X(n49936) );
  inv_x2_sg U75454 ( .A(n30998), .X(n49939) );
  inv_x2_sg U75455 ( .A(n31061), .X(n49307) );
  inv_x2_sg U75456 ( .A(n31067), .X(n49355) );
  inv_x2_sg U75457 ( .A(n31073), .X(n49399) );
  inv_x2_sg U75458 ( .A(n31079), .X(n49445) );
  inv_x2_sg U75459 ( .A(n31085), .X(n49491) );
  inv_x2_sg U75460 ( .A(n31091), .X(n49538) );
  inv_x2_sg U75461 ( .A(n31097), .X(n49585) );
  inv_x2_sg U75462 ( .A(n31103), .X(n49631) );
  inv_x2_sg U75463 ( .A(n31109), .X(n49678) );
  inv_x2_sg U75464 ( .A(n31115), .X(n49725) );
  inv_x2_sg U75465 ( .A(n31121), .X(n49774) );
  inv_x2_sg U75466 ( .A(n31127), .X(n49821) );
  inv_x2_sg U75467 ( .A(n31133), .X(n49869) );
  inv_x2_sg U75468 ( .A(n31145), .X(n49931) );
  inv_x2_sg U75469 ( .A(n45519), .X(n49882) );
  inv_x2_sg U75470 ( .A(n31151), .X(n49924) );
  inv_x2_sg U75471 ( .A(n31157), .X(n49919) );
  inv_x2_sg U75472 ( .A(n31170), .X(n49874) );
  inv_x2_sg U75473 ( .A(n31179), .X(n49881) );
  inv_x2_sg U75474 ( .A(n31192), .X(n49887) );
  inv_x2_sg U75475 ( .A(n31143), .X(n49934) );
  inv_x2_sg U75476 ( .A(n31140), .X(n49937) );
  inv_x2_sg U75477 ( .A(n31205), .X(n49915) );
  inv_x2_sg U75478 ( .A(n25308), .X(n49288) );
  inv_x2_sg U75479 ( .A(n31260), .X(n49309) );
  inv_x2_sg U75480 ( .A(n31264), .X(n49373) );
  inv_x2_sg U75481 ( .A(n31270), .X(n49419) );
  inv_x2_sg U75482 ( .A(n31276), .X(n49465) );
  inv_x2_sg U75483 ( .A(n31282), .X(n49512) );
  inv_x2_sg U75484 ( .A(n31288), .X(n49559) );
  inv_x2_sg U75485 ( .A(n31294), .X(n49605) );
  inv_x2_sg U75486 ( .A(n31300), .X(n49652) );
  inv_x2_sg U75487 ( .A(n31306), .X(n49699) );
  inv_x2_sg U75488 ( .A(n31312), .X(n49748) );
  inv_x2_sg U75489 ( .A(n31318), .X(n49797) );
  inv_x2_sg U75490 ( .A(n31324), .X(n49843) );
  inv_x2_sg U75491 ( .A(n31329), .X(n49890) );
  inv_x2_sg U75492 ( .A(n31335), .X(n49885) );
  inv_x2_sg U75493 ( .A(n45513), .X(n49836) );
  inv_x2_sg U75494 ( .A(n31341), .X(n49878) );
  inv_x2_sg U75495 ( .A(n31162), .X(n49825) );
  inv_x2_sg U75496 ( .A(n31360), .X(n49828) );
  inv_x2_sg U75497 ( .A(n31369), .X(n49835) );
  inv_x2_sg U75498 ( .A(n31382), .X(n49841) );
  inv_x2_sg U75499 ( .A(n31203), .X(n49871) );
  inv_x2_sg U75500 ( .A(n25328), .X(n49287) );
  inv_x2_sg U75501 ( .A(n31440), .X(n49311) );
  inv_x2_sg U75502 ( .A(n31446), .X(n49358) );
  inv_x2_sg U75503 ( .A(n31444), .X(n49372) );
  inv_x2_sg U75504 ( .A(n31452), .X(n49403) );
  inv_x2_sg U75505 ( .A(n31450), .X(n49418) );
  inv_x2_sg U75506 ( .A(n31458), .X(n49448) );
  inv_x2_sg U75507 ( .A(n31456), .X(n49464) );
  inv_x2_sg U75508 ( .A(n31464), .X(n49494) );
  inv_x2_sg U75509 ( .A(n31462), .X(n49511) );
  inv_x2_sg U75510 ( .A(n31470), .X(n49542) );
  inv_x2_sg U75511 ( .A(n31468), .X(n49558) );
  inv_x2_sg U75512 ( .A(n31476), .X(n49588) );
  inv_x2_sg U75513 ( .A(n31474), .X(n49604) );
  inv_x2_sg U75514 ( .A(n31482), .X(n49634) );
  inv_x2_sg U75515 ( .A(n31480), .X(n49651) );
  inv_x2_sg U75516 ( .A(n31488), .X(n49682) );
  inv_x2_sg U75517 ( .A(n31486), .X(n49698) );
  inv_x2_sg U75518 ( .A(n31494), .X(n49728) );
  inv_x2_sg U75519 ( .A(n31492), .X(n49747) );
  inv_x2_sg U75520 ( .A(n31497), .X(n49795) );
  inv_x2_sg U75521 ( .A(n31500), .X(n49778) );
  inv_x2_sg U75522 ( .A(n31506), .X(n49839) );
  inv_x2_sg U75523 ( .A(n45521), .X(n49791) );
  inv_x2_sg U75524 ( .A(n31512), .X(n49832) );
  inv_x2_sg U75525 ( .A(n31518), .X(n49827) );
  inv_x2_sg U75526 ( .A(n31531), .X(n49783) );
  inv_x2_sg U75527 ( .A(n31540), .X(n49790) );
  inv_x2_sg U75528 ( .A(n31553), .X(n49824) );
  inv_x2_sg U75529 ( .A(n25307), .X(n49286) );
  inv_x2_sg U75530 ( .A(n31599), .X(n49327) );
  inv_x2_sg U75531 ( .A(n31605), .X(n49371) );
  inv_x2_sg U75532 ( .A(n31611), .X(n49417) );
  inv_x2_sg U75533 ( .A(n31617), .X(n49463) );
  inv_x2_sg U75534 ( .A(n31623), .X(n49510) );
  inv_x2_sg U75535 ( .A(n31629), .X(n49557) );
  inv_x2_sg U75536 ( .A(n31635), .X(n49603) );
  inv_x2_sg U75537 ( .A(n31641), .X(n49650) );
  inv_x2_sg U75538 ( .A(n31647), .X(n49697) );
  inv_x2_sg U75539 ( .A(n31653), .X(n49746) );
  inv_x2_sg U75540 ( .A(n31659), .X(n49794) );
  inv_x2_sg U75541 ( .A(n45515), .X(n49745) );
  inv_x2_sg U75542 ( .A(n31665), .X(n49787) );
  inv_x2_sg U75543 ( .A(n31523), .X(n49734) );
  inv_x2_sg U75544 ( .A(n31684), .X(n49737) );
  inv_x2_sg U75545 ( .A(n31693), .X(n49744) );
  inv_x2_sg U75546 ( .A(n44621), .X(n49315) );
  inv_x2_sg U75547 ( .A(n31747), .X(n49314) );
  inv_x2_sg U75548 ( .A(n44505), .X(n49363) );
  inv_x2_sg U75549 ( .A(n31754), .X(n49362) );
  inv_x2_sg U75550 ( .A(n44507), .X(n49408) );
  inv_x2_sg U75551 ( .A(n31761), .X(n49407) );
  inv_x2_sg U75552 ( .A(n44509), .X(n49453) );
  inv_x2_sg U75553 ( .A(n31768), .X(n49452) );
  inv_x2_sg U75554 ( .A(n44511), .X(n49499) );
  inv_x2_sg U75555 ( .A(n31775), .X(n49498) );
  inv_x2_sg U75556 ( .A(n44513), .X(n49547) );
  inv_x2_sg U75557 ( .A(n31782), .X(n49546) );
  inv_x2_sg U75558 ( .A(n44515), .X(n49593) );
  inv_x2_sg U75559 ( .A(n31789), .X(n49592) );
  inv_x2_sg U75560 ( .A(n44517), .X(n49639) );
  inv_x2_sg U75561 ( .A(n31796), .X(n49638) );
  inv_x2_sg U75562 ( .A(n44666), .X(n49686) );
  inv_x2_sg U75563 ( .A(n31803), .X(n49685) );
  inv_x2_sg U75564 ( .A(n45523), .X(n49733) );
  inv_x2_sg U75565 ( .A(n31809), .X(n49741) );
  inv_x2_sg U75566 ( .A(n31815), .X(n49736) );
  inv_x2_sg U75567 ( .A(n31828), .X(n49691) );
  inv_x2_sg U75568 ( .A(n31837), .X(n49732) );
  inv_x2_sg U75569 ( .A(n31925), .X(n49695) );
  inv_x2_sg U75570 ( .A(n31820), .X(n49643) );
  inv_x2_sg U75571 ( .A(n31944), .X(n49646) );
  inv_x2_sg U75572 ( .A(n44245), .X(n49319) );
  inv_x2_sg U75573 ( .A(n31988), .X(n49318) );
  inv_x2_sg U75574 ( .A(n31994), .X(n49367) );
  inv_x2_sg U75575 ( .A(n32000), .X(n49412) );
  inv_x2_sg U75576 ( .A(n45489), .X(n49458) );
  inv_x2_sg U75577 ( .A(n32007), .X(n49457) );
  inv_x2_sg U75578 ( .A(n32013), .X(n49503) );
  inv_x2_sg U75579 ( .A(n45491), .X(n49552) );
  inv_x2_sg U75580 ( .A(n32020), .X(n49551) );
  inv_x2_sg U75581 ( .A(n32033), .X(n49645) );
  inv_x2_sg U75582 ( .A(n32036), .X(n49597) );
  inv_x2_sg U75583 ( .A(n32024), .X(n49600) );
  inv_x2_sg U75584 ( .A(n32100), .X(n49506) );
  inv_x2_sg U75585 ( .A(n32111), .X(n49599) );
  inv_x2_sg U75586 ( .A(n32127), .X(n49321) );
  inv_x2_sg U75587 ( .A(n32107), .X(n49505) );
  inv_x2_sg U75588 ( .A(n31504), .X(n49842) );
  inv_x2_sg U75589 ( .A(n21228), .X(n55439) );
  inv_x2_sg U75590 ( .A(n21758), .X(n55448) );
  inv_x2_sg U75591 ( .A(n21767), .X(n55446) );
  inv_x2_sg U75592 ( .A(n21803), .X(n55441) );
  inv_x2_sg U75593 ( .A(n21813), .X(n55404) );
  inv_x2_sg U75594 ( .A(n21815), .X(n55359) );
  inv_x2_sg U75595 ( .A(n21840), .X(n55440) );
  inv_x2_sg U75596 ( .A(n21839), .X(n55418) );
  inv_x2_sg U75597 ( .A(n21691), .X(n55436) );
  inv_x2_sg U75598 ( .A(n21742), .X(n55358) );
  inv_x2_sg U75599 ( .A(n21748), .X(n55371) );
  inv_x2_sg U75600 ( .A(n45415), .X(n55372) );
  inv_x2_sg U75601 ( .A(n21750), .X(n55432) );
  inv_x2_sg U75602 ( .A(n21922), .X(n55431) );
  inv_x2_sg U75603 ( .A(n21232), .X(n55433) );
  inv_x2_sg U75604 ( .A(n21235), .X(n55434) );
  inv_x2_sg U75605 ( .A(n21861), .X(n55382) );
  inv_x2_sg U75606 ( .A(n21773), .X(n55402) );
  inv_x2_sg U75607 ( .A(n21755), .X(n55416) );
  inv_x2_sg U75608 ( .A(n21242), .X(n55437) );
  inv_x2_sg U75609 ( .A(n21631), .X(n55421) );
  inv_x2_sg U75610 ( .A(n21731), .X(n55390) );
  inv_x2_sg U75611 ( .A(n21871), .X(n55259) );
  inv_x2_sg U75612 ( .A(n29528), .X(n55407) );
  inv_x2_sg U75613 ( .A(n21864), .X(n55346) );
  inv_x2_sg U75614 ( .A(n21637), .X(n55420) );
  inv_x2_sg U75615 ( .A(n21213), .X(n55401) );
  inv_x2_sg U75616 ( .A(n21585), .X(n55380) );
  inv_x2_sg U75617 ( .A(n21629), .X(n55395) );
  inv_x2_sg U75618 ( .A(n21720), .X(n55260) );
  inv_x2_sg U75619 ( .A(n21904), .X(n55391) );
  inv_x2_sg U75620 ( .A(n29435), .X(n55385) );
  inv_x2_sg U75621 ( .A(n21905), .X(n55245) );
  inv_x2_sg U75622 ( .A(n21882), .X(n55295) );
  inv_x2_sg U75623 ( .A(n21584), .X(n55398) );
  inv_x2_sg U75624 ( .A(n21685), .X(n55377) );
  inv_x2_sg U75625 ( .A(n21555), .X(n55365) );
  inv_x2_sg U75626 ( .A(n21670), .X(n55258) );
  inv_x2_sg U75627 ( .A(n29441), .X(n55361) );
  inv_x2_sg U75628 ( .A(n21709), .X(n55303) );
  inv_x2_sg U75629 ( .A(n21710), .X(n55330) );
  inv_x2_sg U75630 ( .A(n21647), .X(n55336) );
  inv_x2_sg U75631 ( .A(n21548), .X(n55357) );
  inv_x2_sg U75632 ( .A(n21205), .X(n55356) );
  inv_x2_sg U75633 ( .A(n21574), .X(n55292) );
  inv_x2_sg U75634 ( .A(n29447), .X(n55343) );
  inv_x2_sg U75635 ( .A(n21652), .X(n55347) );
  inv_x2_sg U75636 ( .A(n21610), .X(n55314) );
  inv_x2_sg U75637 ( .A(n21459), .X(n55311) );
  inv_x2_sg U75638 ( .A(n21508), .X(n55301) );
  inv_x2_sg U75639 ( .A(n21488), .X(n55302) );
  inv_x2_sg U75640 ( .A(n21468), .X(n55291) );
  inv_x2_sg U75641 ( .A(n44078), .X(n55312) );
  inv_x2_sg U75642 ( .A(n21534), .X(n55323) );
  inv_x2_sg U75643 ( .A(n29453), .X(n55318) );
  inv_x2_sg U75644 ( .A(n21467), .X(n55325) );
  inv_x2_sg U75645 ( .A(n21252), .X(n55327) );
  inv_x2_sg U75646 ( .A(n21191), .X(n55287) );
  inv_x2_sg U75647 ( .A(n21426), .X(n55309) );
  inv_x2_sg U75648 ( .A(n29459), .X(n55298) );
  inv_x2_sg U75649 ( .A(n21517), .X(n55241) );
  inv_x2_sg U75650 ( .A(n21518), .X(n55230) );
  inv_x2_sg U75651 ( .A(n21476), .X(n55242) );
  inv_x2_sg U75652 ( .A(n21471), .X(n55282) );
  inv_x2_sg U75653 ( .A(n21203), .X(n55310) );
  inv_x2_sg U75654 ( .A(n21373), .X(n55285) );
  inv_x2_sg U75655 ( .A(n21410), .X(n55262) );
  inv_x2_sg U75656 ( .A(n21394), .X(n55261) );
  inv_x2_sg U75657 ( .A(n21422), .X(n55283) );
  inv_x2_sg U75658 ( .A(n21188), .X(n55267) );
  inv_x2_sg U75659 ( .A(n21343), .X(n55252) );
  inv_x2_sg U75660 ( .A(n21372), .X(n55265) );
  inv_x2_sg U75661 ( .A(n29469), .X(n55255) );
  inv_x2_sg U75662 ( .A(n21365), .X(n55209) );
  inv_x2_sg U75663 ( .A(n21409), .X(n55221) );
  inv_x2_sg U75664 ( .A(n21418), .X(n55229) );
  inv_x2_sg U75665 ( .A(n21323), .X(n55249) );
  inv_x2_sg U75666 ( .A(n21354), .X(n55247) );
  inv_x2_sg U75667 ( .A(n21330), .X(n55231) );
  inv_x2_sg U75668 ( .A(n29485), .X(n55226) );
  inv_x2_sg U75669 ( .A(n21324), .X(n55220) );
  inv_x2_sg U75670 ( .A(n21281), .X(n55205) );
  inv_x2_sg U75671 ( .A(n21306), .X(n55216) );
  inv_x2_sg U75672 ( .A(n21305), .X(n55211) );
  inv_x2_sg U75673 ( .A(n29495), .X(n55193) );
  inv_x2_sg U75674 ( .A(n21293), .X(n55203) );
  inv_x2_sg U75675 ( .A(n21271), .X(n55196) );
  inv_x2_sg U75676 ( .A(n29501), .X(n55186) );
  inv_x2_sg U75677 ( .A(n29507), .X(n55180) );
  inv_x2_sg U75678 ( .A(n44267), .X(n55181) );
  inv_x2_sg U75679 ( .A(n46025), .X(n51233) );
  inv_x2_sg U75680 ( .A(n44875), .X(n55175) );
  inv_x2_sg U75681 ( .A(n20455), .X(n55155) );
  inv_x2_sg U75682 ( .A(n20988), .X(n55164) );
  inv_x2_sg U75683 ( .A(n20997), .X(n55162) );
  inv_x2_sg U75684 ( .A(n21032), .X(n55157) );
  inv_x2_sg U75685 ( .A(n21042), .X(n55119) );
  inv_x2_sg U75686 ( .A(n21044), .X(n55061) );
  inv_x2_sg U75687 ( .A(n21069), .X(n55156) );
  inv_x2_sg U75688 ( .A(n21068), .X(n55133) );
  inv_x2_sg U75689 ( .A(n20922), .X(n55151) );
  inv_x2_sg U75690 ( .A(n20972), .X(n55074) );
  inv_x2_sg U75691 ( .A(n20980), .X(n55147) );
  inv_x2_sg U75692 ( .A(n21149), .X(n55146) );
  inv_x2_sg U75693 ( .A(n20459), .X(n55148) );
  inv_x2_sg U75694 ( .A(n20463), .X(n55149) );
  inv_x2_sg U75695 ( .A(n21090), .X(n55097) );
  inv_x2_sg U75696 ( .A(n21003), .X(n55117) );
  inv_x2_sg U75697 ( .A(n20985), .X(n55131) );
  inv_x2_sg U75698 ( .A(n20470), .X(n55152) );
  inv_x2_sg U75699 ( .A(n20862), .X(n55136) );
  inv_x2_sg U75700 ( .A(n20962), .X(n55105) );
  inv_x2_sg U75701 ( .A(n20934), .X(n55056) );
  inv_x2_sg U75702 ( .A(n21100), .X(n54980) );
  inv_x2_sg U75703 ( .A(n21134), .X(n55116) );
  inv_x2_sg U75704 ( .A(n21140), .X(n55127) );
  inv_x2_sg U75705 ( .A(n29250), .X(n55122) );
  inv_x2_sg U75706 ( .A(n21093), .X(n55062) );
  inv_x2_sg U75707 ( .A(n20868), .X(n55135) );
  inv_x2_sg U75708 ( .A(n20440), .X(n55115) );
  inv_x2_sg U75709 ( .A(n20815), .X(n55095) );
  inv_x2_sg U75710 ( .A(n20860), .X(n55109) );
  inv_x2_sg U75711 ( .A(n21132), .X(n55106) );
  inv_x2_sg U75712 ( .A(n29155), .X(n55100) );
  inv_x2_sg U75713 ( .A(n21133), .X(n54973) );
  inv_x2_sg U75714 ( .A(n20951), .X(n55107) );
  inv_x2_sg U75715 ( .A(n20814), .X(n55112) );
  inv_x2_sg U75716 ( .A(n20916), .X(n55092) );
  inv_x2_sg U75717 ( .A(n20785), .X(n55080) );
  inv_x2_sg U75718 ( .A(n20901), .X(n55000) );
  inv_x2_sg U75719 ( .A(n20902), .X(n54979) );
  inv_x2_sg U75720 ( .A(n29161), .X(n55076) );
  inv_x2_sg U75721 ( .A(n20940), .X(n55020) );
  inv_x2_sg U75722 ( .A(n20941), .X(n55037) );
  inv_x2_sg U75723 ( .A(n20878), .X(n55050) );
  inv_x2_sg U75724 ( .A(n20778), .X(n55073) );
  inv_x2_sg U75725 ( .A(n20432), .X(n55072) );
  inv_x2_sg U75726 ( .A(n20804), .X(n55011) );
  inv_x2_sg U75727 ( .A(n29167), .X(n55058) );
  inv_x2_sg U75728 ( .A(n20883), .X(n55063) );
  inv_x2_sg U75729 ( .A(n20841), .X(n55032) );
  inv_x2_sg U75730 ( .A(n20689), .X(n55029) );
  inv_x2_sg U75731 ( .A(n20738), .X(n55018) );
  inv_x2_sg U75732 ( .A(n20718), .X(n55019) );
  inv_x2_sg U75733 ( .A(n20698), .X(n54999) );
  inv_x2_sg U75734 ( .A(n20749), .X(n55030) );
  inv_x2_sg U75735 ( .A(n29173), .X(n55035) );
  inv_x2_sg U75736 ( .A(n20697), .X(n55043) );
  inv_x2_sg U75737 ( .A(n20480), .X(n55045) );
  inv_x2_sg U75738 ( .A(n20418), .X(n55008) );
  inv_x2_sg U75739 ( .A(n20655), .X(n55027) );
  inv_x2_sg U75740 ( .A(n29179), .X(n55015) );
  inv_x2_sg U75741 ( .A(n20747), .X(n54969) );
  inv_x2_sg U75742 ( .A(n20748), .X(n54957) );
  inv_x2_sg U75743 ( .A(n20706), .X(n54970) );
  inv_x2_sg U75744 ( .A(n20701), .X(n55010) );
  inv_x2_sg U75745 ( .A(n20430), .X(n55028) );
  inv_x2_sg U75746 ( .A(n20602), .X(n55006) );
  inv_x2_sg U75747 ( .A(n20639), .X(n54983) );
  inv_x2_sg U75748 ( .A(n20623), .X(n54982) );
  inv_x2_sg U75749 ( .A(n29185), .X(n54994) );
  inv_x2_sg U75750 ( .A(n20652), .X(n55004) );
  inv_x2_sg U75751 ( .A(n20415), .X(n54988) );
  inv_x2_sg U75752 ( .A(n20574), .X(n54967) );
  inv_x2_sg U75753 ( .A(n20601), .X(n54986) );
  inv_x2_sg U75754 ( .A(n29191), .X(n54976) );
  inv_x2_sg U75755 ( .A(n20594), .X(n54929) );
  inv_x2_sg U75756 ( .A(n20638), .X(n54942) );
  inv_x2_sg U75757 ( .A(n20647), .X(n54956) );
  inv_x2_sg U75758 ( .A(n20555), .X(n54964) );
  inv_x2_sg U75759 ( .A(n20576), .X(n54955) );
  inv_x2_sg U75760 ( .A(n20581), .X(n54941) );
  inv_x2_sg U75761 ( .A(n20585), .X(n54962) );
  inv_x2_sg U75762 ( .A(n20549), .X(n54951) );
  inv_x2_sg U75763 ( .A(n29205), .X(n54946) );
  inv_x2_sg U75764 ( .A(n20556), .X(n54940) );
  inv_x2_sg U75765 ( .A(n20511), .X(n54925) );
  inv_x2_sg U75766 ( .A(n20538), .X(n54936) );
  inv_x2_sg U75767 ( .A(n29209), .X(n54934) );
  inv_x2_sg U75768 ( .A(n20537), .X(n54931) );
  inv_x2_sg U75769 ( .A(n29217), .X(n54920) );
  inv_x2_sg U75770 ( .A(n20524), .X(n54923) );
  inv_x2_sg U75771 ( .A(n20489), .X(n54927) );
  inv_x2_sg U75772 ( .A(n29223), .X(n54902) );
  inv_x2_sg U75773 ( .A(n29229), .X(n54896) );
  inv_x2_sg U75774 ( .A(n20386), .X(n54899) );
  inv_x2_sg U75775 ( .A(n44251), .X(n54897) );
  inv_x2_sg U75776 ( .A(n46001), .X(n51214) );
  inv_x2_sg U75777 ( .A(n44827), .X(n54891) );
  inv_x2_sg U75778 ( .A(n19683), .X(n54871) );
  inv_x2_sg U75779 ( .A(n20213), .X(n54880) );
  inv_x2_sg U75780 ( .A(n20222), .X(n54878) );
  inv_x2_sg U75781 ( .A(n20258), .X(n54873) );
  inv_x2_sg U75782 ( .A(n20268), .X(n54836) );
  inv_x2_sg U75783 ( .A(n20270), .X(n54791) );
  inv_x2_sg U75784 ( .A(n20295), .X(n54872) );
  inv_x2_sg U75785 ( .A(n20294), .X(n54850) );
  inv_x2_sg U75786 ( .A(n20146), .X(n54868) );
  inv_x2_sg U75787 ( .A(n20197), .X(n54790) );
  inv_x2_sg U75788 ( .A(n20203), .X(n54803) );
  inv_x2_sg U75789 ( .A(n45417), .X(n54804) );
  inv_x2_sg U75790 ( .A(n20205), .X(n54864) );
  inv_x2_sg U75791 ( .A(n20377), .X(n54863) );
  inv_x2_sg U75792 ( .A(n19687), .X(n54865) );
  inv_x2_sg U75793 ( .A(n19690), .X(n54866) );
  inv_x2_sg U75794 ( .A(n20316), .X(n54814) );
  inv_x2_sg U75795 ( .A(n20228), .X(n54834) );
  inv_x2_sg U75796 ( .A(n20210), .X(n54848) );
  inv_x2_sg U75797 ( .A(n19697), .X(n54869) );
  inv_x2_sg U75798 ( .A(n20086), .X(n54853) );
  inv_x2_sg U75799 ( .A(n20186), .X(n54822) );
  inv_x2_sg U75800 ( .A(n20326), .X(n54691) );
  inv_x2_sg U75801 ( .A(n28967), .X(n54839) );
  inv_x2_sg U75802 ( .A(n20319), .X(n54778) );
  inv_x2_sg U75803 ( .A(n20092), .X(n54852) );
  inv_x2_sg U75804 ( .A(n19668), .X(n54833) );
  inv_x2_sg U75805 ( .A(n20040), .X(n54812) );
  inv_x2_sg U75806 ( .A(n20084), .X(n54827) );
  inv_x2_sg U75807 ( .A(n20175), .X(n54692) );
  inv_x2_sg U75808 ( .A(n20359), .X(n54823) );
  inv_x2_sg U75809 ( .A(n28874), .X(n54817) );
  inv_x2_sg U75810 ( .A(n20360), .X(n54677) );
  inv_x2_sg U75811 ( .A(n20337), .X(n54727) );
  inv_x2_sg U75812 ( .A(n20039), .X(n54830) );
  inv_x2_sg U75813 ( .A(n20140), .X(n54809) );
  inv_x2_sg U75814 ( .A(n20010), .X(n54797) );
  inv_x2_sg U75815 ( .A(n20125), .X(n54690) );
  inv_x2_sg U75816 ( .A(n28880), .X(n54793) );
  inv_x2_sg U75817 ( .A(n20164), .X(n54735) );
  inv_x2_sg U75818 ( .A(n20165), .X(n54762) );
  inv_x2_sg U75819 ( .A(n20102), .X(n54768) );
  inv_x2_sg U75820 ( .A(n20003), .X(n54789) );
  inv_x2_sg U75821 ( .A(n19660), .X(n54788) );
  inv_x2_sg U75822 ( .A(n20029), .X(n54724) );
  inv_x2_sg U75823 ( .A(n28886), .X(n54775) );
  inv_x2_sg U75824 ( .A(n20107), .X(n54779) );
  inv_x2_sg U75825 ( .A(n20065), .X(n54746) );
  inv_x2_sg U75826 ( .A(n19914), .X(n54743) );
  inv_x2_sg U75827 ( .A(n19963), .X(n54733) );
  inv_x2_sg U75828 ( .A(n19943), .X(n54734) );
  inv_x2_sg U75829 ( .A(n19923), .X(n54723) );
  inv_x2_sg U75830 ( .A(n44080), .X(n54744) );
  inv_x2_sg U75831 ( .A(n19989), .X(n54755) );
  inv_x2_sg U75832 ( .A(n28892), .X(n54750) );
  inv_x2_sg U75833 ( .A(n19922), .X(n54757) );
  inv_x2_sg U75834 ( .A(n19707), .X(n54759) );
  inv_x2_sg U75835 ( .A(n19646), .X(n54719) );
  inv_x2_sg U75836 ( .A(n19881), .X(n54741) );
  inv_x2_sg U75837 ( .A(n28898), .X(n54730) );
  inv_x2_sg U75838 ( .A(n19972), .X(n54673) );
  inv_x2_sg U75839 ( .A(n19973), .X(n54662) );
  inv_x2_sg U75840 ( .A(n19931), .X(n54674) );
  inv_x2_sg U75841 ( .A(n19926), .X(n54714) );
  inv_x2_sg U75842 ( .A(n19658), .X(n54742) );
  inv_x2_sg U75843 ( .A(n19828), .X(n54717) );
  inv_x2_sg U75844 ( .A(n19865), .X(n54694) );
  inv_x2_sg U75845 ( .A(n19849), .X(n54693) );
  inv_x2_sg U75846 ( .A(n19877), .X(n54715) );
  inv_x2_sg U75847 ( .A(n19643), .X(n54699) );
  inv_x2_sg U75848 ( .A(n19798), .X(n54684) );
  inv_x2_sg U75849 ( .A(n19827), .X(n54697) );
  inv_x2_sg U75850 ( .A(n28908), .X(n54687) );
  inv_x2_sg U75851 ( .A(n19820), .X(n54641) );
  inv_x2_sg U75852 ( .A(n19864), .X(n54653) );
  inv_x2_sg U75853 ( .A(n19873), .X(n54661) );
  inv_x2_sg U75854 ( .A(n19778), .X(n54681) );
  inv_x2_sg U75855 ( .A(n19809), .X(n54679) );
  inv_x2_sg U75856 ( .A(n19785), .X(n54663) );
  inv_x2_sg U75857 ( .A(n28924), .X(n54658) );
  inv_x2_sg U75858 ( .A(n19779), .X(n54652) );
  inv_x2_sg U75859 ( .A(n19736), .X(n54637) );
  inv_x2_sg U75860 ( .A(n19761), .X(n54648) );
  inv_x2_sg U75861 ( .A(n19760), .X(n54643) );
  inv_x2_sg U75862 ( .A(n28934), .X(n54625) );
  inv_x2_sg U75863 ( .A(n19748), .X(n54635) );
  inv_x2_sg U75864 ( .A(n19726), .X(n54628) );
  inv_x2_sg U75865 ( .A(n28940), .X(n54618) );
  inv_x2_sg U75866 ( .A(n28946), .X(n54612) );
  inv_x2_sg U75867 ( .A(n44263), .X(n54613) );
  inv_x2_sg U75868 ( .A(n46021), .X(n51195) );
  inv_x2_sg U75869 ( .A(n44863), .X(n54607) );
  inv_x2_sg U75870 ( .A(n18911), .X(n54587) );
  inv_x2_sg U75871 ( .A(n19444), .X(n54596) );
  inv_x2_sg U75872 ( .A(n19453), .X(n54594) );
  inv_x2_sg U75873 ( .A(n19488), .X(n54589) );
  inv_x2_sg U75874 ( .A(n19498), .X(n54551) );
  inv_x2_sg U75875 ( .A(n19500), .X(n54493) );
  inv_x2_sg U75876 ( .A(n19525), .X(n54588) );
  inv_x2_sg U75877 ( .A(n19524), .X(n54565) );
  inv_x2_sg U75878 ( .A(n19378), .X(n54583) );
  inv_x2_sg U75879 ( .A(n19428), .X(n54506) );
  inv_x2_sg U75880 ( .A(n19436), .X(n54579) );
  inv_x2_sg U75881 ( .A(n19605), .X(n54578) );
  inv_x2_sg U75882 ( .A(n18915), .X(n54580) );
  inv_x2_sg U75883 ( .A(n18919), .X(n54581) );
  inv_x2_sg U75884 ( .A(n19546), .X(n54529) );
  inv_x2_sg U75885 ( .A(n19459), .X(n54549) );
  inv_x2_sg U75886 ( .A(n19441), .X(n54563) );
  inv_x2_sg U75887 ( .A(n18926), .X(n54584) );
  inv_x2_sg U75888 ( .A(n19318), .X(n54568) );
  inv_x2_sg U75889 ( .A(n19418), .X(n54537) );
  inv_x2_sg U75890 ( .A(n19390), .X(n54488) );
  inv_x2_sg U75891 ( .A(n19556), .X(n54412) );
  inv_x2_sg U75892 ( .A(n19590), .X(n54548) );
  inv_x2_sg U75893 ( .A(n19596), .X(n54559) );
  inv_x2_sg U75894 ( .A(n28689), .X(n54554) );
  inv_x2_sg U75895 ( .A(n19549), .X(n54494) );
  inv_x2_sg U75896 ( .A(n19324), .X(n54567) );
  inv_x2_sg U75897 ( .A(n18896), .X(n54547) );
  inv_x2_sg U75898 ( .A(n19271), .X(n54527) );
  inv_x2_sg U75899 ( .A(n19316), .X(n54541) );
  inv_x2_sg U75900 ( .A(n19588), .X(n54538) );
  inv_x2_sg U75901 ( .A(n28594), .X(n54532) );
  inv_x2_sg U75902 ( .A(n19589), .X(n54405) );
  inv_x2_sg U75903 ( .A(n19407), .X(n54539) );
  inv_x2_sg U75904 ( .A(n19270), .X(n54544) );
  inv_x2_sg U75905 ( .A(n19372), .X(n54524) );
  inv_x2_sg U75906 ( .A(n19241), .X(n54512) );
  inv_x2_sg U75907 ( .A(n19357), .X(n54432) );
  inv_x2_sg U75908 ( .A(n19358), .X(n54411) );
  inv_x2_sg U75909 ( .A(n28600), .X(n54508) );
  inv_x2_sg U75910 ( .A(n19396), .X(n54452) );
  inv_x2_sg U75911 ( .A(n19397), .X(n54469) );
  inv_x2_sg U75912 ( .A(n19334), .X(n54482) );
  inv_x2_sg U75913 ( .A(n19234), .X(n54505) );
  inv_x2_sg U75914 ( .A(n18888), .X(n54504) );
  inv_x2_sg U75915 ( .A(n19260), .X(n54443) );
  inv_x2_sg U75916 ( .A(n28606), .X(n54490) );
  inv_x2_sg U75917 ( .A(n19339), .X(n54495) );
  inv_x2_sg U75918 ( .A(n19297), .X(n54464) );
  inv_x2_sg U75919 ( .A(n19145), .X(n54461) );
  inv_x2_sg U75920 ( .A(n19194), .X(n54450) );
  inv_x2_sg U75921 ( .A(n19174), .X(n54451) );
  inv_x2_sg U75922 ( .A(n19154), .X(n54431) );
  inv_x2_sg U75923 ( .A(n19205), .X(n54462) );
  inv_x2_sg U75924 ( .A(n28612), .X(n54467) );
  inv_x2_sg U75925 ( .A(n19153), .X(n54475) );
  inv_x2_sg U75926 ( .A(n18936), .X(n54477) );
  inv_x2_sg U75927 ( .A(n18874), .X(n54440) );
  inv_x2_sg U75928 ( .A(n19111), .X(n54459) );
  inv_x2_sg U75929 ( .A(n28618), .X(n54447) );
  inv_x2_sg U75930 ( .A(n19203), .X(n54401) );
  inv_x2_sg U75931 ( .A(n19204), .X(n54389) );
  inv_x2_sg U75932 ( .A(n19162), .X(n54402) );
  inv_x2_sg U75933 ( .A(n19157), .X(n54442) );
  inv_x2_sg U75934 ( .A(n18886), .X(n54460) );
  inv_x2_sg U75935 ( .A(n19058), .X(n54438) );
  inv_x2_sg U75936 ( .A(n19095), .X(n54415) );
  inv_x2_sg U75937 ( .A(n19079), .X(n54414) );
  inv_x2_sg U75938 ( .A(n28624), .X(n54426) );
  inv_x2_sg U75939 ( .A(n19108), .X(n54436) );
  inv_x2_sg U75940 ( .A(n18871), .X(n54420) );
  inv_x2_sg U75941 ( .A(n19030), .X(n54399) );
  inv_x2_sg U75942 ( .A(n19057), .X(n54418) );
  inv_x2_sg U75943 ( .A(n28630), .X(n54408) );
  inv_x2_sg U75944 ( .A(n19050), .X(n54361) );
  inv_x2_sg U75945 ( .A(n19094), .X(n54374) );
  inv_x2_sg U75946 ( .A(n19103), .X(n54388) );
  inv_x2_sg U75947 ( .A(n19011), .X(n54396) );
  inv_x2_sg U75948 ( .A(n19032), .X(n54387) );
  inv_x2_sg U75949 ( .A(n19037), .X(n54373) );
  inv_x2_sg U75950 ( .A(n19041), .X(n54394) );
  inv_x2_sg U75951 ( .A(n19005), .X(n54383) );
  inv_x2_sg U75952 ( .A(n28644), .X(n54378) );
  inv_x2_sg U75953 ( .A(n19012), .X(n54372) );
  inv_x2_sg U75954 ( .A(n18967), .X(n54357) );
  inv_x2_sg U75955 ( .A(n18994), .X(n54368) );
  inv_x2_sg U75956 ( .A(n28648), .X(n54366) );
  inv_x2_sg U75957 ( .A(n18993), .X(n54363) );
  inv_x2_sg U75958 ( .A(n28656), .X(n54352) );
  inv_x2_sg U75959 ( .A(n18980), .X(n54355) );
  inv_x2_sg U75960 ( .A(n18945), .X(n54359) );
  inv_x2_sg U75961 ( .A(n28662), .X(n54334) );
  inv_x2_sg U75962 ( .A(n28668), .X(n54328) );
  inv_x2_sg U75963 ( .A(n18842), .X(n54331) );
  inv_x2_sg U75964 ( .A(n44253), .X(n54329) );
  inv_x2_sg U75965 ( .A(n46003), .X(n51176) );
  inv_x2_sg U75966 ( .A(n44829), .X(n54323) );
  inv_x2_sg U75967 ( .A(n18138), .X(n54303) );
  inv_x2_sg U75968 ( .A(n18668), .X(n54312) );
  inv_x2_sg U75969 ( .A(n18677), .X(n54310) );
  inv_x2_sg U75970 ( .A(n18712), .X(n54305) );
  inv_x2_sg U75971 ( .A(n18722), .X(n54269) );
  inv_x2_sg U75972 ( .A(n18724), .X(n54224) );
  inv_x2_sg U75973 ( .A(n18749), .X(n54304) );
  inv_x2_sg U75974 ( .A(n18748), .X(n54283) );
  inv_x2_sg U75975 ( .A(n18600), .X(n54300) );
  inv_x2_sg U75976 ( .A(n18658), .X(n54238) );
  inv_x2_sg U75977 ( .A(n44329), .X(n54239) );
  inv_x2_sg U75978 ( .A(n18660), .X(n54296) );
  inv_x2_sg U75979 ( .A(n18832), .X(n54295) );
  inv_x2_sg U75980 ( .A(n18142), .X(n54297) );
  inv_x2_sg U75981 ( .A(n18145), .X(n54298) );
  inv_x2_sg U75982 ( .A(n18683), .X(n54267) );
  inv_x2_sg U75983 ( .A(n18779), .X(n54246) );
  inv_x2_sg U75984 ( .A(n18790), .X(n54253) );
  inv_x2_sg U75985 ( .A(n18665), .X(n54281) );
  inv_x2_sg U75986 ( .A(n18152), .X(n54301) );
  inv_x2_sg U75987 ( .A(n18541), .X(n54285) );
  inv_x2_sg U75988 ( .A(n18640), .X(n54255) );
  inv_x2_sg U75989 ( .A(n18798), .X(n54254) );
  inv_x2_sg U75990 ( .A(n18599), .X(n54279) );
  inv_x2_sg U75991 ( .A(n28410), .X(n54272) );
  inv_x2_sg U75992 ( .A(n18547), .X(n54284) );
  inv_x2_sg U75993 ( .A(n18123), .X(n54266) );
  inv_x2_sg U75994 ( .A(n18495), .X(n54244) );
  inv_x2_sg U75995 ( .A(n18539), .X(n54260) );
  inv_x2_sg U75996 ( .A(n18629), .X(n54129) );
  inv_x2_sg U75997 ( .A(n18814), .X(n54256) );
  inv_x2_sg U75998 ( .A(n28317), .X(n54249) );
  inv_x2_sg U75999 ( .A(n18815), .X(n54114) );
  inv_x2_sg U76000 ( .A(n18793), .X(n54161) );
  inv_x2_sg U76001 ( .A(n18494), .X(n54263) );
  inv_x2_sg U76002 ( .A(n18465), .X(n54232) );
  inv_x2_sg U76003 ( .A(n18579), .X(n54127) );
  inv_x2_sg U76004 ( .A(n28323), .X(n54228) );
  inv_x2_sg U76005 ( .A(n18618), .X(n54169) );
  inv_x2_sg U76006 ( .A(n18619), .X(n54195) );
  inv_x2_sg U76007 ( .A(n18458), .X(n54222) );
  inv_x2_sg U76008 ( .A(n18115), .X(n54219) );
  inv_x2_sg U76009 ( .A(n18484), .X(n54159) );
  inv_x2_sg U76010 ( .A(n18487), .X(n54211) );
  inv_x2_sg U76011 ( .A(n28329), .X(n54208) );
  inv_x2_sg U76012 ( .A(n18467), .X(n54212) );
  inv_x2_sg U76013 ( .A(n18520), .X(n54179) );
  inv_x2_sg U76014 ( .A(n18369), .X(n54176) );
  inv_x2_sg U76015 ( .A(n18418), .X(n54167) );
  inv_x2_sg U76016 ( .A(n18398), .X(n54168) );
  inv_x2_sg U76017 ( .A(n18378), .X(n54158) );
  inv_x2_sg U76018 ( .A(n18429), .X(n54177) );
  inv_x2_sg U76019 ( .A(n18444), .X(n54188) );
  inv_x2_sg U76020 ( .A(n28335), .X(n54183) );
  inv_x2_sg U76021 ( .A(n18377), .X(n54190) );
  inv_x2_sg U76022 ( .A(n18162), .X(n54192) );
  inv_x2_sg U76023 ( .A(n18101), .X(n54154) );
  inv_x2_sg U76024 ( .A(n18336), .X(n54175) );
  inv_x2_sg U76025 ( .A(n28341), .X(n54164) );
  inv_x2_sg U76026 ( .A(n18427), .X(n54110) );
  inv_x2_sg U76027 ( .A(n18428), .X(n54106) );
  inv_x2_sg U76028 ( .A(n18386), .X(n54111) );
  inv_x2_sg U76029 ( .A(n18381), .X(n54149) );
  inv_x2_sg U76030 ( .A(n18282), .X(n54152) );
  inv_x2_sg U76031 ( .A(n18321), .X(n54131) );
  inv_x2_sg U76032 ( .A(n18332), .X(n54150) );
  inv_x2_sg U76033 ( .A(n18098), .X(n54135) );
  inv_x2_sg U76034 ( .A(n18253), .X(n54121) );
  inv_x2_sg U76035 ( .A(n28351), .X(n54123) );
  inv_x2_sg U76036 ( .A(n18319), .X(n54077) );
  inv_x2_sg U76037 ( .A(n18320), .X(n54091) );
  inv_x2_sg U76038 ( .A(n18232), .X(n54118) );
  inv_x2_sg U76039 ( .A(n18264), .X(n54116) );
  inv_x2_sg U76040 ( .A(n18240), .X(n54099) );
  inv_x2_sg U76041 ( .A(n45983), .X(n51163) );
  inv_x2_sg U76042 ( .A(n28365), .X(n54096) );
  inv_x2_sg U76043 ( .A(n18233), .X(n54089) );
  inv_x2_sg U76044 ( .A(n18189), .X(n54073) );
  inv_x2_sg U76045 ( .A(n18215), .X(n54085) );
  inv_x2_sg U76046 ( .A(n28371), .X(n54067) );
  inv_x2_sg U76047 ( .A(n28373), .X(n54082) );
  inv_x2_sg U76048 ( .A(n18214), .X(n54079) );
  inv_x2_sg U76049 ( .A(n28377), .X(n54058) );
  inv_x2_sg U76050 ( .A(n45987), .X(n51161) );
  inv_x2_sg U76051 ( .A(n18201), .X(n54071) );
  inv_x2_sg U76052 ( .A(n18180), .X(n54060) );
  inv_x2_sg U76053 ( .A(n28381), .X(n54059) );
  inv_x2_sg U76054 ( .A(n46193), .X(n51159) );
  inv_x2_sg U76055 ( .A(n28395), .X(n54049) );
  inv_x2_sg U76056 ( .A(n45985), .X(n51158) );
  inv_x2_sg U76057 ( .A(n44815), .X(n54042) );
  inv_x2_sg U76058 ( .A(n17366), .X(n54022) );
  inv_x2_sg U76059 ( .A(n17899), .X(n54031) );
  inv_x2_sg U76060 ( .A(n17908), .X(n54029) );
  inv_x2_sg U76061 ( .A(n17943), .X(n54024) );
  inv_x2_sg U76062 ( .A(n17953), .X(n53986) );
  inv_x2_sg U76063 ( .A(n17955), .X(n53928) );
  inv_x2_sg U76064 ( .A(n17980), .X(n54023) );
  inv_x2_sg U76065 ( .A(n17979), .X(n54000) );
  inv_x2_sg U76066 ( .A(n17833), .X(n54018) );
  inv_x2_sg U76067 ( .A(n17883), .X(n53941) );
  inv_x2_sg U76068 ( .A(n17891), .X(n54014) );
  inv_x2_sg U76069 ( .A(n18060), .X(n54013) );
  inv_x2_sg U76070 ( .A(n17370), .X(n54015) );
  inv_x2_sg U76071 ( .A(n17374), .X(n54016) );
  inv_x2_sg U76072 ( .A(n18001), .X(n53964) );
  inv_x2_sg U76073 ( .A(n17914), .X(n53984) );
  inv_x2_sg U76074 ( .A(n17896), .X(n53998) );
  inv_x2_sg U76075 ( .A(n17381), .X(n54019) );
  inv_x2_sg U76076 ( .A(n17773), .X(n54003) );
  inv_x2_sg U76077 ( .A(n17873), .X(n53972) );
  inv_x2_sg U76078 ( .A(n17845), .X(n53923) );
  inv_x2_sg U76079 ( .A(n18011), .X(n53847) );
  inv_x2_sg U76080 ( .A(n18045), .X(n53983) );
  inv_x2_sg U76081 ( .A(n18051), .X(n53994) );
  inv_x2_sg U76082 ( .A(n28131), .X(n53989) );
  inv_x2_sg U76083 ( .A(n18004), .X(n53929) );
  inv_x2_sg U76084 ( .A(n17779), .X(n54002) );
  inv_x2_sg U76085 ( .A(n17351), .X(n53982) );
  inv_x2_sg U76086 ( .A(n17726), .X(n53962) );
  inv_x2_sg U76087 ( .A(n17771), .X(n53976) );
  inv_x2_sg U76088 ( .A(n18043), .X(n53973) );
  inv_x2_sg U76089 ( .A(n28036), .X(n53967) );
  inv_x2_sg U76090 ( .A(n18044), .X(n53840) );
  inv_x2_sg U76091 ( .A(n17862), .X(n53974) );
  inv_x2_sg U76092 ( .A(n17725), .X(n53979) );
  inv_x2_sg U76093 ( .A(n17827), .X(n53959) );
  inv_x2_sg U76094 ( .A(n17696), .X(n53947) );
  inv_x2_sg U76095 ( .A(n17812), .X(n53867) );
  inv_x2_sg U76096 ( .A(n17813), .X(n53846) );
  inv_x2_sg U76097 ( .A(n28042), .X(n53943) );
  inv_x2_sg U76098 ( .A(n17851), .X(n53887) );
  inv_x2_sg U76099 ( .A(n17852), .X(n53904) );
  inv_x2_sg U76100 ( .A(n17789), .X(n53917) );
  inv_x2_sg U76101 ( .A(n17689), .X(n53940) );
  inv_x2_sg U76102 ( .A(n17343), .X(n53939) );
  inv_x2_sg U76103 ( .A(n17715), .X(n53878) );
  inv_x2_sg U76104 ( .A(n28048), .X(n53925) );
  inv_x2_sg U76105 ( .A(n17794), .X(n53930) );
  inv_x2_sg U76106 ( .A(n17752), .X(n53899) );
  inv_x2_sg U76107 ( .A(n17600), .X(n53896) );
  inv_x2_sg U76108 ( .A(n17649), .X(n53885) );
  inv_x2_sg U76109 ( .A(n17629), .X(n53886) );
  inv_x2_sg U76110 ( .A(n17609), .X(n53866) );
  inv_x2_sg U76111 ( .A(n17660), .X(n53897) );
  inv_x2_sg U76112 ( .A(n28054), .X(n53902) );
  inv_x2_sg U76113 ( .A(n17608), .X(n53910) );
  inv_x2_sg U76114 ( .A(n17391), .X(n53912) );
  inv_x2_sg U76115 ( .A(n17329), .X(n53875) );
  inv_x2_sg U76116 ( .A(n17566), .X(n53894) );
  inv_x2_sg U76117 ( .A(n28060), .X(n53882) );
  inv_x2_sg U76118 ( .A(n17658), .X(n53836) );
  inv_x2_sg U76119 ( .A(n17659), .X(n53824) );
  inv_x2_sg U76120 ( .A(n17617), .X(n53837) );
  inv_x2_sg U76121 ( .A(n17612), .X(n53877) );
  inv_x2_sg U76122 ( .A(n17341), .X(n53895) );
  inv_x2_sg U76123 ( .A(n17513), .X(n53873) );
  inv_x2_sg U76124 ( .A(n17550), .X(n53850) );
  inv_x2_sg U76125 ( .A(n17534), .X(n53849) );
  inv_x2_sg U76126 ( .A(n28066), .X(n53861) );
  inv_x2_sg U76127 ( .A(n17563), .X(n53871) );
  inv_x2_sg U76128 ( .A(n17326), .X(n53855) );
  inv_x2_sg U76129 ( .A(n17485), .X(n53834) );
  inv_x2_sg U76130 ( .A(n17512), .X(n53853) );
  inv_x2_sg U76131 ( .A(n28072), .X(n53843) );
  inv_x2_sg U76132 ( .A(n17505), .X(n53796) );
  inv_x2_sg U76133 ( .A(n17549), .X(n53809) );
  inv_x2_sg U76134 ( .A(n17558), .X(n53823) );
  inv_x2_sg U76135 ( .A(n17466), .X(n53831) );
  inv_x2_sg U76136 ( .A(n17487), .X(n53822) );
  inv_x2_sg U76137 ( .A(n17492), .X(n53808) );
  inv_x2_sg U76138 ( .A(n17496), .X(n53829) );
  inv_x2_sg U76139 ( .A(n17460), .X(n53818) );
  inv_x2_sg U76140 ( .A(n28086), .X(n53813) );
  inv_x2_sg U76141 ( .A(n17467), .X(n53807) );
  inv_x2_sg U76142 ( .A(n17422), .X(n53792) );
  inv_x2_sg U76143 ( .A(n17449), .X(n53803) );
  inv_x2_sg U76144 ( .A(n28090), .X(n53801) );
  inv_x2_sg U76145 ( .A(n17448), .X(n53798) );
  inv_x2_sg U76146 ( .A(n28098), .X(n53787) );
  inv_x2_sg U76147 ( .A(n17435), .X(n53790) );
  inv_x2_sg U76148 ( .A(n17400), .X(n53794) );
  inv_x2_sg U76149 ( .A(n28104), .X(n53769) );
  inv_x2_sg U76150 ( .A(n28110), .X(n53763) );
  inv_x2_sg U76151 ( .A(n17297), .X(n53766) );
  inv_x2_sg U76152 ( .A(n44255), .X(n53764) );
  inv_x2_sg U76153 ( .A(n46005), .X(n51139) );
  inv_x2_sg U76154 ( .A(n44831), .X(n53758) );
  inv_x2_sg U76155 ( .A(n16583), .X(n53740) );
  inv_x2_sg U76156 ( .A(n17126), .X(n53747) );
  inv_x2_sg U76157 ( .A(n17135), .X(n53745) );
  inv_x2_sg U76158 ( .A(n17163), .X(n53686) );
  inv_x2_sg U76159 ( .A(n17170), .X(n53735) );
  inv_x2_sg U76160 ( .A(n17182), .X(n53655) );
  inv_x2_sg U76161 ( .A(n17207), .X(n53734) );
  inv_x2_sg U76162 ( .A(n17206), .X(n53720) );
  inv_x2_sg U76163 ( .A(n17060), .X(n53736) );
  inv_x2_sg U76164 ( .A(n17110), .X(n53660) );
  inv_x2_sg U76165 ( .A(n17179), .X(n53712) );
  inv_x2_sg U76166 ( .A(n17124), .X(n53718) );
  inv_x2_sg U76167 ( .A(n16598), .X(n53737) );
  inv_x2_sg U76168 ( .A(n17002), .X(n53722) );
  inv_x2_sg U76169 ( .A(n17092), .X(n53679) );
  inv_x2_sg U76170 ( .A(n17059), .X(n53715) );
  inv_x2_sg U76171 ( .A(n17268), .X(n53704) );
  inv_x2_sg U76172 ( .A(n17274), .X(n53713) );
  inv_x2_sg U76173 ( .A(n27850), .X(n53709) );
  inv_x2_sg U76174 ( .A(n17008), .X(n53721) );
  inv_x2_sg U76175 ( .A(n16568), .X(n53703) );
  inv_x2_sg U76176 ( .A(n16954), .X(n53678) );
  inv_x2_sg U76177 ( .A(n17000), .X(n53696) );
  inv_x2_sg U76178 ( .A(n17267), .X(n53693) );
  inv_x2_sg U76179 ( .A(n17089), .X(n53694) );
  inv_x2_sg U76180 ( .A(n16953), .X(n53700) );
  inv_x2_sg U76181 ( .A(n16564), .X(n53670) );
  inv_x2_sg U76182 ( .A(n44142), .X(n53659) );
  inv_x2_sg U76183 ( .A(n17041), .X(n53589) );
  inv_x2_sg U76184 ( .A(n17042), .X(n53567) );
  inv_x2_sg U76185 ( .A(n27761), .X(n53662) );
  inv_x2_sg U76186 ( .A(n17078), .X(n53609) );
  inv_x2_sg U76187 ( .A(n17079), .X(n53620) );
  inv_x2_sg U76188 ( .A(n16996), .X(n53664) );
  inv_x2_sg U76189 ( .A(n45405), .X(n53665) );
  inv_x2_sg U76190 ( .A(n16921), .X(n53666) );
  inv_x2_sg U76191 ( .A(n16912), .X(n53667) );
  inv_x2_sg U76192 ( .A(n16560), .X(n53650) );
  inv_x2_sg U76193 ( .A(n16943), .X(n53594) );
  inv_x2_sg U76194 ( .A(n27767), .X(n53640) );
  inv_x2_sg U76195 ( .A(n16939), .X(n53645) );
  inv_x2_sg U76196 ( .A(n16979), .X(n53615) );
  inv_x2_sg U76197 ( .A(n16824), .X(n53608) );
  inv_x2_sg U76198 ( .A(n16875), .X(n53606) );
  inv_x2_sg U76199 ( .A(n16833), .X(n53588) );
  inv_x2_sg U76200 ( .A(n27773), .X(n53618) );
  inv_x2_sg U76201 ( .A(n16832), .X(n53626) );
  inv_x2_sg U76202 ( .A(n16607), .X(n53628) );
  inv_x2_sg U76203 ( .A(n16546), .X(n53584) );
  inv_x2_sg U76204 ( .A(n16837), .X(n53600) );
  inv_x2_sg U76205 ( .A(n16838), .X(n53593) );
  inv_x2_sg U76206 ( .A(n27779), .X(n53597) );
  inv_x2_sg U76207 ( .A(n16885), .X(n53558) );
  inv_x2_sg U76208 ( .A(n16886), .X(n53545) );
  inv_x2_sg U76209 ( .A(n16843), .X(n53599) );
  inv_x2_sg U76210 ( .A(n16789), .X(n53602) );
  inv_x2_sg U76211 ( .A(n16557), .X(n53603) );
  inv_x2_sg U76212 ( .A(n16558), .X(n53604) );
  inv_x2_sg U76213 ( .A(n16735), .X(n53582) );
  inv_x2_sg U76214 ( .A(n16799), .X(n53569) );
  inv_x2_sg U76215 ( .A(n27785), .X(n53578) );
  inv_x2_sg U76216 ( .A(n16543), .X(n53575) );
  inv_x2_sg U76217 ( .A(n16707), .X(n53555) );
  inv_x2_sg U76218 ( .A(n16734), .X(n53573) );
  inv_x2_sg U76219 ( .A(n27791), .X(n53564) );
  inv_x2_sg U76220 ( .A(n16741), .X(n53557) );
  inv_x2_sg U76221 ( .A(n16686), .X(n53552) );
  inv_x2_sg U76222 ( .A(n16709), .X(n53544) );
  inv_x2_sg U76223 ( .A(n16718), .X(n53550) );
  inv_x2_sg U76224 ( .A(n16680), .X(n53540) );
  inv_x2_sg U76225 ( .A(n43837), .X(n53516) );
  inv_x2_sg U76226 ( .A(n16667), .X(n53526) );
  inv_x2_sg U76227 ( .A(n16643), .X(n53501) );
  inv_x2_sg U76228 ( .A(n27817), .X(n53508) );
  inv_x2_sg U76229 ( .A(n16658), .X(n53511) );
  inv_x2_sg U76230 ( .A(n16617), .X(n53495) );
  inv_x2_sg U76231 ( .A(n27823), .X(n53489) );
  inv_x2_sg U76232 ( .A(n27829), .X(n53485) );
  inv_x2_sg U76233 ( .A(n44271), .X(n53486) );
  inv_x2_sg U76234 ( .A(n16514), .X(n53487) );
  inv_x2_sg U76235 ( .A(n46007), .X(n51120) );
  inv_x2_sg U76236 ( .A(n44841), .X(n53480) );
  inv_x2_sg U76237 ( .A(n15802), .X(n53462) );
  inv_x2_sg U76238 ( .A(n16345), .X(n53468) );
  inv_x2_sg U76239 ( .A(n16358), .X(n53466) );
  inv_x2_sg U76240 ( .A(n16372), .X(n53409) );
  inv_x2_sg U76241 ( .A(n16371), .X(n53431) );
  inv_x2_sg U76242 ( .A(n16390), .X(n53450) );
  inv_x2_sg U76243 ( .A(n16395), .X(n53426) );
  inv_x2_sg U76244 ( .A(n16397), .X(n53381) );
  inv_x2_sg U76245 ( .A(n16389), .X(n53433) );
  inv_x2_sg U76246 ( .A(n16222), .X(n53459) );
  inv_x2_sg U76247 ( .A(n16325), .X(n53380) );
  inv_x2_sg U76248 ( .A(n15806), .X(n53455) );
  inv_x2_sg U76249 ( .A(n15810), .X(n53456) );
  inv_x2_sg U76250 ( .A(n16338), .X(n53439) );
  inv_x2_sg U76251 ( .A(n16217), .X(n53443) );
  inv_x2_sg U76252 ( .A(n16315), .X(n53412) );
  inv_x2_sg U76253 ( .A(n16312), .X(n53393) );
  inv_x2_sg U76254 ( .A(n16461), .X(n53394) );
  inv_x2_sg U76255 ( .A(n16452), .X(n53285) );
  inv_x2_sg U76256 ( .A(n16275), .X(n53437) );
  inv_x2_sg U76257 ( .A(n16487), .X(n53423) );
  inv_x2_sg U76258 ( .A(n16493), .X(n53435) );
  inv_x2_sg U76259 ( .A(n27571), .X(n53429) );
  inv_x2_sg U76260 ( .A(n16477), .X(n53360) );
  inv_x2_sg U76261 ( .A(n16223), .X(n53442) );
  inv_x2_sg U76262 ( .A(n15786), .X(n53422) );
  inv_x2_sg U76263 ( .A(n16169), .X(n53399) );
  inv_x2_sg U76264 ( .A(n16215), .X(n53416) );
  inv_x2_sg U76265 ( .A(n27476), .X(n53407) );
  inv_x2_sg U76266 ( .A(n16486), .X(n53413) );
  inv_x2_sg U76267 ( .A(n16305), .X(n53414) );
  inv_x2_sg U76268 ( .A(n16168), .X(n53419) );
  inv_x2_sg U76269 ( .A(n16258), .X(n53379) );
  inv_x2_sg U76270 ( .A(n16270), .X(n53396) );
  inv_x2_sg U76271 ( .A(n15782), .X(n53391) );
  inv_x2_sg U76272 ( .A(n16256), .X(n53309) );
  inv_x2_sg U76273 ( .A(n16257), .X(n53284) );
  inv_x2_sg U76274 ( .A(n27482), .X(n53383) );
  inv_x2_sg U76275 ( .A(n16294), .X(n53330) );
  inv_x2_sg U76276 ( .A(n16295), .X(n53341) );
  inv_x2_sg U76277 ( .A(n16136), .X(n53387) );
  inv_x2_sg U76278 ( .A(n16127), .X(n53388) );
  inv_x2_sg U76279 ( .A(n16233), .X(n53354) );
  inv_x2_sg U76280 ( .A(n15778), .X(n53372) );
  inv_x2_sg U76281 ( .A(n16158), .X(n53314) );
  inv_x2_sg U76282 ( .A(n27488), .X(n53362) );
  inv_x2_sg U76283 ( .A(n16238), .X(n53364) );
  inv_x2_sg U76284 ( .A(n16194), .X(n53336) );
  inv_x2_sg U76285 ( .A(n16039), .X(n53329) );
  inv_x2_sg U76286 ( .A(n16090), .X(n53327) );
  inv_x2_sg U76287 ( .A(n16048), .X(n53308) );
  inv_x2_sg U76288 ( .A(n27494), .X(n53339) );
  inv_x2_sg U76289 ( .A(n16047), .X(n53347) );
  inv_x2_sg U76290 ( .A(n15825), .X(n53349) );
  inv_x2_sg U76291 ( .A(n15764), .X(n53304) );
  inv_x2_sg U76292 ( .A(n16052), .X(n53321) );
  inv_x2_sg U76293 ( .A(n16053), .X(n53313) );
  inv_x2_sg U76294 ( .A(n27500), .X(n53318) );
  inv_x2_sg U76295 ( .A(n16100), .X(n53276) );
  inv_x2_sg U76296 ( .A(n16101), .X(n53254) );
  inv_x2_sg U76297 ( .A(n16058), .X(n53320) );
  inv_x2_sg U76298 ( .A(n16004), .X(n53323) );
  inv_x2_sg U76299 ( .A(n15775), .X(n53324) );
  inv_x2_sg U76300 ( .A(n15776), .X(n53325) );
  inv_x2_sg U76301 ( .A(n15949), .X(n53302) );
  inv_x2_sg U76302 ( .A(n15941), .X(n53248) );
  inv_x2_sg U76303 ( .A(n16014), .X(n53293) );
  inv_x2_sg U76304 ( .A(n27506), .X(n53297) );
  inv_x2_sg U76305 ( .A(n15761), .X(n53291) );
  inv_x2_sg U76306 ( .A(n15918), .X(n53273) );
  inv_x2_sg U76307 ( .A(n15948), .X(n53289) );
  inv_x2_sg U76308 ( .A(n27512), .X(n53281) );
  inv_x2_sg U76309 ( .A(n15955), .X(n53275) );
  inv_x2_sg U76310 ( .A(n15898), .X(n53270) );
  inv_x2_sg U76311 ( .A(n15930), .X(n53268) );
  inv_x2_sg U76312 ( .A(n15903), .X(n53255) );
  inv_x2_sg U76313 ( .A(n27528), .X(n53251) );
  inv_x2_sg U76314 ( .A(n15911), .X(n53232) );
  inv_x2_sg U76315 ( .A(n15893), .X(n53257) );
  inv_x2_sg U76316 ( .A(n15862), .X(n53231) );
  inv_x2_sg U76317 ( .A(n15881), .X(n53241) );
  inv_x2_sg U76318 ( .A(n27530), .X(n53239) );
  inv_x2_sg U76319 ( .A(n15880), .X(n53235) );
  inv_x2_sg U76320 ( .A(n15851), .X(n53224) );
  inv_x2_sg U76321 ( .A(n15856), .X(n53221) );
  inv_x2_sg U76322 ( .A(n27538), .X(n53219) );
  inv_x2_sg U76323 ( .A(n15872), .X(n53228) );
  inv_x2_sg U76324 ( .A(n15844), .X(n53223) );
  inv_x2_sg U76325 ( .A(n27544), .X(n53211) );
  inv_x2_sg U76326 ( .A(n27550), .X(n53205) );
  inv_x2_sg U76327 ( .A(n44261), .X(n53206) );
  inv_x2_sg U76328 ( .A(n46013), .X(n51101) );
  inv_x2_sg U76329 ( .A(n44847), .X(n53200) );
  inv_x2_sg U76330 ( .A(n15017), .X(n53182) );
  inv_x2_sg U76331 ( .A(n15560), .X(n53189) );
  inv_x2_sg U76332 ( .A(n15569), .X(n53187) );
  inv_x2_sg U76333 ( .A(n15597), .X(n53128) );
  inv_x2_sg U76334 ( .A(n15604), .X(n53177) );
  inv_x2_sg U76335 ( .A(n15616), .X(n53097) );
  inv_x2_sg U76336 ( .A(n15641), .X(n53176) );
  inv_x2_sg U76337 ( .A(n15640), .X(n53162) );
  inv_x2_sg U76338 ( .A(n15494), .X(n53178) );
  inv_x2_sg U76339 ( .A(n15544), .X(n53102) );
  inv_x2_sg U76340 ( .A(n15613), .X(n53154) );
  inv_x2_sg U76341 ( .A(n15558), .X(n53160) );
  inv_x2_sg U76342 ( .A(n15032), .X(n53179) );
  inv_x2_sg U76343 ( .A(n15436), .X(n53164) );
  inv_x2_sg U76344 ( .A(n15526), .X(n53121) );
  inv_x2_sg U76345 ( .A(n15493), .X(n53157) );
  inv_x2_sg U76346 ( .A(n15702), .X(n53146) );
  inv_x2_sg U76347 ( .A(n15708), .X(n53155) );
  inv_x2_sg U76348 ( .A(n27292), .X(n53151) );
  inv_x2_sg U76349 ( .A(n15442), .X(n53163) );
  inv_x2_sg U76350 ( .A(n15002), .X(n53145) );
  inv_x2_sg U76351 ( .A(n15388), .X(n53120) );
  inv_x2_sg U76352 ( .A(n15434), .X(n53138) );
  inv_x2_sg U76353 ( .A(n15701), .X(n53135) );
  inv_x2_sg U76354 ( .A(n15523), .X(n53136) );
  inv_x2_sg U76355 ( .A(n15387), .X(n53142) );
  inv_x2_sg U76356 ( .A(n14998), .X(n53112) );
  inv_x2_sg U76357 ( .A(n44144), .X(n53101) );
  inv_x2_sg U76358 ( .A(n15475), .X(n53031) );
  inv_x2_sg U76359 ( .A(n15476), .X(n53009) );
  inv_x2_sg U76360 ( .A(n27203), .X(n53104) );
  inv_x2_sg U76361 ( .A(n15512), .X(n53051) );
  inv_x2_sg U76362 ( .A(n15513), .X(n53062) );
  inv_x2_sg U76363 ( .A(n15430), .X(n53106) );
  inv_x2_sg U76364 ( .A(n45407), .X(n53107) );
  inv_x2_sg U76365 ( .A(n15355), .X(n53108) );
  inv_x2_sg U76366 ( .A(n15346), .X(n53109) );
  inv_x2_sg U76367 ( .A(n14994), .X(n53092) );
  inv_x2_sg U76368 ( .A(n15377), .X(n53036) );
  inv_x2_sg U76369 ( .A(n27209), .X(n53082) );
  inv_x2_sg U76370 ( .A(n15373), .X(n53087) );
  inv_x2_sg U76371 ( .A(n15413), .X(n53057) );
  inv_x2_sg U76372 ( .A(n15258), .X(n53050) );
  inv_x2_sg U76373 ( .A(n15309), .X(n53048) );
  inv_x2_sg U76374 ( .A(n15267), .X(n53030) );
  inv_x2_sg U76375 ( .A(n27215), .X(n53060) );
  inv_x2_sg U76376 ( .A(n15266), .X(n53068) );
  inv_x2_sg U76377 ( .A(n15041), .X(n53070) );
  inv_x2_sg U76378 ( .A(n14980), .X(n53026) );
  inv_x2_sg U76379 ( .A(n15271), .X(n53042) );
  inv_x2_sg U76380 ( .A(n15272), .X(n53035) );
  inv_x2_sg U76381 ( .A(n27221), .X(n53039) );
  inv_x2_sg U76382 ( .A(n15319), .X(n53000) );
  inv_x2_sg U76383 ( .A(n15320), .X(n52987) );
  inv_x2_sg U76384 ( .A(n15277), .X(n53041) );
  inv_x2_sg U76385 ( .A(n15223), .X(n53044) );
  inv_x2_sg U76386 ( .A(n14991), .X(n53045) );
  inv_x2_sg U76387 ( .A(n14992), .X(n53046) );
  inv_x2_sg U76388 ( .A(n15169), .X(n53024) );
  inv_x2_sg U76389 ( .A(n15233), .X(n53011) );
  inv_x2_sg U76390 ( .A(n27227), .X(n53020) );
  inv_x2_sg U76391 ( .A(n14977), .X(n53017) );
  inv_x2_sg U76392 ( .A(n15141), .X(n52997) );
  inv_x2_sg U76393 ( .A(n15168), .X(n53015) );
  inv_x2_sg U76394 ( .A(n27233), .X(n53006) );
  inv_x2_sg U76395 ( .A(n15175), .X(n52999) );
  inv_x2_sg U76396 ( .A(n15120), .X(n52994) );
  inv_x2_sg U76397 ( .A(n15143), .X(n52986) );
  inv_x2_sg U76398 ( .A(n15152), .X(n52992) );
  inv_x2_sg U76399 ( .A(n15114), .X(n52982) );
  inv_x2_sg U76400 ( .A(n43839), .X(n52958) );
  inv_x2_sg U76401 ( .A(n15101), .X(n52968) );
  inv_x2_sg U76402 ( .A(n15077), .X(n52943) );
  inv_x2_sg U76403 ( .A(n27259), .X(n52950) );
  inv_x2_sg U76404 ( .A(n15092), .X(n52953) );
  inv_x2_sg U76405 ( .A(n15051), .X(n52937) );
  inv_x2_sg U76406 ( .A(n27265), .X(n52931) );
  inv_x2_sg U76407 ( .A(n27271), .X(n52927) );
  inv_x2_sg U76408 ( .A(n44273), .X(n52928) );
  inv_x2_sg U76409 ( .A(n14948), .X(n52929) );
  inv_x2_sg U76410 ( .A(n46009), .X(n51082) );
  inv_x2_sg U76411 ( .A(n44843), .X(n52922) );
  inv_x2_sg U76412 ( .A(n14247), .X(n52902) );
  inv_x2_sg U76413 ( .A(n14778), .X(n52911) );
  inv_x2_sg U76414 ( .A(n14787), .X(n52909) );
  inv_x2_sg U76415 ( .A(n14822), .X(n52904) );
  inv_x2_sg U76416 ( .A(n14832), .X(n52866) );
  inv_x2_sg U76417 ( .A(n14834), .X(n52808) );
  inv_x2_sg U76418 ( .A(n14859), .X(n52903) );
  inv_x2_sg U76419 ( .A(n14858), .X(n52880) );
  inv_x2_sg U76420 ( .A(n14712), .X(n52898) );
  inv_x2_sg U76421 ( .A(n14762), .X(n52821) );
  inv_x2_sg U76422 ( .A(n14770), .X(n52894) );
  inv_x2_sg U76423 ( .A(n14939), .X(n52893) );
  inv_x2_sg U76424 ( .A(n14251), .X(n52895) );
  inv_x2_sg U76425 ( .A(n14255), .X(n52896) );
  inv_x2_sg U76426 ( .A(n14880), .X(n52844) );
  inv_x2_sg U76427 ( .A(n14793), .X(n52864) );
  inv_x2_sg U76428 ( .A(n14775), .X(n52878) );
  inv_x2_sg U76429 ( .A(n14262), .X(n52899) );
  inv_x2_sg U76430 ( .A(n14652), .X(n52883) );
  inv_x2_sg U76431 ( .A(n14752), .X(n52852) );
  inv_x2_sg U76432 ( .A(n14890), .X(n52727) );
  inv_x2_sg U76433 ( .A(n14924), .X(n52863) );
  inv_x2_sg U76434 ( .A(n14930), .X(n52874) );
  inv_x2_sg U76435 ( .A(n27012), .X(n52869) );
  inv_x2_sg U76436 ( .A(n14883), .X(n52809) );
  inv_x2_sg U76437 ( .A(n14658), .X(n52882) );
  inv_x2_sg U76438 ( .A(n14232), .X(n52862) );
  inv_x2_sg U76439 ( .A(n14605), .X(n52842) );
  inv_x2_sg U76440 ( .A(n14650), .X(n52856) );
  inv_x2_sg U76441 ( .A(n14922), .X(n52853) );
  inv_x2_sg U76442 ( .A(n26917), .X(n52847) );
  inv_x2_sg U76443 ( .A(n14923), .X(n52713) );
  inv_x2_sg U76444 ( .A(n14741), .X(n52854) );
  inv_x2_sg U76445 ( .A(n14604), .X(n52859) );
  inv_x2_sg U76446 ( .A(n14706), .X(n52839) );
  inv_x2_sg U76447 ( .A(n14575), .X(n52827) );
  inv_x2_sg U76448 ( .A(n14691), .X(n52747) );
  inv_x2_sg U76449 ( .A(n14692), .X(n52726) );
  inv_x2_sg U76450 ( .A(n26923), .X(n52823) );
  inv_x2_sg U76451 ( .A(n14730), .X(n52767) );
  inv_x2_sg U76452 ( .A(n14731), .X(n52784) );
  inv_x2_sg U76453 ( .A(n14668), .X(n52796) );
  inv_x2_sg U76454 ( .A(n14568), .X(n52820) );
  inv_x2_sg U76455 ( .A(n14224), .X(n52819) );
  inv_x2_sg U76456 ( .A(n14594), .X(n52758) );
  inv_x2_sg U76457 ( .A(n26929), .X(n52805) );
  inv_x2_sg U76458 ( .A(n14673), .X(n52810) );
  inv_x2_sg U76459 ( .A(n14631), .X(n52779) );
  inv_x2_sg U76460 ( .A(n14479), .X(n52776) );
  inv_x2_sg U76461 ( .A(n14528), .X(n52765) );
  inv_x2_sg U76462 ( .A(n14508), .X(n52766) );
  inv_x2_sg U76463 ( .A(n14488), .X(n52746) );
  inv_x2_sg U76464 ( .A(n14539), .X(n52777) );
  inv_x2_sg U76465 ( .A(n26935), .X(n52782) );
  inv_x2_sg U76466 ( .A(n14487), .X(n52790) );
  inv_x2_sg U76467 ( .A(n14272), .X(n52792) );
  inv_x2_sg U76468 ( .A(n14210), .X(n52755) );
  inv_x2_sg U76469 ( .A(n14446), .X(n52774) );
  inv_x2_sg U76470 ( .A(n26941), .X(n52762) );
  inv_x2_sg U76471 ( .A(n14537), .X(n52709) );
  inv_x2_sg U76472 ( .A(n14538), .X(n52697) );
  inv_x2_sg U76473 ( .A(n14496), .X(n52710) );
  inv_x2_sg U76474 ( .A(n14491), .X(n52757) );
  inv_x2_sg U76475 ( .A(n14222), .X(n52775) );
  inv_x2_sg U76476 ( .A(n14392), .X(n52753) );
  inv_x2_sg U76477 ( .A(n14431), .X(n52730) );
  inv_x2_sg U76478 ( .A(n14414), .X(n52729) );
  inv_x2_sg U76479 ( .A(n26947), .X(n52741) );
  inv_x2_sg U76480 ( .A(n14443), .X(n52751) );
  inv_x2_sg U76481 ( .A(n14207), .X(n52735) );
  inv_x2_sg U76482 ( .A(n14363), .X(n52720) );
  inv_x2_sg U76483 ( .A(n14391), .X(n52733) );
  inv_x2_sg U76484 ( .A(n26953), .X(n52723) );
  inv_x2_sg U76485 ( .A(n14430), .X(n52677) );
  inv_x2_sg U76486 ( .A(n14429), .X(n52689) );
  inv_x2_sg U76487 ( .A(n14439), .X(n52696) );
  inv_x2_sg U76488 ( .A(n14343), .X(n52717) );
  inv_x2_sg U76489 ( .A(n14374), .X(n52715) );
  inv_x2_sg U76490 ( .A(n14347), .X(n52698) );
  inv_x2_sg U76491 ( .A(n26973), .X(n52668) );
  inv_x2_sg U76492 ( .A(n26969), .X(n52693) );
  inv_x2_sg U76493 ( .A(n14344), .X(n52688) );
  inv_x2_sg U76494 ( .A(n14301), .X(n52673) );
  inv_x2_sg U76495 ( .A(n14326), .X(n52684) );
  inv_x2_sg U76496 ( .A(n14325), .X(n52679) );
  inv_x2_sg U76497 ( .A(n26979), .X(n52660) );
  inv_x2_sg U76498 ( .A(n14313), .X(n52671) );
  inv_x2_sg U76499 ( .A(n14291), .X(n52663) );
  inv_x2_sg U76500 ( .A(n26985), .X(n52652) );
  inv_x2_sg U76501 ( .A(n26991), .X(n52646) );
  inv_x2_sg U76502 ( .A(n44265), .X(n52647) );
  inv_x2_sg U76503 ( .A(n46023), .X(n51063) );
  inv_x2_sg U76504 ( .A(n44867), .X(n52641) );
  inv_x2_sg U76505 ( .A(n13468), .X(n52623) );
  inv_x2_sg U76506 ( .A(n14007), .X(n52630) );
  inv_x2_sg U76507 ( .A(n14016), .X(n52628) );
  inv_x2_sg U76508 ( .A(n14044), .X(n52569) );
  inv_x2_sg U76509 ( .A(n14051), .X(n52618) );
  inv_x2_sg U76510 ( .A(n14063), .X(n52539) );
  inv_x2_sg U76511 ( .A(n14088), .X(n52617) );
  inv_x2_sg U76512 ( .A(n14087), .X(n52603) );
  inv_x2_sg U76513 ( .A(n13941), .X(n52619) );
  inv_x2_sg U76514 ( .A(n14060), .X(n52595) );
  inv_x2_sg U76515 ( .A(n14005), .X(n52601) );
  inv_x2_sg U76516 ( .A(n13483), .X(n52620) );
  inv_x2_sg U76517 ( .A(n13883), .X(n52605) );
  inv_x2_sg U76518 ( .A(n13973), .X(n52562) );
  inv_x2_sg U76519 ( .A(n13940), .X(n52598) );
  inv_x2_sg U76520 ( .A(n14149), .X(n52587) );
  inv_x2_sg U76521 ( .A(n14155), .X(n52596) );
  inv_x2_sg U76522 ( .A(n26733), .X(n52592) );
  inv_x2_sg U76523 ( .A(n13889), .X(n52604) );
  inv_x2_sg U76524 ( .A(n13453), .X(n52586) );
  inv_x2_sg U76525 ( .A(n13835), .X(n52561) );
  inv_x2_sg U76526 ( .A(n13881), .X(n52579) );
  inv_x2_sg U76527 ( .A(n14148), .X(n52576) );
  inv_x2_sg U76528 ( .A(n13970), .X(n52577) );
  inv_x2_sg U76529 ( .A(n13834), .X(n52583) );
  inv_x2_sg U76530 ( .A(n13449), .X(n52553) );
  inv_x2_sg U76531 ( .A(n44146), .X(n52543) );
  inv_x2_sg U76532 ( .A(n13922), .X(n52474) );
  inv_x2_sg U76533 ( .A(n13923), .X(n52450) );
  inv_x2_sg U76534 ( .A(n26644), .X(n52545) );
  inv_x2_sg U76535 ( .A(n13959), .X(n52494) );
  inv_x2_sg U76536 ( .A(n13960), .X(n52505) );
  inv_x2_sg U76537 ( .A(n13877), .X(n52547) );
  inv_x2_sg U76538 ( .A(n45409), .X(n52548) );
  inv_x2_sg U76539 ( .A(n13802), .X(n52549) );
  inv_x2_sg U76540 ( .A(n13793), .X(n52550) );
  inv_x2_sg U76541 ( .A(n13445), .X(n52534) );
  inv_x2_sg U76542 ( .A(n13824), .X(n52479) );
  inv_x2_sg U76543 ( .A(n26650), .X(n52524) );
  inv_x2_sg U76544 ( .A(n13820), .X(n52529) );
  inv_x2_sg U76545 ( .A(n13860), .X(n52500) );
  inv_x2_sg U76546 ( .A(n13705), .X(n52493) );
  inv_x2_sg U76547 ( .A(n13756), .X(n52491) );
  inv_x2_sg U76548 ( .A(n13714), .X(n52473) );
  inv_x2_sg U76549 ( .A(n26656), .X(n52503) );
  inv_x2_sg U76550 ( .A(n13713), .X(n52511) );
  inv_x2_sg U76551 ( .A(n13492), .X(n52513) );
  inv_x2_sg U76552 ( .A(n13431), .X(n52469) );
  inv_x2_sg U76553 ( .A(n13718), .X(n52485) );
  inv_x2_sg U76554 ( .A(n13719), .X(n52478) );
  inv_x2_sg U76555 ( .A(n26662), .X(n52482) );
  inv_x2_sg U76556 ( .A(n13766), .X(n52440) );
  inv_x2_sg U76557 ( .A(n13767), .X(n52419) );
  inv_x2_sg U76558 ( .A(n13724), .X(n52484) );
  inv_x2_sg U76559 ( .A(n13670), .X(n52487) );
  inv_x2_sg U76560 ( .A(n13442), .X(n52488) );
  inv_x2_sg U76561 ( .A(n13443), .X(n52489) );
  inv_x2_sg U76562 ( .A(n13615), .X(n52467) );
  inv_x2_sg U76563 ( .A(n13680), .X(n52452) );
  inv_x2_sg U76564 ( .A(n13624), .X(n52438) );
  inv_x2_sg U76565 ( .A(n26668), .X(n52462) );
  inv_x2_sg U76566 ( .A(n13428), .X(n52459) );
  inv_x2_sg U76567 ( .A(n13584), .X(n52437) );
  inv_x2_sg U76568 ( .A(n13614), .X(n52457) );
  inv_x2_sg U76569 ( .A(n26674), .X(n52446) );
  inv_x2_sg U76570 ( .A(n13626), .X(n52439) );
  inv_x2_sg U76571 ( .A(n13564), .X(n52434) );
  inv_x2_sg U76572 ( .A(n13589), .X(n52432) );
  inv_x2_sg U76573 ( .A(n13569), .X(n52420) );
  inv_x2_sg U76574 ( .A(n26690), .X(n52417) );
  inv_x2_sg U76575 ( .A(n13577), .X(n52398) );
  inv_x2_sg U76576 ( .A(n13559), .X(n52422) );
  inv_x2_sg U76577 ( .A(n43936), .X(n52397) );
  inv_x2_sg U76578 ( .A(n13547), .X(n52407) );
  inv_x2_sg U76579 ( .A(n13546), .X(n52401) );
  inv_x2_sg U76580 ( .A(n13517), .X(n52388) );
  inv_x2_sg U76581 ( .A(n13522), .X(n52385) );
  inv_x2_sg U76582 ( .A(n26700), .X(n52383) );
  inv_x2_sg U76583 ( .A(n13538), .X(n52392) );
  inv_x2_sg U76584 ( .A(n44325), .X(n52394) );
  inv_x2_sg U76585 ( .A(n13511), .X(n52387) );
  inv_x2_sg U76586 ( .A(n26706), .X(n52375) );
  inv_x2_sg U76587 ( .A(n26712), .X(n52370) );
  inv_x2_sg U76588 ( .A(n44269), .X(n52371) );
  inv_x2_sg U76589 ( .A(n46015), .X(n51044) );
  inv_x2_sg U76590 ( .A(n44855), .X(n52365) );
  inv_x2_sg U76591 ( .A(n12684), .X(n52348) );
  inv_x2_sg U76592 ( .A(n13227), .X(n52355) );
  inv_x2_sg U76593 ( .A(n13236), .X(n52353) );
  inv_x2_sg U76594 ( .A(n13264), .X(n52294) );
  inv_x2_sg U76595 ( .A(n13271), .X(n52343) );
  inv_x2_sg U76596 ( .A(n13283), .X(n52263) );
  inv_x2_sg U76597 ( .A(n13308), .X(n52342) );
  inv_x2_sg U76598 ( .A(n13307), .X(n52328) );
  inv_x2_sg U76599 ( .A(n13161), .X(n52344) );
  inv_x2_sg U76600 ( .A(n13211), .X(n52268) );
  inv_x2_sg U76601 ( .A(n13280), .X(n52320) );
  inv_x2_sg U76602 ( .A(n13225), .X(n52326) );
  inv_x2_sg U76603 ( .A(n12699), .X(n52345) );
  inv_x2_sg U76604 ( .A(n13103), .X(n52330) );
  inv_x2_sg U76605 ( .A(n13193), .X(n52287) );
  inv_x2_sg U76606 ( .A(n13160), .X(n52323) );
  inv_x2_sg U76607 ( .A(n13369), .X(n52312) );
  inv_x2_sg U76608 ( .A(n13375), .X(n52321) );
  inv_x2_sg U76609 ( .A(n26455), .X(n52317) );
  inv_x2_sg U76610 ( .A(n13109), .X(n52329) );
  inv_x2_sg U76611 ( .A(n12669), .X(n52311) );
  inv_x2_sg U76612 ( .A(n13055), .X(n52286) );
  inv_x2_sg U76613 ( .A(n13101), .X(n52304) );
  inv_x2_sg U76614 ( .A(n13368), .X(n52301) );
  inv_x2_sg U76615 ( .A(n13190), .X(n52302) );
  inv_x2_sg U76616 ( .A(n13054), .X(n52308) );
  inv_x2_sg U76617 ( .A(n12665), .X(n52278) );
  inv_x2_sg U76618 ( .A(n44148), .X(n52267) );
  inv_x2_sg U76619 ( .A(n13142), .X(n52197) );
  inv_x2_sg U76620 ( .A(n13143), .X(n52175) );
  inv_x2_sg U76621 ( .A(n26366), .X(n52270) );
  inv_x2_sg U76622 ( .A(n13179), .X(n52217) );
  inv_x2_sg U76623 ( .A(n13180), .X(n52228) );
  inv_x2_sg U76624 ( .A(n13097), .X(n52272) );
  inv_x2_sg U76625 ( .A(n45411), .X(n52273) );
  inv_x2_sg U76626 ( .A(n13022), .X(n52274) );
  inv_x2_sg U76627 ( .A(n13013), .X(n52275) );
  inv_x2_sg U76628 ( .A(n12661), .X(n52258) );
  inv_x2_sg U76629 ( .A(n13044), .X(n52202) );
  inv_x2_sg U76630 ( .A(n26372), .X(n52248) );
  inv_x2_sg U76631 ( .A(n13040), .X(n52253) );
  inv_x2_sg U76632 ( .A(n13080), .X(n52223) );
  inv_x2_sg U76633 ( .A(n12925), .X(n52216) );
  inv_x2_sg U76634 ( .A(n12976), .X(n52214) );
  inv_x2_sg U76635 ( .A(n12934), .X(n52196) );
  inv_x2_sg U76636 ( .A(n26378), .X(n52226) );
  inv_x2_sg U76637 ( .A(n12933), .X(n52234) );
  inv_x2_sg U76638 ( .A(n12708), .X(n52236) );
  inv_x2_sg U76639 ( .A(n12647), .X(n52192) );
  inv_x2_sg U76640 ( .A(n12938), .X(n52208) );
  inv_x2_sg U76641 ( .A(n12939), .X(n52201) );
  inv_x2_sg U76642 ( .A(n26384), .X(n52205) );
  inv_x2_sg U76643 ( .A(n12986), .X(n52166) );
  inv_x2_sg U76644 ( .A(n12987), .X(n52153) );
  inv_x2_sg U76645 ( .A(n12944), .X(n52207) );
  inv_x2_sg U76646 ( .A(n12890), .X(n52210) );
  inv_x2_sg U76647 ( .A(n12658), .X(n52211) );
  inv_x2_sg U76648 ( .A(n12659), .X(n52212) );
  inv_x2_sg U76649 ( .A(n12836), .X(n52190) );
  inv_x2_sg U76650 ( .A(n12900), .X(n52177) );
  inv_x2_sg U76651 ( .A(n26390), .X(n52186) );
  inv_x2_sg U76652 ( .A(n12644), .X(n52183) );
  inv_x2_sg U76653 ( .A(n12808), .X(n52163) );
  inv_x2_sg U76654 ( .A(n12835), .X(n52181) );
  inv_x2_sg U76655 ( .A(n26396), .X(n52172) );
  inv_x2_sg U76656 ( .A(n12842), .X(n52165) );
  inv_x2_sg U76657 ( .A(n12787), .X(n52160) );
  inv_x2_sg U76658 ( .A(n12810), .X(n52152) );
  inv_x2_sg U76659 ( .A(n12819), .X(n52158) );
  inv_x2_sg U76660 ( .A(n12781), .X(n52148) );
  inv_x2_sg U76661 ( .A(n43841), .X(n52124) );
  inv_x2_sg U76662 ( .A(n12768), .X(n52134) );
  inv_x2_sg U76663 ( .A(n12744), .X(n52109) );
  inv_x2_sg U76664 ( .A(n26422), .X(n52116) );
  inv_x2_sg U76665 ( .A(n12759), .X(n52119) );
  inv_x2_sg U76666 ( .A(n12718), .X(n52103) );
  inv_x2_sg U76667 ( .A(n26428), .X(n52097) );
  inv_x2_sg U76668 ( .A(n26434), .X(n52093) );
  inv_x2_sg U76669 ( .A(n44275), .X(n52094) );
  inv_x2_sg U76670 ( .A(n12615), .X(n52095) );
  inv_x2_sg U76671 ( .A(n46011), .X(n51024) );
  inv_x2_sg U76672 ( .A(n44845), .X(n52088) );
  inv_x2_sg U76673 ( .A(n11906), .X(n52070) );
  inv_x2_sg U76674 ( .A(n12446), .X(n52077) );
  inv_x2_sg U76675 ( .A(n12455), .X(n52075) );
  inv_x2_sg U76676 ( .A(n12483), .X(n52018) );
  inv_x2_sg U76677 ( .A(n12490), .X(n52066) );
  inv_x2_sg U76678 ( .A(n12502), .X(n51992) );
  inv_x2_sg U76679 ( .A(n12527), .X(n52065) );
  inv_x2_sg U76680 ( .A(n12526), .X(n52051) );
  inv_x2_sg U76681 ( .A(n12381), .X(n52067) );
  inv_x2_sg U76682 ( .A(n12430), .X(n51991) );
  inv_x2_sg U76683 ( .A(n12499), .X(n52044) );
  inv_x2_sg U76684 ( .A(n12444), .X(n52049) );
  inv_x2_sg U76685 ( .A(n11921), .X(n52068) );
  inv_x2_sg U76686 ( .A(n12322), .X(n52053) );
  inv_x2_sg U76687 ( .A(n12386), .X(n52024) );
  inv_x2_sg U76688 ( .A(n12380), .X(n52047) );
  inv_x2_sg U76689 ( .A(n12593), .X(n52045) );
  inv_x2_sg U76690 ( .A(n26176), .X(n52041) );
  inv_x2_sg U76691 ( .A(n12328), .X(n52052) );
  inv_x2_sg U76692 ( .A(n11891), .X(n52036) );
  inv_x2_sg U76693 ( .A(n12274), .X(n52008) );
  inv_x2_sg U76694 ( .A(n12320), .X(n52029) );
  inv_x2_sg U76695 ( .A(n12410), .X(n51901) );
  inv_x2_sg U76696 ( .A(n12586), .X(n52025) );
  inv_x2_sg U76697 ( .A(n12273), .X(n52033) );
  inv_x2_sg U76698 ( .A(n12363), .X(n51988) );
  inv_x2_sg U76699 ( .A(n11887), .X(n52002) );
  inv_x2_sg U76700 ( .A(n12361), .X(n51922) );
  inv_x2_sg U76701 ( .A(n12362), .X(n51898) );
  inv_x2_sg U76702 ( .A(n26087), .X(n51994) );
  inv_x2_sg U76703 ( .A(n12399), .X(n51942) );
  inv_x2_sg U76704 ( .A(n12400), .X(n51953) );
  inv_x2_sg U76705 ( .A(n12241), .X(n51998) );
  inv_x2_sg U76706 ( .A(n12232), .X(n51999) );
  inv_x2_sg U76707 ( .A(n12338), .X(n51965) );
  inv_x2_sg U76708 ( .A(n11883), .X(n51983) );
  inv_x2_sg U76709 ( .A(n12263), .X(n51926) );
  inv_x2_sg U76710 ( .A(n26093), .X(n51973) );
  inv_x2_sg U76711 ( .A(n12343), .X(n51975) );
  inv_x2_sg U76712 ( .A(n12299), .X(n51948) );
  inv_x2_sg U76713 ( .A(n12144), .X(n51941) );
  inv_x2_sg U76714 ( .A(n12195), .X(n51939) );
  inv_x2_sg U76715 ( .A(n12153), .X(n51921) );
  inv_x2_sg U76716 ( .A(n26099), .X(n51951) );
  inv_x2_sg U76717 ( .A(n12152), .X(n51959) );
  inv_x2_sg U76718 ( .A(n11930), .X(n51961) );
  inv_x2_sg U76719 ( .A(n11869), .X(n51917) );
  inv_x2_sg U76720 ( .A(n12157), .X(n51933) );
  inv_x2_sg U76721 ( .A(n12158), .X(n51925) );
  inv_x2_sg U76722 ( .A(n26105), .X(n51930) );
  inv_x2_sg U76723 ( .A(n12205), .X(n51889) );
  inv_x2_sg U76724 ( .A(n12206), .X(n51867) );
  inv_x2_sg U76725 ( .A(n12163), .X(n51932) );
  inv_x2_sg U76726 ( .A(n12109), .X(n51935) );
  inv_x2_sg U76727 ( .A(n11880), .X(n51936) );
  inv_x2_sg U76728 ( .A(n11881), .X(n51937) );
  inv_x2_sg U76729 ( .A(n12054), .X(n51915) );
  inv_x2_sg U76730 ( .A(n12119), .X(n51900) );
  inv_x2_sg U76731 ( .A(n26111), .X(n51910) );
  inv_x2_sg U76732 ( .A(n11866), .X(n51906) );
  inv_x2_sg U76733 ( .A(n12023), .X(n51886) );
  inv_x2_sg U76734 ( .A(n12053), .X(n51904) );
  inv_x2_sg U76735 ( .A(n26117), .X(n51895) );
  inv_x2_sg U76736 ( .A(n12060), .X(n51888) );
  inv_x2_sg U76737 ( .A(n12003), .X(n51883) );
  inv_x2_sg U76738 ( .A(n12035), .X(n51881) );
  inv_x2_sg U76739 ( .A(n12008), .X(n51868) );
  inv_x2_sg U76740 ( .A(n26133), .X(n51865) );
  inv_x2_sg U76741 ( .A(n12016), .X(n51846) );
  inv_x2_sg U76742 ( .A(n11998), .X(n51870) );
  inv_x2_sg U76743 ( .A(n43938), .X(n51845) );
  inv_x2_sg U76744 ( .A(n11986), .X(n51855) );
  inv_x2_sg U76745 ( .A(n26135), .X(n51853) );
  inv_x2_sg U76746 ( .A(n11985), .X(n51849) );
  inv_x2_sg U76747 ( .A(n11956), .X(n51836) );
  inv_x2_sg U76748 ( .A(n11961), .X(n51833) );
  inv_x2_sg U76749 ( .A(n26143), .X(n51831) );
  inv_x2_sg U76750 ( .A(n11977), .X(n51840) );
  inv_x2_sg U76751 ( .A(n44327), .X(n51842) );
  inv_x2_sg U76752 ( .A(n11949), .X(n51835) );
  inv_x2_sg U76753 ( .A(n26149), .X(n51823) );
  inv_x2_sg U76754 ( .A(n26155), .X(n51817) );
  inv_x2_sg U76755 ( .A(n44277), .X(n51818) );
  inv_x2_sg U76756 ( .A(n46017), .X(n51005) );
  inv_x2_sg U76757 ( .A(n44857), .X(n51812) );
  inv_x2_sg U76758 ( .A(n11123), .X(n51792) );
  inv_x2_sg U76759 ( .A(n11666), .X(n51801) );
  inv_x2_sg U76760 ( .A(n11675), .X(n51799) );
  inv_x2_sg U76761 ( .A(n11710), .X(n51794) );
  inv_x2_sg U76762 ( .A(n11720), .X(n51757) );
  inv_x2_sg U76763 ( .A(n11722), .X(n51707) );
  inv_x2_sg U76764 ( .A(n11747), .X(n51793) );
  inv_x2_sg U76765 ( .A(n11746), .X(n51771) );
  inv_x2_sg U76766 ( .A(n11600), .X(n51788) );
  inv_x2_sg U76767 ( .A(n11650), .X(n51712) );
  inv_x2_sg U76768 ( .A(n11827), .X(n51783) );
  inv_x2_sg U76769 ( .A(n11660), .X(n51784) );
  inv_x2_sg U76770 ( .A(n11127), .X(n51785) );
  inv_x2_sg U76771 ( .A(n11131), .X(n51786) );
  inv_x2_sg U76772 ( .A(n11681), .X(n51755) );
  inv_x2_sg U76773 ( .A(n11787), .X(n51741) );
  inv_x2_sg U76774 ( .A(n11663), .X(n51769) );
  inv_x2_sg U76775 ( .A(n11138), .X(n51789) );
  inv_x2_sg U76776 ( .A(n11542), .X(n51773) );
  inv_x2_sg U76777 ( .A(n11640), .X(n51743) );
  inv_x2_sg U76778 ( .A(n11795), .X(n51742) );
  inv_x2_sg U76779 ( .A(n11599), .X(n51767) );
  inv_x2_sg U76780 ( .A(n11812), .X(n51754) );
  inv_x2_sg U76781 ( .A(n11818), .X(n51765) );
  inv_x2_sg U76782 ( .A(n25896), .X(n51760) );
  inv_x2_sg U76783 ( .A(n11805), .X(n51731) );
  inv_x2_sg U76784 ( .A(n11548), .X(n51772) );
  inv_x2_sg U76785 ( .A(n11108), .X(n51753) );
  inv_x2_sg U76786 ( .A(n11494), .X(n51730) );
  inv_x2_sg U76787 ( .A(n11540), .X(n51747) );
  inv_x2_sg U76788 ( .A(n25801), .X(n51737) );
  inv_x2_sg U76789 ( .A(n11811), .X(n51744) );
  inv_x2_sg U76790 ( .A(n11629), .X(n51745) );
  inv_x2_sg U76791 ( .A(n11493), .X(n51750) );
  inv_x2_sg U76792 ( .A(n11104), .X(n51724) );
  inv_x2_sg U76793 ( .A(n44150), .X(n51711) );
  inv_x2_sg U76794 ( .A(n11581), .X(n51641) );
  inv_x2_sg U76795 ( .A(n11582), .X(n51617) );
  inv_x2_sg U76796 ( .A(n25807), .X(n51716) );
  inv_x2_sg U76797 ( .A(n11618), .X(n51661) );
  inv_x2_sg U76798 ( .A(n11619), .X(n51672) );
  inv_x2_sg U76799 ( .A(n11536), .X(n51718) );
  inv_x2_sg U76800 ( .A(n45413), .X(n51719) );
  inv_x2_sg U76801 ( .A(n11461), .X(n51720) );
  inv_x2_sg U76802 ( .A(n11452), .X(n51721) );
  inv_x2_sg U76803 ( .A(n11100), .X(n51702) );
  inv_x2_sg U76804 ( .A(n11483), .X(n51646) );
  inv_x2_sg U76805 ( .A(n25813), .X(n51692) );
  inv_x2_sg U76806 ( .A(n11479), .X(n51697) );
  inv_x2_sg U76807 ( .A(n11519), .X(n51667) );
  inv_x2_sg U76808 ( .A(n11364), .X(n51660) );
  inv_x2_sg U76809 ( .A(n11415), .X(n51658) );
  inv_x2_sg U76810 ( .A(n11373), .X(n51640) );
  inv_x2_sg U76811 ( .A(n25819), .X(n51670) );
  inv_x2_sg U76812 ( .A(n11372), .X(n51678) );
  inv_x2_sg U76813 ( .A(n11147), .X(n51680) );
  inv_x2_sg U76814 ( .A(n11086), .X(n51636) );
  inv_x2_sg U76815 ( .A(n11377), .X(n51652) );
  inv_x2_sg U76816 ( .A(n11378), .X(n51645) );
  inv_x2_sg U76817 ( .A(n25825), .X(n51649) );
  inv_x2_sg U76818 ( .A(n11425), .X(n51608) );
  inv_x2_sg U76819 ( .A(n11426), .X(n51595) );
  inv_x2_sg U76820 ( .A(n11383), .X(n51651) );
  inv_x2_sg U76821 ( .A(n11329), .X(n51654) );
  inv_x2_sg U76822 ( .A(n11097), .X(n51655) );
  inv_x2_sg U76823 ( .A(n11098), .X(n51656) );
  inv_x2_sg U76824 ( .A(n11275), .X(n51634) );
  inv_x2_sg U76825 ( .A(n11267), .X(n51581) );
  inv_x2_sg U76826 ( .A(n11339), .X(n51626) );
  inv_x2_sg U76827 ( .A(n25831), .X(n51629) );
  inv_x2_sg U76828 ( .A(n11083), .X(n51624) );
  inv_x2_sg U76829 ( .A(n11247), .X(n51605) );
  inv_x2_sg U76830 ( .A(n11274), .X(n51622) );
  inv_x2_sg U76831 ( .A(n25837), .X(n51614) );
  inv_x2_sg U76832 ( .A(n11281), .X(n51607) );
  inv_x2_sg U76833 ( .A(n11226), .X(n51602) );
  inv_x2_sg U76834 ( .A(n11249), .X(n51594) );
  inv_x2_sg U76835 ( .A(n11258), .X(n51600) );
  inv_x2_sg U76836 ( .A(n11220), .X(n51590) );
  inv_x2_sg U76837 ( .A(n43843), .X(n51567) );
  inv_x2_sg U76838 ( .A(n11207), .X(n51576) );
  inv_x2_sg U76839 ( .A(n11183), .X(n51552) );
  inv_x2_sg U76840 ( .A(n25863), .X(n51559) );
  inv_x2_sg U76841 ( .A(n11198), .X(n51562) );
  inv_x2_sg U76842 ( .A(n11157), .X(n51546) );
  inv_x2_sg U76843 ( .A(n25869), .X(n51540) );
  inv_x2_sg U76844 ( .A(n25875), .X(n51535) );
  inv_x2_sg U76845 ( .A(n44259), .X(n51536) );
  inv_x2_sg U76846 ( .A(n11054), .X(n51538) );
  inv_x2_sg U76847 ( .A(n46019), .X(n50986) );
  inv_x2_sg U76848 ( .A(n44835), .X(n51530) );
  inv_x2_sg U76849 ( .A(n10356), .X(n51512) );
  inv_x2_sg U76850 ( .A(n10890), .X(n51519) );
  inv_x2_sg U76851 ( .A(n44249), .X(n51516) );
  inv_x2_sg U76852 ( .A(n10903), .X(n51517) );
  inv_x2_sg U76853 ( .A(n10913), .X(n51475) );
  inv_x2_sg U76854 ( .A(n10912), .X(n51482) );
  inv_x2_sg U76855 ( .A(n10932), .X(n51502) );
  inv_x2_sg U76856 ( .A(n10937), .X(n51477) );
  inv_x2_sg U76857 ( .A(n10939), .X(n51432) );
  inv_x2_sg U76858 ( .A(n10931), .X(n51484) );
  inv_x2_sg U76859 ( .A(n10765), .X(n51509) );
  inv_x2_sg U76860 ( .A(n10870), .X(n51431) );
  inv_x2_sg U76861 ( .A(n11043), .X(n51503) );
  inv_x2_sg U76862 ( .A(n10880), .X(n51504) );
  inv_x2_sg U76863 ( .A(n10360), .X(n51505) );
  inv_x2_sg U76864 ( .A(n10364), .X(n51506) );
  inv_x2_sg U76865 ( .A(n10883), .X(n51490) );
  inv_x2_sg U76866 ( .A(n10860), .X(n51462) );
  inv_x2_sg U76867 ( .A(n10994), .X(n51459) );
  inv_x2_sg U76868 ( .A(n11011), .X(n51461) );
  inv_x2_sg U76869 ( .A(n10819), .X(n51488) );
  inv_x2_sg U76870 ( .A(n25615), .X(n51480) );
  inv_x2_sg U76871 ( .A(n10766), .X(n51493) );
  inv_x2_sg U76872 ( .A(n10340), .X(n51473) );
  inv_x2_sg U76873 ( .A(n10713), .X(n51451) );
  inv_x2_sg U76874 ( .A(n10758), .X(n51467) );
  inv_x2_sg U76875 ( .A(n10849), .X(n51338) );
  inv_x2_sg U76876 ( .A(n11027), .X(n51463) );
  inv_x2_sg U76877 ( .A(n25522), .X(n51457) );
  inv_x2_sg U76878 ( .A(n11028), .X(n51323) );
  inv_x2_sg U76879 ( .A(n10712), .X(n51470) );
  inv_x2_sg U76880 ( .A(n10683), .X(n51438) );
  inv_x2_sg U76881 ( .A(n10799), .X(n51336) );
  inv_x2_sg U76882 ( .A(n25528), .X(n51434) );
  inv_x2_sg U76883 ( .A(n10838), .X(n51381) );
  inv_x2_sg U76884 ( .A(n10676), .X(n51430) );
  inv_x2_sg U76885 ( .A(n10332), .X(n51429) );
  inv_x2_sg U76886 ( .A(n10702), .X(n51370) );
  inv_x2_sg U76887 ( .A(n25534), .X(n51417) );
  inv_x2_sg U76888 ( .A(n10781), .X(n51420) );
  inv_x2_sg U76889 ( .A(n10739), .X(n51390) );
  inv_x2_sg U76890 ( .A(n10587), .X(n51388) );
  inv_x2_sg U76891 ( .A(n10636), .X(n51379) );
  inv_x2_sg U76892 ( .A(n10616), .X(n51380) );
  inv_x2_sg U76893 ( .A(n10596), .X(n51369) );
  inv_x2_sg U76894 ( .A(n44082), .X(n51389) );
  inv_x2_sg U76895 ( .A(n10662), .X(n51399) );
  inv_x2_sg U76896 ( .A(n10595), .X(n51401) );
  inv_x2_sg U76897 ( .A(n10380), .X(n51403) );
  inv_x2_sg U76898 ( .A(n10318), .X(n51365) );
  inv_x2_sg U76899 ( .A(n10554), .X(n51387) );
  inv_x2_sg U76900 ( .A(n25546), .X(n51376) );
  inv_x2_sg U76901 ( .A(n10645), .X(n51319) );
  inv_x2_sg U76902 ( .A(n10646), .X(n51308) );
  inv_x2_sg U76903 ( .A(n10604), .X(n51320) );
  inv_x2_sg U76904 ( .A(n10599), .X(n51360) );
  inv_x2_sg U76905 ( .A(n10501), .X(n51363) );
  inv_x2_sg U76906 ( .A(n10538), .X(n51340) );
  inv_x2_sg U76907 ( .A(n10522), .X(n51339) );
  inv_x2_sg U76908 ( .A(n10550), .X(n51361) );
  inv_x2_sg U76909 ( .A(n10315), .X(n51345) );
  inv_x2_sg U76910 ( .A(n10471), .X(n51330) );
  inv_x2_sg U76911 ( .A(n10500), .X(n51343) );
  inv_x2_sg U76912 ( .A(n25556), .X(n51333) );
  inv_x2_sg U76913 ( .A(n10493), .X(n51287) );
  inv_x2_sg U76914 ( .A(n10537), .X(n51299) );
  inv_x2_sg U76915 ( .A(n10451), .X(n51327) );
  inv_x2_sg U76916 ( .A(n10482), .X(n51325) );
  inv_x2_sg U76917 ( .A(n10458), .X(n51309) );
  inv_x2_sg U76918 ( .A(n25572), .X(n51304) );
  inv_x2_sg U76919 ( .A(n10452), .X(n51298) );
  inv_x2_sg U76920 ( .A(n10409), .X(n51283) );
  inv_x2_sg U76921 ( .A(n10434), .X(n51294) );
  inv_x2_sg U76922 ( .A(n25574), .X(n51292) );
  inv_x2_sg U76923 ( .A(n10433), .X(n51289) );
  inv_x2_sg U76924 ( .A(n10425), .X(n51269) );
  inv_x2_sg U76925 ( .A(n25582), .X(n51271) );
  inv_x2_sg U76926 ( .A(n10421), .X(n51281) );
  inv_x2_sg U76927 ( .A(n10399), .X(n51274) );
  inv_x2_sg U76928 ( .A(n25588), .X(n51264) );
  inv_x2_sg U76929 ( .A(n25594), .X(n51259) );
  inv_x2_sg U76930 ( .A(n44257), .X(n51260) );
  inv_x2_sg U76931 ( .A(n46027), .X(n50967) );
  inv_x2_sg U76932 ( .A(n44865), .X(n51254) );
  inv_x2_sg U76933 ( .A(n10230), .X(n50125) );
  inv_x2_sg U76934 ( .A(n44070), .X(n50158) );
  inv_x2_sg U76935 ( .A(n22066), .X(n50157) );
  inv_x2_sg U76936 ( .A(n44577), .X(n50201) );
  inv_x2_sg U76937 ( .A(n22073), .X(n50200) );
  inv_x2_sg U76938 ( .A(n44579), .X(n50245) );
  inv_x2_sg U76939 ( .A(n22080), .X(n50244) );
  inv_x2_sg U76940 ( .A(n44581), .X(n50291) );
  inv_x2_sg U76941 ( .A(n22087), .X(n50290) );
  inv_x2_sg U76942 ( .A(n44585), .X(n50337) );
  inv_x2_sg U76943 ( .A(n22094), .X(n50336) );
  inv_x2_sg U76944 ( .A(n44587), .X(n50384) );
  inv_x2_sg U76945 ( .A(n22101), .X(n50383) );
  inv_x2_sg U76946 ( .A(n44591), .X(n50431) );
  inv_x2_sg U76947 ( .A(n22108), .X(n50430) );
  inv_x2_sg U76948 ( .A(n44595), .X(n50477) );
  inv_x2_sg U76949 ( .A(n22115), .X(n50476) );
  inv_x2_sg U76950 ( .A(n44599), .X(n50524) );
  inv_x2_sg U76951 ( .A(n22122), .X(n50523) );
  inv_x2_sg U76952 ( .A(n44603), .X(n50571) );
  inv_x2_sg U76953 ( .A(n22129), .X(n50570) );
  inv_x2_sg U76954 ( .A(n44607), .X(n50620) );
  inv_x2_sg U76955 ( .A(n22136), .X(n50619) );
  inv_x2_sg U76956 ( .A(n44609), .X(n50667) );
  inv_x2_sg U76957 ( .A(n22143), .X(n50666) );
  inv_x2_sg U76958 ( .A(n44613), .X(n50715) );
  inv_x2_sg U76959 ( .A(n22150), .X(n50714) );
  inv_x2_sg U76960 ( .A(n44617), .X(n50762) );
  inv_x2_sg U76961 ( .A(n22157), .X(n50761) );
  inv_x2_sg U76962 ( .A(n44619), .X(n50810) );
  inv_x2_sg U76963 ( .A(n22164), .X(n50809) );
  inv_x2_sg U76964 ( .A(n44655), .X(n50854) );
  inv_x2_sg U76965 ( .A(n22171), .X(n50853) );
  inv_x2_sg U76966 ( .A(n44653), .X(n50904) );
  inv_x2_sg U76967 ( .A(n22183), .X(n50906) );
  inv_x2_sg U76968 ( .A(n22192), .X(n50903) );
  inv_x2_sg U76969 ( .A(n22343), .X(n50897) );
  inv_x2_sg U76970 ( .A(n22349), .X(n50858) );
  inv_x2_sg U76971 ( .A(n22412), .X(n50160) );
  inv_x2_sg U76972 ( .A(n22418), .X(n50205) );
  inv_x2_sg U76973 ( .A(n22424), .X(n50249) );
  inv_x2_sg U76974 ( .A(n22430), .X(n50295) );
  inv_x2_sg U76975 ( .A(n22436), .X(n50341) );
  inv_x2_sg U76976 ( .A(n22442), .X(n50388) );
  inv_x2_sg U76977 ( .A(n22448), .X(n50435) );
  inv_x2_sg U76978 ( .A(n22454), .X(n50481) );
  inv_x2_sg U76979 ( .A(n22460), .X(n50528) );
  inv_x2_sg U76980 ( .A(n22466), .X(n50575) );
  inv_x2_sg U76981 ( .A(n22472), .X(n50624) );
  inv_x2_sg U76982 ( .A(n22478), .X(n50671) );
  inv_x2_sg U76983 ( .A(n22484), .X(n50719) );
  inv_x2_sg U76984 ( .A(n22490), .X(n50766) );
  inv_x2_sg U76985 ( .A(n22496), .X(n50814) );
  inv_x2_sg U76986 ( .A(n22571), .X(n50923) );
  inv_x2_sg U76987 ( .A(n22578), .X(n50951) );
  inv_x2_sg U76988 ( .A(n22586), .X(n50928) );
  inv_x2_sg U76989 ( .A(n22614), .X(n50950) );
  inv_x2_sg U76990 ( .A(n10213), .X(n50151) );
  inv_x2_sg U76991 ( .A(n22679), .X(n50192) );
  inv_x2_sg U76992 ( .A(n22685), .X(n50236) );
  inv_x2_sg U76993 ( .A(n22691), .X(n50282) );
  inv_x2_sg U76994 ( .A(n22697), .X(n50328) );
  inv_x2_sg U76995 ( .A(n22703), .X(n50375) );
  inv_x2_sg U76996 ( .A(n22709), .X(n50422) );
  inv_x2_sg U76997 ( .A(n22715), .X(n50468) );
  inv_x2_sg U76998 ( .A(n22721), .X(n50515) );
  inv_x2_sg U76999 ( .A(n22727), .X(n50562) );
  inv_x2_sg U77000 ( .A(n22733), .X(n50611) );
  inv_x2_sg U77001 ( .A(n22739), .X(n50659) );
  inv_x2_sg U77002 ( .A(n22745), .X(n50706) );
  inv_x2_sg U77003 ( .A(n22751), .X(n50753) );
  inv_x2_sg U77004 ( .A(n22757), .X(n50801) );
  inv_x2_sg U77005 ( .A(n22763), .X(n50846) );
  inv_x2_sg U77006 ( .A(n22769), .X(n50893) );
  inv_x2_sg U77007 ( .A(n22775), .X(n50938) );
  inv_x2_sg U77008 ( .A(n44633), .X(n50892) );
  inv_x2_sg U77009 ( .A(n22790), .X(n50924) );
  inv_x2_sg U77010 ( .A(n22793), .X(n50921) );
  inv_x2_sg U77011 ( .A(n45525), .X(n50875) );
  inv_x2_sg U77012 ( .A(n22799), .X(n50915) );
  inv_x2_sg U77013 ( .A(n44647), .X(n50868) );
  inv_x2_sg U77014 ( .A(n22806), .X(n50909) );
  inv_x2_sg U77015 ( .A(n22814), .X(n50867) );
  inv_x2_sg U77016 ( .A(n22818), .X(n50866) );
  inv_x2_sg U77017 ( .A(n22827), .X(n50874) );
  inv_x2_sg U77018 ( .A(n22840), .X(n50880) );
  inv_x2_sg U77019 ( .A(n22788), .X(n50926) );
  inv_x2_sg U77020 ( .A(n22851), .X(n50886) );
  inv_x2_sg U77021 ( .A(n22863), .X(n50891) );
  inv_x2_sg U77022 ( .A(n44072), .X(n50164) );
  inv_x2_sg U77023 ( .A(n22934), .X(n50163) );
  inv_x2_sg U77024 ( .A(n44651), .X(n50210) );
  inv_x2_sg U77025 ( .A(n22941), .X(n50209) );
  inv_x2_sg U77026 ( .A(n44641), .X(n50254) );
  inv_x2_sg U77027 ( .A(n22948), .X(n50253) );
  inv_x2_sg U77028 ( .A(n44583), .X(n50300) );
  inv_x2_sg U77029 ( .A(n22955), .X(n50299) );
  inv_x2_sg U77030 ( .A(n44643), .X(n50346) );
  inv_x2_sg U77031 ( .A(n22962), .X(n50345) );
  inv_x2_sg U77032 ( .A(n44589), .X(n50393) );
  inv_x2_sg U77033 ( .A(n22969), .X(n50392) );
  inv_x2_sg U77034 ( .A(n44593), .X(n50440) );
  inv_x2_sg U77035 ( .A(n22976), .X(n50439) );
  inv_x2_sg U77036 ( .A(n44597), .X(n50486) );
  inv_x2_sg U77037 ( .A(n22983), .X(n50485) );
  inv_x2_sg U77038 ( .A(n44601), .X(n50533) );
  inv_x2_sg U77039 ( .A(n22990), .X(n50532) );
  inv_x2_sg U77040 ( .A(n44605), .X(n50580) );
  inv_x2_sg U77041 ( .A(n22997), .X(n50579) );
  inv_x2_sg U77042 ( .A(n44645), .X(n50629) );
  inv_x2_sg U77043 ( .A(n23004), .X(n50628) );
  inv_x2_sg U77044 ( .A(n44611), .X(n50676) );
  inv_x2_sg U77045 ( .A(n23011), .X(n50675) );
  inv_x2_sg U77046 ( .A(n44615), .X(n50724) );
  inv_x2_sg U77047 ( .A(n23018), .X(n50723) );
  inv_x2_sg U77048 ( .A(n23024), .X(n50770) );
  inv_x2_sg U77049 ( .A(n23030), .X(n50818) );
  inv_x2_sg U77050 ( .A(n23048), .X(n50878) );
  inv_x2_sg U77051 ( .A(n45503), .X(n50831) );
  inv_x2_sg U77052 ( .A(n23054), .X(n50871) );
  inv_x2_sg U77053 ( .A(n23060), .X(n50865) );
  inv_x2_sg U77054 ( .A(n23073), .X(n50823) );
  inv_x2_sg U77055 ( .A(n23082), .X(n50830) );
  inv_x2_sg U77056 ( .A(n23095), .X(n50836) );
  inv_x2_sg U77057 ( .A(n23046), .X(n50881) );
  inv_x2_sg U77058 ( .A(n23043), .X(n50884) );
  inv_x2_sg U77059 ( .A(n23108), .X(n50841) );
  inv_x2_sg U77060 ( .A(n23120), .X(n50862) );
  inv_x2_sg U77061 ( .A(n23268), .X(n50839) );
  inv_x2_sg U77062 ( .A(n23274), .X(n50834) );
  inv_x2_sg U77063 ( .A(n45497), .X(n50787) );
  inv_x2_sg U77064 ( .A(n23280), .X(n50827) );
  inv_x2_sg U77065 ( .A(n23065), .X(n50776) );
  inv_x2_sg U77066 ( .A(n23299), .X(n50779) );
  inv_x2_sg U77067 ( .A(n23308), .X(n50786) );
  inv_x2_sg U77068 ( .A(n23321), .X(n50792) );
  inv_x2_sg U77069 ( .A(n23106), .X(n50795) );
  inv_x2_sg U77070 ( .A(n23332), .X(n50798) );
  inv_x2_sg U77071 ( .A(n23395), .X(n50166) );
  inv_x2_sg U77072 ( .A(n23401), .X(n50214) );
  inv_x2_sg U77073 ( .A(n23407), .X(n50258) );
  inv_x2_sg U77074 ( .A(n23413), .X(n50304) );
  inv_x2_sg U77075 ( .A(n23419), .X(n50350) );
  inv_x2_sg U77076 ( .A(n23425), .X(n50397) );
  inv_x2_sg U77077 ( .A(n23431), .X(n50444) );
  inv_x2_sg U77078 ( .A(n23437), .X(n50490) );
  inv_x2_sg U77079 ( .A(n23443), .X(n50537) );
  inv_x2_sg U77080 ( .A(n23449), .X(n50584) );
  inv_x2_sg U77081 ( .A(n23455), .X(n50633) );
  inv_x2_sg U77082 ( .A(n23461), .X(n50680) );
  inv_x2_sg U77083 ( .A(n23467), .X(n50728) );
  inv_x2_sg U77084 ( .A(n23479), .X(n50790) );
  inv_x2_sg U77085 ( .A(n45505), .X(n50741) );
  inv_x2_sg U77086 ( .A(n23485), .X(n50783) );
  inv_x2_sg U77087 ( .A(n23491), .X(n50778) );
  inv_x2_sg U77088 ( .A(n23504), .X(n50733) );
  inv_x2_sg U77089 ( .A(n23513), .X(n50740) );
  inv_x2_sg U77090 ( .A(n23526), .X(n50746) );
  inv_x2_sg U77091 ( .A(n23477), .X(n50793) );
  inv_x2_sg U77092 ( .A(n23474), .X(n50796) );
  inv_x2_sg U77093 ( .A(n23539), .X(n50774) );
  inv_x2_sg U77094 ( .A(n10197), .X(n50147) );
  inv_x2_sg U77095 ( .A(n23594), .X(n50168) );
  inv_x2_sg U77096 ( .A(n23598), .X(n50232) );
  inv_x2_sg U77097 ( .A(n23604), .X(n50278) );
  inv_x2_sg U77098 ( .A(n23610), .X(n50324) );
  inv_x2_sg U77099 ( .A(n23616), .X(n50371) );
  inv_x2_sg U77100 ( .A(n23622), .X(n50418) );
  inv_x2_sg U77101 ( .A(n23628), .X(n50464) );
  inv_x2_sg U77102 ( .A(n23634), .X(n50511) );
  inv_x2_sg U77103 ( .A(n23640), .X(n50558) );
  inv_x2_sg U77104 ( .A(n23646), .X(n50607) );
  inv_x2_sg U77105 ( .A(n23652), .X(n50656) );
  inv_x2_sg U77106 ( .A(n23658), .X(n50702) );
  inv_x2_sg U77107 ( .A(n23663), .X(n50749) );
  inv_x2_sg U77108 ( .A(n23669), .X(n50744) );
  inv_x2_sg U77109 ( .A(n45499), .X(n50695) );
  inv_x2_sg U77110 ( .A(n23675), .X(n50737) );
  inv_x2_sg U77111 ( .A(n23496), .X(n50684) );
  inv_x2_sg U77112 ( .A(n23694), .X(n50687) );
  inv_x2_sg U77113 ( .A(n23703), .X(n50694) );
  inv_x2_sg U77114 ( .A(n23716), .X(n50700) );
  inv_x2_sg U77115 ( .A(n23537), .X(n50730) );
  inv_x2_sg U77116 ( .A(n10220), .X(n50146) );
  inv_x2_sg U77117 ( .A(n23774), .X(n50170) );
  inv_x2_sg U77118 ( .A(n23780), .X(n50217) );
  inv_x2_sg U77119 ( .A(n23778), .X(n50231) );
  inv_x2_sg U77120 ( .A(n23786), .X(n50262) );
  inv_x2_sg U77121 ( .A(n23784), .X(n50277) );
  inv_x2_sg U77122 ( .A(n23792), .X(n50307) );
  inv_x2_sg U77123 ( .A(n23790), .X(n50323) );
  inv_x2_sg U77124 ( .A(n23798), .X(n50353) );
  inv_x2_sg U77125 ( .A(n23796), .X(n50370) );
  inv_x2_sg U77126 ( .A(n23804), .X(n50401) );
  inv_x2_sg U77127 ( .A(n23802), .X(n50417) );
  inv_x2_sg U77128 ( .A(n23810), .X(n50447) );
  inv_x2_sg U77129 ( .A(n23808), .X(n50463) );
  inv_x2_sg U77130 ( .A(n23816), .X(n50493) );
  inv_x2_sg U77131 ( .A(n23814), .X(n50510) );
  inv_x2_sg U77132 ( .A(n23822), .X(n50541) );
  inv_x2_sg U77133 ( .A(n23820), .X(n50557) );
  inv_x2_sg U77134 ( .A(n23828), .X(n50587) );
  inv_x2_sg U77135 ( .A(n23826), .X(n50606) );
  inv_x2_sg U77136 ( .A(n23831), .X(n50654) );
  inv_x2_sg U77137 ( .A(n23834), .X(n50637) );
  inv_x2_sg U77138 ( .A(n23840), .X(n50698) );
  inv_x2_sg U77139 ( .A(n45507), .X(n50650) );
  inv_x2_sg U77140 ( .A(n23846), .X(n50691) );
  inv_x2_sg U77141 ( .A(n23852), .X(n50686) );
  inv_x2_sg U77142 ( .A(n23865), .X(n50642) );
  inv_x2_sg U77143 ( .A(n23874), .X(n50649) );
  inv_x2_sg U77144 ( .A(n23887), .X(n50683) );
  inv_x2_sg U77145 ( .A(n10200), .X(n50145) );
  inv_x2_sg U77146 ( .A(n23933), .X(n50186) );
  inv_x2_sg U77147 ( .A(n23939), .X(n50230) );
  inv_x2_sg U77148 ( .A(n23945), .X(n50276) );
  inv_x2_sg U77149 ( .A(n23951), .X(n50322) );
  inv_x2_sg U77150 ( .A(n23957), .X(n50369) );
  inv_x2_sg U77151 ( .A(n23963), .X(n50416) );
  inv_x2_sg U77152 ( .A(n23969), .X(n50462) );
  inv_x2_sg U77153 ( .A(n23975), .X(n50509) );
  inv_x2_sg U77154 ( .A(n23981), .X(n50556) );
  inv_x2_sg U77155 ( .A(n23987), .X(n50605) );
  inv_x2_sg U77156 ( .A(n23993), .X(n50653) );
  inv_x2_sg U77157 ( .A(n45501), .X(n50604) );
  inv_x2_sg U77158 ( .A(n23999), .X(n50646) );
  inv_x2_sg U77159 ( .A(n23857), .X(n50593) );
  inv_x2_sg U77160 ( .A(n24018), .X(n50596) );
  inv_x2_sg U77161 ( .A(n24027), .X(n50603) );
  inv_x2_sg U77162 ( .A(n44519), .X(n50174) );
  inv_x2_sg U77163 ( .A(n24081), .X(n50173) );
  inv_x2_sg U77164 ( .A(n44625), .X(n50222) );
  inv_x2_sg U77165 ( .A(n24088), .X(n50221) );
  inv_x2_sg U77166 ( .A(n44627), .X(n50267) );
  inv_x2_sg U77167 ( .A(n24095), .X(n50266) );
  inv_x2_sg U77168 ( .A(n44521), .X(n50312) );
  inv_x2_sg U77169 ( .A(n24102), .X(n50311) );
  inv_x2_sg U77170 ( .A(n44629), .X(n50358) );
  inv_x2_sg U77171 ( .A(n24109), .X(n50357) );
  inv_x2_sg U77172 ( .A(n44523), .X(n50406) );
  inv_x2_sg U77173 ( .A(n24116), .X(n50405) );
  inv_x2_sg U77174 ( .A(n44525), .X(n50452) );
  inv_x2_sg U77175 ( .A(n24123), .X(n50451) );
  inv_x2_sg U77176 ( .A(n44527), .X(n50498) );
  inv_x2_sg U77177 ( .A(n24130), .X(n50497) );
  inv_x2_sg U77178 ( .A(n44657), .X(n50545) );
  inv_x2_sg U77179 ( .A(n24137), .X(n50544) );
  inv_x2_sg U77180 ( .A(n45509), .X(n50592) );
  inv_x2_sg U77181 ( .A(n24143), .X(n50600) );
  inv_x2_sg U77182 ( .A(n24149), .X(n50595) );
  inv_x2_sg U77183 ( .A(n24162), .X(n50550) );
  inv_x2_sg U77184 ( .A(n24171), .X(n50591) );
  inv_x2_sg U77185 ( .A(n24259), .X(n50554) );
  inv_x2_sg U77186 ( .A(n24154), .X(n50502) );
  inv_x2_sg U77187 ( .A(n24278), .X(n50505) );
  inv_x2_sg U77188 ( .A(n44247), .X(n50178) );
  inv_x2_sg U77189 ( .A(n24322), .X(n50177) );
  inv_x2_sg U77190 ( .A(n24328), .X(n50226) );
  inv_x2_sg U77191 ( .A(n24334), .X(n50271) );
  inv_x2_sg U77192 ( .A(n45495), .X(n50317) );
  inv_x2_sg U77193 ( .A(n24341), .X(n50316) );
  inv_x2_sg U77194 ( .A(n24347), .X(n50362) );
  inv_x2_sg U77195 ( .A(n45493), .X(n50411) );
  inv_x2_sg U77196 ( .A(n24354), .X(n50410) );
  inv_x2_sg U77197 ( .A(n24367), .X(n50504) );
  inv_x2_sg U77198 ( .A(n24370), .X(n50456) );
  inv_x2_sg U77199 ( .A(n24358), .X(n50459) );
  inv_x2_sg U77200 ( .A(n24434), .X(n50365) );
  inv_x2_sg U77201 ( .A(n24445), .X(n50458) );
  inv_x2_sg U77202 ( .A(n24461), .X(n50180) );
  inv_x2_sg U77203 ( .A(n24441), .X(n50364) );
  inv_x2_sg U77204 ( .A(n23838), .X(n50701) );
  inv_x2_sg U77205 ( .A(reset), .X(n55511) );
endmodule

