
module pooling ( clk, reset, .im({\im[3][19] , \im[3][18] , \im[3][17] , 
        \im[3][16] , \im[3][15] , \im[3][14] , \im[3][13] , \im[3][12] , 
        \im[3][11] , \im[3][10] , \im[3][9] , \im[3][8] , \im[3][7] , 
        \im[3][6] , \im[3][5] , \im[3][4] , \im[3][3] , \im[3][2] , \im[3][1] , 
        \im[3][0] , \im[2][19] , \im[2][18] , \im[2][17] , \im[2][16] , 
        \im[2][15] , \im[2][14] , \im[2][13] , \im[2][12] , \im[2][11] , 
        \im[2][10] , \im[2][9] , \im[2][8] , \im[2][7] , \im[2][6] , 
        \im[2][5] , \im[2][4] , \im[2][3] , \im[2][2] , \im[2][1] , \im[2][0] , 
        \im[1][19] , \im[1][18] , \im[1][17] , \im[1][16] , \im[1][15] , 
        \im[1][14] , \im[1][13] , \im[1][12] , \im[1][11] , \im[1][10] , 
        \im[1][9] , \im[1][8] , \im[1][7] , \im[1][6] , \im[1][5] , \im[1][4] , 
        \im[1][3] , \im[1][2] , \im[1][1] , \im[1][0] , \im[0][19] , 
        \im[0][18] , \im[0][17] , \im[0][16] , \im[0][15] , \im[0][14] , 
        \im[0][13] , \im[0][12] , \im[0][11] , \im[0][10] , \im[0][9] , 
        \im[0][8] , \im[0][7] , \im[0][6] , \im[0][5] , \im[0][4] , \im[0][3] , 
        \im[0][2] , \im[0][1] , \im[0][0] }), input_ready, output_taken, mode, 
        om, state );
  input [1:0] mode;
  output [19:0] om;
  output [1:0] state;
  input clk, reset, \im[3][19] , \im[3][18] , \im[3][17] , \im[3][16] ,
         \im[3][15] , \im[3][14] , \im[3][13] , \im[3][12] , \im[3][11] ,
         \im[3][10] , \im[3][9] , \im[3][8] , \im[3][7] , \im[3][6] ,
         \im[3][5] , \im[3][4] , \im[3][3] , \im[3][2] , \im[3][1] ,
         \im[3][0] , \im[2][19] , \im[2][18] , \im[2][17] , \im[2][16] ,
         \im[2][15] , \im[2][14] , \im[2][13] , \im[2][12] , \im[2][11] ,
         \im[2][10] , \im[2][9] , \im[2][8] , \im[2][7] , \im[2][6] ,
         \im[2][5] , \im[2][4] , \im[2][3] , \im[2][2] , \im[2][1] ,
         \im[2][0] , \im[1][19] , \im[1][18] , \im[1][17] , \im[1][16] ,
         \im[1][15] , \im[1][14] , \im[1][13] , \im[1][12] , \im[1][11] ,
         \im[1][10] , \im[1][9] , \im[1][8] , \im[1][7] , \im[1][6] ,
         \im[1][5] , \im[1][4] , \im[1][3] , \im[1][2] , \im[1][1] ,
         \im[1][0] , \im[0][19] , \im[0][18] , \im[0][17] , \im[0][16] ,
         \im[0][15] , \im[0][14] , \im[0][13] , \im[0][12] , \im[0][11] ,
         \im[0][10] , \im[0][9] , \im[0][8] , \im[0][7] , \im[0][6] ,
         \im[0][5] , \im[0][4] , \im[0][3] , \im[0][2] , \im[0][1] ,
         \im[0][0] , input_ready, output_taken;
  wire   \reg_im[3][19] , \reg_im[3][18] , \reg_im[3][17] , \reg_im[3][16] ,
         \reg_im[3][15] , \reg_im[3][14] , \reg_im[3][13] , \reg_im[3][12] ,
         \reg_im[3][11] , \reg_im[3][10] , \reg_im[3][9] , \reg_im[3][8] ,
         \reg_im[3][7] , \reg_im[3][6] , \reg_im[3][5] , \reg_im[3][4] ,
         \reg_im[3][3] , \reg_im[3][2] , \reg_im[3][1] , \reg_im[3][0] ,
         \reg_im[2][19] , \reg_im[2][18] , \reg_im[2][17] , \reg_im[2][16] ,
         \reg_im[2][15] , \reg_im[2][14] , \reg_im[2][13] , \reg_im[2][12] ,
         \reg_im[2][11] , \reg_im[2][10] , \reg_im[2][9] , \reg_im[2][8] ,
         \reg_im[2][7] , \reg_im[2][6] , \reg_im[2][5] , \reg_im[2][4] ,
         \reg_im[2][3] , \reg_im[2][2] , \reg_im[2][1] , \reg_im[2][0] ,
         \reg_im[1][19] , \reg_im[1][18] , \reg_im[1][17] , \reg_im[1][16] ,
         \reg_im[1][15] , \reg_im[1][14] , \reg_im[1][13] , \reg_im[1][12] ,
         \reg_im[1][11] , \reg_im[1][10] , \reg_im[1][9] , \reg_im[1][8] ,
         \reg_im[1][7] , \reg_im[1][6] , \reg_im[1][5] , \reg_im[1][4] ,
         \reg_im[1][3] , \reg_im[1][2] , \reg_im[1][1] , \reg_im[1][0] ,
         \reg_im[0][19] , \reg_im[0][18] , \reg_im[0][17] , \reg_im[0][16] ,
         \reg_im[0][15] , \reg_im[0][14] , \reg_im[0][13] , \reg_im[0][12] ,
         \reg_im[0][11] , \reg_im[0][10] , \reg_im[0][9] , \reg_im[0][8] ,
         \reg_im[0][7] , \reg_im[0][6] , \reg_im[0][5] , \reg_im[0][4] ,
         \reg_im[0][3] , \reg_im[0][2] , \reg_im[0][1] , \reg_im[0][0] , N112,
         reg_input_ready, n472, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n5053, n5054,
         \max_pooling_0/n821 , \max_pooling_0/n820 , \max_pooling_0/n819 ,
         \max_pooling_0/n818 , \max_pooling_0/n817 , \max_pooling_0/n816 ,
         \max_pooling_0/n815 , \max_pooling_0/n814 , \max_pooling_0/n813 ,
         \max_pooling_0/n812 , \max_pooling_0/n811 , \max_pooling_0/n810 ,
         \max_pooling_0/n809 , \max_pooling_0/n808 , \max_pooling_0/n807 ,
         \max_pooling_0/n806 , \max_pooling_0/n805 , \max_pooling_0/n804 ,
         \max_pooling_0/n803 , \max_pooling_0/n802 , \max_pooling_0/N4 ,
         \max_pooling_0/N3 , \mean_pooling_0/n212 , \mean_pooling_0/n211 ,
         \mean_pooling_0/n210 , \mean_pooling_0/n209 , \mean_pooling_0/n208 ,
         \mean_pooling_0/n194 , \mean_pooling_0/n193 , \mean_pooling_0/n192 ,
         \mean_pooling_0/n191 , \mean_pooling_0/n190 , \mean_pooling_0/n189 ,
         \mean_pooling_0/n179 , \mean_pooling_0/n178 , \mean_pooling_0/n2 ,
         \mean_pooling_0/n159 , \mean_pooling_0/n687 , \mean_pooling_0/n686 ,
         \mean_pooling_0/n685 , \mean_pooling_0/n684 , \mean_pooling_0/n683 ,
         \mean_pooling_0/n682 , \mean_pooling_0/n681 , \mean_pooling_0/n680 ,
         \mean_pooling_0/n679 , \mean_pooling_0/n678 , \mean_pooling_0/n677 ,
         \mean_pooling_0/n676 , \mean_pooling_0/n675 , \mean_pooling_0/n674 ,
         \mean_pooling_0/n673 , \mean_pooling_0/n672 , \mean_pooling_0/n671 ,
         \mean_pooling_0/n670 , \mean_pooling_0/N5 , \mean_pooling_0/N4 ,
         \min_pooling_0/n452 , \min_pooling_0/n451 , \min_pooling_0/n450 ,
         \min_pooling_0/n449 , \min_pooling_0/n448 , \min_pooling_0/n447 ,
         \min_pooling_0/n446 , \min_pooling_0/n445 , \min_pooling_0/n444 ,
         \min_pooling_0/n443 , \min_pooling_0/n442 , \min_pooling_0/n441 ,
         \min_pooling_0/n440 , \min_pooling_0/n439 , \min_pooling_0/n438 ,
         \min_pooling_0/n437 , \min_pooling_0/n436 , \min_pooling_0/n435 ,
         \min_pooling_0/n434 , \min_pooling_0/n433 , \min_pooling_0/n306 ,
         \min_pooling_0/n305 , \min_pooling_0/n304 , \min_pooling_0/n303 ,
         \min_pooling_0/n302 , \min_pooling_0/n301 , \min_pooling_0/n300 ,
         \min_pooling_0/n299 , \min_pooling_0/n298 , \min_pooling_0/n297 ,
         \min_pooling_0/n296 , \min_pooling_0/n295 , \min_pooling_0/n294 ,
         \min_pooling_0/n293 , \min_pooling_0/n292 , \min_pooling_0/n291 ,
         \min_pooling_0/n290 , \min_pooling_0/n289 , \min_pooling_0/n288 ,
         \min_pooling_0/n287 , \min_pooling_0/n873 , \min_pooling_0/n872 ,
         \min_pooling_0/n871 , \min_pooling_0/n870 , \min_pooling_0/n869 ,
         \min_pooling_0/n868 , \min_pooling_0/n867 , \min_pooling_0/n866 ,
         \min_pooling_0/n865 , \min_pooling_0/n864 , \min_pooling_0/n863 ,
         \min_pooling_0/n862 , \min_pooling_0/n861 , \min_pooling_0/n860 ,
         \min_pooling_0/n859 , \min_pooling_0/n858 , \min_pooling_0/n857 ,
         \min_pooling_0/n856 , \min_pooling_0/n855 , \min_pooling_0/n854 ,
         \min_pooling_0/N4 , \min_pooling_0/N3 , n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n470, n469, n466, n465, n462, n461, n458, n457, n454, n453,
         n450, n449, n446, n445, n442, n441, n438, n437, n434, n433, n430,
         n429, n426, n425, n422, n421, n418, n417, n414, n413, n410, n409,
         n406, n405, n402, n401, n398, n397, n394, n393, n390, n386, n385,
         n382, n381, n378, n377, n2756, n2755, n2754, n2753, n2752, n2751,
         n2750, n2749, n2748, n2747, n2746, n2745, n2744, n2743, n2742, n2741,
         n2740, n2739, n2738, n2737, n2736, n2735, n2734, n2733, n2732, n2731,
         n2730, n2729, n2728, n2727, n2726, n2725, n2724, n2723, n2722, n2721,
         n2720, n2719, n2718, n2717, n2716, n2715, n2714, n2713, n2712, n2711,
         n2710, n2709, n2708, n2707, n2706, n2705, n2704, n2703, n2702, n2701,
         n2700, n2699, n2698, n2697, n2696, n2695, n2694, n2693, n2692, n2691,
         n2690, n2689, n2688, n2687, n2686, n2685, n2684, n2683, n2682, n2681,
         n2680, n2679, n2678, n2677, n2676, n2675, n2674, n2673, n2672, n2671,
         n2670, n2669, n2668, n2667, n2666, n2665, n2664, n2663, n2662, n2661,
         n2660, n2659, n2658, n2657, n2656, n2655, n2654, n2653, n2652, n2651,
         n2650, n2649, n2648, n2647, n2646, n2645, n2644, n2643, n2642, n2641,
         n2640, n2639, n2638, n2637, n2636, n2635, n2634, n2633, n2632, n2631,
         n2630, n2629, n2628, n2627, n2626, n2625, n2624, n2623, n2622, n2621,
         n2620, n2619, n2618, n2617, n2616, n2615, n2614, n2613, n2612, n2611,
         n2610, n2609, n2608, n2607, n2606, n2605, n2604, n2603, n2602, n2601,
         n2600, n2599, n2598, n2597, n2596, n2595, n2594, n2593, n2592, n2591,
         n2590, n2589, n2588, n2587, n2586, n2585, n2584, n2583, n2582, n2581,
         n2580, n2579, n2578, n2577, n2576, n2575, n2574, n2573, n2572, n2571,
         n2570, n2569, n2568, n2567, n2566, n2565, n2564, n2563, n2562, n2561,
         n2560, n2559, n2558, n2557, n2556, n2555, n2554, n2553, n2552, n2551,
         n2550, n2549, n2548, n2547, n2546, n2545, n2544, n2543, n2542, n2541,
         n2540, n2539, n2538, n2537, n2536, n2535, n2534, n2533, n2532, n2531,
         n2530, n2529, n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521,
         n2520, n2519, n2518, n2517, n2516, n2515, n2514, n2513, n2512, n2511,
         n2510, n2509, n2508, n2507, n2506, n2505, n2504, n2503, n2502, n2501,
         n2500, n2499, n2498, n2497, n2496, n2495, n2494, n2493, n2492, n2491,
         n2490, n2489, n2488, n2487, n2486, n2485, n2484, n2483, n2482, n2481,
         n2480, n2479, n2478, n2477, n2476, n2475, n2474, n2473, n2472, n2471,
         n2470, n2469, n2468, n2467, n2466, n2465, n2464, n2463, n2462, n2461,
         n2460, n2459, n2458, n2457, n2456, n2455, n2454, n2453, n2452, n2451,
         n2450, n2449, n2448, n2447, n2446, n2445, n2444, n2443, n2442, n2441,
         n2440, n2439, n2438, n2437, n2436, n2435, n2434, n2433, n2432, n2431,
         n2430, n2429, n2428, n2427, n2426, n2425, n2424, n2423, n2422, n2421,
         n2420, n2419, n2418, n2417, n2416, n2415, n2414, n2413, n2412, n2411,
         n2410, n2409, n2408, n2407, n2406, n2405, n2404, n2403, n2402, n2401,
         n2400, n2399, n2398, n2397, n2396, n2395, n2394, n2393, n2392, n2391,
         n2390, n2389, n2388, n2387, n2386, n2385, n2384, n2383, n2382, n2381,
         n2380, n2379, n2378, n2377, n2376, n2375, n2374, n2373, n2372, n2371,
         n2370, n2369, n2368, n2367, n2366, n2365, n2364, n2363, n2362, n2361,
         n2360, n2359, n2358, n2357, n2356, n2355, n2354, n2353, n2352, n2351,
         n2350, n2349, n2348, n2347, n2346, n2345, n2344, n2343, n2342, n2341,
         n2340, n2339, n2338, n2337, n2336, n2335, n2334, n2333, n2332, n2331,
         n2330, n2329, n2328, n2327, n2326, n2325, n2324, n2323, n2322, n2321,
         n2320, n2319, n2318, n2317, n2316, n2315, n2314, n2313, n2312, n2311,
         n2310, n2309, n2308, n2307, n2306, n2305, n2304, n2303, n2302, n2301,
         n2300, n2299, n2298, n2297, n2296, n2295, n2294, n2293, n2292, n2291,
         n2290, n2289, n2288, n2287, n2286, n2285, n2284, n2283, n2282, n2281,
         n2280, n2279, n2278, n2277, n2276, n2275, n2274, n2273, n2272, n2271,
         n2270, n2269, n2268, n2267, n2266, n2265, n2264, n2263, n2262, n2261,
         n2260, n2259, n2258, n2257, n2256, n2255, n2254, n2253, n2252, n2251,
         n2250, n2249, n2248, n2247, n2246, n2245, n2244, n2243, n2242, n2241,
         n2240, n2239, n2238, n2237, n2236, n2235, n2234, n2233, n2232, n2231,
         n2230, n2229, n2228, n2227, n2226, n2225, n2224, n2223, n2222, n2221,
         n2220, n2219, n2218, n2217, n2216, n2215, n2214, n2213, n2212, n2211,
         n2210, n2209, n2208, n2207, n2206, n2205, n2204, n2203, n2202, n2201,
         n2200, n2199, n2198, n2197, n2196, n2195, n2194, n2193, n2192, n2191,
         n2190, n2189, n2188, n2187, n2186, n2185, n2184, n2183, n2182, n2181,
         n2180, n2179, n2178, n2177, n2176, n2175, n2174, n2173, n2172, n2171,
         n2170, n2169, n2168, n2167, n2166, n2165, n2164, n2163, n2162, n2161,
         n2160, n2159, n2158, n2157, n2156, n2155, n2154, n2153, n2152, n2151,
         n2150, n2149, n2148, n2147, n2146, n2145, n2144, n2143, n2142, n2141,
         n2140, n2139, n2138, n2137, n2136, n2135, n2134, n2133, n2132, n2131,
         n2130, n2129, n2128, n2127, n2126, n2125, n2124, n2123, n2122, n2121,
         n2120, n2119, n2118, n2117, n2116, n2115, n2114, n2113, n2112, n2111,
         n2110, n2109, n2108, n2107, n2106, n2105, n2104, n2103, n2102, n2101,
         n2100, n2099, n2098, n2097, n2096, n2095, n2094, n2093, n2092, n2091,
         n2090, n2089, n2088, n2087, n2086, n2085, n2084, n2083, n2082, n2081,
         n2080, n2079, n2078, n2077, n2076, n2075, n2074, n2073, n2072, n2071,
         n2070, n2069, n2068, n2067, n2066, n2065, n2064, n2063, n2062, n2061,
         n2060, n2059, n2058, n2057, n2056, n2055, n2054, n2053, n2052, n2051,
         n2050, n2049, n2048, n2047, n2046, n2045, n2044, n2043, n2042, n2041,
         n2040, n2039, n2038, n2037, n2036, n2035, n2034, n2033, n2032, n2031,
         n2030, n2029, n2028, n2027, n2026, n2025, n2024, n2023, n2022, n2021,
         n2020, n2019, n2018, n2017, n2016, n2015, n2014, n2013, n2012, n2011,
         n2010, n2009, n2008, n2007, n2006, n2005, n2004, n2003, n2002, n2001,
         n2000, n1999, n1998, n1997, n1996, n1995, n1994, n1993, n1992, n1991,
         n1990, n1989, n1988, n1987, n1986, n1985, n1984, n1983, n1982, n1981,
         n1980, n1979, n1978, n1977, n1976, n1975, n1974, n1973, n1972, n1971,
         n1970, n1969, n1968, n1967, n1966, n1965, n1964, n1963, n1962, n1961,
         n1960, n1959, n1958, n1957, n1956, n1955, n1954, n1953, n1952, n1951,
         n1950, n1949, n1948, n1947, n1946, n1945, n1944, n1943, n1942, n1941,
         n1940, n1939, n1938, n1937, n1936, n1935, n1934, n1933, n1932, n1931,
         n1930, n1929, n1928, n1927, n1926, n1925, n1924, n1923, n1922, n1921,
         n1920, n1919, n1918, n1917, n1916, n1915, n1914, n1913, n1912, n1911,
         n1910, n1909, n1908, n1907, n1906, n1905, n1904, n1903, n1902, n1901,
         n1900, n1899, n1898, n1897, n1896, n1895, n1894, n1893, n1892, n1891,
         n1890, n1889, n1888, n1887, n1886, n1885, n1884, n1883, n1882, n1881,
         n1880, n1879, n1878, n1877, n1876, n1875, n1874, n1873, n1872, n1871,
         n1870, n1869, n1868, n1867, n1866, n1865, n1864, n1863, n1862, n1861,
         n1860, n1859, n1858, n1857, n1856, n1855, n1854, n1853, n1852, n1851,
         n1850, n1849, n1848, n1847, n1846, n1845, n1844, n1843, n1842, n1841,
         n1840, n1839, n1838, n1837, n1836, n1835, n1834, n1833, n1832, n1831,
         n1830, n1829, n1828, n1827, n1826, n1825, n1824, n1823, n1822, n1821,
         n1820, n1819, n1818, n1817, n1816, n1815, n1814, n1813, n1812, n1811,
         n1810, n1809, n1808, n1807, n1806, n1805, n1804, n1803, n1802, n1801,
         n1800, n1799, n1798, n1797, n1796, n1795, n1794, n1793, n1792, n1791,
         n1790, n1789, n1788, n1787, n1786, n1785, n1784, n1783, n1782, n1781,
         n1780, n1779, n1778, n1777, n1776, n1775, n1774, n1773, n1772, n1771,
         n1770, n1769, n1768, n1767, n1766, n1765, n1764, n1763, n1762, n1761,
         n1760, n1759, n1758, n1757, n1756, n1755, n1754, n1753, n1752, n1751,
         n1750, n1749, n1748, n1747, n1746, n1745, n1744, n1743, n1742, n1741,
         n1740, n1739, n1738, n1737, n1736, n1735, n1734, n1733, n1732, n1731,
         n1730, n1729, n1728, n1727, n1726, n1725, n1724, n1723, n1722, n1721,
         n1720, n1719, n1718, n1717, n1716, n1715, n1714, n1713, n1712, n1711,
         n1710, n1709, n1708, n1707, n1706, n1705, n1704, n1703, n1702, n1701,
         n1700, n1699, n1698, n1697, n1696, n1695, n1694, n1693, n1692, n1691,
         n1690, n1689, n1688, n1687, n1686, n1685, n1684, n1683, n1682, n1681,
         n1680, n1679, n1678, n1677, n1676, n1675, n1674, n1673, n1672, n1671,
         n1670, n1669, n1668, n1667, n1666, n1665, n1664, n1663, n1662, n1661,
         n1660, n1659, n1658, n1657, n1656, n1655, n1654, n1653, n1652, n1651,
         n1650, n1649, n1648, n1647, n1646, n1645, n1644, n1643, n1642, n1641,
         n1640, n1639, n1638, n1637, n1636, n1635, n1634, n1633, n1632, n1631,
         n1630, n1629, n1628, n1627, n1626, n1625, n1624, n1623, n1622, n1621,
         n1620, n1619, n1618, n1617, n1616, n1615, n1614, n1613, n1612, n1611,
         n1610, n1609, n1608, n1607, n1606, n1605, n1604, n1603, n1602, n1601,
         n1600, n1599, n1598, n1597, n1596, n1595, n1594, n1593, n1592, n1591,
         n1590, n1589, n1588, n1587, n1586, \min_pooling_0/n355 ,
         \min_pooling_0/n354 , \mean_pooling_0/n302 , \mean_pooling_0/n298 ,
         \mean_pooling_0/n294 , \mean_pooling_0/n290 , \mean_pooling_0/n286 ,
         \mean_pooling_0/n282 , \mean_pooling_0/n278 , \mean_pooling_0/n274 ,
         \mean_pooling_0/n270 , \mean_pooling_0/n266 , \mean_pooling_0/n262 ,
         \mean_pooling_0/n258 , \mean_pooling_0/n254 , \mean_pooling_0/n250 ,
         \mean_pooling_0/n246 , \mean_pooling_0/n242 , \mean_pooling_0/n238 ,
         \mean_pooling_0/n234 , \mean_pooling_0/n230 , \mean_pooling_0/n226 ,
         \mean_pooling_0/n225 , \mean_pooling_0/n222 , \mean_pooling_0/n175 ,
         \mean_pooling_0/n172 , \mean_pooling_0/n169 , \mean_pooling_0/n166 ,
         \max_pooling_0/n314 , \max_pooling_0/n313 , done_min, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052;

  dff_sg \state_reg[1]  ( .D(n3436), .CP(clk), .Q(n5053) );
  dff_sg \state_reg[0]  ( .D(n3437), .CP(clk), .Q(n5054) );
  dff_sg reg_input_ready_reg ( .D(N112), .CP(clk), .Q(reg_input_ready) );
  dff_sg \reg_im_reg[3][19]  ( .D(n475), .CP(clk), .Q(\reg_im[3][19] ) );
  dff_sg \reg_im_reg[3][18]  ( .D(n476), .CP(clk), .Q(\reg_im[3][18] ) );
  dff_sg \reg_im_reg[3][17]  ( .D(n477), .CP(clk), .Q(\reg_im[3][17] ) );
  dff_sg \reg_im_reg[3][16]  ( .D(n478), .CP(clk), .Q(\reg_im[3][16] ) );
  dff_sg \reg_im_reg[3][15]  ( .D(n479), .CP(clk), .Q(\reg_im[3][15] ) );
  dff_sg \reg_im_reg[3][14]  ( .D(n480), .CP(clk), .Q(\reg_im[3][14] ) );
  dff_sg \reg_im_reg[3][13]  ( .D(n481), .CP(clk), .Q(\reg_im[3][13] ) );
  dff_sg \reg_im_reg[3][12]  ( .D(n482), .CP(clk), .Q(\reg_im[3][12] ) );
  dff_sg \reg_im_reg[3][11]  ( .D(n483), .CP(clk), .Q(\reg_im[3][11] ) );
  dff_sg \reg_im_reg[3][10]  ( .D(n484), .CP(clk), .Q(\reg_im[3][10] ) );
  dff_sg \reg_im_reg[3][9]  ( .D(n485), .CP(clk), .Q(\reg_im[3][9] ) );
  dff_sg \reg_im_reg[3][8]  ( .D(n486), .CP(clk), .Q(\reg_im[3][8] ) );
  dff_sg \reg_im_reg[3][7]  ( .D(n487), .CP(clk), .Q(\reg_im[3][7] ) );
  dff_sg \reg_im_reg[3][6]  ( .D(n488), .CP(clk), .Q(\reg_im[3][6] ) );
  dff_sg \reg_im_reg[3][5]  ( .D(n489), .CP(clk), .Q(\reg_im[3][5] ) );
  dff_sg \reg_im_reg[3][4]  ( .D(n490), .CP(clk), .Q(\reg_im[3][4] ) );
  dff_sg \reg_im_reg[3][3]  ( .D(n491), .CP(clk), .Q(\reg_im[3][3] ) );
  dff_sg \reg_im_reg[3][2]  ( .D(n492), .CP(clk), .Q(\reg_im[3][2] ) );
  dff_sg \reg_im_reg[3][1]  ( .D(n493), .CP(clk), .Q(\reg_im[3][1] ) );
  dff_sg \reg_im_reg[3][0]  ( .D(n494), .CP(clk), .Q(\reg_im[3][0] ) );
  dff_sg \reg_im_reg[2][19]  ( .D(n495), .CP(clk), .Q(\reg_im[2][19] ) );
  dff_sg \reg_im_reg[2][18]  ( .D(n496), .CP(clk), .Q(\reg_im[2][18] ) );
  dff_sg \reg_im_reg[2][17]  ( .D(n497), .CP(clk), .Q(\reg_im[2][17] ) );
  dff_sg \reg_im_reg[2][16]  ( .D(n498), .CP(clk), .Q(\reg_im[2][16] ) );
  dff_sg \reg_im_reg[2][15]  ( .D(n499), .CP(clk), .Q(\reg_im[2][15] ) );
  dff_sg \reg_im_reg[2][14]  ( .D(n500), .CP(clk), .Q(\reg_im[2][14] ) );
  dff_sg \reg_im_reg[2][13]  ( .D(n501), .CP(clk), .Q(\reg_im[2][13] ) );
  dff_sg \reg_im_reg[2][12]  ( .D(n502), .CP(clk), .Q(\reg_im[2][12] ) );
  dff_sg \reg_im_reg[2][11]  ( .D(n503), .CP(clk), .Q(\reg_im[2][11] ) );
  dff_sg \reg_im_reg[2][10]  ( .D(n504), .CP(clk), .Q(\reg_im[2][10] ) );
  dff_sg \reg_im_reg[2][9]  ( .D(n505), .CP(clk), .Q(\reg_im[2][9] ) );
  dff_sg \reg_im_reg[2][8]  ( .D(n506), .CP(clk), .Q(\reg_im[2][8] ) );
  dff_sg \reg_im_reg[2][7]  ( .D(n507), .CP(clk), .Q(\reg_im[2][7] ) );
  dff_sg \reg_im_reg[2][6]  ( .D(n508), .CP(clk), .Q(\reg_im[2][6] ) );
  dff_sg \reg_im_reg[2][5]  ( .D(n509), .CP(clk), .Q(\reg_im[2][5] ) );
  dff_sg \reg_im_reg[2][4]  ( .D(n510), .CP(clk), .Q(\reg_im[2][4] ) );
  dff_sg \reg_im_reg[2][3]  ( .D(n511), .CP(clk), .Q(\reg_im[2][3] ) );
  dff_sg \reg_im_reg[2][2]  ( .D(n512), .CP(clk), .Q(\reg_im[2][2] ) );
  dff_sg \reg_im_reg[2][1]  ( .D(n513), .CP(clk), .Q(\reg_im[2][1] ) );
  dff_sg \reg_im_reg[2][0]  ( .D(n514), .CP(clk), .Q(\reg_im[2][0] ) );
  dff_sg \reg_im_reg[1][19]  ( .D(n515), .CP(clk), .Q(\reg_im[1][19] ) );
  dff_sg \reg_im_reg[1][18]  ( .D(n516), .CP(clk), .Q(\reg_im[1][18] ) );
  dff_sg \reg_im_reg[1][17]  ( .D(n517), .CP(clk), .Q(\reg_im[1][17] ) );
  dff_sg \reg_im_reg[1][16]  ( .D(n518), .CP(clk), .Q(\reg_im[1][16] ) );
  dff_sg \reg_im_reg[1][15]  ( .D(n519), .CP(clk), .Q(\reg_im[1][15] ) );
  dff_sg \reg_im_reg[1][14]  ( .D(n520), .CP(clk), .Q(\reg_im[1][14] ) );
  dff_sg \reg_im_reg[1][13]  ( .D(n521), .CP(clk), .Q(\reg_im[1][13] ) );
  dff_sg \reg_im_reg[1][12]  ( .D(n522), .CP(clk), .Q(\reg_im[1][12] ) );
  dff_sg \reg_im_reg[1][11]  ( .D(n523), .CP(clk), .Q(\reg_im[1][11] ) );
  dff_sg \reg_im_reg[1][10]  ( .D(n524), .CP(clk), .Q(\reg_im[1][10] ) );
  dff_sg \reg_im_reg[1][9]  ( .D(n525), .CP(clk), .Q(\reg_im[1][9] ) );
  dff_sg \reg_im_reg[1][8]  ( .D(n526), .CP(clk), .Q(\reg_im[1][8] ) );
  dff_sg \reg_im_reg[1][7]  ( .D(n527), .CP(clk), .Q(\reg_im[1][7] ) );
  dff_sg \reg_im_reg[1][6]  ( .D(n528), .CP(clk), .Q(\reg_im[1][6] ) );
  dff_sg \reg_im_reg[1][5]  ( .D(n529), .CP(clk), .Q(\reg_im[1][5] ) );
  dff_sg \reg_im_reg[1][4]  ( .D(n530), .CP(clk), .Q(\reg_im[1][4] ) );
  dff_sg \reg_im_reg[1][3]  ( .D(n531), .CP(clk), .Q(\reg_im[1][3] ) );
  dff_sg \reg_im_reg[1][2]  ( .D(n532), .CP(clk), .Q(\reg_im[1][2] ) );
  dff_sg \reg_im_reg[1][1]  ( .D(n533), .CP(clk), .Q(\reg_im[1][1] ) );
  dff_sg \reg_im_reg[1][0]  ( .D(n534), .CP(clk), .Q(\reg_im[1][0] ) );
  dff_sg \reg_im_reg[0][19]  ( .D(n535), .CP(clk), .Q(\reg_im[0][19] ) );
  dff_sg \reg_im_reg[0][18]  ( .D(n536), .CP(clk), .Q(\reg_im[0][18] ) );
  dff_sg \reg_im_reg[0][17]  ( .D(n537), .CP(clk), .Q(\reg_im[0][17] ) );
  dff_sg \reg_im_reg[0][16]  ( .D(n538), .CP(clk), .Q(\reg_im[0][16] ) );
  dff_sg \reg_im_reg[0][15]  ( .D(n539), .CP(clk), .Q(\reg_im[0][15] ) );
  dff_sg \reg_im_reg[0][14]  ( .D(n540), .CP(clk), .Q(\reg_im[0][14] ) );
  dff_sg \reg_im_reg[0][13]  ( .D(n541), .CP(clk), .Q(\reg_im[0][13] ) );
  dff_sg \reg_im_reg[0][12]  ( .D(n542), .CP(clk), .Q(\reg_im[0][12] ) );
  dff_sg \reg_im_reg[0][11]  ( .D(n543), .CP(clk), .Q(\reg_im[0][11] ) );
  dff_sg \reg_im_reg[0][10]  ( .D(n544), .CP(clk), .Q(\reg_im[0][10] ) );
  dff_sg \reg_im_reg[0][9]  ( .D(n545), .CP(clk), .Q(\reg_im[0][9] ) );
  dff_sg \reg_im_reg[0][8]  ( .D(n546), .CP(clk), .Q(\reg_im[0][8] ) );
  dff_sg \reg_im_reg[0][7]  ( .D(n547), .CP(clk), .Q(\reg_im[0][7] ) );
  dff_sg \reg_im_reg[0][6]  ( .D(n548), .CP(clk), .Q(\reg_im[0][6] ) );
  dff_sg \reg_im_reg[0][5]  ( .D(n549), .CP(clk), .Q(\reg_im[0][5] ) );
  dff_sg \reg_im_reg[0][4]  ( .D(n550), .CP(clk), .Q(\reg_im[0][4] ) );
  dff_sg \reg_im_reg[0][3]  ( .D(n551), .CP(clk), .Q(\reg_im[0][3] ) );
  dff_sg \reg_im_reg[0][2]  ( .D(n552), .CP(clk), .Q(\reg_im[0][2] ) );
  dff_sg \reg_im_reg[0][1]  ( .D(n553), .CP(clk), .Q(\reg_im[0][1] ) );
  dff_sg \reg_im_reg[0][0]  ( .D(n554), .CP(clk), .Q(\reg_im[0][0] ) );
  dff_sg \max_pooling_0/om_reg[19]  ( .D(n3442), .CP(clk), .Q(
        \max_pooling_0/n802 ) );
  dff_sg \max_pooling_0/om_reg[18]  ( .D(n3460), .CP(clk), .Q(
        \max_pooling_0/n803 ) );
  dff_sg \max_pooling_0/om_reg[17]  ( .D(n3455), .CP(clk), .Q(
        \max_pooling_0/n804 ) );
  dff_sg \max_pooling_0/om_reg[16]  ( .D(n3457), .CP(clk), .Q(
        \max_pooling_0/n805 ) );
  dff_sg \max_pooling_0/om_reg[15]  ( .D(n3454), .CP(clk), .Q(
        \max_pooling_0/n806 ) );
  dff_sg \max_pooling_0/om_reg[14]  ( .D(n3456), .CP(clk), .Q(
        \max_pooling_0/n807 ) );
  dff_sg \max_pooling_0/om_reg[13]  ( .D(n3453), .CP(clk), .Q(
        \max_pooling_0/n808 ) );
  dff_sg \max_pooling_0/om_reg[12]  ( .D(n3443), .CP(clk), .Q(
        \max_pooling_0/n809 ) );
  dff_sg \max_pooling_0/om_reg[11]  ( .D(n3458), .CP(clk), .Q(
        \max_pooling_0/n810 ) );
  dff_sg \max_pooling_0/om_reg[10]  ( .D(n3450), .CP(clk), .Q(
        \max_pooling_0/n811 ) );
  dff_sg \max_pooling_0/om_reg[9]  ( .D(n3459), .CP(clk), .Q(
        \max_pooling_0/n812 ) );
  dff_sg \max_pooling_0/om_reg[8]  ( .D(n3452), .CP(clk), .Q(
        \max_pooling_0/n813 ) );
  dff_sg \max_pooling_0/om_reg[7]  ( .D(n3447), .CP(clk), .Q(
        \max_pooling_0/n814 ) );
  dff_sg \max_pooling_0/om_reg[6]  ( .D(n3448), .CP(clk), .Q(
        \max_pooling_0/n815 ) );
  dff_sg \max_pooling_0/om_reg[5]  ( .D(n3446), .CP(clk), .Q(
        \max_pooling_0/n816 ) );
  dff_sg \max_pooling_0/om_reg[4]  ( .D(n3444), .CP(clk), .Q(
        \max_pooling_0/n817 ) );
  dff_sg \max_pooling_0/om_reg[3]  ( .D(n3441), .CP(clk), .Q(
        \max_pooling_0/n818 ) );
  dff_sg \max_pooling_0/om_reg[2]  ( .D(n3461), .CP(clk), .Q(
        \max_pooling_0/n819 ) );
  dff_sg \max_pooling_0/om_reg[1]  ( .D(n3445), .CP(clk), .Q(
        \max_pooling_0/n820 ) );
  dff_sg \max_pooling_0/om_reg[0]  ( .D(n3449), .CP(clk), .Q(
        \max_pooling_0/n821 ) );
  dff_sg \max_pooling_0/pointer_reg[1]  ( .D(n3440), .CP(clk), .Q(
        \max_pooling_0/N4 ) );
  dff_sg \max_pooling_0/pointer_reg[0]  ( .D(n3451), .CP(clk), .Q(
        \max_pooling_0/N3 ) );
  dff_sg \mean_pooling_0/om_reg[17]  ( .D(n3472), .CP(clk), .Q(
        \mean_pooling_0/n670 ) );
  dff_sg \mean_pooling_0/om_reg[16]  ( .D(n3473), .CP(clk), .Q(
        \mean_pooling_0/n671 ) );
  dff_sg \mean_pooling_0/om_reg[15]  ( .D(n3479), .CP(clk), .Q(
        \mean_pooling_0/n672 ) );
  dff_sg \mean_pooling_0/om_reg[14]  ( .D(n3465), .CP(clk), .Q(
        \mean_pooling_0/n673 ) );
  dff_sg \mean_pooling_0/om_reg[13]  ( .D(n3478), .CP(clk), .Q(
        \mean_pooling_0/n674 ) );
  dff_sg \mean_pooling_0/om_reg[12]  ( .D(n3468), .CP(clk), .Q(
        \mean_pooling_0/n675 ) );
  dff_sg \mean_pooling_0/om_reg[11]  ( .D(n3474), .CP(clk), .Q(
        \mean_pooling_0/n676 ) );
  dff_sg \mean_pooling_0/om_reg[10]  ( .D(n3466), .CP(clk), .Q(
        \mean_pooling_0/n677 ) );
  dff_sg \mean_pooling_0/om_reg[9]  ( .D(n3470), .CP(clk), .Q(
        \mean_pooling_0/n678 ) );
  dff_sg \mean_pooling_0/om_reg[8]  ( .D(n3464), .CP(clk), .Q(
        \mean_pooling_0/n679 ) );
  dff_sg \mean_pooling_0/om_reg[7]  ( .D(n3475), .CP(clk), .Q(
        \mean_pooling_0/n680 ) );
  dff_sg \mean_pooling_0/om_reg[6]  ( .D(n3467), .CP(clk), .Q(
        \mean_pooling_0/n681 ) );
  dff_sg \mean_pooling_0/om_reg[5]  ( .D(n3471), .CP(clk), .Q(
        \mean_pooling_0/n682 ) );
  dff_sg \mean_pooling_0/om_reg[4]  ( .D(n3462), .CP(clk), .Q(
        \mean_pooling_0/n683 ) );
  dff_sg \mean_pooling_0/om_reg[3]  ( .D(n3476), .CP(clk), .Q(
        \mean_pooling_0/n684 ) );
  dff_sg \mean_pooling_0/om_reg[2]  ( .D(n3469), .CP(clk), .Q(
        \mean_pooling_0/n685 ) );
  dff_sg \mean_pooling_0/om_reg[1]  ( .D(n3477), .CP(clk), .Q(
        \mean_pooling_0/n686 ) );
  dff_sg \mean_pooling_0/om_reg[0]  ( .D(n3463), .CP(clk), .Q(
        \mean_pooling_0/n687 ) );
  dff_sg \mean_pooling_0/pointer_reg[1]  ( .D(n3481), .CP(clk), .Q(
        \mean_pooling_0/N5 ) );
  dff_sg \mean_pooling_0/pointer_reg[0]  ( .D(n3480), .CP(clk), .Q(
        \mean_pooling_0/N4 ) );
  dff_sg \min_pooling_0/om_reg[19]  ( .D(\min_pooling_0/n433 ), .CP(clk), .Q(
        \min_pooling_0/n854 ) );
  dff_sg \min_pooling_0/om_reg[18]  ( .D(\min_pooling_0/n434 ), .CP(clk), .Q(
        \min_pooling_0/n855 ) );
  dff_sg \min_pooling_0/om_reg[17]  ( .D(\min_pooling_0/n435 ), .CP(clk), .Q(
        \min_pooling_0/n856 ) );
  dff_sg \min_pooling_0/om_reg[16]  ( .D(\min_pooling_0/n436 ), .CP(clk), .Q(
        \min_pooling_0/n857 ) );
  dff_sg \min_pooling_0/om_reg[15]  ( .D(\min_pooling_0/n437 ), .CP(clk), .Q(
        \min_pooling_0/n858 ) );
  dff_sg \min_pooling_0/om_reg[14]  ( .D(\min_pooling_0/n438 ), .CP(clk), .Q(
        \min_pooling_0/n859 ) );
  dff_sg \min_pooling_0/om_reg[13]  ( .D(\min_pooling_0/n439 ), .CP(clk), .Q(
        \min_pooling_0/n860 ) );
  dff_sg \min_pooling_0/om_reg[12]  ( .D(\min_pooling_0/n440 ), .CP(clk), .Q(
        \min_pooling_0/n861 ) );
  dff_sg \min_pooling_0/om_reg[11]  ( .D(\min_pooling_0/n441 ), .CP(clk), .Q(
        \min_pooling_0/n862 ) );
  dff_sg \min_pooling_0/om_reg[10]  ( .D(\min_pooling_0/n442 ), .CP(clk), .Q(
        \min_pooling_0/n863 ) );
  dff_sg \min_pooling_0/om_reg[9]  ( .D(\min_pooling_0/n443 ), .CP(clk), .Q(
        \min_pooling_0/n864 ) );
  dff_sg \min_pooling_0/om_reg[8]  ( .D(\min_pooling_0/n444 ), .CP(clk), .Q(
        \min_pooling_0/n865 ) );
  dff_sg \min_pooling_0/om_reg[7]  ( .D(\min_pooling_0/n445 ), .CP(clk), .Q(
        \min_pooling_0/n866 ) );
  dff_sg \min_pooling_0/om_reg[6]  ( .D(\min_pooling_0/n446 ), .CP(clk), .Q(
        \min_pooling_0/n867 ) );
  dff_sg \min_pooling_0/om_reg[5]  ( .D(\min_pooling_0/n447 ), .CP(clk), .Q(
        \min_pooling_0/n868 ) );
  dff_sg \min_pooling_0/om_reg[4]  ( .D(\min_pooling_0/n448 ), .CP(clk), .Q(
        \min_pooling_0/n869 ) );
  dff_sg \min_pooling_0/om_reg[3]  ( .D(\min_pooling_0/n449 ), .CP(clk), .Q(
        \min_pooling_0/n870 ) );
  dff_sg \min_pooling_0/om_reg[2]  ( .D(\min_pooling_0/n450 ), .CP(clk), .Q(
        \min_pooling_0/n871 ) );
  dff_sg \min_pooling_0/om_reg[1]  ( .D(\min_pooling_0/n451 ), .CP(clk), .Q(
        \min_pooling_0/n872 ) );
  dff_sg \min_pooling_0/om_reg[0]  ( .D(\min_pooling_0/n452 ), .CP(clk), .Q(
        \min_pooling_0/n873 ) );
  dff_sg \min_pooling_0/pointer_reg[1]  ( .D(n3438), .CP(clk), .Q(
        \min_pooling_0/N4 ) );
  dff_sg \min_pooling_0/pointer_reg[0]  ( .D(n3439), .CP(clk), .Q(
        \min_pooling_0/N3 ) );
  nor_x2_sg U2449 ( .A(n4433), .B(n3061), .X(n3060) );
  nor_x2_sg U2450 ( .A(n3062), .B(n4425), .X(n3059) );
  nor_x2_sg U2457 ( .A(n4433), .B(n3070), .X(n3069) );
  nor_x2_sg U2458 ( .A(n5029), .B(n3071), .X(n3068) );
  nor_x2_sg U2579 ( .A(n3435), .B(\mean_pooling_0/n159 ), .X(n3153) );
  nor_x2_sg U2586 ( .A(n4433), .B(n3162), .X(n3161) );
  nor_x2_sg U2587 ( .A(n4415), .B(n3163), .X(n3160) );
  nor_x2_sg U2829 ( .A(n3326), .B(n3327), .X(n3167) );
  nand_x8_sg U2832 ( .A(n3328), .B(n5023), .X(n3054) );
  nor_x2_sg U2838 ( .A(n4425), .B(\min_pooling_0/n306 ), .X(n3333) );
  nor_x2_sg U2843 ( .A(n4425), .B(\min_pooling_0/n305 ), .X(n3338) );
  nor_x2_sg U2848 ( .A(n4425), .B(\min_pooling_0/n304 ), .X(n3342) );
  nor_x2_sg U2853 ( .A(n4425), .B(\min_pooling_0/n303 ), .X(n3346) );
  nor_x2_sg U2858 ( .A(n4425), .B(\min_pooling_0/n302 ), .X(n3350) );
  nor_x2_sg U2863 ( .A(n4425), .B(\min_pooling_0/n301 ), .X(n3354) );
  nor_x2_sg U2868 ( .A(n4425), .B(\min_pooling_0/n300 ), .X(n3358) );
  nor_x2_sg U2873 ( .A(n4425), .B(\min_pooling_0/n299 ), .X(n3362) );
  nor_x2_sg U2878 ( .A(n4425), .B(\min_pooling_0/n298 ), .X(n3366) );
  nor_x2_sg U2883 ( .A(n4425), .B(\min_pooling_0/n297 ), .X(n3370) );
  nor_x2_sg U2888 ( .A(n4425), .B(\min_pooling_0/n296 ), .X(n3374) );
  nor_x2_sg U2893 ( .A(n4425), .B(\min_pooling_0/n295 ), .X(n3378) );
  nor_x2_sg U2898 ( .A(n4425), .B(\min_pooling_0/n294 ), .X(n3382) );
  nor_x2_sg U2903 ( .A(n4425), .B(\min_pooling_0/n293 ), .X(n3386) );
  nor_x2_sg U2908 ( .A(n4425), .B(\min_pooling_0/n292 ), .X(n3390) );
  nor_x2_sg U2913 ( .A(n4425), .B(\min_pooling_0/n291 ), .X(n3394) );
  nor_x2_sg U2918 ( .A(n4425), .B(\min_pooling_0/n290 ), .X(n3398) );
  nor_x2_sg U2923 ( .A(n4425), .B(\min_pooling_0/n289 ), .X(n3402) );
  nor_x2_sg U2928 ( .A(n4425), .B(\min_pooling_0/n288 ), .X(n3406) );
  nor_x2_sg U2933 ( .A(n4425), .B(\min_pooling_0/n287 ), .X(n3410) );
  nand_x8_sg U2936 ( .A(n4433), .B(n3486), .X(n3334) );
  \**FFGEN**  \om_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n377), .force_10(n378), .force_11(1'b0), .Q(om[0]) );
  \**FFGEN**  \om_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n469), .force_10(n470), .force_11(1'b0), .Q(om[1]) );
  \**FFGEN**  \om_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n465), .force_10(n466), .force_11(1'b0), .Q(om[2]) );
  \**FFGEN**  \om_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n461), .force_10(n462), .force_11(1'b0), .Q(om[3]) );
  \**FFGEN**  \om_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n457), .force_10(n458), .force_11(1'b0), .Q(om[4]) );
  \**FFGEN**  \om_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n453), .force_10(n454), .force_11(1'b0), .Q(om[5]) );
  \**FFGEN**  \om_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n449), .force_10(n450), .force_11(1'b0), .Q(om[6]) );
  \**FFGEN**  \om_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n445), .force_10(n446), .force_11(1'b0), .Q(om[7]) );
  \**FFGEN**  \om_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n441), .force_10(n442), .force_11(1'b0), .Q(om[8]) );
  \**FFGEN**  \om_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n437), .force_10(n438), .force_11(1'b0), .Q(om[9]) );
  \**FFGEN**  \om_reg[10]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n433), .force_10(n434), .force_11(1'b0), .Q(om[10])
         );
  \**FFGEN**  \om_reg[11]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n429), .force_10(n430), .force_11(1'b0), .Q(om[11])
         );
  \**FFGEN**  \om_reg[12]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n425), .force_10(n426), .force_11(1'b0), .Q(om[12])
         );
  \**FFGEN**  \om_reg[13]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n421), .force_10(n422), .force_11(1'b0), .Q(om[13])
         );
  \**FFGEN**  \om_reg[14]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n417), .force_10(n418), .force_11(1'b0), .Q(om[14])
         );
  \**FFGEN**  \om_reg[15]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n413), .force_10(n414), .force_11(1'b0), .Q(om[15])
         );
  \**FFGEN**  \om_reg[16]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n409), .force_10(n410), .force_11(1'b0), .Q(om[16])
         );
  \**FFGEN**  \om_reg[17]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n405), .force_10(n406), .force_11(1'b0), .Q(om[17])
         );
  \**FFGEN**  \om_reg[18]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n401), .force_10(n402), .force_11(1'b0), .Q(om[18])
         );
  \**FFGEN**  \om_reg[19]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n397), .force_10(n398), .force_11(1'b0), .Q(om[19])
         );
  \**FFGEN**  en_mean_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n393), .force_10(n394), .force_11(1'b0), .Q(n3485), 
        .QN(n3435) );
  \**FFGEN**  en_max_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n1686), .force_10(n390), .force_11(1'b0), .QN(n3434)
         );
  \**FFGEN**  en_min_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n385), .force_10(n386), .force_11(1'b0), .Q(n3486), 
        .QN(n3433) );
  \**FFGEN**  done_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), 
        .force_01(n381), .force_10(n382), .force_11(1'b0), .Q(n472) );
  \**FFGEN**  \max_pooling_0/done_reg  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\max_pooling_0/n313 ), .force_10(
        \max_pooling_0/n314 ), .force_11(1'b0), .QN(n1689) );
  \**FFGEN**  \max_pooling_0/max_num_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1614), .force_10(n1611), .force_11(
        1'b0), .Q(n3413) );
  \**FFGEN**  \max_pooling_0/max_num_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1605), .force_10(n1602), .force_11(
        1'b0), .Q(n3414) );
  \**FFGEN**  \max_pooling_0/max_num_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1617), .force_10(n1616), .force_11(
        1'b0), .Q(n3415) );
  \**FFGEN**  \max_pooling_0/max_num_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1619), .force_10(n1618), .force_11(
        1'b0), .Q(n3416) );
  \**FFGEN**  \max_pooling_0/max_num_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1622), .force_10(n1621), .force_11(
        1'b0), .Q(n3417) );
  \**FFGEN**  \max_pooling_0/max_num_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1599), .force_10(n1596), .force_11(
        1'b0), .Q(n3418) );
  \**FFGEN**  \max_pooling_0/max_num_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1624), .force_10(n1593), .force_11(
        1'b0), .Q(n3419) );
  \**FFGEN**  \max_pooling_0/max_num_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1598), .force_10(n1597), .force_11(
        1'b0), .Q(n3420) );
  \**FFGEN**  \max_pooling_0/max_num_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1601), .force_10(n1600), .force_11(
        1'b0), .Q(n3421) );
  \**FFGEN**  \max_pooling_0/max_num_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1592), .force_10(n1591), .force_11(
        1'b0), .Q(n3422) );
  \**FFGEN**  \max_pooling_0/max_num_reg[10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1595), .force_10(n1594), 
        .force_11(1'b0), .Q(n3423) );
  \**FFGEN**  \max_pooling_0/max_num_reg[11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1610), .force_10(n1609), 
        .force_11(1'b0), .Q(n3424) );
  \**FFGEN**  \max_pooling_0/max_num_reg[12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1613), .force_10(n1612), 
        .force_11(1'b0), .Q(n3425) );
  \**FFGEN**  \max_pooling_0/max_num_reg[13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1604), .force_10(n1603), 
        .force_11(1'b0), .Q(n3426) );
  \**FFGEN**  \max_pooling_0/max_num_reg[14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1607), .force_10(n1606), 
        .force_11(1'b0), .Q(n3427) );
  \**FFGEN**  \max_pooling_0/max_num_reg[15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1625), .force_10(n1623), 
        .force_11(1'b0), .Q(n3428) );
  \**FFGEN**  \max_pooling_0/max_num_reg[16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1590), .force_10(n1589), 
        .force_11(1'b0), .Q(n3429) );
  \**FFGEN**  \max_pooling_0/max_num_reg[17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1586), .force_10(n1620), 
        .force_11(1'b0), .Q(n3430) );
  \**FFGEN**  \max_pooling_0/max_num_reg[18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1588), .force_10(n1587), 
        .force_11(1'b0), .Q(n3431) );
  \**FFGEN**  \max_pooling_0/max_num_reg[19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1615), .force_10(n1608), 
        .force_11(1'b0), .Q(n3432) );
  \**FFGEN**  \mean_pooling_0/done_reg  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\mean_pooling_0/n225 ), .force_10(
        \mean_pooling_0/n226 ), .force_11(1'b0), .QN(\mean_pooling_0/n159 ) );
  \**FFGEN**  \mean_pooling_0/sum_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1676), .force_10(
        \mean_pooling_0/n230 ), .force_11(1'b0), .QN(n1687) );
  \**FFGEN**  \mean_pooling_0/sum_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1682), .force_10(
        \mean_pooling_0/n234 ), .force_11(1'b0), .Q(n3503), .QN(n1688) );
  \**FFGEN**  \mean_pooling_0/sum_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1678), .force_10(
        \mean_pooling_0/n238 ), .force_11(1'b0), .Q(\mean_pooling_0/n179 ), 
        .QN(n3501) );
  \**FFGEN**  \mean_pooling_0/sum_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1669), .force_10(
        \mean_pooling_0/n242 ), .force_11(1'b0), .Q(\mean_pooling_0/n194 ), 
        .QN(n3499) );
  \**FFGEN**  \mean_pooling_0/sum_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1684), .force_10(
        \mean_pooling_0/n246 ), .force_11(1'b0), .Q(\mean_pooling_0/n212 ), 
        .QN(n3498) );
  \**FFGEN**  \mean_pooling_0/sum_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1677), .force_10(
        \mean_pooling_0/n250 ), .force_11(1'b0), .Q(\mean_pooling_0/n178 ), 
        .QN(n3488) );
  \**FFGEN**  \mean_pooling_0/sum_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1680), .force_10(
        \mean_pooling_0/n254 ), .force_11(1'b0), .Q(\mean_pooling_0/n193 ), 
        .QN(n3494) );
  \**FFGEN**  \mean_pooling_0/sum_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1666), .force_10(
        \mean_pooling_0/n258 ), .force_11(1'b0), .Q(\mean_pooling_0/n211 ), 
        .QN(n3493) );
  \**FFGEN**  \mean_pooling_0/sum_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1673), .force_10(
        \mean_pooling_0/n262 ), .force_11(1'b0), .Q(n3497), .QN(
        \mean_pooling_0/n166 ) );
  \**FFGEN**  \mean_pooling_0/sum_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1679), .force_10(
        \mean_pooling_0/n266 ), .force_11(1'b0), .Q(\mean_pooling_0/n192 ), 
        .QN(n3492) );
  \**FFGEN**  \mean_pooling_0/sum_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1675), .force_10(
        \mean_pooling_0/n270 ), .force_11(1'b0), .Q(\mean_pooling_0/n210 ), 
        .QN(n3491) );
  \**FFGEN**  \mean_pooling_0/sum_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1674), .force_10(
        \mean_pooling_0/n274 ), .force_11(1'b0), .Q(n3496), .QN(
        \mean_pooling_0/n169 ) );
  \**FFGEN**  \mean_pooling_0/sum_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1668), .force_10(
        \mean_pooling_0/n278 ), .force_11(1'b0), .Q(\mean_pooling_0/n191 ), 
        .QN(n3490) );
  \**FFGEN**  \mean_pooling_0/sum_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1681), .force_10(
        \mean_pooling_0/n282 ), .force_11(1'b0), .Q(\mean_pooling_0/n209 ), 
        .QN(n3489) );
  \**FFGEN**  \mean_pooling_0/sum_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1671), .force_10(
        \mean_pooling_0/n286 ), .force_11(1'b0), .Q(n3495), .QN(
        \mean_pooling_0/n172 ) );
  \**FFGEN**  \mean_pooling_0/sum_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1685), .force_10(
        \mean_pooling_0/n290 ), .force_11(1'b0), .Q(\mean_pooling_0/n190 ), 
        .QN(n3487) );
  \**FFGEN**  \mean_pooling_0/sum_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1667), .force_10(
        \mean_pooling_0/n294 ), .force_11(1'b0), .Q(\mean_pooling_0/n208 ) );
  \**FFGEN**  \mean_pooling_0/sum_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1670), .force_10(
        \mean_pooling_0/n298 ), .force_11(1'b0), .Q(n3500), .QN(
        \mean_pooling_0/n175 ) );
  \**FFGEN**  \mean_pooling_0/sum_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1683), .force_10(
        \mean_pooling_0/n302 ), .force_11(1'b0), .Q(\mean_pooling_0/n189 ), 
        .QN(n3502) );
  \**FFGEN**  \mean_pooling_0/sum_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1672), .force_10(
        \mean_pooling_0/n222 ), .force_11(1'b0), .Q(\mean_pooling_0/n2 ) );
  \**FFGEN**  \min_pooling_0/done_reg  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\min_pooling_0/n354 ), .force_10(
        \min_pooling_0/n355 ), .force_11(1'b0), .Q(done_min) );
  \**FFGEN**  \min_pooling_0/min_num_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1654), .force_10(n1651), .force_11(
        1'b0), .QN(\min_pooling_0/n306 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1645), .force_10(n1642), .force_11(
        1'b0), .QN(\min_pooling_0/n305 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1657), .force_10(n1656), .force_11(
        1'b0), .QN(\min_pooling_0/n304 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1659), .force_10(n1658), .force_11(
        1'b0), .QN(\min_pooling_0/n303 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1662), .force_10(n1661), .force_11(
        1'b0), .QN(\min_pooling_0/n302 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1639), .force_10(n1636), .force_11(
        1'b0), .QN(\min_pooling_0/n301 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1664), .force_10(n1633), .force_11(
        1'b0), .QN(\min_pooling_0/n300 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1638), .force_10(n1637), .force_11(
        1'b0), .QN(\min_pooling_0/n299 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1641), .force_10(n1640), .force_11(
        1'b0), .QN(\min_pooling_0/n298 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n1632), .force_10(n1631), .force_11(
        1'b0), .QN(\min_pooling_0/n297 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1635), .force_10(n1634), 
        .force_11(1'b0), .QN(\min_pooling_0/n296 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1650), .force_10(n1649), 
        .force_11(1'b0), .QN(\min_pooling_0/n295 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1653), .force_10(n1652), 
        .force_11(1'b0), .QN(\min_pooling_0/n294 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1644), .force_10(n1643), 
        .force_11(1'b0), .QN(\min_pooling_0/n293 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1647), .force_10(n1646), 
        .force_11(1'b0), .QN(\min_pooling_0/n292 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1665), .force_10(n1663), 
        .force_11(1'b0), .QN(\min_pooling_0/n291 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1630), .force_10(n1629), 
        .force_11(1'b0), .QN(\min_pooling_0/n290 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1626), .force_10(n1660), 
        .force_11(1'b0), .QN(\min_pooling_0/n289 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1628), .force_10(n1627), 
        .force_11(1'b0), .QN(\min_pooling_0/n288 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n1655), .force_10(n1648), 
        .force_11(1'b0), .QN(\min_pooling_0/n287 ) );
  nor_x2_sg U1299 ( .A(n2011), .B(n2012), .X(n1835) );
  nor_x2_sg U1298 ( .A(n2019), .B(n2020), .X(n2011) );
  nor_x2_sg U1297 ( .A(n2021), .B(n1840), .X(n2019) );
  nor_x2_sg U1296 ( .A(n2030), .B(n2031), .X(n2021) );
  nand_x8_sg U1294 ( .A(n3915), .B(n3975), .X(n1745) );
  nand_x8_sg U1291 ( .A(n4102), .B(n5052), .X(n3061) );
  nand_x8_sg U1286 ( .A(n5052), .B(n4801), .X(n1905) );
  nand_x8_sg U1283 ( .A(n4112), .B(n4801), .X(n3062) );
  nand_x8_sg U1280 ( .A(n3917), .B(n3977), .X(n1821) );
  nand_x8_sg U1269 ( .A(n3913), .B(n3973), .X(n1826) );
  nor_x2_sg U1251 ( .A(n1837), .B(n1838), .X(n1836) );
  nor_x2_sg U1247 ( .A(n1857), .B(n1858), .X(n1855) );
  nand_x8_sg U1234 ( .A(n3921), .B(n3945), .X(n1786) );
  nand_x8_sg U1222 ( .A(n3919), .B(n3943), .X(n1732) );
  nor_x2_sg U1184 ( .A(n1864), .B(n1865), .X(n1863) );
  nor_x2_sg U1183 ( .A(n4092), .B(n1869), .X(n1864) );
  nand_x8_sg U1168 ( .A(n3923), .B(n3947), .X(n1793) );
  nor_x2_sg U1159 ( .A(n1876), .B(n1877), .X(n1874) );
  nor_x2_sg U1127 ( .A(n1938), .B(n1939), .X(n1880) );
  nand_x8_sg U1112 ( .A(n3925), .B(n3969), .X(n1750) );
  nand_x8_sg U1088 ( .A(n3927), .B(n3979), .X(n1783) );
  nor_x2_sg U1047 ( .A(n1847), .B(n1848), .X(n1846) );
  nor_x2_sg U1046 ( .A(n1849), .B(n1850), .X(n1847) );
  nand_x8_sg U1780 ( .A(n4433), .B(n3485), .X(n3154) );
  nor_x2_sg U1325 ( .A(n2750), .B(\mean_pooling_0/n2 ), .X(n2748) );
  nand_x8_sg U1770 ( .A(n4104), .B(n5051), .X(n3162) );
  nand_x8_sg U1765 ( .A(n5051), .B(n4815), .X(n2637) );
  nand_x8_sg U1762 ( .A(n4114), .B(n4815), .X(n3163) );
  nand_x8_sg U1341 ( .A(n3889), .B(n3949), .X(n2449) );
  nand_x8_sg U1364 ( .A(n3881), .B(n3933), .X(n2455) );
  nand_x8_sg U1396 ( .A(n2587), .B(n2588), .X(n2466) );
  nand_x8_sg U1413 ( .A(n3891), .B(n3941), .X(n2470) );
  nand_x8_sg U1436 ( .A(n3883), .B(n3935), .X(n2476) );
  nand_x8_sg U1461 ( .A(n3893), .B(n3951), .X(n2484) );
  nand_x8_sg U1485 ( .A(n3895), .B(n3953), .X(n2491) );
  nand_x8_sg U1508 ( .A(n3885), .B(n3937), .X(n2497) );
  nand_x8_sg U1533 ( .A(n3897), .B(n3955), .X(n2505) );
  nand_x8_sg U1557 ( .A(n3899), .B(n3957), .X(n2512) );
  nand_x8_sg U1580 ( .A(n3887), .B(n3939), .X(n2518) );
  nand_x8_sg U1605 ( .A(n3901), .B(n3959), .X(n2526) );
  nand_x8_sg U1629 ( .A(n3903), .B(n3961), .X(n2533) );
  nand_x8_sg U1653 ( .A(n3905), .B(n3963), .X(n2540) );
  nand_x8_sg U1677 ( .A(n3907), .B(n3965), .X(n2547) );
  nand_x8_sg U1701 ( .A(n3909), .B(n3967), .X(n2554) );
  nand_x8_sg U1747 ( .A(n3911), .B(n3983), .X(n2568) );
  nor_x2_sg U1313 ( .A(n5013), .B(\mean_pooling_0/n189 ), .X(n2579) );
  nor_x2_sg U1357 ( .A(n2454), .B(n2455), .X(n2453) );
  nor_x2_sg U1398 ( .A(n2464), .B(n4994), .X(n2462) );
  nor_x2_sg U1397 ( .A(n2466), .B(\mean_pooling_0/n208 ), .X(n2464) );
  nor_x2_sg U1429 ( .A(n2475), .B(n2476), .X(n2474) );
  nor_x2_sg U1501 ( .A(n2496), .B(n2497), .X(n2495) );
  nor_x2_sg U1573 ( .A(n2517), .B(n2518), .X(n2516) );
  nor_x2_sg U1733 ( .A(n2562), .B(n2563), .X(n2560) );
  nor_x2_sg U1740 ( .A(n2567), .B(n2568), .X(n2566) );
  nor_x2_sg U2246 ( .A(n2324), .B(n2325), .X(n2149) );
  nor_x2_sg U2245 ( .A(n2332), .B(n2333), .X(n2324) );
  nor_x2_sg U2244 ( .A(n2334), .B(n2154), .X(n2332) );
  nor_x2_sg U2243 ( .A(n2343), .B(n2344), .X(n2334) );
  nand_x8_sg U2237 ( .A(n4100), .B(n5050), .X(n3070) );
  nand_x8_sg U2229 ( .A(n5050), .B(n4834), .X(n2218) );
  nand_x8_sg U2226 ( .A(n4110), .B(n4834), .X(n3071) );
  nand_x8_sg U2193 ( .A(n3929), .B(n3971), .X(n2090) );
  nor_x2_sg U2182 ( .A(n2151), .B(n2152), .X(n2150) );
  nor_x2_sg U2178 ( .A(n2171), .B(n2172), .X(n2169) );
  nand_x8_sg U2147 ( .A(n3931), .B(n3981), .X(n2093) );
  nor_x2_sg U2122 ( .A(n4965), .B(n2285), .X(n2176) );
  nor_x2_sg U2095 ( .A(n2178), .B(n2179), .X(n2177) );
  nor_x2_sg U2094 ( .A(n2182), .B(n2183), .X(n2178) );
  nor_x2_sg U2062 ( .A(n2190), .B(n2191), .X(n2188) );
  nor_x2_sg U2002 ( .A(n2205), .B(n2206), .X(n2204) );
  nor_x2_sg U1984 ( .A(n2224), .B(n2225), .X(n2222) );
  nor_x2_sg U1921 ( .A(n2161), .B(n4991), .X(n2160) );
  nor_x2_sg U1920 ( .A(n2163), .B(n2164), .X(n2161) );
  nor_x2_sg U1919 ( .A(n4978), .B(n2165), .X(n2163) );
  nor_x2_sg U2258 ( .A(n1689), .B(n4410), .X(n2439) );
  nor_x2_sg U2257 ( .A(\mean_pooling_0/n159 ), .B(n4408), .X(n2440) );
  nand_x8_sg U2420 ( .A(mode[1]), .B(n5020), .X(n2436) );
  nor_x2_sg U2284 ( .A(n4833), .B(n4408), .X(n2425) );
  nor_x2_sg U2292 ( .A(n4832), .B(n4408), .X(n2421) );
  nor_x2_sg U2300 ( .A(n4831), .B(n4408), .X(n2417) );
  nor_x2_sg U2308 ( .A(n4830), .B(n4408), .X(n2413) );
  nor_x2_sg U2316 ( .A(n4829), .B(n4408), .X(n2409) );
  nor_x2_sg U2324 ( .A(n4828), .B(n4408), .X(n2405) );
  nor_x2_sg U2332 ( .A(n4827), .B(n4408), .X(n2401) );
  nor_x2_sg U2340 ( .A(n4826), .B(n4408), .X(n2397) );
  nor_x2_sg U2348 ( .A(n4825), .B(n4408), .X(n2393) );
  nor_x2_sg U2356 ( .A(n4824), .B(n4408), .X(n2389) );
  nor_x2_sg U2364 ( .A(n4823), .B(n4408), .X(n2385) );
  nor_x2_sg U2372 ( .A(n4822), .B(n4408), .X(n2381) );
  nor_x2_sg U2380 ( .A(n4821), .B(n4408), .X(n2377) );
  nor_x2_sg U2388 ( .A(n4820), .B(n4408), .X(n2373) );
  nor_x2_sg U2396 ( .A(n4819), .B(n4408), .X(n2369) );
  nor_x2_sg U2404 ( .A(n4818), .B(n4408), .X(n2365) );
  nor_x2_sg U2412 ( .A(n4817), .B(n4408), .X(n2361) );
  nor_x2_sg U2427 ( .A(n4816), .B(n4408), .X(n2445) );
  nor_x1_sg U2947 ( .A(n2585), .B(\mean_pooling_0/n208 ), .X(n2584) );
  nand_x1_sg U2948 ( .A(n4999), .B(n2466), .X(n2586) );
  nand_x4_sg U2949 ( .A(n2586), .B(n4097), .X(n3482) );
  inv_x8_sg U2950 ( .A(n3482), .X(n2459) );
  inv_x2_sg U2951 ( .A(n2584), .X(n4097) );
  nor_x1_sg U2952 ( .A(n2628), .B(\mean_pooling_0/n179 ), .X(n2627) );
  inv_x1_sg U2953 ( .A(n2626), .X(n4096) );
  nor_x1_sg U2954 ( .A(n2561), .B(n2564), .X(n2626) );
  nand_x4_sg U2955 ( .A(n4096), .B(n4095), .X(n3483) );
  inv_x8_sg U2956 ( .A(n3483), .X(n2557) );
  inv_x2_sg U2957 ( .A(n2627), .X(n4095) );
  nand_x4_sg U2958 ( .A(n4083), .B(n4084), .X(n3484) );
  inv_x8_sg U2959 ( .A(n3484), .X(n2564) );
  inv_x4_sg U2960 ( .A(n1733), .X(n4435) );
  inv_x4_sg U2961 ( .A(n2046), .X(n4437) );
  inv_x4_sg U2962 ( .A(n4440), .X(n4439) );
  inv_x4_sg U2963 ( .A(n4447), .X(n4446) );
  inv_x4_sg U2964 ( .A(n4451), .X(n4450) );
  inv_x4_sg U2965 ( .A(n4444), .X(n4443) );
  inv_x2_sg U2966 ( .A(n2167), .X(n4093) );
  nor_x1_sg U2967 ( .A(n2052), .B(n4850), .X(n2167) );
  inv_x1_sg U2968 ( .A(n2630), .X(n4084) );
  inv_x1_sg U2969 ( .A(n2629), .X(n4083) );
  inv_x2_sg U2970 ( .A(n2576), .X(n4085) );
  nor_x1_sg U2971 ( .A(n2748), .B(n5018), .X(n2576) );
  inv_x2_sg U2972 ( .A(n2575), .X(n4080) );
  nor_x1_sg U2973 ( .A(n2578), .B(n2579), .X(n2575) );
  inv_x2_sg U2974 ( .A(n4802), .X(n4087) );
  inv_x1_sg U2975 ( .A(n4340), .X(n4802) );
  inv_x2_sg U2976 ( .A(n1697), .X(n4076) );
  nor_x1_sg U2977 ( .A(n2565), .B(n2566), .X(n1697) );
  inv_x2_sg U2978 ( .A(n4902), .X(n4089) );
  inv_x1_sg U2979 ( .A(n2105), .X(n4902) );
  inv_x2_sg U2980 ( .A(n2428), .X(n5021) );
  nor_x2_sg U2981 ( .A(n2441), .B(n2434), .X(n2357) );
  nand_x2_sg U2982 ( .A(n2436), .B(n4410), .X(n2441) );
  inv_x2_sg U2983 ( .A(n4281), .X(n4282) );
  inv_x1_sg U2984 ( .A(reg_input_ready), .X(n4281) );
  inv_x2_sg U2985 ( .A(n3166), .X(n4452) );
  nor_x1_sg U2986 ( .A(n3054), .B(n4447), .X(n3166) );
  inv_x4_sg U2987 ( .A(n4452), .X(n4451) );
  inv_x4_sg U2988 ( .A(n4282), .X(n4432) );
  inv_x4_sg U2989 ( .A(n4280), .X(n4428) );
  inv_x4_sg U2990 ( .A(n5021), .X(n4409) );
  inv_x4_sg U2991 ( .A(n2357), .X(n4405) );
  inv_x4_sg U2992 ( .A(n4375), .X(n4376) );
  inv_x4_sg U2993 ( .A(n4373), .X(n4374) );
  inv_x2_sg U2994 ( .A(n2047), .X(n4441) );
  inv_x1_sg U2995 ( .A(n1853), .X(n3504) );
  inv_x2_sg U2996 ( .A(n3504), .X(n3505) );
  inv_x1_sg U2997 ( .A(n2250), .X(n3506) );
  inv_x2_sg U2998 ( .A(n3506), .X(n3507) );
  inv_x1_sg U2999 ( .A(n2416), .X(n3508) );
  inv_x2_sg U3000 ( .A(n3508), .X(n3509) );
  inv_x1_sg U3001 ( .A(n2360), .X(n3510) );
  inv_x2_sg U3002 ( .A(n3510), .X(n3511) );
  inv_x1_sg U3003 ( .A(n1922), .X(n3512) );
  inv_x2_sg U3004 ( .A(n3512), .X(n3513) );
  inv_x1_sg U3005 ( .A(n1924), .X(n3514) );
  inv_x2_sg U3006 ( .A(n3514), .X(n3515) );
  inv_x1_sg U3007 ( .A(n2235), .X(n3516) );
  inv_x2_sg U3008 ( .A(n3516), .X(n3517) );
  inv_x1_sg U3009 ( .A(n2237), .X(n3518) );
  inv_x2_sg U3010 ( .A(n3518), .X(n3519) );
  inv_x1_sg U3011 ( .A(n1904), .X(n3520) );
  inv_x2_sg U3012 ( .A(n3520), .X(n3521) );
  inv_x1_sg U3013 ( .A(n1907), .X(n3522) );
  inv_x2_sg U3014 ( .A(n3522), .X(n3523) );
  inv_x1_sg U3015 ( .A(n2217), .X(n3524) );
  inv_x2_sg U3016 ( .A(n3524), .X(n3525) );
  inv_x1_sg U3017 ( .A(n2220), .X(n3526) );
  inv_x2_sg U3018 ( .A(n3526), .X(n3527) );
  inv_x1_sg U3019 ( .A(n1950), .X(n3528) );
  inv_x2_sg U3020 ( .A(n3528), .X(n3529) );
  inv_x1_sg U3021 ( .A(n1952), .X(n3530) );
  inv_x2_sg U3022 ( .A(n3530), .X(n3531) );
  inv_x1_sg U3023 ( .A(n2256), .X(n3532) );
  inv_x2_sg U3024 ( .A(n3532), .X(n3533) );
  inv_x1_sg U3025 ( .A(n2258), .X(n3534) );
  inv_x2_sg U3026 ( .A(n3534), .X(n3535) );
  inv_x1_sg U3027 ( .A(n2241), .X(n3536) );
  inv_x2_sg U3028 ( .A(n3536), .X(n3537) );
  inv_x1_sg U3029 ( .A(n2243), .X(n3538) );
  inv_x2_sg U3030 ( .A(n3538), .X(n3539) );
  inv_x1_sg U3031 ( .A(n2247), .X(n3540) );
  inv_x2_sg U3032 ( .A(n3540), .X(n3541) );
  inv_x1_sg U3033 ( .A(n2249), .X(n3542) );
  inv_x2_sg U3034 ( .A(n3542), .X(n3543) );
  inv_x1_sg U3035 ( .A(n1928), .X(n3544) );
  inv_x2_sg U3036 ( .A(n3544), .X(n3545) );
  inv_x1_sg U3037 ( .A(n1930), .X(n3546) );
  inv_x2_sg U3038 ( .A(n3546), .X(n3547) );
  inv_x1_sg U3039 ( .A(n1943), .X(n3548) );
  inv_x2_sg U3040 ( .A(n3548), .X(n3549) );
  inv_x1_sg U3041 ( .A(n1945), .X(n3550) );
  inv_x2_sg U3042 ( .A(n3550), .X(n3551) );
  inv_x1_sg U3043 ( .A(n2269), .X(n3552) );
  inv_x2_sg U3044 ( .A(n3552), .X(n3553) );
  inv_x1_sg U3045 ( .A(n2271), .X(n3554) );
  inv_x2_sg U3046 ( .A(n3554), .X(n3555) );
  inv_x1_sg U3047 ( .A(n2263), .X(n3556) );
  inv_x2_sg U3048 ( .A(n3556), .X(n3557) );
  inv_x1_sg U3049 ( .A(n2265), .X(n3558) );
  inv_x2_sg U3050 ( .A(n3558), .X(n3559) );
  inv_x1_sg U3051 ( .A(n2276), .X(n3560) );
  inv_x2_sg U3052 ( .A(n3560), .X(n3561) );
  inv_x1_sg U3053 ( .A(n2278), .X(n3562) );
  inv_x2_sg U3054 ( .A(n3562), .X(n3563) );
  inv_x1_sg U3055 ( .A(n2282), .X(n3564) );
  inv_x2_sg U3056 ( .A(n3564), .X(n3565) );
  inv_x1_sg U3057 ( .A(n2284), .X(n3566) );
  inv_x2_sg U3058 ( .A(n3566), .X(n3567) );
  inv_x1_sg U3059 ( .A(n2289), .X(n3568) );
  inv_x2_sg U3060 ( .A(n3568), .X(n3569) );
  inv_x1_sg U3061 ( .A(n2291), .X(n3570) );
  inv_x2_sg U3062 ( .A(n3570), .X(n3571) );
  inv_x1_sg U3063 ( .A(n1969), .X(n3572) );
  inv_x2_sg U3064 ( .A(n3572), .X(n3573) );
  inv_x1_sg U3065 ( .A(n1971), .X(n3574) );
  inv_x2_sg U3066 ( .A(n3574), .X(n3575) );
  inv_x1_sg U3067 ( .A(n1976), .X(n3576) );
  inv_x2_sg U3068 ( .A(n3576), .X(n3577) );
  inv_x1_sg U3069 ( .A(n1978), .X(n3578) );
  inv_x2_sg U3070 ( .A(n3578), .X(n3579) );
  inv_x1_sg U3071 ( .A(n1982), .X(n3580) );
  inv_x2_sg U3072 ( .A(n3580), .X(n3581) );
  inv_x1_sg U3073 ( .A(n1984), .X(n3582) );
  inv_x2_sg U3074 ( .A(n3582), .X(n3583) );
  inv_x1_sg U3075 ( .A(n2008), .X(n3584) );
  inv_x2_sg U3076 ( .A(n3584), .X(n3585) );
  inv_x1_sg U3077 ( .A(n2010), .X(n3586) );
  inv_x2_sg U3078 ( .A(n3586), .X(n3587) );
  inv_x1_sg U3079 ( .A(n1989), .X(n3588) );
  inv_x2_sg U3080 ( .A(n3588), .X(n3589) );
  inv_x1_sg U3081 ( .A(n1991), .X(n3590) );
  inv_x2_sg U3082 ( .A(n3590), .X(n3591) );
  inv_x1_sg U3083 ( .A(n2295), .X(n3592) );
  inv_x2_sg U3084 ( .A(n3592), .X(n3593) );
  inv_x1_sg U3085 ( .A(n2297), .X(n3594) );
  inv_x2_sg U3086 ( .A(n3594), .X(n3595) );
  inv_x1_sg U3087 ( .A(n2315), .X(n3596) );
  inv_x2_sg U3088 ( .A(n3596), .X(n3597) );
  inv_x1_sg U3089 ( .A(n2317), .X(n3598) );
  inv_x2_sg U3090 ( .A(n3598), .X(n3599) );
  inv_x1_sg U3091 ( .A(n2321), .X(n3600) );
  inv_x2_sg U3092 ( .A(n3600), .X(n3601) );
  inv_x1_sg U3093 ( .A(n2323), .X(n3602) );
  inv_x2_sg U3094 ( .A(n3602), .X(n3603) );
  inv_x1_sg U3095 ( .A(n2302), .X(n3604) );
  inv_x2_sg U3096 ( .A(n3604), .X(n3605) );
  inv_x1_sg U3097 ( .A(n2304), .X(n3606) );
  inv_x2_sg U3098 ( .A(n3606), .X(n3607) );
  inv_x1_sg U3099 ( .A(n2354), .X(n3608) );
  inv_x2_sg U3100 ( .A(n3608), .X(n3609) );
  inv_x1_sg U3101 ( .A(n2356), .X(n3610) );
  inv_x2_sg U3102 ( .A(n3610), .X(n3611) );
  inv_x1_sg U3103 ( .A(n2348), .X(n3612) );
  inv_x2_sg U3104 ( .A(n3612), .X(n3613) );
  inv_x1_sg U3105 ( .A(n2350), .X(n3614) );
  inv_x2_sg U3106 ( .A(n3614), .X(n3615) );
  inv_x1_sg U3107 ( .A(n2016), .X(n3616) );
  inv_x2_sg U3108 ( .A(n3616), .X(n3617) );
  inv_x1_sg U3109 ( .A(n2018), .X(n3618) );
  inv_x2_sg U3110 ( .A(n3618), .X(n3619) );
  inv_x1_sg U3111 ( .A(n2636), .X(n3620) );
  inv_x2_sg U3112 ( .A(n3620), .X(n3621) );
  inv_x1_sg U3113 ( .A(n2639), .X(n3622) );
  inv_x2_sg U3114 ( .A(n3622), .X(n3623) );
  inv_x1_sg U3115 ( .A(n2638), .X(n3624) );
  inv_x2_sg U3116 ( .A(n3624), .X(n3625) );
  inv_x1_sg U3117 ( .A(n2329), .X(n3626) );
  inv_x2_sg U3118 ( .A(n3626), .X(n3627) );
  inv_x1_sg U3119 ( .A(n2331), .X(n3628) );
  inv_x2_sg U3120 ( .A(n3628), .X(n3629) );
  inv_x1_sg U3121 ( .A(n2649), .X(n3630) );
  inv_x2_sg U3122 ( .A(n3630), .X(n3631) );
  inv_x1_sg U3123 ( .A(n2651), .X(n3632) );
  inv_x2_sg U3124 ( .A(n3632), .X(n3633) );
  inv_x1_sg U3125 ( .A(n2643), .X(n3634) );
  inv_x2_sg U3126 ( .A(n3634), .X(n3635) );
  inv_x1_sg U3127 ( .A(n2645), .X(n3636) );
  inv_x2_sg U3128 ( .A(n3636), .X(n3637) );
  inv_x1_sg U3129 ( .A(n2754), .X(n3638) );
  inv_x2_sg U3130 ( .A(n3638), .X(n3639) );
  inv_x1_sg U3131 ( .A(n2756), .X(n3640) );
  inv_x2_sg U3132 ( .A(n3640), .X(n3641) );
  inv_x1_sg U3133 ( .A(n2745), .X(n3642) );
  inv_x2_sg U3134 ( .A(n3642), .X(n3643) );
  inv_x1_sg U3135 ( .A(n2747), .X(n3644) );
  inv_x2_sg U3136 ( .A(n3644), .X(n3645) );
  inv_x1_sg U3137 ( .A(n2733), .X(n3646) );
  inv_x2_sg U3138 ( .A(n3646), .X(n3647) );
  inv_x1_sg U3139 ( .A(n2735), .X(n3648) );
  inv_x2_sg U3140 ( .A(n3648), .X(n3649) );
  inv_x1_sg U3141 ( .A(n2727), .X(n3650) );
  inv_x2_sg U3142 ( .A(n3650), .X(n3651) );
  inv_x1_sg U3143 ( .A(n2729), .X(n3652) );
  inv_x2_sg U3144 ( .A(n3652), .X(n3653) );
  inv_x1_sg U3145 ( .A(n2715), .X(n3654) );
  inv_x2_sg U3146 ( .A(n3654), .X(n3655) );
  inv_x1_sg U3147 ( .A(n2717), .X(n3656) );
  inv_x2_sg U3148 ( .A(n3656), .X(n3657) );
  inv_x1_sg U3149 ( .A(n2709), .X(n3658) );
  inv_x2_sg U3150 ( .A(n3658), .X(n3659) );
  inv_x1_sg U3151 ( .A(n2711), .X(n3660) );
  inv_x2_sg U3152 ( .A(n3660), .X(n3661) );
  inv_x1_sg U3153 ( .A(n2697), .X(n3662) );
  inv_x2_sg U3154 ( .A(n3662), .X(n3663) );
  inv_x1_sg U3155 ( .A(n2699), .X(n3664) );
  inv_x2_sg U3156 ( .A(n3664), .X(n3665) );
  inv_x1_sg U3157 ( .A(n2691), .X(n3666) );
  inv_x2_sg U3158 ( .A(n3666), .X(n3667) );
  inv_x1_sg U3159 ( .A(n2693), .X(n3668) );
  inv_x2_sg U3160 ( .A(n3668), .X(n3669) );
  inv_x1_sg U3161 ( .A(n2679), .X(n3670) );
  inv_x2_sg U3162 ( .A(n3670), .X(n3671) );
  inv_x1_sg U3163 ( .A(n2681), .X(n3672) );
  inv_x2_sg U3164 ( .A(n3672), .X(n3673) );
  inv_x1_sg U3165 ( .A(n2673), .X(n3674) );
  inv_x2_sg U3166 ( .A(n3674), .X(n3675) );
  inv_x1_sg U3167 ( .A(n2675), .X(n3676) );
  inv_x2_sg U3168 ( .A(n3676), .X(n3677) );
  inv_x1_sg U3169 ( .A(n2667), .X(n3678) );
  inv_x2_sg U3170 ( .A(n3678), .X(n3679) );
  inv_x1_sg U3171 ( .A(n2669), .X(n3680) );
  inv_x2_sg U3172 ( .A(n3680), .X(n3681) );
  inv_x1_sg U3173 ( .A(n2661), .X(n3682) );
  inv_x2_sg U3174 ( .A(n3682), .X(n3683) );
  inv_x1_sg U3175 ( .A(n2663), .X(n3684) );
  inv_x2_sg U3176 ( .A(n3684), .X(n3685) );
  inv_x1_sg U3177 ( .A(n2655), .X(n3686) );
  inv_x2_sg U3178 ( .A(n3686), .X(n3687) );
  inv_x1_sg U3179 ( .A(n2657), .X(n3688) );
  inv_x2_sg U3180 ( .A(n3688), .X(n3689) );
  inv_x1_sg U3181 ( .A(n1956), .X(n3690) );
  inv_x2_sg U3182 ( .A(n3690), .X(n3691) );
  inv_x1_sg U3183 ( .A(n1958), .X(n3692) );
  inv_x2_sg U3184 ( .A(n3692), .X(n3693) );
  inv_x1_sg U3185 ( .A(n1934), .X(n3694) );
  inv_x2_sg U3186 ( .A(n3694), .X(n3695) );
  inv_x1_sg U3187 ( .A(n1936), .X(n3696) );
  inv_x2_sg U3188 ( .A(n3696), .X(n3697) );
  inv_x1_sg U3189 ( .A(n2739), .X(n3698) );
  inv_x2_sg U3190 ( .A(n3698), .X(n3699) );
  inv_x1_sg U3191 ( .A(n2741), .X(n3700) );
  inv_x2_sg U3192 ( .A(n3700), .X(n3701) );
  inv_x1_sg U3193 ( .A(n2721), .X(n3702) );
  inv_x2_sg U3194 ( .A(n3702), .X(n3703) );
  inv_x1_sg U3195 ( .A(n2723), .X(n3704) );
  inv_x2_sg U3196 ( .A(n3704), .X(n3705) );
  inv_x1_sg U3197 ( .A(n2703), .X(n3706) );
  inv_x2_sg U3198 ( .A(n3706), .X(n3707) );
  inv_x1_sg U3199 ( .A(n2705), .X(n3708) );
  inv_x2_sg U3200 ( .A(n3708), .X(n3709) );
  inv_x1_sg U3201 ( .A(n2685), .X(n3710) );
  inv_x2_sg U3202 ( .A(n3710), .X(n3711) );
  inv_x1_sg U3203 ( .A(n2687), .X(n3712) );
  inv_x2_sg U3204 ( .A(n3712), .X(n3713) );
  inv_x1_sg U3205 ( .A(n2340), .X(n3714) );
  inv_x2_sg U3206 ( .A(n3714), .X(n3715) );
  inv_x1_sg U3207 ( .A(n2342), .X(n3716) );
  inv_x2_sg U3208 ( .A(n3716), .X(n3717) );
  inv_x1_sg U3209 ( .A(n2027), .X(n3718) );
  inv_x2_sg U3210 ( .A(n3718), .X(n3719) );
  inv_x1_sg U3211 ( .A(n2029), .X(n3720) );
  inv_x2_sg U3212 ( .A(n3720), .X(n3721) );
  inv_x1_sg U3213 ( .A(n2041), .X(n3722) );
  inv_x2_sg U3214 ( .A(n3722), .X(n3723) );
  inv_x1_sg U3215 ( .A(n2043), .X(n3724) );
  inv_x2_sg U3216 ( .A(n3724), .X(n3725) );
  inv_x1_sg U3217 ( .A(n2035), .X(n3726) );
  inv_x2_sg U3218 ( .A(n3726), .X(n3727) );
  inv_x1_sg U3219 ( .A(n2037), .X(n3728) );
  inv_x2_sg U3220 ( .A(n3728), .X(n3729) );
  inv_x1_sg U3221 ( .A(n1995), .X(n3730) );
  inv_x2_sg U3222 ( .A(n3730), .X(n3731) );
  inv_x1_sg U3223 ( .A(n1997), .X(n3732) );
  inv_x2_sg U3224 ( .A(n3732), .X(n3733) );
  inv_x1_sg U3225 ( .A(n2002), .X(n3734) );
  inv_x2_sg U3226 ( .A(n3734), .X(n3735) );
  inv_x1_sg U3227 ( .A(n2004), .X(n3736) );
  inv_x2_sg U3228 ( .A(n3736), .X(n3737) );
  inv_x1_sg U3229 ( .A(n1963), .X(n3738) );
  inv_x2_sg U3230 ( .A(n3738), .X(n3739) );
  inv_x1_sg U3231 ( .A(n1965), .X(n3740) );
  inv_x2_sg U3232 ( .A(n3740), .X(n3741) );
  inv_x1_sg U3233 ( .A(n1916), .X(n3742) );
  inv_x2_sg U3234 ( .A(n3742), .X(n3743) );
  inv_x1_sg U3235 ( .A(n1918), .X(n3744) );
  inv_x2_sg U3236 ( .A(n3744), .X(n3745) );
  inv_x1_sg U3237 ( .A(n2308), .X(n3746) );
  inv_x2_sg U3238 ( .A(n3746), .X(n3747) );
  inv_x1_sg U3239 ( .A(n2310), .X(n3748) );
  inv_x2_sg U3240 ( .A(n3748), .X(n3749) );
  inv_x1_sg U3241 ( .A(n2229), .X(n3750) );
  inv_x2_sg U3242 ( .A(n3750), .X(n3751) );
  inv_x1_sg U3243 ( .A(n2231), .X(n3752) );
  inv_x2_sg U3244 ( .A(n3752), .X(n3753) );
  inv_x1_sg U3245 ( .A(n2159), .X(n3754) );
  inv_x2_sg U3246 ( .A(n3754), .X(n3755) );
  inv_x1_sg U3247 ( .A(n2746), .X(n3756) );
  inv_x2_sg U3248 ( .A(n3756), .X(n3757) );
  inv_x1_sg U3249 ( .A(n2716), .X(n3758) );
  inv_x2_sg U3250 ( .A(n3758), .X(n3759) );
  inv_x1_sg U3251 ( .A(n2710), .X(n3760) );
  inv_x2_sg U3252 ( .A(n3760), .X(n3761) );
  inv_x1_sg U3253 ( .A(n2698), .X(n3762) );
  inv_x2_sg U3254 ( .A(n3762), .X(n3763) );
  inv_x1_sg U3255 ( .A(n2692), .X(n3764) );
  inv_x2_sg U3256 ( .A(n3764), .X(n3765) );
  inv_x1_sg U3257 ( .A(n2680), .X(n3766) );
  inv_x2_sg U3258 ( .A(n3766), .X(n3767) );
  inv_x1_sg U3259 ( .A(n2674), .X(n3768) );
  inv_x2_sg U3260 ( .A(n3768), .X(n3769) );
  inv_x1_sg U3261 ( .A(n2668), .X(n3770) );
  inv_x2_sg U3262 ( .A(n3770), .X(n3771) );
  inv_x1_sg U3263 ( .A(n2662), .X(n3772) );
  inv_x2_sg U3264 ( .A(n3772), .X(n3773) );
  inv_x1_sg U3265 ( .A(n2656), .X(n3774) );
  inv_x2_sg U3266 ( .A(n3774), .X(n3775) );
  inv_x1_sg U3267 ( .A(n2740), .X(n3776) );
  inv_x2_sg U3268 ( .A(n3776), .X(n3777) );
  inv_x1_sg U3269 ( .A(n2722), .X(n3778) );
  inv_x2_sg U3270 ( .A(n3778), .X(n3779) );
  inv_x1_sg U3271 ( .A(n2704), .X(n3780) );
  inv_x2_sg U3272 ( .A(n3780), .X(n3781) );
  inv_x1_sg U3273 ( .A(n2686), .X(n3782) );
  inv_x2_sg U3274 ( .A(n3782), .X(n3783) );
  inv_x1_sg U3275 ( .A(n1929), .X(n3784) );
  inv_x2_sg U3276 ( .A(n3784), .X(n3785) );
  inv_x1_sg U3277 ( .A(n2330), .X(n3786) );
  inv_x2_sg U3278 ( .A(n3786), .X(n3787) );
  inv_x1_sg U3279 ( .A(n2728), .X(n3788) );
  inv_x2_sg U3280 ( .A(n3788), .X(n3789) );
  inv_x1_sg U3281 ( .A(n2028), .X(n3790) );
  inv_x2_sg U3282 ( .A(n3790), .X(n3791) );
  inv_x1_sg U3283 ( .A(n2042), .X(n3792) );
  inv_x2_sg U3284 ( .A(n3792), .X(n3793) );
  inv_x1_sg U3285 ( .A(n2036), .X(n3794) );
  inv_x2_sg U3286 ( .A(n3794), .X(n3795) );
  inv_x1_sg U3287 ( .A(n1996), .X(n3796) );
  inv_x2_sg U3288 ( .A(n3796), .X(n3797) );
  inv_x1_sg U3289 ( .A(n2003), .X(n3798) );
  inv_x2_sg U3290 ( .A(n3798), .X(n3799) );
  inv_x1_sg U3291 ( .A(n1964), .X(n3800) );
  inv_x2_sg U3292 ( .A(n3800), .X(n3801) );
  inv_x1_sg U3293 ( .A(n1917), .X(n3802) );
  inv_x2_sg U3294 ( .A(n3802), .X(n3803) );
  inv_x1_sg U3295 ( .A(n2309), .X(n3804) );
  inv_x2_sg U3296 ( .A(n3804), .X(n3805) );
  inv_x1_sg U3297 ( .A(n2213), .X(n3806) );
  inv_x2_sg U3298 ( .A(n3806), .X(n3807) );
  inv_x1_sg U3299 ( .A(n1845), .X(n3808) );
  inv_x2_sg U3300 ( .A(n3808), .X(n3809) );
  inv_x1_sg U3301 ( .A(n2644), .X(n3810) );
  inv_x2_sg U3302 ( .A(n3810), .X(n3811) );
  inv_x1_sg U3303 ( .A(n2236), .X(n3812) );
  inv_x2_sg U3304 ( .A(n3812), .X(n3813) );
  inv_x1_sg U3305 ( .A(n1906), .X(n3814) );
  inv_x2_sg U3306 ( .A(n3814), .X(n3815) );
  inv_x1_sg U3307 ( .A(n2219), .X(n3816) );
  inv_x2_sg U3308 ( .A(n3816), .X(n3817) );
  inv_x1_sg U3309 ( .A(n1951), .X(n3818) );
  inv_x2_sg U3310 ( .A(n3818), .X(n3819) );
  inv_x1_sg U3311 ( .A(n2257), .X(n3820) );
  inv_x2_sg U3312 ( .A(n3820), .X(n3821) );
  inv_x1_sg U3313 ( .A(n1944), .X(n3822) );
  inv_x2_sg U3314 ( .A(n3822), .X(n3823) );
  inv_x1_sg U3315 ( .A(n1970), .X(n3824) );
  inv_x2_sg U3316 ( .A(n3824), .X(n3825) );
  inv_x1_sg U3317 ( .A(n2303), .X(n3826) );
  inv_x2_sg U3318 ( .A(n3826), .X(n3827) );
  inv_x1_sg U3319 ( .A(n2650), .X(n3828) );
  inv_x2_sg U3320 ( .A(n3828), .X(n3829) );
  inv_x1_sg U3321 ( .A(n2248), .X(n3830) );
  inv_x2_sg U3322 ( .A(n3830), .X(n3831) );
  inv_x1_sg U3323 ( .A(n2264), .X(n3832) );
  inv_x2_sg U3324 ( .A(n3832), .X(n3833) );
  inv_x1_sg U3325 ( .A(n2290), .X(n3834) );
  inv_x2_sg U3326 ( .A(n3834), .X(n3835) );
  inv_x1_sg U3327 ( .A(n1977), .X(n3836) );
  inv_x2_sg U3328 ( .A(n3836), .X(n3837) );
  inv_x1_sg U3329 ( .A(n1983), .X(n3838) );
  inv_x2_sg U3330 ( .A(n3838), .X(n3839) );
  inv_x1_sg U3331 ( .A(n2009), .X(n3840) );
  inv_x2_sg U3332 ( .A(n3840), .X(n3841) );
  inv_x1_sg U3333 ( .A(n1990), .X(n3842) );
  inv_x2_sg U3334 ( .A(n3842), .X(n3843) );
  inv_x1_sg U3335 ( .A(n2296), .X(n3844) );
  inv_x2_sg U3336 ( .A(n3844), .X(n3845) );
  inv_x1_sg U3337 ( .A(n2322), .X(n3846) );
  inv_x2_sg U3338 ( .A(n3846), .X(n3847) );
  inv_x1_sg U3339 ( .A(n2017), .X(n3848) );
  inv_x2_sg U3340 ( .A(n3848), .X(n3849) );
  inv_x1_sg U3341 ( .A(n2230), .X(n3850) );
  inv_x2_sg U3342 ( .A(n3850), .X(n3851) );
  inv_x1_sg U3343 ( .A(n2755), .X(n3852) );
  inv_x2_sg U3344 ( .A(n3852), .X(n3853) );
  inv_x1_sg U3345 ( .A(n1923), .X(n3854) );
  inv_x2_sg U3346 ( .A(n3854), .X(n3855) );
  inv_x1_sg U3347 ( .A(n2242), .X(n3856) );
  inv_x2_sg U3348 ( .A(n3856), .X(n3857) );
  inv_x1_sg U3349 ( .A(n2270), .X(n3858) );
  inv_x2_sg U3350 ( .A(n3858), .X(n3859) );
  inv_x1_sg U3351 ( .A(n2277), .X(n3860) );
  inv_x2_sg U3352 ( .A(n3860), .X(n3861) );
  inv_x1_sg U3353 ( .A(n2283), .X(n3862) );
  inv_x2_sg U3354 ( .A(n3862), .X(n3863) );
  inv_x1_sg U3355 ( .A(n2316), .X(n3864) );
  inv_x2_sg U3356 ( .A(n3864), .X(n3865) );
  inv_x1_sg U3357 ( .A(n2355), .X(n3866) );
  inv_x2_sg U3358 ( .A(n3866), .X(n3867) );
  inv_x1_sg U3359 ( .A(n2349), .X(n3868) );
  inv_x2_sg U3360 ( .A(n3868), .X(n3869) );
  inv_x1_sg U3361 ( .A(n2734), .X(n3870) );
  inv_x2_sg U3362 ( .A(n3870), .X(n3871) );
  inv_x1_sg U3363 ( .A(n1957), .X(n3872) );
  inv_x2_sg U3364 ( .A(n3872), .X(n3873) );
  inv_x1_sg U3365 ( .A(n1935), .X(n3874) );
  inv_x2_sg U3366 ( .A(n3874), .X(n3875) );
  inv_x1_sg U3367 ( .A(n2341), .X(n3876) );
  inv_x2_sg U3368 ( .A(n3876), .X(n3877) );
  inv_x1_sg U3369 ( .A(n4937), .X(n3878) );
  inv_x2_sg U3370 ( .A(n3878), .X(n3879) );
  inv_x1_sg U3371 ( .A(n2736), .X(n3880) );
  inv_x2_sg U3372 ( .A(n3880), .X(n3881) );
  inv_x1_sg U3373 ( .A(n2718), .X(n3882) );
  inv_x2_sg U3374 ( .A(n3882), .X(n3883) );
  inv_x1_sg U3375 ( .A(n2700), .X(n3884) );
  inv_x2_sg U3376 ( .A(n3884), .X(n3885) );
  inv_x1_sg U3377 ( .A(n2682), .X(n3886) );
  inv_x2_sg U3378 ( .A(n3886), .X(n3887) );
  inv_x1_sg U3379 ( .A(n2742), .X(n3888) );
  inv_x2_sg U3380 ( .A(n3888), .X(n3889) );
  inv_x1_sg U3381 ( .A(n2724), .X(n3890) );
  inv_x2_sg U3382 ( .A(n3890), .X(n3891) );
  inv_x1_sg U3383 ( .A(n2712), .X(n3892) );
  inv_x2_sg U3384 ( .A(n3892), .X(n3893) );
  inv_x1_sg U3385 ( .A(n2706), .X(n3894) );
  inv_x2_sg U3386 ( .A(n3894), .X(n3895) );
  inv_x1_sg U3387 ( .A(n2694), .X(n3896) );
  inv_x2_sg U3388 ( .A(n3896), .X(n3897) );
  inv_x1_sg U3389 ( .A(n2688), .X(n3898) );
  inv_x2_sg U3390 ( .A(n3898), .X(n3899) );
  inv_x1_sg U3391 ( .A(n2676), .X(n3900) );
  inv_x2_sg U3392 ( .A(n3900), .X(n3901) );
  inv_x1_sg U3393 ( .A(n2670), .X(n3902) );
  inv_x2_sg U3394 ( .A(n3902), .X(n3903) );
  inv_x1_sg U3395 ( .A(n2664), .X(n3904) );
  inv_x2_sg U3396 ( .A(n3904), .X(n3905) );
  inv_x1_sg U3397 ( .A(n2658), .X(n3906) );
  inv_x2_sg U3398 ( .A(n3906), .X(n3907) );
  inv_x1_sg U3399 ( .A(n2652), .X(n3908) );
  inv_x2_sg U3400 ( .A(n3908), .X(n3909) );
  inv_x1_sg U3401 ( .A(n2640), .X(n3910) );
  inv_x2_sg U3402 ( .A(n3910), .X(n3911) );
  inv_x1_sg U3403 ( .A(n2024), .X(n3912) );
  inv_x2_sg U3404 ( .A(n3912), .X(n3913) );
  inv_x1_sg U3405 ( .A(n2038), .X(n3914) );
  inv_x2_sg U3406 ( .A(n3914), .X(n3915) );
  inv_x1_sg U3407 ( .A(n2032), .X(n3916) );
  inv_x2_sg U3408 ( .A(n3916), .X(n3917) );
  inv_x1_sg U3409 ( .A(n1992), .X(n3918) );
  inv_x2_sg U3410 ( .A(n3918), .X(n3919) );
  inv_x1_sg U3411 ( .A(n1999), .X(n3920) );
  inv_x2_sg U3412 ( .A(n3920), .X(n3921) );
  inv_x1_sg U3413 ( .A(n1960), .X(n3922) );
  inv_x2_sg U3414 ( .A(n3922), .X(n3923) );
  inv_x1_sg U3415 ( .A(n1925), .X(n3924) );
  inv_x2_sg U3416 ( .A(n3924), .X(n3925) );
  inv_x1_sg U3417 ( .A(n1913), .X(n3926) );
  inv_x2_sg U3418 ( .A(n3926), .X(n3927) );
  inv_x1_sg U3419 ( .A(n2326), .X(n3928) );
  inv_x2_sg U3420 ( .A(n3928), .X(n3929) );
  inv_x1_sg U3421 ( .A(n2305), .X(n3930) );
  inv_x2_sg U3422 ( .A(n3930), .X(n3931) );
  inv_x1_sg U3423 ( .A(n2737), .X(n3932) );
  inv_x2_sg U3424 ( .A(n3932), .X(n3933) );
  inv_x1_sg U3425 ( .A(n2719), .X(n3934) );
  inv_x2_sg U3426 ( .A(n3934), .X(n3935) );
  inv_x1_sg U3427 ( .A(n2701), .X(n3936) );
  inv_x2_sg U3428 ( .A(n3936), .X(n3937) );
  inv_x1_sg U3429 ( .A(n2683), .X(n3938) );
  inv_x2_sg U3430 ( .A(n3938), .X(n3939) );
  inv_x1_sg U3431 ( .A(n2725), .X(n3940) );
  inv_x2_sg U3432 ( .A(n3940), .X(n3941) );
  inv_x1_sg U3433 ( .A(n1993), .X(n3942) );
  inv_x2_sg U3434 ( .A(n3942), .X(n3943) );
  inv_x1_sg U3435 ( .A(n2000), .X(n3944) );
  inv_x2_sg U3436 ( .A(n3944), .X(n3945) );
  inv_x1_sg U3437 ( .A(n1961), .X(n3946) );
  inv_x2_sg U3438 ( .A(n3946), .X(n3947) );
  inv_x1_sg U3439 ( .A(n2743), .X(n3948) );
  inv_x2_sg U3440 ( .A(n3948), .X(n3949) );
  inv_x1_sg U3441 ( .A(n2713), .X(n3950) );
  inv_x2_sg U3442 ( .A(n3950), .X(n3951) );
  inv_x1_sg U3443 ( .A(n2707), .X(n3952) );
  inv_x2_sg U3444 ( .A(n3952), .X(n3953) );
  inv_x1_sg U3445 ( .A(n2695), .X(n3954) );
  inv_x2_sg U3446 ( .A(n3954), .X(n3955) );
  inv_x1_sg U3447 ( .A(n2689), .X(n3956) );
  inv_x2_sg U3448 ( .A(n3956), .X(n3957) );
  inv_x1_sg U3449 ( .A(n2677), .X(n3958) );
  inv_x2_sg U3450 ( .A(n3958), .X(n3959) );
  inv_x1_sg U3451 ( .A(n2671), .X(n3960) );
  inv_x2_sg U3452 ( .A(n3960), .X(n3961) );
  inv_x1_sg U3453 ( .A(n2665), .X(n3962) );
  inv_x2_sg U3454 ( .A(n3962), .X(n3963) );
  inv_x1_sg U3455 ( .A(n2659), .X(n3964) );
  inv_x2_sg U3456 ( .A(n3964), .X(n3965) );
  inv_x1_sg U3457 ( .A(n2653), .X(n3966) );
  inv_x2_sg U3458 ( .A(n3966), .X(n3967) );
  inv_x1_sg U3459 ( .A(n1926), .X(n3968) );
  inv_x2_sg U3460 ( .A(n3968), .X(n3969) );
  inv_x1_sg U3461 ( .A(n2327), .X(n3970) );
  inv_x2_sg U3462 ( .A(n3970), .X(n3971) );
  inv_x1_sg U3463 ( .A(n2025), .X(n3972) );
  inv_x2_sg U3464 ( .A(n3972), .X(n3973) );
  inv_x1_sg U3465 ( .A(n2039), .X(n3974) );
  inv_x2_sg U3466 ( .A(n3974), .X(n3975) );
  inv_x1_sg U3467 ( .A(n2033), .X(n3976) );
  inv_x2_sg U3468 ( .A(n3976), .X(n3977) );
  inv_x1_sg U3469 ( .A(n1914), .X(n3978) );
  inv_x2_sg U3470 ( .A(n3978), .X(n3979) );
  inv_x1_sg U3471 ( .A(n2306), .X(n3980) );
  inv_x2_sg U3472 ( .A(n3980), .X(n3981) );
  inv_x1_sg U3473 ( .A(n2641), .X(n3982) );
  inv_x2_sg U3474 ( .A(n3982), .X(n3983) );
  inv_x1_sg U3475 ( .A(\min_pooling_0/N3 ), .X(n3984) );
  inv_x2_sg U3476 ( .A(n3984), .X(n3985) );
  inv_x1_sg U3477 ( .A(\min_pooling_0/N4 ), .X(n3986) );
  inv_x2_sg U3478 ( .A(n3986), .X(n3987) );
  inv_x1_sg U3479 ( .A(\min_pooling_0/n872 ), .X(n3988) );
  inv_x2_sg U3480 ( .A(n3988), .X(n3989) );
  inv_x1_sg U3481 ( .A(\min_pooling_0/n871 ), .X(n3990) );
  inv_x2_sg U3482 ( .A(n3990), .X(n3991) );
  inv_x1_sg U3483 ( .A(\min_pooling_0/n870 ), .X(n3992) );
  inv_x2_sg U3484 ( .A(n3992), .X(n3993) );
  inv_x1_sg U3485 ( .A(\min_pooling_0/n869 ), .X(n3994) );
  inv_x2_sg U3486 ( .A(n3994), .X(n3995) );
  inv_x1_sg U3487 ( .A(\min_pooling_0/n868 ), .X(n3996) );
  inv_x2_sg U3488 ( .A(n3996), .X(n3997) );
  inv_x1_sg U3489 ( .A(\min_pooling_0/n867 ), .X(n3998) );
  inv_x2_sg U3490 ( .A(n3998), .X(n3999) );
  inv_x1_sg U3491 ( .A(\min_pooling_0/n866 ), .X(n4000) );
  inv_x2_sg U3492 ( .A(n4000), .X(n4001) );
  inv_x1_sg U3493 ( .A(\min_pooling_0/n865 ), .X(n4002) );
  inv_x2_sg U3494 ( .A(n4002), .X(n4003) );
  inv_x1_sg U3495 ( .A(\min_pooling_0/n864 ), .X(n4004) );
  inv_x2_sg U3496 ( .A(n4004), .X(n4005) );
  inv_x1_sg U3497 ( .A(\min_pooling_0/n863 ), .X(n4006) );
  inv_x2_sg U3498 ( .A(n4006), .X(n4007) );
  inv_x1_sg U3499 ( .A(\min_pooling_0/n862 ), .X(n4008) );
  inv_x2_sg U3500 ( .A(n4008), .X(n4009) );
  inv_x1_sg U3501 ( .A(\min_pooling_0/n861 ), .X(n4010) );
  inv_x2_sg U3502 ( .A(n4010), .X(n4011) );
  inv_x1_sg U3503 ( .A(\min_pooling_0/n860 ), .X(n4012) );
  inv_x2_sg U3504 ( .A(n4012), .X(n4013) );
  inv_x1_sg U3505 ( .A(\min_pooling_0/n859 ), .X(n4014) );
  inv_x2_sg U3506 ( .A(n4014), .X(n4015) );
  inv_x1_sg U3507 ( .A(\min_pooling_0/n858 ), .X(n4016) );
  inv_x2_sg U3508 ( .A(n4016), .X(n4017) );
  inv_x1_sg U3509 ( .A(\min_pooling_0/n857 ), .X(n4018) );
  inv_x2_sg U3510 ( .A(n4018), .X(n4019) );
  inv_x1_sg U3511 ( .A(\min_pooling_0/n856 ), .X(n4020) );
  inv_x2_sg U3512 ( .A(n4020), .X(n4021) );
  inv_x1_sg U3513 ( .A(\min_pooling_0/n855 ), .X(n4022) );
  inv_x2_sg U3514 ( .A(n4022), .X(n4023) );
  inv_x1_sg U3515 ( .A(\min_pooling_0/n854 ), .X(n4024) );
  inv_x2_sg U3516 ( .A(n4024), .X(n4025) );
  inv_x1_sg U3517 ( .A(\mean_pooling_0/N4 ), .X(n4026) );
  inv_x2_sg U3518 ( .A(n4026), .X(n4027) );
  inv_x1_sg U3519 ( .A(\mean_pooling_0/N5 ), .X(n4028) );
  inv_x2_sg U3520 ( .A(n4028), .X(n4029) );
  inv_x1_sg U3521 ( .A(\max_pooling_0/N3 ), .X(n4030) );
  inv_x2_sg U3522 ( .A(n4030), .X(n4031) );
  inv_x1_sg U3523 ( .A(\max_pooling_0/N4 ), .X(n4032) );
  inv_x2_sg U3524 ( .A(n4032), .X(n4033) );
  inv_x1_sg U3525 ( .A(\max_pooling_0/n820 ), .X(n4034) );
  inv_x2_sg U3526 ( .A(n4034), .X(n4035) );
  inv_x1_sg U3527 ( .A(\max_pooling_0/n819 ), .X(n4036) );
  inv_x2_sg U3528 ( .A(n4036), .X(n4037) );
  inv_x1_sg U3529 ( .A(\max_pooling_0/n818 ), .X(n4038) );
  inv_x2_sg U3530 ( .A(n4038), .X(n4039) );
  inv_x1_sg U3531 ( .A(\max_pooling_0/n817 ), .X(n4040) );
  inv_x2_sg U3532 ( .A(n4040), .X(n4041) );
  inv_x1_sg U3533 ( .A(\max_pooling_0/n816 ), .X(n4042) );
  inv_x2_sg U3534 ( .A(n4042), .X(n4043) );
  inv_x1_sg U3535 ( .A(\max_pooling_0/n815 ), .X(n4044) );
  inv_x2_sg U3536 ( .A(n4044), .X(n4045) );
  inv_x1_sg U3537 ( .A(\max_pooling_0/n814 ), .X(n4046) );
  inv_x2_sg U3538 ( .A(n4046), .X(n4047) );
  inv_x1_sg U3539 ( .A(\max_pooling_0/n813 ), .X(n4048) );
  inv_x2_sg U3540 ( .A(n4048), .X(n4049) );
  inv_x1_sg U3541 ( .A(\max_pooling_0/n812 ), .X(n4050) );
  inv_x2_sg U3542 ( .A(n4050), .X(n4051) );
  inv_x1_sg U3543 ( .A(\max_pooling_0/n811 ), .X(n4052) );
  inv_x2_sg U3544 ( .A(n4052), .X(n4053) );
  inv_x1_sg U3545 ( .A(\max_pooling_0/n810 ), .X(n4054) );
  inv_x2_sg U3546 ( .A(n4054), .X(n4055) );
  inv_x1_sg U3547 ( .A(\max_pooling_0/n809 ), .X(n4056) );
  inv_x2_sg U3548 ( .A(n4056), .X(n4057) );
  inv_x1_sg U3549 ( .A(\max_pooling_0/n808 ), .X(n4058) );
  inv_x2_sg U3550 ( .A(n4058), .X(n4059) );
  inv_x1_sg U3551 ( .A(\max_pooling_0/n807 ), .X(n4060) );
  inv_x2_sg U3552 ( .A(n4060), .X(n4061) );
  inv_x1_sg U3553 ( .A(\max_pooling_0/n806 ), .X(n4062) );
  inv_x2_sg U3554 ( .A(n4062), .X(n4063) );
  inv_x1_sg U3555 ( .A(\max_pooling_0/n805 ), .X(n4064) );
  inv_x2_sg U3556 ( .A(n4064), .X(n4065) );
  inv_x1_sg U3557 ( .A(\max_pooling_0/n804 ), .X(n4066) );
  inv_x2_sg U3558 ( .A(n4066), .X(n4067) );
  inv_x1_sg U3559 ( .A(\max_pooling_0/n803 ), .X(n4068) );
  inv_x2_sg U3560 ( .A(n4068), .X(n4069) );
  inv_x1_sg U3561 ( .A(\max_pooling_0/n802 ), .X(n4070) );
  inv_x2_sg U3562 ( .A(n4070), .X(n4071) );
  inv_x1_sg U3563 ( .A(n5054), .X(n4072) );
  inv_x2_sg U3564 ( .A(n4072), .X(n4073) );
  inv_x1_sg U3565 ( .A(n5053), .X(n4074) );
  inv_x2_sg U3566 ( .A(n4074), .X(n4075) );
  nor_x2_sg U3567 ( .A(n5030), .B(n4426), .X(n3409) );
  nor_x2_sg U3568 ( .A(n5038), .B(n3334), .X(n3377) );
  nor_x2_sg U3569 ( .A(n4370), .B(n4078), .X(n2170) );
  nor_x2_sg U3570 ( .A(n5041), .B(n3334), .X(n3365) );
  nor_x2_sg U3571 ( .A(n5045), .B(n4426), .X(n3349) );
  inv_x4_sg U3572 ( .A(n4076), .X(n4077) );
  inv_x4_sg U3573 ( .A(n2052), .X(n4078) );
  inv_x4_sg U3574 ( .A(n4378), .X(n4805) );
  nor_x2_sg U3575 ( .A(n4904), .B(n4079), .X(n2628) );
  nor_x2_sg U3576 ( .A(n5042), .B(n4426), .X(n3361) );
  nor_x2_sg U3577 ( .A(n5040), .B(n4427), .X(n3369) );
  nor_x2_sg U3578 ( .A(n4416), .B(n5045), .X(n2660) );
  nor_x2_sg U3579 ( .A(n4417), .B(n5043), .X(n2672) );
  nor_x2_sg U3580 ( .A(n5041), .B(n1905), .X(n1962) );
  nor_x2_sg U3581 ( .A(n2637), .B(n5038), .X(n2702) );
  nor_x2_sg U3582 ( .A(n1909), .B(n1910), .X(n1899) );
  nor_x2_sg U3583 ( .A(n4088), .B(n1911), .X(n1909) );
  nor_x2_sg U3584 ( .A(n2222), .B(n2223), .X(n2212) );
  nor_x2_sg U3585 ( .A(n4090), .B(n4366), .X(n2223) );
  inv_x4_sg U3586 ( .A(n2561), .X(n4079) );
  inv_x4_sg U3587 ( .A(n4080), .X(n4081) );
  inv_x1_sg U3588 ( .A(n1868), .X(n4091) );
  nor_x1_sg U3589 ( .A(n2298), .B(n4094), .X(n4082) );
  nor_x1_sg U3590 ( .A(n2298), .B(n4094), .X(n2162) );
  nor_x4_sg U3591 ( .A(n2093), .B(n4849), .X(n2298) );
  nor_x2_sg U3592 ( .A(n3501), .B(n2564), .X(n2563) );
  nor_x2_sg U3593 ( .A(n5047), .B(n3334), .X(n3341) );
  nor_x2_sg U3594 ( .A(n5043), .B(n4427), .X(n3357) );
  nor_x2_sg U3595 ( .A(n4416), .B(n5042), .X(n2678) );
  nor_x2_sg U3596 ( .A(n4417), .B(n5040), .X(n2690) );
  nor_x2_sg U3597 ( .A(n1732), .B(n4810), .X(n1856) );
  nor_x2_sg U3598 ( .A(n5030), .B(n4411), .X(n2328) );
  nor_x2_sg U3599 ( .A(n1891), .B(n1892), .X(n1890) );
  nor_x2_sg U3600 ( .A(n1750), .B(n4804), .X(n1891) );
  nor_x2_sg U3601 ( .A(n2637), .B(n5041), .X(n2684) );
  nor_x2_sg U3602 ( .A(n4396), .B(n4917), .X(n1937) );
  inv_x4_sg U3603 ( .A(n1742), .X(n4917) );
  inv_x4_sg U3604 ( .A(n4085), .X(n4086) );
  inv_x4_sg U3605 ( .A(n4087), .X(n4088) );
  inv_x4_sg U3606 ( .A(n4089), .X(n4090) );
  nor_x2_sg U3607 ( .A(n4904), .B(\mean_pooling_0/n179 ), .X(n2562) );
  inv_x2_sg U3608 ( .A(n4091), .X(n4092) );
  nor_x2_sg U3609 ( .A(n4899), .B(n4903), .X(n2565) );
  nor_x2_sg U3610 ( .A(n4898), .B(n4903), .X(n2631) );
  inv_x4_sg U3611 ( .A(n2568), .X(n4903) );
  inv_x4_sg U3612 ( .A(n4093), .X(n4094) );
  nor_x4_sg U3613 ( .A(n4278), .B(n4923), .X(n1885) );
  inv_x8_sg U3614 ( .A(n1805), .X(n4923) );
  nor_x4_sg U3615 ( .A(n4398), .B(n4936), .X(n1938) );
  inv_x8_sg U3616 ( .A(n1802), .X(n4936) );
  inv_x4_sg U3617 ( .A(n2564), .X(n4904) );
  nand_x1_sg U3618 ( .A(n1897), .B(n1898), .X(n1893) );
  nor_x1_sg U3619 ( .A(n1899), .B(n1900), .X(n1897) );
  nand_x1_sg U3620 ( .A(n2209), .B(n2210), .X(n2208) );
  inv_x1_sg U3621 ( .A(n1880), .X(n4937) );
  inv_x2_sg U3622 ( .A(n2198), .X(n4105) );
  nand_x1_sg U3623 ( .A(n4924), .B(n4360), .X(n2198) );
  nand_x1_sg U3624 ( .A(n2211), .B(n2210), .X(n2207) );
  nand_x1_sg U3625 ( .A(n1882), .B(n1883), .X(n1881) );
  nand_x1_sg U3626 ( .A(n1888), .B(n1889), .X(n1887) );
  nand_x1_sg U3627 ( .A(n4939), .B(n2194), .X(n2193) );
  inv_x1_sg U3628 ( .A(n2199), .X(n4939) );
  nand_x1_sg U3629 ( .A(n2195), .B(n2196), .X(n2194) );
  nand_x1_sg U3630 ( .A(n2202), .B(n2203), .X(n2201) );
  nand_x1_sg U3631 ( .A(n1872), .B(n1873), .X(n1871) );
  nand_x1_sg U3632 ( .A(n1793), .B(n4373), .X(n1873) );
  nand_x1_sg U3633 ( .A(n2186), .B(n2187), .X(n2185) );
  nand_x1_sg U3634 ( .A(n1860), .B(n1861), .X(n1859) );
  inv_x1_sg U3635 ( .A(n1848), .X(n4990) );
  nand_x1_sg U3636 ( .A(n2174), .B(n2175), .X(n2173) );
  inv_x1_sg U3637 ( .A(n1840), .X(n5009) );
  nand_x1_sg U3638 ( .A(n1775), .B(n4814), .X(n1842) );
  inv_x1_sg U3639 ( .A(n2154), .X(n5011) );
  nand_x1_sg U3640 ( .A(n1843), .B(n1844), .X(n1841) );
  nand_x1_sg U3641 ( .A(n2157), .B(n2158), .X(n2155) );
  inv_x1_sg U3642 ( .A(n2470), .X(n4992) );
  inv_x1_sg U3643 ( .A(n2595), .X(n4980) );
  nand_x1_sg U3644 ( .A(n2594), .B(n3489), .X(n2593) );
  inv_x1_sg U3645 ( .A(n2604), .X(n4960) );
  nand_x1_sg U3646 ( .A(n2603), .B(n3491), .X(n2602) );
  inv_x1_sg U3647 ( .A(n2613), .X(n4941) );
  nand_x1_sg U3648 ( .A(n2612), .B(n3493), .X(n2611) );
  inv_x1_sg U3649 ( .A(n2583), .X(n5005) );
  nand_x1_sg U3650 ( .A(\mean_pooling_0/n175 ), .B(n2582), .X(n2581) );
  nor_x1_sg U3651 ( .A(n3777), .B(n3701), .X(n2736) );
  inv_x1_sg U3652 ( .A(n2458), .X(n5000) );
  nand_x1_sg U3653 ( .A(n4987), .B(n2470), .X(n2589) );
  inv_x1_sg U3654 ( .A(n2592), .X(n4986) );
  nand_x1_sg U3655 ( .A(\mean_pooling_0/n172 ), .B(n2591), .X(n2590) );
  nor_x1_sg U3656 ( .A(n3779), .B(n3705), .X(n2718) );
  nand_x1_sg U3657 ( .A(\mean_pooling_0/n172 ), .B(n2480), .X(n2479) );
  inv_x1_sg U3658 ( .A(n2598), .X(n4973) );
  nand_x1_sg U3659 ( .A(n2597), .B(n3490), .X(n2596) );
  inv_x1_sg U3660 ( .A(n2601), .X(n4967) );
  nand_x1_sg U3661 ( .A(\mean_pooling_0/n169 ), .B(n2600), .X(n2599) );
  nor_x1_sg U3662 ( .A(n3781), .B(n3709), .X(n2700) );
  nand_x1_sg U3663 ( .A(\mean_pooling_0/n169 ), .B(n2501), .X(n2500) );
  inv_x1_sg U3664 ( .A(n2607), .X(n4954) );
  nand_x1_sg U3665 ( .A(n2606), .B(n3492), .X(n2605) );
  inv_x1_sg U3666 ( .A(n2610), .X(n4947) );
  nand_x1_sg U3667 ( .A(\mean_pooling_0/n166 ), .B(n2609), .X(n2608) );
  nor_x1_sg U3668 ( .A(n3783), .B(n3713), .X(n2682) );
  nand_x1_sg U3669 ( .A(\mean_pooling_0/n166 ), .B(n2522), .X(n2521) );
  inv_x1_sg U3670 ( .A(n2616), .X(n4933) );
  nand_x1_sg U3671 ( .A(n2615), .B(n3494), .X(n2614) );
  inv_x1_sg U3672 ( .A(n2619), .X(n4927) );
  nand_x1_sg U3673 ( .A(n2618), .B(n3488), .X(n2617) );
  inv_x1_sg U3674 ( .A(n2622), .X(n4920) );
  nand_x1_sg U3675 ( .A(n2621), .B(n3498), .X(n2620) );
  inv_x1_sg U3676 ( .A(n2625), .X(n4914) );
  nor_x1_sg U3677 ( .A(n2146), .B(n3434), .X(n2047) );
  nand_x1_sg U3678 ( .A(\mean_pooling_0/n2 ), .B(n2750), .X(n2749) );
  nand_x1_sg U3679 ( .A(\mean_pooling_0/n189 ), .B(n2452), .X(n2451) );
  nor_x1_sg U3680 ( .A(n3757), .B(n3645), .X(n2742) );
  nand_x1_sg U3681 ( .A(n2454), .B(n2455), .X(n2456) );
  nand_x1_sg U3682 ( .A(\mean_pooling_0/n208 ), .B(n2466), .X(n2465) );
  nand_x1_sg U3683 ( .A(\mean_pooling_0/n190 ), .B(n2473), .X(n2472) );
  nor_x1_sg U3684 ( .A(n3789), .B(n3653), .X(n2724) );
  nand_x1_sg U3685 ( .A(n2475), .B(n2476), .X(n2477) );
  nand_x1_sg U3686 ( .A(\mean_pooling_0/n209 ), .B(n2487), .X(n2486) );
  nor_x1_sg U3687 ( .A(n3759), .B(n3657), .X(n2712) );
  nand_x1_sg U3688 ( .A(\mean_pooling_0/n191 ), .B(n2494), .X(n2493) );
  nor_x1_sg U3689 ( .A(n3761), .B(n3661), .X(n2706) );
  nand_x1_sg U3690 ( .A(n2496), .B(n2497), .X(n2498) );
  nand_x1_sg U3691 ( .A(\mean_pooling_0/n210 ), .B(n2508), .X(n2507) );
  nor_x1_sg U3692 ( .A(n3763), .B(n3665), .X(n2694) );
  nand_x1_sg U3693 ( .A(\mean_pooling_0/n192 ), .B(n2515), .X(n2514) );
  nor_x1_sg U3694 ( .A(n3765), .B(n3669), .X(n2688) );
  nand_x1_sg U3695 ( .A(n2517), .B(n2518), .X(n2519) );
  nand_x1_sg U3696 ( .A(\mean_pooling_0/n211 ), .B(n2529), .X(n2528) );
  nor_x1_sg U3697 ( .A(n3767), .B(n3673), .X(n2676) );
  nand_x1_sg U3698 ( .A(\mean_pooling_0/n193 ), .B(n2536), .X(n2535) );
  nor_x1_sg U3699 ( .A(n3769), .B(n3677), .X(n2670) );
  nand_x1_sg U3700 ( .A(\mean_pooling_0/n178 ), .B(n2543), .X(n2542) );
  nor_x1_sg U3701 ( .A(n3771), .B(n3681), .X(n2664) );
  nand_x1_sg U3702 ( .A(\mean_pooling_0/n212 ), .B(n2550), .X(n2549) );
  nor_x1_sg U3703 ( .A(n3773), .B(n3685), .X(n2658) );
  inv_x1_sg U3704 ( .A(n2556), .X(n4909) );
  nor_x1_sg U3705 ( .A(n3775), .B(n3689), .X(n2652) );
  nor_x1_sg U3706 ( .A(n3811), .B(n3637), .X(n2640) );
  inv_x2_sg U3707 ( .A(n3118), .X(n4279) );
  nor_x1_sg U3708 ( .A(n3153), .B(n5028), .X(n3118) );
  nor_x1_sg U3709 ( .A(n3791), .B(n3721), .X(n2024) );
  nor_x1_sg U3710 ( .A(n3793), .B(n3725), .X(n2038) );
  nor_x1_sg U3711 ( .A(n3795), .B(n3729), .X(n2032) );
  nor_x1_sg U3712 ( .A(n3797), .B(n3733), .X(n1992) );
  nor_x1_sg U3713 ( .A(n3799), .B(n3737), .X(n1999) );
  nor_x1_sg U3714 ( .A(n3801), .B(n3741), .X(n1960) );
  nor_x1_sg U3715 ( .A(n3785), .B(n3547), .X(n1925) );
  nor_x1_sg U3716 ( .A(n3803), .B(n3745), .X(n1913) );
  inv_x1_sg U3717 ( .A(n2577), .X(n5019) );
  inv_x1_sg U3718 ( .A(n2447), .X(n5012) );
  nand_x1_sg U3719 ( .A(n2448), .B(n2449), .X(n2446) );
  inv_x2_sg U3720 ( .A(n1721), .X(n4119) );
  nor_x1_sg U3721 ( .A(n5004), .B(n2453), .X(n1721) );
  nand_x1_sg U3722 ( .A(n4995), .B(n2463), .X(n2460) );
  inv_x1_sg U3723 ( .A(n2468), .X(n4993) );
  nand_x1_sg U3724 ( .A(n2469), .B(n2470), .X(n2467) );
  inv_x2_sg U3725 ( .A(n1719), .X(n4117) );
  nor_x1_sg U3726 ( .A(n4985), .B(n2474), .X(n1719) );
  inv_x1_sg U3727 ( .A(n2482), .X(n4979) );
  nand_x1_sg U3728 ( .A(n2483), .B(n2484), .X(n2481) );
  inv_x1_sg U3729 ( .A(n2489), .X(n4972) );
  nand_x1_sg U3730 ( .A(n2490), .B(n2491), .X(n2488) );
  inv_x2_sg U3731 ( .A(n1713), .X(n4107) );
  nor_x1_sg U3732 ( .A(n4966), .B(n2495), .X(n1713) );
  inv_x1_sg U3733 ( .A(n2503), .X(n4959) );
  nand_x1_sg U3734 ( .A(n2504), .B(n2505), .X(n2502) );
  inv_x1_sg U3735 ( .A(n2510), .X(n4953) );
  nand_x1_sg U3736 ( .A(n2511), .B(n2512), .X(n2509) );
  inv_x2_sg U3737 ( .A(n1715), .X(n4115) );
  nor_x1_sg U3738 ( .A(n4946), .B(n2516), .X(n1715) );
  inv_x1_sg U3739 ( .A(n2524), .X(n4940) );
  nand_x1_sg U3740 ( .A(n2525), .B(n2526), .X(n2523) );
  inv_x1_sg U3741 ( .A(n2531), .X(n4932) );
  nand_x1_sg U3742 ( .A(n2532), .B(n2533), .X(n2530) );
  inv_x1_sg U3743 ( .A(n2538), .X(n4926) );
  nand_x1_sg U3744 ( .A(n2539), .B(n2540), .X(n2537) );
  inv_x1_sg U3745 ( .A(n2545), .X(n4919) );
  nand_x1_sg U3746 ( .A(n2546), .B(n2547), .X(n2544) );
  inv_x1_sg U3747 ( .A(n2552), .X(n4913) );
  nand_x1_sg U3748 ( .A(n2553), .B(n2554), .X(n2551) );
  nand_x1_sg U3749 ( .A(n4905), .B(n2561), .X(n2558) );
  inv_x1_sg U3750 ( .A(n2560), .X(n4905) );
  nor_x1_sg U3751 ( .A(n3787), .B(n3629), .X(n2326) );
  nor_x1_sg U3752 ( .A(n3805), .B(n3749), .X(n2305) );
  inv_x2_sg U3753 ( .A(n2087), .X(n4964) );
  nand_x1_sg U3754 ( .A(n1773), .B(n1774), .X(n1648) );
  nand_x1_sg U3755 ( .A(n4442), .B(n1775), .X(n1774) );
  nand_x1_sg U3756 ( .A(n1756), .B(n1757), .X(n1655) );
  nand_x1_sg U3757 ( .A(n1827), .B(n1828), .X(n1627) );
  nand_x1_sg U3758 ( .A(n4442), .B(n1826), .X(n1828) );
  nand_x1_sg U3759 ( .A(n1824), .B(n1825), .X(n1628) );
  nand_x1_sg U3760 ( .A(n4442), .B(n5008), .X(n1825) );
  inv_x1_sg U3761 ( .A(n1826), .X(n5008) );
  nand_x1_sg U3762 ( .A(n1743), .B(n1744), .X(n1660) );
  nand_x1_sg U3763 ( .A(n4444), .B(n1745), .X(n1744) );
  nand_x1_sg U3764 ( .A(n1829), .B(n1830), .X(n1626) );
  nand_x1_sg U3765 ( .A(n4442), .B(n5002), .X(n1830) );
  inv_x1_sg U3766 ( .A(n1745), .X(n5002) );
  nand_x1_sg U3767 ( .A(n1822), .B(n1823), .X(n1629) );
  nand_x1_sg U3768 ( .A(n4442), .B(n1821), .X(n1823) );
  nand_x1_sg U3769 ( .A(n1819), .B(n1820), .X(n1630) );
  nand_x1_sg U3770 ( .A(n4442), .B(n4997), .X(n1820) );
  inv_x1_sg U3771 ( .A(n1821), .X(n4997) );
  nand_x1_sg U3772 ( .A(n1736), .B(n1737), .X(n1663) );
  nand_x1_sg U3773 ( .A(n4442), .B(n1732), .X(n1737) );
  nand_x1_sg U3774 ( .A(n1730), .B(n1731), .X(n1665) );
  nand_x1_sg U3775 ( .A(n4442), .B(n4989), .X(n1731) );
  inv_x1_sg U3776 ( .A(n1732), .X(n4989) );
  nand_x1_sg U3777 ( .A(n1778), .B(n1779), .X(n1646) );
  nand_x1_sg U3778 ( .A(n4442), .B(n1780), .X(n1779) );
  nand_x1_sg U3779 ( .A(n1776), .B(n1777), .X(n1647) );
  nand_x1_sg U3780 ( .A(n1787), .B(n1788), .X(n1643) );
  nand_x1_sg U3781 ( .A(n4442), .B(n1786), .X(n1788) );
  nand_x1_sg U3782 ( .A(n1784), .B(n1785), .X(n1644) );
  nand_x1_sg U3783 ( .A(n4442), .B(n4976), .X(n1785) );
  inv_x1_sg U3784 ( .A(n1786), .X(n4976) );
  nand_x1_sg U3785 ( .A(n1762), .B(n1763), .X(n1652) );
  nand_x1_sg U3786 ( .A(n4442), .B(n1764), .X(n1763) );
  nand_x1_sg U3787 ( .A(n1760), .B(n1761), .X(n1653) );
  nand_x1_sg U3788 ( .A(n1770), .B(n1771), .X(n1649) );
  nand_x1_sg U3789 ( .A(n4442), .B(n1772), .X(n1771) );
  nand_x1_sg U3790 ( .A(n1768), .B(n1769), .X(n1650) );
  nand_x1_sg U3791 ( .A(n4442), .B(n4963), .X(n1769) );
  nand_x1_sg U3792 ( .A(n1808), .B(n1809), .X(n1634) );
  nand_x1_sg U3793 ( .A(n4442), .B(n1810), .X(n1809) );
  nand_x1_sg U3794 ( .A(n1806), .B(n1807), .X(n1635) );
  nand_x1_sg U3795 ( .A(n1816), .B(n1817), .X(n1631) );
  nand_x1_sg U3796 ( .A(n1814), .B(n1815), .X(n1632) );
  nand_x1_sg U3797 ( .A(n1794), .B(n1795), .X(n1640) );
  nand_x1_sg U3798 ( .A(n4442), .B(n1793), .X(n1795) );
  nand_x1_sg U3799 ( .A(n1791), .B(n1792), .X(n1641) );
  nand_x1_sg U3800 ( .A(n4442), .B(n4944), .X(n1792) );
  inv_x1_sg U3801 ( .A(n1793), .X(n4944) );
  nand_x1_sg U3802 ( .A(n1800), .B(n1801), .X(n1637) );
  nand_x1_sg U3803 ( .A(n4442), .B(n1802), .X(n1801) );
  nand_x1_sg U3804 ( .A(n1798), .B(n1799), .X(n1638) );
  nand_x1_sg U3805 ( .A(n4434), .B(n4397), .X(n1798) );
  nand_x1_sg U3806 ( .A(n1811), .B(n1812), .X(n1633) );
  nand_x1_sg U3807 ( .A(n1734), .B(n1735), .X(n1664) );
  nand_x1_sg U3808 ( .A(n4434), .B(n4399), .X(n1734) );
  nand_x1_sg U3809 ( .A(n1803), .B(n1804), .X(n1636) );
  nand_x1_sg U3810 ( .A(n4442), .B(n1805), .X(n1804) );
  nand_x1_sg U3811 ( .A(n1796), .B(n1797), .X(n1639) );
  nand_x1_sg U3812 ( .A(n4434), .B(n4277), .X(n1796) );
  nand_x1_sg U3813 ( .A(n1740), .B(n1741), .X(n1661) );
  nand_x1_sg U3814 ( .A(n4442), .B(n1742), .X(n1741) );
  nand_x1_sg U3815 ( .A(n1738), .B(n1739), .X(n1662) );
  nand_x1_sg U3816 ( .A(n4434), .B(n4395), .X(n1738) );
  nand_x1_sg U3817 ( .A(n1748), .B(n1749), .X(n1658) );
  nand_x1_sg U3818 ( .A(n4442), .B(n1750), .X(n1749) );
  nand_x1_sg U3819 ( .A(n1746), .B(n1747), .X(n1659) );
  nand_x1_sg U3820 ( .A(n1753), .B(n1754), .X(n1656) );
  nand_x1_sg U3821 ( .A(n1751), .B(n1752), .X(n1657) );
  nand_x1_sg U3822 ( .A(n4434), .B(n4393), .X(n1751) );
  nand_x1_sg U3823 ( .A(n1789), .B(n1790), .X(n1642) );
  nand_x1_sg U3824 ( .A(n4442), .B(n1783), .X(n1790) );
  nand_x1_sg U3825 ( .A(n1781), .B(n1782), .X(n1645) );
  nand_x1_sg U3826 ( .A(n4442), .B(n4901), .X(n1782) );
  inv_x1_sg U3827 ( .A(n1783), .X(n4901) );
  nand_x1_sg U3828 ( .A(n1765), .B(n1766), .X(n1651) );
  nand_x1_sg U3829 ( .A(n4442), .B(n1767), .X(n1766) );
  nand_x1_sg U3830 ( .A(n1758), .B(n1759), .X(n1654) );
  nand_x1_sg U3831 ( .A(n4420), .B(n1716), .X(n1672) );
  nand_x1_sg U3832 ( .A(n1717), .B(n3485), .X(n1716) );
  nand_x1_sg U3833 ( .A(n4420), .B(n1694), .X(n1683) );
  nand_x1_sg U3834 ( .A(n1695), .B(n3485), .X(n1694) );
  nand_x1_sg U3835 ( .A(n4420), .B(n1720), .X(n1670) );
  nand_x1_sg U3836 ( .A(n3154), .B(n1726), .X(n1667) );
  nand_x1_sg U3837 ( .A(n1727), .B(n3485), .X(n1726) );
  nand_x1_sg U3838 ( .A(n3154), .B(n1690), .X(n1685) );
  nand_x1_sg U3839 ( .A(n1691), .B(n3485), .X(n1690) );
  nand_x1_sg U3840 ( .A(n3154), .B(n1718), .X(n1671) );
  nand_x1_sg U3841 ( .A(n4420), .B(n1698), .X(n1681) );
  nand_x1_sg U3842 ( .A(n1699), .B(n3485), .X(n1698) );
  nand_x1_sg U3843 ( .A(n4420), .B(n1724), .X(n1668) );
  nand_x1_sg U3844 ( .A(n1725), .B(n3485), .X(n1724) );
  nand_x1_sg U3845 ( .A(n4420), .B(n1712), .X(n1674) );
  nand_x1_sg U3846 ( .A(n4420), .B(n1710), .X(n1675) );
  nand_x1_sg U3847 ( .A(n1711), .B(n3485), .X(n1710) );
  nand_x1_sg U3848 ( .A(n4420), .B(n1702), .X(n1679) );
  nand_x1_sg U3849 ( .A(n1703), .B(n3485), .X(n1702) );
  nand_x1_sg U3850 ( .A(n3154), .B(n1714), .X(n1673) );
  nand_x1_sg U3851 ( .A(n4420), .B(n1728), .X(n1666) );
  nand_x1_sg U3852 ( .A(n1729), .B(n3485), .X(n1728) );
  nand_x1_sg U3853 ( .A(n4420), .B(n1700), .X(n1680) );
  nand_x1_sg U3854 ( .A(n1701), .B(n3485), .X(n1700) );
  nand_x1_sg U3855 ( .A(n4420), .B(n1706), .X(n1677) );
  nand_x1_sg U3856 ( .A(n1707), .B(n3485), .X(n1706) );
  nand_x1_sg U3857 ( .A(n3154), .B(n1692), .X(n1684) );
  nand_x1_sg U3858 ( .A(n1693), .B(n3485), .X(n1692) );
  nand_x1_sg U3859 ( .A(n3154), .B(n1722), .X(n1669) );
  nand_x1_sg U3860 ( .A(n1723), .B(n3485), .X(n1722) );
  nand_x1_sg U3861 ( .A(n4420), .B(n1704), .X(n1678) );
  nand_x1_sg U3862 ( .A(n1705), .B(n3485), .X(n1704) );
  nand_x1_sg U3863 ( .A(n4420), .B(n1696), .X(n1682) );
  nand_x1_sg U3864 ( .A(n4420), .B(n1708), .X(n1676) );
  nand_x1_sg U3865 ( .A(n2088), .B(n2089), .X(n1608) );
  nand_x1_sg U3866 ( .A(n4436), .B(n2090), .X(n2089) );
  nand_x1_sg U3867 ( .A(n2071), .B(n2072), .X(n1615) );
  nand_x1_sg U3868 ( .A(n4436), .B(n5016), .X(n2072) );
  nand_x1_sg U3869 ( .A(n2141), .B(n2142), .X(n1587) );
  nand_x1_sg U3870 ( .A(n2046), .B(n2143), .X(n2142) );
  nand_x1_sg U3871 ( .A(n2139), .B(n2140), .X(n1588) );
  nand_x1_sg U3872 ( .A(n4440), .B(n4391), .X(n2139) );
  nand_x1_sg U3873 ( .A(n2058), .B(n2059), .X(n1620) );
  nand_x1_sg U3874 ( .A(n4436), .B(n2060), .X(n2059) );
  nand_x1_sg U3875 ( .A(n2144), .B(n2145), .X(n1586) );
  nand_x1_sg U3876 ( .A(n2136), .B(n2137), .X(n1589) );
  nand_x1_sg U3877 ( .A(n4436), .B(n2138), .X(n2137) );
  nand_x1_sg U3878 ( .A(n2134), .B(n2135), .X(n1590) );
  nand_x1_sg U3879 ( .A(n2050), .B(n2051), .X(n1623) );
  nand_x1_sg U3880 ( .A(n4436), .B(n2052), .X(n2051) );
  nand_x1_sg U3881 ( .A(n2044), .B(n2045), .X(n1625) );
  nand_x1_sg U3882 ( .A(n2094), .B(n2095), .X(n1606) );
  nand_x1_sg U3883 ( .A(n4436), .B(n2093), .X(n2095) );
  nand_x1_sg U3884 ( .A(n2091), .B(n2092), .X(n1607) );
  nand_x1_sg U3885 ( .A(n4436), .B(n4984), .X(n2092) );
  inv_x1_sg U3886 ( .A(n2093), .X(n4984) );
  nand_x1_sg U3887 ( .A(n2100), .B(n2101), .X(n1603) );
  nand_x1_sg U3888 ( .A(n4436), .B(n2102), .X(n2101) );
  nand_x1_sg U3889 ( .A(n2098), .B(n2099), .X(n1604) );
  nand_x1_sg U3890 ( .A(n2078), .B(n2079), .X(n1612) );
  nand_x1_sg U3891 ( .A(n4436), .B(n2080), .X(n2079) );
  nand_x1_sg U3892 ( .A(n2076), .B(n2077), .X(n1613) );
  nand_x1_sg U3893 ( .A(n4436), .B(n4971), .X(n2077) );
  nand_x1_sg U3894 ( .A(n2085), .B(n2086), .X(n1609) );
  nand_x1_sg U3895 ( .A(n4436), .B(n2087), .X(n2086) );
  nand_x1_sg U3896 ( .A(n2083), .B(n2084), .X(n1610) );
  nand_x1_sg U3897 ( .A(n4436), .B(n4964), .X(n2084) );
  nand_x1_sg U3898 ( .A(n2123), .B(n2124), .X(n1594) );
  nand_x1_sg U3899 ( .A(n4436), .B(n2125), .X(n2124) );
  nand_x1_sg U3900 ( .A(n2121), .B(n2122), .X(n1595) );
  nand_x1_sg U3901 ( .A(n4436), .B(n4958), .X(n2122) );
  nand_x1_sg U3902 ( .A(n2131), .B(n2132), .X(n1591) );
  nand_x1_sg U3903 ( .A(n4436), .B(n2133), .X(n2132) );
  nand_x1_sg U3904 ( .A(n2129), .B(n2130), .X(n1592) );
  nand_x1_sg U3905 ( .A(n2108), .B(n2109), .X(n1600) );
  nand_x1_sg U3906 ( .A(n4436), .B(n2110), .X(n2109) );
  nand_x1_sg U3907 ( .A(n2106), .B(n2107), .X(n1601) );
  nand_x1_sg U3908 ( .A(n2115), .B(n2116), .X(n1597) );
  nand_x1_sg U3909 ( .A(n4436), .B(n2117), .X(n2116) );
  nand_x1_sg U3910 ( .A(n2113), .B(n2114), .X(n1598) );
  nand_x1_sg U3911 ( .A(n4436), .B(n4938), .X(n2114) );
  nand_x1_sg U3912 ( .A(n2126), .B(n2127), .X(n1593) );
  nand_x1_sg U3913 ( .A(n4436), .B(n2128), .X(n2127) );
  nand_x1_sg U3914 ( .A(n2048), .B(n2049), .X(n1624) );
  nand_x1_sg U3915 ( .A(n2118), .B(n2119), .X(n1596) );
  nand_x1_sg U3916 ( .A(n4436), .B(n2120), .X(n2119) );
  nand_x1_sg U3917 ( .A(n2111), .B(n2112), .X(n1599) );
  nand_x1_sg U3918 ( .A(n4436), .B(n4924), .X(n2112) );
  nand_x1_sg U3919 ( .A(n2055), .B(n2056), .X(n1621) );
  nand_x1_sg U3920 ( .A(n2053), .B(n2054), .X(n1622) );
  nand_x1_sg U3921 ( .A(n2063), .B(n2064), .X(n1618) );
  nand_x1_sg U3922 ( .A(n4436), .B(n2065), .X(n2064) );
  nand_x1_sg U3923 ( .A(n2061), .B(n2062), .X(n1619) );
  nand_x1_sg U3924 ( .A(n2068), .B(n2069), .X(n1616) );
  nand_x1_sg U3925 ( .A(n2066), .B(n2067), .X(n1617) );
  nand_x1_sg U3926 ( .A(n2103), .B(n2104), .X(n1602) );
  nand_x1_sg U3927 ( .A(n4436), .B(n2105), .X(n2104) );
  nand_x1_sg U3928 ( .A(n2096), .B(n2097), .X(n1605) );
  nand_x1_sg U3929 ( .A(n2081), .B(n2082), .X(n1611) );
  nand_x1_sg U3930 ( .A(n4436), .B(n2075), .X(n2082) );
  nand_x1_sg U3931 ( .A(n2073), .B(n2074), .X(n1614) );
  nand_x1_sg U3932 ( .A(n4896), .B(n4436), .X(n2074) );
  inv_x1_sg U3933 ( .A(n2075), .X(n4896) );
  nand_x1_sg U3934 ( .A(n4407), .B(done_min), .X(n2438) );
  nand_x1_sg U3935 ( .A(n3063), .B(n3064), .X(n3439) );
  nand_x1_sg U3936 ( .A(n3057), .B(n3058), .X(n3438) );
  nand_x1_sg U3937 ( .A(n3330), .B(n3331), .X(\min_pooling_0/n452 ) );
  nand_x1_sg U3938 ( .A(n3335), .B(n3336), .X(\min_pooling_0/n451 ) );
  nand_x1_sg U3939 ( .A(n3339), .B(n3340), .X(\min_pooling_0/n450 ) );
  nand_x1_sg U3940 ( .A(n3343), .B(n3344), .X(\min_pooling_0/n449 ) );
  nand_x1_sg U3941 ( .A(n3347), .B(n3348), .X(\min_pooling_0/n448 ) );
  nand_x1_sg U3942 ( .A(n3351), .B(n3352), .X(\min_pooling_0/n447 ) );
  nand_x1_sg U3943 ( .A(n3355), .B(n3356), .X(\min_pooling_0/n446 ) );
  nand_x1_sg U3944 ( .A(n3359), .B(n3360), .X(\min_pooling_0/n445 ) );
  nand_x1_sg U3945 ( .A(n3363), .B(n3364), .X(\min_pooling_0/n444 ) );
  nand_x1_sg U3946 ( .A(n3367), .B(n3368), .X(\min_pooling_0/n443 ) );
  nand_x1_sg U3947 ( .A(n3371), .B(n3372), .X(\min_pooling_0/n442 ) );
  nand_x1_sg U3948 ( .A(n3375), .B(n3376), .X(\min_pooling_0/n441 ) );
  nand_x1_sg U3949 ( .A(n3379), .B(n3380), .X(\min_pooling_0/n440 ) );
  nand_x1_sg U3950 ( .A(n3383), .B(n3384), .X(\min_pooling_0/n439 ) );
  nand_x1_sg U3951 ( .A(n3387), .B(n3388), .X(\min_pooling_0/n438 ) );
  nand_x1_sg U3952 ( .A(n3391), .B(n3392), .X(\min_pooling_0/n437 ) );
  nand_x1_sg U3953 ( .A(n3395), .B(n3396), .X(\min_pooling_0/n436 ) );
  nand_x1_sg U3954 ( .A(n3399), .B(n3400), .X(\min_pooling_0/n435 ) );
  nand_x1_sg U3955 ( .A(n3403), .B(n3404), .X(\min_pooling_0/n434 ) );
  nand_x1_sg U3956 ( .A(n3407), .B(n3408), .X(\min_pooling_0/n433 ) );
  nand_x1_sg U3957 ( .A(n3155), .B(n3156), .X(n3480) );
  nand_x1_sg U3958 ( .A(n3158), .B(n3159), .X(n3481) );
  nand_x1_sg U3959 ( .A(n3119), .B(n3120), .X(n3463) );
  nand_x1_sg U3960 ( .A(\mean_pooling_0/n179 ), .B(n3117), .X(n3120) );
  nand_x1_sg U3961 ( .A(n3147), .B(n3148), .X(n3477) );
  nand_x1_sg U3962 ( .A(\mean_pooling_0/n194 ), .B(n3117), .X(n3148) );
  nand_x1_sg U3963 ( .A(n3131), .B(n3132), .X(n3469) );
  nand_x1_sg U3964 ( .A(\mean_pooling_0/n212 ), .B(n3117), .X(n3132) );
  nand_x1_sg U3965 ( .A(n3145), .B(n3146), .X(n3476) );
  nand_x1_sg U3966 ( .A(\mean_pooling_0/n178 ), .B(n3117), .X(n3146) );
  nand_x1_sg U3967 ( .A(n3115), .B(n3116), .X(n3462) );
  nand_x1_sg U3968 ( .A(\mean_pooling_0/n193 ), .B(n3117), .X(n3116) );
  nand_x1_sg U3969 ( .A(n3135), .B(n3136), .X(n3471) );
  nand_x1_sg U3970 ( .A(\mean_pooling_0/n211 ), .B(n3117), .X(n3136) );
  nand_x1_sg U3971 ( .A(n3127), .B(n3128), .X(n3467) );
  nand_x1_sg U3972 ( .A(n3117), .B(n3497), .X(n3128) );
  nand_x1_sg U3973 ( .A(n3143), .B(n3144), .X(n3475) );
  nand_x1_sg U3974 ( .A(\mean_pooling_0/n192 ), .B(n3117), .X(n3144) );
  nand_x1_sg U3975 ( .A(n3121), .B(n3122), .X(n3464) );
  nand_x1_sg U3976 ( .A(\mean_pooling_0/n210 ), .B(n3117), .X(n3122) );
  nand_x1_sg U3977 ( .A(n3133), .B(n3134), .X(n3470) );
  nand_x1_sg U3978 ( .A(n3117), .B(n3496), .X(n3134) );
  nand_x1_sg U3979 ( .A(n3125), .B(n3126), .X(n3466) );
  nand_x1_sg U3980 ( .A(\mean_pooling_0/n191 ), .B(n3117), .X(n3126) );
  nand_x1_sg U3981 ( .A(n3141), .B(n3142), .X(n3474) );
  nand_x1_sg U3982 ( .A(\mean_pooling_0/n209 ), .B(n3117), .X(n3142) );
  nand_x1_sg U3983 ( .A(n3129), .B(n3130), .X(n3468) );
  nand_x1_sg U3984 ( .A(n3117), .B(n3495), .X(n3130) );
  nand_x1_sg U3985 ( .A(n3149), .B(n3150), .X(n3478) );
  nand_x1_sg U3986 ( .A(\mean_pooling_0/n190 ), .B(n3117), .X(n3150) );
  nand_x1_sg U3987 ( .A(n3123), .B(n3124), .X(n3465) );
  nand_x1_sg U3988 ( .A(\mean_pooling_0/n208 ), .B(n3117), .X(n3124) );
  nand_x1_sg U3989 ( .A(n3151), .B(n3152), .X(n3479) );
  nand_x1_sg U3990 ( .A(n3139), .B(n3140), .X(n3473) );
  nand_x1_sg U3991 ( .A(\mean_pooling_0/n189 ), .B(n3117), .X(n3140) );
  nand_x1_sg U3992 ( .A(n3137), .B(n3138), .X(n3472) );
  nand_x1_sg U3993 ( .A(\mean_pooling_0/n2 ), .B(n3117), .X(n3138) );
  nand_x1_sg U3994 ( .A(n3093), .B(n3094), .X(n3451) );
  nand_x1_sg U3995 ( .A(n3066), .B(n3067), .X(n3440) );
  nand_x1_sg U3996 ( .A(n3089), .B(n3090), .X(n3449) );
  nand_x1_sg U3997 ( .A(n3413), .B(n4430), .X(n3090) );
  nand_x1_sg U3998 ( .A(n3081), .B(n3082), .X(n3445) );
  nand_x1_sg U3999 ( .A(n3414), .B(n4431), .X(n3082) );
  nand_x1_sg U4000 ( .A(n3113), .B(n3114), .X(n3461) );
  nand_x1_sg U4001 ( .A(n3415), .B(n4430), .X(n3114) );
  nand_x1_sg U4002 ( .A(n3073), .B(n3074), .X(n3441) );
  nand_x1_sg U4003 ( .A(n3416), .B(n3072), .X(n3074) );
  nand_x1_sg U4004 ( .A(n3079), .B(n3080), .X(n3444) );
  nand_x1_sg U4005 ( .A(n3417), .B(n3072), .X(n3080) );
  nand_x1_sg U4006 ( .A(n3083), .B(n3084), .X(n3446) );
  nand_x1_sg U4007 ( .A(n3418), .B(n4430), .X(n3084) );
  nand_x1_sg U4008 ( .A(n3087), .B(n3088), .X(n3448) );
  nand_x1_sg U4009 ( .A(n3419), .B(n4431), .X(n3088) );
  nand_x1_sg U4010 ( .A(n3085), .B(n3086), .X(n3447) );
  nand_x1_sg U4011 ( .A(n3420), .B(n3072), .X(n3086) );
  nand_x1_sg U4012 ( .A(n3095), .B(n3096), .X(n3452) );
  nand_x1_sg U4013 ( .A(n3421), .B(n4430), .X(n3096) );
  nand_x1_sg U4014 ( .A(n3109), .B(n3110), .X(n3459) );
  nand_x1_sg U4015 ( .A(n3422), .B(n3072), .X(n3110) );
  nand_x1_sg U4016 ( .A(n3091), .B(n3092), .X(n3450) );
  nand_x1_sg U4017 ( .A(n3423), .B(n3072), .X(n3092) );
  nand_x1_sg U4018 ( .A(n3107), .B(n3108), .X(n3458) );
  nand_x1_sg U4019 ( .A(n3424), .B(n4430), .X(n3108) );
  nand_x1_sg U4020 ( .A(n3077), .B(n3078), .X(n3443) );
  nand_x1_sg U4021 ( .A(n3425), .B(n4430), .X(n3078) );
  nand_x1_sg U4022 ( .A(n3097), .B(n3098), .X(n3453) );
  nand_x1_sg U4023 ( .A(n3426), .B(n3072), .X(n3098) );
  nand_x1_sg U4024 ( .A(n3103), .B(n3104), .X(n3456) );
  nand_x1_sg U4025 ( .A(n3427), .B(n3072), .X(n3104) );
  nand_x1_sg U4026 ( .A(n3099), .B(n3100), .X(n3454) );
  nand_x1_sg U4027 ( .A(n3428), .B(n4431), .X(n3100) );
  nand_x1_sg U4028 ( .A(n3105), .B(n3106), .X(n3457) );
  nand_x1_sg U4029 ( .A(n3429), .B(n4431), .X(n3106) );
  nand_x1_sg U4030 ( .A(n3101), .B(n3102), .X(n3455) );
  nand_x1_sg U4031 ( .A(n3430), .B(n4430), .X(n3102) );
  nand_x1_sg U4032 ( .A(n3111), .B(n3112), .X(n3460) );
  nand_x1_sg U4033 ( .A(n3431), .B(n4431), .X(n3112) );
  nand_x1_sg U4034 ( .A(n3075), .B(n3076), .X(n3442) );
  nand_x1_sg U4035 ( .A(n3432), .B(n4431), .X(n3076) );
  nand_x1_sg U4036 ( .A(n3164), .B(n3165), .X(n554) );
  nand_x1_sg U4037 ( .A(\im[0][0] ), .B(n4445), .X(n3164) );
  nand_x1_sg U4038 ( .A(n3168), .B(n3169), .X(n553) );
  nand_x1_sg U4039 ( .A(\im[0][1] ), .B(n4445), .X(n3168) );
  nand_x1_sg U4040 ( .A(n3170), .B(n3171), .X(n552) );
  nand_x1_sg U4041 ( .A(\im[0][2] ), .B(n4445), .X(n3170) );
  nand_x1_sg U4042 ( .A(n3172), .B(n3173), .X(n551) );
  nand_x1_sg U4043 ( .A(\im[0][3] ), .B(n4445), .X(n3172) );
  nand_x1_sg U4044 ( .A(n3174), .B(n3175), .X(n550) );
  nand_x1_sg U4045 ( .A(\im[0][4] ), .B(n4445), .X(n3174) );
  nand_x1_sg U4046 ( .A(n3176), .B(n3177), .X(n549) );
  nand_x1_sg U4047 ( .A(\im[0][5] ), .B(n4445), .X(n3176) );
  nand_x1_sg U4048 ( .A(n3178), .B(n3179), .X(n548) );
  nand_x1_sg U4049 ( .A(\im[0][6] ), .B(n4445), .X(n3178) );
  nand_x1_sg U4050 ( .A(n3180), .B(n3181), .X(n547) );
  nand_x1_sg U4051 ( .A(\im[0][7] ), .B(n4445), .X(n3180) );
  nand_x1_sg U4052 ( .A(n3182), .B(n3183), .X(n546) );
  nand_x1_sg U4053 ( .A(\im[0][8] ), .B(n4445), .X(n3182) );
  nand_x1_sg U4054 ( .A(n3184), .B(n3185), .X(n545) );
  nand_x1_sg U4055 ( .A(\im[0][9] ), .B(n4445), .X(n3184) );
  nand_x1_sg U4056 ( .A(n3186), .B(n3187), .X(n544) );
  nand_x1_sg U4057 ( .A(\im[0][10] ), .B(n4445), .X(n3186) );
  nand_x1_sg U4058 ( .A(n3188), .B(n3189), .X(n543) );
  nand_x1_sg U4059 ( .A(\im[0][11] ), .B(n4445), .X(n3188) );
  nand_x1_sg U4060 ( .A(n3190), .B(n3191), .X(n542) );
  nand_x1_sg U4061 ( .A(\im[0][12] ), .B(n4445), .X(n3190) );
  nand_x1_sg U4062 ( .A(n3192), .B(n3193), .X(n541) );
  nand_x1_sg U4063 ( .A(\im[0][13] ), .B(n4445), .X(n3192) );
  nand_x1_sg U4064 ( .A(n3194), .B(n3195), .X(n540) );
  nand_x1_sg U4065 ( .A(\im[0][14] ), .B(n4447), .X(n3194) );
  nand_x1_sg U4066 ( .A(n3196), .B(n3197), .X(n539) );
  nand_x1_sg U4067 ( .A(\im[0][15] ), .B(n4447), .X(n3196) );
  nand_x1_sg U4068 ( .A(n3198), .B(n3199), .X(n538) );
  nand_x1_sg U4069 ( .A(\im[0][16] ), .B(n4447), .X(n3198) );
  nand_x1_sg U4070 ( .A(n3200), .B(n3201), .X(n537) );
  nand_x1_sg U4071 ( .A(\im[0][17] ), .B(n4445), .X(n3200) );
  nand_x1_sg U4072 ( .A(n3202), .B(n3203), .X(n536) );
  nand_x1_sg U4073 ( .A(\im[0][18] ), .B(n4445), .X(n3202) );
  nand_x1_sg U4074 ( .A(n3204), .B(n3205), .X(n535) );
  nand_x1_sg U4075 ( .A(\im[0][19] ), .B(n4445), .X(n3204) );
  nand_x1_sg U4076 ( .A(n3206), .B(n3207), .X(n534) );
  nand_x1_sg U4077 ( .A(\im[1][0] ), .B(n4445), .X(n3206) );
  nand_x1_sg U4078 ( .A(n3208), .B(n3209), .X(n533) );
  nand_x1_sg U4079 ( .A(\im[1][1] ), .B(n4445), .X(n3208) );
  nand_x1_sg U4080 ( .A(n3210), .B(n3211), .X(n532) );
  nand_x1_sg U4081 ( .A(\im[1][2] ), .B(n4445), .X(n3210) );
  nand_x1_sg U4082 ( .A(n3212), .B(n3213), .X(n531) );
  nand_x1_sg U4083 ( .A(\im[1][3] ), .B(n4445), .X(n3212) );
  nand_x1_sg U4084 ( .A(n3214), .B(n3215), .X(n530) );
  nand_x1_sg U4085 ( .A(\im[1][4] ), .B(n4445), .X(n3214) );
  nand_x1_sg U4086 ( .A(n3216), .B(n3217), .X(n529) );
  nand_x1_sg U4087 ( .A(\im[1][5] ), .B(n4445), .X(n3216) );
  nand_x1_sg U4088 ( .A(n3218), .B(n3219), .X(n528) );
  nand_x1_sg U4089 ( .A(\im[1][6] ), .B(n4445), .X(n3218) );
  nand_x1_sg U4090 ( .A(n3220), .B(n3221), .X(n527) );
  nand_x1_sg U4091 ( .A(\im[1][7] ), .B(n4445), .X(n3220) );
  nand_x1_sg U4092 ( .A(n3222), .B(n3223), .X(n526) );
  nand_x1_sg U4093 ( .A(\im[1][8] ), .B(n4445), .X(n3222) );
  nand_x1_sg U4094 ( .A(n3224), .B(n3225), .X(n525) );
  nand_x1_sg U4095 ( .A(\im[1][9] ), .B(n4445), .X(n3224) );
  nand_x1_sg U4096 ( .A(n3226), .B(n3227), .X(n524) );
  nand_x1_sg U4097 ( .A(\im[1][10] ), .B(n4445), .X(n3226) );
  nand_x1_sg U4098 ( .A(n3228), .B(n3229), .X(n523) );
  nand_x1_sg U4099 ( .A(\im[1][11] ), .B(n4445), .X(n3228) );
  nand_x1_sg U4100 ( .A(n3230), .B(n3231), .X(n522) );
  nand_x1_sg U4101 ( .A(\im[1][12] ), .B(n4445), .X(n3230) );
  nand_x1_sg U4102 ( .A(n3232), .B(n3233), .X(n521) );
  nand_x1_sg U4103 ( .A(\im[1][13] ), .B(n4445), .X(n3232) );
  nand_x1_sg U4104 ( .A(n3234), .B(n3235), .X(n520) );
  nand_x1_sg U4105 ( .A(\im[1][14] ), .B(n4445), .X(n3234) );
  nand_x1_sg U4106 ( .A(n3236), .B(n3237), .X(n519) );
  nand_x1_sg U4107 ( .A(\im[1][15] ), .B(n4445), .X(n3236) );
  nand_x1_sg U4108 ( .A(n3238), .B(n3239), .X(n518) );
  nand_x1_sg U4109 ( .A(\im[1][16] ), .B(n4445), .X(n3238) );
  nand_x1_sg U4110 ( .A(n3240), .B(n3241), .X(n517) );
  nand_x1_sg U4111 ( .A(\im[1][17] ), .B(n4445), .X(n3240) );
  nand_x1_sg U4112 ( .A(n3242), .B(n3243), .X(n516) );
  nand_x1_sg U4113 ( .A(\im[1][18] ), .B(n4445), .X(n3242) );
  nand_x1_sg U4114 ( .A(n3244), .B(n3245), .X(n515) );
  nand_x1_sg U4115 ( .A(\im[1][19] ), .B(n4445), .X(n3244) );
  nand_x1_sg U4116 ( .A(n3246), .B(n3247), .X(n514) );
  nand_x1_sg U4117 ( .A(\im[2][0] ), .B(n4445), .X(n3246) );
  nand_x1_sg U4118 ( .A(n3248), .B(n3249), .X(n513) );
  nand_x1_sg U4119 ( .A(\im[2][1] ), .B(n4445), .X(n3248) );
  nand_x1_sg U4120 ( .A(n3250), .B(n3251), .X(n512) );
  nand_x1_sg U4121 ( .A(\im[2][2] ), .B(n4445), .X(n3250) );
  nand_x1_sg U4122 ( .A(n3252), .B(n3253), .X(n511) );
  nand_x1_sg U4123 ( .A(\im[2][3] ), .B(n4445), .X(n3252) );
  nand_x1_sg U4124 ( .A(n3254), .B(n3255), .X(n510) );
  nand_x1_sg U4125 ( .A(\im[2][4] ), .B(n4445), .X(n3254) );
  nand_x1_sg U4126 ( .A(n3256), .B(n3257), .X(n509) );
  nand_x1_sg U4127 ( .A(\im[2][5] ), .B(n4445), .X(n3256) );
  nand_x1_sg U4128 ( .A(n3258), .B(n3259), .X(n508) );
  nand_x1_sg U4129 ( .A(\im[2][6] ), .B(n4445), .X(n3258) );
  nand_x1_sg U4130 ( .A(n3260), .B(n3261), .X(n507) );
  nand_x1_sg U4131 ( .A(\im[2][7] ), .B(n4445), .X(n3260) );
  nand_x1_sg U4132 ( .A(n3262), .B(n3263), .X(n506) );
  nand_x1_sg U4133 ( .A(\im[2][8] ), .B(n4445), .X(n3262) );
  nand_x1_sg U4134 ( .A(n3264), .B(n3265), .X(n505) );
  nand_x1_sg U4135 ( .A(\im[2][9] ), .B(n4445), .X(n3264) );
  nand_x1_sg U4136 ( .A(n3266), .B(n3267), .X(n504) );
  nand_x1_sg U4137 ( .A(\im[2][10] ), .B(n4445), .X(n3266) );
  nand_x1_sg U4138 ( .A(n3268), .B(n3269), .X(n503) );
  nand_x1_sg U4139 ( .A(\im[2][11] ), .B(n4445), .X(n3268) );
  nand_x1_sg U4140 ( .A(n3270), .B(n3271), .X(n502) );
  nand_x1_sg U4141 ( .A(\im[2][12] ), .B(n4445), .X(n3270) );
  nand_x1_sg U4142 ( .A(n3272), .B(n3273), .X(n501) );
  nand_x1_sg U4143 ( .A(\im[2][13] ), .B(n4445), .X(n3272) );
  nand_x1_sg U4144 ( .A(n3274), .B(n3275), .X(n500) );
  nand_x1_sg U4145 ( .A(\im[2][14] ), .B(n4447), .X(n3274) );
  nand_x1_sg U4146 ( .A(n3276), .B(n3277), .X(n499) );
  nand_x1_sg U4147 ( .A(\im[2][15] ), .B(n4447), .X(n3276) );
  nand_x1_sg U4148 ( .A(n3278), .B(n3279), .X(n498) );
  nand_x1_sg U4149 ( .A(\im[2][16] ), .B(n4447), .X(n3278) );
  nand_x1_sg U4150 ( .A(n3280), .B(n3281), .X(n497) );
  nand_x1_sg U4151 ( .A(\im[2][17] ), .B(n4447), .X(n3280) );
  nand_x1_sg U4152 ( .A(n3282), .B(n3283), .X(n496) );
  nand_x1_sg U4153 ( .A(\im[2][18] ), .B(n4445), .X(n3282) );
  nand_x1_sg U4154 ( .A(n3284), .B(n3285), .X(n495) );
  nand_x1_sg U4155 ( .A(\im[2][19] ), .B(n4445), .X(n3284) );
  nand_x1_sg U4156 ( .A(n3286), .B(n3287), .X(n494) );
  nand_x1_sg U4157 ( .A(\im[3][0] ), .B(n4445), .X(n3286) );
  nand_x1_sg U4158 ( .A(n3288), .B(n3289), .X(n493) );
  nand_x1_sg U4159 ( .A(\im[3][1] ), .B(n4445), .X(n3288) );
  nand_x1_sg U4160 ( .A(n3290), .B(n3291), .X(n492) );
  nand_x1_sg U4161 ( .A(\im[3][2] ), .B(n4445), .X(n3290) );
  nand_x1_sg U4162 ( .A(n3292), .B(n3293), .X(n491) );
  nand_x1_sg U4163 ( .A(\im[3][3] ), .B(n4445), .X(n3292) );
  nand_x1_sg U4164 ( .A(n3294), .B(n3295), .X(n490) );
  nand_x1_sg U4165 ( .A(\im[3][4] ), .B(n4445), .X(n3294) );
  nand_x1_sg U4166 ( .A(n3296), .B(n3297), .X(n489) );
  nand_x1_sg U4167 ( .A(\im[3][5] ), .B(n4445), .X(n3296) );
  nand_x1_sg U4168 ( .A(n3298), .B(n3299), .X(n488) );
  nand_x1_sg U4169 ( .A(\im[3][6] ), .B(n4445), .X(n3298) );
  nand_x1_sg U4170 ( .A(n3300), .B(n3301), .X(n487) );
  nand_x1_sg U4171 ( .A(\im[3][7] ), .B(n4445), .X(n3300) );
  nand_x1_sg U4172 ( .A(n3302), .B(n3303), .X(n486) );
  nand_x1_sg U4173 ( .A(\im[3][8] ), .B(n4445), .X(n3302) );
  nand_x1_sg U4174 ( .A(n3304), .B(n3305), .X(n485) );
  nand_x1_sg U4175 ( .A(\im[3][9] ), .B(n4445), .X(n3304) );
  nand_x1_sg U4176 ( .A(n3306), .B(n3307), .X(n484) );
  nand_x1_sg U4177 ( .A(\im[3][10] ), .B(n4445), .X(n3306) );
  nand_x1_sg U4178 ( .A(n3308), .B(n3309), .X(n483) );
  nand_x1_sg U4179 ( .A(\im[3][11] ), .B(n4445), .X(n3308) );
  nand_x1_sg U4180 ( .A(n3310), .B(n3311), .X(n482) );
  nand_x1_sg U4181 ( .A(\im[3][12] ), .B(n4445), .X(n3310) );
  nand_x1_sg U4182 ( .A(n3312), .B(n3313), .X(n481) );
  nand_x1_sg U4183 ( .A(\im[3][13] ), .B(n4445), .X(n3312) );
  nand_x1_sg U4184 ( .A(n3314), .B(n3315), .X(n480) );
  nand_x1_sg U4185 ( .A(\im[3][14] ), .B(n4445), .X(n3314) );
  nand_x1_sg U4186 ( .A(n3316), .B(n3317), .X(n479) );
  nand_x1_sg U4187 ( .A(\im[3][15] ), .B(n4445), .X(n3316) );
  nand_x1_sg U4188 ( .A(n3318), .B(n3319), .X(n478) );
  nand_x1_sg U4189 ( .A(\im[3][16] ), .B(n4445), .X(n3318) );
  nand_x1_sg U4190 ( .A(n3320), .B(n3321), .X(n477) );
  nand_x1_sg U4191 ( .A(\im[3][17] ), .B(n4445), .X(n3320) );
  nand_x1_sg U4192 ( .A(n3322), .B(n3323), .X(n476) );
  nand_x1_sg U4193 ( .A(\im[3][18] ), .B(n4445), .X(n3322) );
  nand_x1_sg U4194 ( .A(n3324), .B(n3325), .X(n475) );
  nand_x1_sg U4195 ( .A(\im[3][19] ), .B(n4445), .X(n3324) );
  nand_x1_sg U4196 ( .A(n3050), .B(n3051), .X(n3437) );
  nand_x1_sg U4197 ( .A(n3047), .B(n3048), .X(n3436) );
  nor_x2_sg U4198 ( .A(n4837), .B(n4410), .X(n2364) );
  nor_x2_sg U4199 ( .A(n5030), .B(n4421), .X(n2015) );
  nor_x2_sg U4200 ( .A(n5038), .B(n2218), .X(n2294) );
  nor_x2_sg U4201 ( .A(n5047), .B(n4412), .X(n2216) );
  nor_x2_sg U4202 ( .A(n5043), .B(n4422), .X(n1949) );
  nor_x2_sg U4203 ( .A(n4835), .B(n4410), .X(n2444) );
  nor_x2_sg U4204 ( .A(n4840), .B(n4410), .X(n2376) );
  nand_x1_sg U4205 ( .A(n4442), .B(n1755), .X(n1754) );
  inv_x1_sg U4206 ( .A(n3053), .X(n4098) );
  nand_x4_sg U4207 ( .A(n5025), .B(n472), .X(n3053) );
  nand_x2_sg U4208 ( .A(n2093), .B(n4849), .X(n2168) );
  nor_x2_sg U4209 ( .A(n5040), .B(n4412), .X(n2281) );
  nor_x2_sg U4210 ( .A(n5041), .B(n2218), .X(n2275) );
  nor_x2_sg U4211 ( .A(n5047), .B(n4422), .X(n1903) );
  nor_x2_sg U4212 ( .A(n5045), .B(n1905), .X(n1942) );
  nor_x2_sg U4213 ( .A(n5042), .B(n4421), .X(n1955) );
  nor_x2_sg U4214 ( .A(n4839), .B(n4410), .X(n2372) );
  nor_x2_sg U4215 ( .A(n4846), .B(n4410), .X(n2400) );
  nand_x4_sg U4216 ( .A(n2433), .B(n5025), .X(n1686) );
  nand_x1_sg U4217 ( .A(n4442), .B(n1813), .X(n1812) );
  nand_x1_sg U4218 ( .A(n4436), .B(n2057), .X(n2056) );
  nand_x1_sg U4219 ( .A(n4442), .B(n1818), .X(n1817) );
  nand_x1_sg U4220 ( .A(n4436), .B(n2070), .X(n2069) );
  nor_x2_sg U4221 ( .A(n4852), .B(n4410), .X(n2424) );
  inv_x4_sg U4222 ( .A(n4274), .X(n4852) );
  nor_x2_sg U4223 ( .A(n4853), .B(n2090), .X(n2325) );
  nor_x4_sg U4224 ( .A(n1832), .B(n3433), .X(n1733) );
  inv_x4_sg U4225 ( .A(n3054), .X(n5022) );
  inv_x4_sg U4226 ( .A(n4033), .X(n4099) );
  inv_x8_sg U4227 ( .A(n4099), .X(n4100) );
  nand_x4_sg U4228 ( .A(n4100), .B(n4110), .X(n2221) );
  inv_x4_sg U4229 ( .A(n3987), .X(n4101) );
  inv_x8_sg U4230 ( .A(n4101), .X(n4102) );
  nand_x4_sg U4231 ( .A(n4102), .B(n4112), .X(n1908) );
  inv_x4_sg U4232 ( .A(n4029), .X(n4103) );
  inv_x8_sg U4233 ( .A(n4103), .X(n4104) );
  nand_x4_sg U4234 ( .A(n4104), .B(n4114), .X(n2573) );
  nand_x2_sg U4235 ( .A(input_ready), .B(n5026), .X(n3412) );
  nor_x2_sg U4236 ( .A(n4416), .B(n5030), .X(n2753) );
  nor_x2_sg U4237 ( .A(n2637), .B(n5047), .X(n2648) );
  nor_x2_sg U4238 ( .A(n5038), .B(n4421), .X(n1975) );
  nor_x2_sg U4239 ( .A(n5040), .B(n4422), .X(n1968) );
  nor_x2_sg U4240 ( .A(n5042), .B(n4412), .X(n2262) );
  nor_x2_sg U4241 ( .A(n5045), .B(n2218), .X(n2255) );
  nor_x2_sg U4242 ( .A(n5043), .B(n4411), .X(n2268) );
  nor_x2_sg U4243 ( .A(n4842), .B(n4410), .X(n2384) );
  nor_x2_sg U4244 ( .A(n4849), .B(n4410), .X(n2412) );
  nor_x4_sg U4245 ( .A(n2436), .B(n2432), .X(n386) );
  inv_x4_sg U4246 ( .A(n4105), .X(n4106) );
  nor_x2_sg U4247 ( .A(n4838), .B(n4410), .X(n2368) );
  inv_x4_sg U4248 ( .A(n4388), .X(n4838) );
  nor_x2_sg U4249 ( .A(n4841), .B(n4410), .X(n2380) );
  inv_x4_sg U4250 ( .A(n4382), .X(n4841) );
  nor_x2_sg U4251 ( .A(n4843), .B(n4410), .X(n2388) );
  inv_x4_sg U4252 ( .A(n4380), .X(n4843) );
  nor_x2_sg U4253 ( .A(n4844), .B(n4410), .X(n2392) );
  inv_x4_sg U4254 ( .A(n4390), .X(n4844) );
  nor_x2_sg U4255 ( .A(n4848), .B(n4410), .X(n2408) );
  inv_x4_sg U4256 ( .A(n4386), .X(n4848) );
  nor_x2_sg U4257 ( .A(n4276), .B(n4911), .X(n1896) );
  inv_x4_sg U4258 ( .A(n1750), .X(n4911) );
  nor_x2_sg U4259 ( .A(n4394), .B(n4907), .X(n1900) );
  inv_x4_sg U4260 ( .A(n1755), .X(n4907) );
  inv_x4_sg U4261 ( .A(n4107), .X(n4108) );
  nand_x4_sg U4262 ( .A(n4898), .B(n2572), .X(n1709) );
  inv_x4_sg U4263 ( .A(n2571), .X(n4898) );
  inv_x2_sg U4264 ( .A(\mean_pooling_0/n672 ), .X(n4121) );
  inv_x2_sg U4265 ( .A(\reg_im[1][7] ), .X(n4123) );
  inv_x2_sg U4266 ( .A(\reg_im[1][6] ), .X(n4125) );
  inv_x2_sg U4267 ( .A(\reg_im[3][18] ), .X(n4127) );
  inv_x2_sg U4268 ( .A(\reg_im[3][17] ), .X(n4129) );
  inv_x2_sg U4269 ( .A(\reg_im[3][15] ), .X(n4131) );
  inv_x2_sg U4270 ( .A(\reg_im[3][14] ), .X(n4133) );
  inv_x2_sg U4271 ( .A(\reg_im[3][13] ), .X(n4135) );
  inv_x2_sg U4272 ( .A(\reg_im[3][8] ), .X(n4137) );
  inv_x2_sg U4273 ( .A(\reg_im[3][3] ), .X(n4139) );
  inv_x2_sg U4274 ( .A(\reg_im[3][1] ), .X(n4141) );
  inv_x2_sg U4275 ( .A(\reg_im[1][5] ), .X(n4143) );
  inv_x2_sg U4276 ( .A(\reg_im[0][18] ), .X(n4243) );
  inv_x2_sg U4277 ( .A(\reg_im[0][17] ), .X(n4245) );
  inv_x2_sg U4278 ( .A(\reg_im[0][15] ), .X(n4247) );
  inv_x2_sg U4279 ( .A(\reg_im[0][14] ), .X(n4249) );
  inv_x2_sg U4280 ( .A(\reg_im[0][13] ), .X(n4251) );
  inv_x2_sg U4281 ( .A(\reg_im[0][3] ), .X(n4253) );
  inv_x2_sg U4282 ( .A(\reg_im[0][1] ), .X(n4255) );
  inv_x2_sg U4283 ( .A(\reg_im[3][16] ), .X(n4145) );
  inv_x2_sg U4284 ( .A(\reg_im[3][12] ), .X(n4147) );
  inv_x2_sg U4285 ( .A(\reg_im[3][11] ), .X(n4149) );
  inv_x2_sg U4286 ( .A(\reg_im[3][10] ), .X(n4151) );
  inv_x2_sg U4287 ( .A(\reg_im[3][9] ), .X(n4153) );
  inv_x2_sg U4288 ( .A(\reg_im[3][5] ), .X(n4155) );
  inv_x2_sg U4289 ( .A(\reg_im[3][0] ), .X(n4157) );
  inv_x2_sg U4290 ( .A(\reg_im[0][16] ), .X(n4257) );
  inv_x2_sg U4291 ( .A(\reg_im[0][12] ), .X(n4259) );
  inv_x2_sg U4292 ( .A(\reg_im[0][10] ), .X(n4261) );
  inv_x2_sg U4293 ( .A(\reg_im[0][5] ), .X(n4263) );
  inv_x2_sg U4294 ( .A(\reg_im[0][0] ), .X(n4265) );
  inv_x2_sg U4295 ( .A(\reg_im[3][19] ), .X(n4159) );
  inv_x2_sg U4296 ( .A(\reg_im[3][7] ), .X(n4161) );
  inv_x2_sg U4297 ( .A(\reg_im[3][4] ), .X(n4163) );
  inv_x2_sg U4298 ( .A(\reg_im[3][6] ), .X(n4165) );
  inv_x2_sg U4299 ( .A(\reg_im[3][2] ), .X(n4167) );
  inv_x2_sg U4300 ( .A(\reg_im[1][2] ), .X(n4169) );
  inv_x2_sg U4301 ( .A(\reg_im[2][2] ), .X(n4171) );
  inv_x2_sg U4302 ( .A(\reg_im[1][0] ), .X(n4173) );
  inv_x2_sg U4303 ( .A(\reg_im[2][0] ), .X(n4175) );
  inv_x2_sg U4304 ( .A(\reg_im[1][4] ), .X(n4177) );
  inv_x2_sg U4305 ( .A(\reg_im[1][19] ), .X(n4179) );
  inv_x2_sg U4306 ( .A(\reg_im[1][16] ), .X(n4181) );
  inv_x2_sg U4307 ( .A(\reg_im[1][12] ), .X(n4183) );
  inv_x2_sg U4308 ( .A(\reg_im[1][11] ), .X(n4185) );
  inv_x2_sg U4309 ( .A(\reg_im[1][10] ), .X(n4187) );
  inv_x2_sg U4310 ( .A(\reg_im[1][9] ), .X(n4189) );
  inv_x2_sg U4311 ( .A(\reg_im[2][19] ), .X(n4191) );
  inv_x2_sg U4312 ( .A(\reg_im[2][16] ), .X(n4193) );
  inv_x2_sg U4313 ( .A(\reg_im[2][12] ), .X(n4195) );
  inv_x2_sg U4314 ( .A(\reg_im[2][11] ), .X(n4197) );
  inv_x2_sg U4315 ( .A(\reg_im[2][10] ), .X(n4199) );
  inv_x2_sg U4316 ( .A(\reg_im[2][9] ), .X(n4201) );
  inv_x2_sg U4317 ( .A(\reg_im[2][7] ), .X(n4203) );
  inv_x2_sg U4318 ( .A(\reg_im[2][6] ), .X(n4205) );
  inv_x2_sg U4319 ( .A(\reg_im[2][5] ), .X(n4207) );
  inv_x2_sg U4320 ( .A(\reg_im[2][4] ), .X(n4209) );
  inv_x2_sg U4321 ( .A(\reg_im[1][18] ), .X(n4211) );
  inv_x2_sg U4322 ( .A(\reg_im[1][17] ), .X(n4213) );
  inv_x2_sg U4323 ( .A(\reg_im[1][15] ), .X(n4215) );
  inv_x2_sg U4324 ( .A(\reg_im[1][14] ), .X(n4217) );
  inv_x2_sg U4325 ( .A(\reg_im[1][13] ), .X(n4219) );
  inv_x2_sg U4326 ( .A(\reg_im[1][8] ), .X(n4221) );
  inv_x2_sg U4327 ( .A(\reg_im[1][3] ), .X(n4223) );
  inv_x2_sg U4328 ( .A(\reg_im[1][1] ), .X(n4225) );
  inv_x2_sg U4329 ( .A(\reg_im[2][18] ), .X(n4227) );
  inv_x2_sg U4330 ( .A(\reg_im[2][17] ), .X(n4229) );
  inv_x2_sg U4331 ( .A(\reg_im[2][15] ), .X(n4231) );
  inv_x2_sg U4332 ( .A(\reg_im[2][14] ), .X(n4233) );
  inv_x2_sg U4333 ( .A(\reg_im[2][13] ), .X(n4235) );
  inv_x2_sg U4334 ( .A(\reg_im[2][8] ), .X(n4237) );
  inv_x2_sg U4335 ( .A(\reg_im[2][3] ), .X(n4239) );
  inv_x2_sg U4336 ( .A(\reg_im[2][1] ), .X(n4241) );
  nor_x2_sg U4337 ( .A(n1826), .B(n4813), .X(n2020) );
  nor_x4_sg U4338 ( .A(n3054), .B(n3055), .X(n3049) );
  nor_x4_sg U4339 ( .A(state[1]), .B(n3056), .X(n3055) );
  nor_x4_sg U4340 ( .A(input_ready), .B(state[0]), .X(n3056) );
  nor_x2_sg U4341 ( .A(n4998), .B(n4384), .X(n2344) );
  inv_x4_sg U4342 ( .A(n2138), .X(n4998) );
  nor_x2_sg U4343 ( .A(n5003), .B(n4274), .X(n2343) );
  inv_x4_sg U4344 ( .A(n2060), .X(n5003) );
  inv_x4_sg U4345 ( .A(n4031), .X(n4109) );
  inv_x8_sg U4346 ( .A(n4109), .X(n4110) );
  inv_x4_sg U4347 ( .A(n3985), .X(n4111) );
  inv_x8_sg U4348 ( .A(n4111), .X(n4112) );
  inv_x4_sg U4349 ( .A(n4027), .X(n4113) );
  inv_x8_sg U4350 ( .A(n4113), .X(n4114) );
  nor_x2_sg U4351 ( .A(n4806), .B(n1972), .X(n1862) );
  nor_x2_sg U4352 ( .A(n4845), .B(n4410), .X(n2396) );
  nor_x2_sg U4353 ( .A(n4847), .B(n4410), .X(n2404) );
  nor_x4_sg U4354 ( .A(n4408), .B(n2432), .X(n394) );
  nor_x2_sg U4355 ( .A(n4851), .B(n4410), .X(n2420) );
  inv_x4_sg U4356 ( .A(n4384), .X(n4851) );
  inv_x4_sg U4357 ( .A(n2057), .X(n4918) );
  inv_x4_sg U4358 ( .A(n2070), .X(n4908) );
  nor_x2_sg U4359 ( .A(n4930), .B(n4400), .X(n1939) );
  inv_x4_sg U4360 ( .A(n1813), .X(n4930) );
  inv_x4_sg U4361 ( .A(n4115), .X(n4116) );
  inv_x4_sg U4362 ( .A(n4117), .X(n4118) );
  inv_x4_sg U4363 ( .A(n4119), .X(n4120) );
  nand_x4_sg U4364 ( .A(n4964), .B(n4364), .X(n2181) );
  inv_x2_sg U4365 ( .A(\mean_pooling_0/n670 ), .X(n4283) );
  inv_x2_sg U4366 ( .A(\mean_pooling_0/n671 ), .X(n4285) );
  inv_x2_sg U4367 ( .A(\mean_pooling_0/n673 ), .X(n4287) );
  inv_x2_sg U4368 ( .A(\mean_pooling_0/n674 ), .X(n4289) );
  inv_x2_sg U4369 ( .A(\mean_pooling_0/n675 ), .X(n4291) );
  inv_x2_sg U4370 ( .A(\mean_pooling_0/n676 ), .X(n4293) );
  inv_x2_sg U4371 ( .A(\mean_pooling_0/n677 ), .X(n4295) );
  inv_x2_sg U4372 ( .A(\mean_pooling_0/n678 ), .X(n4297) );
  inv_x2_sg U4373 ( .A(\mean_pooling_0/n679 ), .X(n4299) );
  inv_x2_sg U4374 ( .A(\mean_pooling_0/n680 ), .X(n4301) );
  inv_x2_sg U4375 ( .A(\mean_pooling_0/n681 ), .X(n4303) );
  inv_x2_sg U4376 ( .A(\mean_pooling_0/n682 ), .X(n4305) );
  inv_x2_sg U4377 ( .A(\mean_pooling_0/n683 ), .X(n4307) );
  inv_x2_sg U4378 ( .A(\mean_pooling_0/n684 ), .X(n4309) );
  inv_x2_sg U4379 ( .A(\mean_pooling_0/n685 ), .X(n4311) );
  inv_x2_sg U4380 ( .A(\mean_pooling_0/n686 ), .X(n4313) );
  inv_x2_sg U4381 ( .A(\mean_pooling_0/n687 ), .X(n4315) );
  inv_x2_sg U4382 ( .A(\min_pooling_0/n873 ), .X(n4339) );
  inv_x2_sg U4383 ( .A(\max_pooling_0/n821 ), .X(n4333) );
  inv_x2_sg U4384 ( .A(\reg_im[0][8] ), .X(n4317) );
  inv_x2_sg U4385 ( .A(\reg_im[0][11] ), .X(n4319) );
  inv_x2_sg U4386 ( .A(\reg_im[0][9] ), .X(n4321) );
  inv_x2_sg U4387 ( .A(\reg_im[0][19] ), .X(n4323) );
  inv_x2_sg U4388 ( .A(\reg_im[0][7] ), .X(n4325) );
  inv_x2_sg U4389 ( .A(\reg_im[0][4] ), .X(n4327) );
  inv_x2_sg U4390 ( .A(\reg_im[0][6] ), .X(n4329) );
  inv_x2_sg U4391 ( .A(\reg_im[0][2] ), .X(n4331) );
  nor_x2_sg U4392 ( .A(n5010), .B(n4392), .X(n2333) );
  inv_x4_sg U4393 ( .A(n2143), .X(n5010) );
  nor_x2_sg U4394 ( .A(n4836), .B(n2105), .X(n2224) );
  nor_x2_sg U4395 ( .A(n1786), .B(n4808), .X(n1850) );
  nor_x2_sg U4396 ( .A(n1783), .B(n4803), .X(n1910) );
  nor_x2_sg U4397 ( .A(n1745), .B(n4812), .X(n2030) );
  nor_x2_sg U4398 ( .A(n1821), .B(n4811), .X(n2031) );
  inv_x4_sg U4399 ( .A(reset), .X(n5023) );
  nand_x2_sg U4400 ( .A(n5027), .B(n5023), .X(n3411) );
  nor_x4_sg U4401 ( .A(n1687), .B(n4897), .X(n2571) );
  inv_x4_sg U4402 ( .A(n2632), .X(n4897) );
  inv_x4_sg U4403 ( .A(n4121), .X(n4122) );
  inv_x4_sg U4404 ( .A(n2432), .X(n5025) );
  nand_x8_sg U4405 ( .A(state[0]), .B(n5026), .X(n2432) );
  nor_x4_sg U4406 ( .A(n4378), .B(n4950), .X(n1875) );
  inv_x4_sg U4407 ( .A(n1818), .X(n4950) );
  inv_x4_sg U4408 ( .A(n2110), .X(n4945) );
  nor_x2_sg U4409 ( .A(n4402), .B(n5015), .X(n2012) );
  inv_x4_sg U4410 ( .A(n1775), .X(n5015) );
  nor_x2_sg U4411 ( .A(n2466), .B(n4999), .X(n2585) );
  inv_x4_sg U4412 ( .A(n2463), .X(n4999) );
  inv_x4_sg U4413 ( .A(n2128), .X(n4931) );
  inv_x4_sg U4414 ( .A(n2487), .X(n4974) );
  inv_x4_sg U4415 ( .A(n2501), .X(n4961) );
  inv_x4_sg U4416 ( .A(n2515), .X(n4948) );
  inv_x4_sg U4417 ( .A(n2529), .X(n4934) );
  inv_x4_sg U4418 ( .A(n2543), .X(n4921) );
  inv_x4_sg U4419 ( .A(n4123), .X(n4124) );
  inv_x4_sg U4420 ( .A(n4125), .X(n4126) );
  inv_x4_sg U4421 ( .A(n4127), .X(n4128) );
  inv_x4_sg U4422 ( .A(n4129), .X(n4130) );
  inv_x4_sg U4423 ( .A(n4131), .X(n4132) );
  inv_x4_sg U4424 ( .A(n4133), .X(n4134) );
  inv_x4_sg U4425 ( .A(n4135), .X(n4136) );
  inv_x4_sg U4426 ( .A(n4137), .X(n4138) );
  inv_x4_sg U4427 ( .A(n4139), .X(n4140) );
  inv_x4_sg U4428 ( .A(n4141), .X(n4142) );
  inv_x4_sg U4429 ( .A(n4143), .X(n4144) );
  inv_x4_sg U4430 ( .A(n4145), .X(n4146) );
  inv_x4_sg U4431 ( .A(n4147), .X(n4148) );
  inv_x4_sg U4432 ( .A(n4149), .X(n4150) );
  inv_x4_sg U4433 ( .A(n4151), .X(n4152) );
  inv_x4_sg U4434 ( .A(n4153), .X(n4154) );
  inv_x4_sg U4435 ( .A(n4155), .X(n4156) );
  inv_x4_sg U4436 ( .A(n4157), .X(n4158) );
  inv_x4_sg U4437 ( .A(n4159), .X(n4160) );
  inv_x4_sg U4438 ( .A(n4161), .X(n4162) );
  inv_x4_sg U4439 ( .A(n4163), .X(n4164) );
  inv_x4_sg U4440 ( .A(n4165), .X(n4166) );
  inv_x4_sg U4441 ( .A(n4167), .X(n4168) );
  inv_x4_sg U4442 ( .A(n4169), .X(n4170) );
  inv_x4_sg U4443 ( .A(n4171), .X(n4172) );
  inv_x4_sg U4444 ( .A(n4173), .X(n4174) );
  inv_x4_sg U4445 ( .A(n4175), .X(n4176) );
  inv_x4_sg U4446 ( .A(n4177), .X(n4178) );
  inv_x4_sg U4447 ( .A(n4179), .X(n4180) );
  inv_x4_sg U4448 ( .A(n4181), .X(n4182) );
  inv_x4_sg U4449 ( .A(n4183), .X(n4184) );
  inv_x4_sg U4450 ( .A(n4185), .X(n4186) );
  inv_x4_sg U4451 ( .A(n4187), .X(n4188) );
  inv_x4_sg U4452 ( .A(n4189), .X(n4190) );
  inv_x4_sg U4453 ( .A(n4191), .X(n4192) );
  inv_x4_sg U4454 ( .A(n4193), .X(n4194) );
  inv_x4_sg U4455 ( .A(n4195), .X(n4196) );
  inv_x4_sg U4456 ( .A(n4197), .X(n4198) );
  inv_x4_sg U4457 ( .A(n4199), .X(n4200) );
  inv_x4_sg U4458 ( .A(n4201), .X(n4202) );
  inv_x4_sg U4459 ( .A(n4203), .X(n4204) );
  inv_x4_sg U4460 ( .A(n4205), .X(n4206) );
  inv_x4_sg U4461 ( .A(n4207), .X(n4208) );
  inv_x4_sg U4462 ( .A(n4209), .X(n4210) );
  inv_x4_sg U4463 ( .A(n4211), .X(n4212) );
  inv_x4_sg U4464 ( .A(n4213), .X(n4214) );
  inv_x4_sg U4465 ( .A(n4215), .X(n4216) );
  inv_x4_sg U4466 ( .A(n4217), .X(n4218) );
  inv_x4_sg U4467 ( .A(n4219), .X(n4220) );
  inv_x4_sg U4468 ( .A(n4221), .X(n4222) );
  inv_x4_sg U4469 ( .A(n4223), .X(n4224) );
  inv_x4_sg U4470 ( .A(n4225), .X(n4226) );
  inv_x4_sg U4471 ( .A(n4227), .X(n4228) );
  inv_x4_sg U4472 ( .A(n4229), .X(n4230) );
  inv_x4_sg U4473 ( .A(n4231), .X(n4232) );
  inv_x4_sg U4474 ( .A(n4233), .X(n4234) );
  inv_x4_sg U4475 ( .A(n4235), .X(n4236) );
  inv_x4_sg U4476 ( .A(n4237), .X(n4238) );
  inv_x4_sg U4477 ( .A(n4239), .X(n4240) );
  inv_x4_sg U4478 ( .A(n4241), .X(n4242) );
  nor_x2_sg U4479 ( .A(n4390), .B(n4951), .X(n2182) );
  nand_x4_sg U4480 ( .A(n4951), .B(n4390), .X(n2189) );
  inv_x4_sg U4481 ( .A(n2133), .X(n4951) );
  nor_x2_sg U4482 ( .A(n4912), .B(n4388), .X(n2205) );
  inv_x4_sg U4483 ( .A(n2065), .X(n4912) );
  nor_x2_sg U4484 ( .A(n4386), .B(n4977), .X(n2164) );
  nand_x4_sg U4485 ( .A(n4977), .B(n4386), .X(n2166) );
  inv_x4_sg U4486 ( .A(n2102), .X(n4977) );
  inv_x4_sg U4487 ( .A(n4243), .X(n4244) );
  inv_x4_sg U4488 ( .A(n4245), .X(n4246) );
  inv_x4_sg U4489 ( .A(n4247), .X(n4248) );
  inv_x4_sg U4490 ( .A(n4249), .X(n4250) );
  inv_x4_sg U4491 ( .A(n4251), .X(n4252) );
  inv_x4_sg U4492 ( .A(n4253), .X(n4254) );
  inv_x4_sg U4493 ( .A(n4255), .X(n4256) );
  inv_x4_sg U4494 ( .A(n4257), .X(n4258) );
  inv_x4_sg U4495 ( .A(n4259), .X(n4260) );
  inv_x4_sg U4496 ( .A(n4261), .X(n4262) );
  inv_x4_sg U4497 ( .A(n4263), .X(n4264) );
  inv_x4_sg U4498 ( .A(n4265), .X(n4266) );
  inv_x4_sg U4499 ( .A(n4023), .X(n4267) );
  inv_x8_sg U4500 ( .A(n4267), .X(n4268) );
  inv_x4_sg U4501 ( .A(n4268), .X(n4813) );
  inv_x4_sg U4502 ( .A(n4075), .X(n4269) );
  inv_x8_sg U4503 ( .A(n4269), .X(state[1]) );
  inv_x8_sg U4504 ( .A(state[1]), .X(n5026) );
  inv_x8_sg U4505 ( .A(n4100), .X(n4834) );
  inv_x8_sg U4506 ( .A(n4102), .X(n4801) );
  inv_x8_sg U4507 ( .A(n4104), .X(n4815) );
  inv_x4_sg U4508 ( .A(n4071), .X(n4271) );
  inv_x8_sg U4509 ( .A(n4271), .X(n4272) );
  inv_x4_sg U4510 ( .A(n4272), .X(n4853) );
  inv_x4_sg U4511 ( .A(n4067), .X(n4273) );
  inv_x8_sg U4512 ( .A(n4273), .X(n4274) );
  inv_x4_sg U4513 ( .A(n3993), .X(n4275) );
  inv_x8_sg U4514 ( .A(n4275), .X(n4276) );
  inv_x4_sg U4515 ( .A(n4276), .X(n4804) );
  inv_x4_sg U4516 ( .A(n3997), .X(n4277) );
  inv_x8_sg U4517 ( .A(n4277), .X(n4278) );
  inv_x1_sg U4518 ( .A(n2462), .X(n4995) );
  nor_x2_sg U4519 ( .A(n4807), .B(n1851), .X(n1849) );
  inv_x4_sg U4520 ( .A(n4279), .X(n4280) );
  nor_x4_sg U4521 ( .A(n3433), .B(n4433), .X(n3065) );
  nor_x4_sg U4522 ( .A(n3435), .B(n4433), .X(n3157) );
  nor_x4_sg U4523 ( .A(n3434), .B(n5017), .X(n2046) );
  inv_x4_sg U4524 ( .A(n2146), .X(n5017) );
  nor_x4_sg U4525 ( .A(mode[0]), .B(mode[1]), .X(n2428) );
  inv_x4_sg U4526 ( .A(n4283), .X(n4284) );
  inv_x4_sg U4527 ( .A(n4285), .X(n4286) );
  inv_x4_sg U4528 ( .A(n4287), .X(n4288) );
  inv_x4_sg U4529 ( .A(n4289), .X(n4290) );
  inv_x4_sg U4530 ( .A(n4291), .X(n4292) );
  inv_x4_sg U4531 ( .A(n4293), .X(n4294) );
  inv_x4_sg U4532 ( .A(n4295), .X(n4296) );
  inv_x4_sg U4533 ( .A(n4297), .X(n4298) );
  inv_x4_sg U4534 ( .A(n4299), .X(n4300) );
  inv_x4_sg U4535 ( .A(n4301), .X(n4302) );
  inv_x4_sg U4536 ( .A(n4303), .X(n4304) );
  inv_x4_sg U4537 ( .A(n4305), .X(n4306) );
  inv_x4_sg U4538 ( .A(n4307), .X(n4308) );
  inv_x4_sg U4539 ( .A(n4309), .X(n4310) );
  inv_x4_sg U4540 ( .A(n4311), .X(n4312) );
  inv_x4_sg U4541 ( .A(n4313), .X(n4314) );
  inv_x4_sg U4542 ( .A(n4315), .X(n4316) );
  inv_x4_sg U4543 ( .A(n4317), .X(n4318) );
  inv_x8_sg U4544 ( .A(n4318), .X(n5041) );
  inv_x4_sg U4545 ( .A(n4319), .X(n4320) );
  inv_x8_sg U4546 ( .A(n4320), .X(n5038) );
  inv_x4_sg U4547 ( .A(n4321), .X(n4322) );
  inv_x8_sg U4548 ( .A(n4322), .X(n5040) );
  inv_x4_sg U4549 ( .A(n4323), .X(n4324) );
  inv_x8_sg U4550 ( .A(n4324), .X(n5030) );
  inv_x4_sg U4551 ( .A(n4325), .X(n4326) );
  inv_x8_sg U4552 ( .A(n4326), .X(n5042) );
  inv_x4_sg U4553 ( .A(n4327), .X(n4328) );
  inv_x8_sg U4554 ( .A(n4328), .X(n5045) );
  inv_x4_sg U4555 ( .A(n4329), .X(n4330) );
  inv_x8_sg U4556 ( .A(n4330), .X(n5043) );
  inv_x4_sg U4557 ( .A(n4331), .X(n4332) );
  inv_x8_sg U4558 ( .A(n4332), .X(n5047) );
  nor_x2_sg U4559 ( .A(n2449), .B(n5006), .X(n2578) );
  inv_x4_sg U4560 ( .A(n2452), .X(n5006) );
  inv_x4_sg U4561 ( .A(n2480), .X(n4981) );
  inv_x4_sg U4562 ( .A(n2494), .X(n4968) );
  inv_x4_sg U4563 ( .A(n2508), .X(n4955) );
  inv_x4_sg U4564 ( .A(n2522), .X(n4942) );
  inv_x4_sg U4565 ( .A(n2536), .X(n4928) );
  inv_x4_sg U4566 ( .A(n2550), .X(n4915) );
  inv_x4_sg U4567 ( .A(n4128), .X(n5007) );
  inv_x4_sg U4568 ( .A(n4138), .X(n4943) );
  inv_x4_sg U4569 ( .A(n4130), .X(n5001) );
  inv_x4_sg U4570 ( .A(n4156), .X(n4922) );
  inv_x4_sg U4571 ( .A(n4144), .X(n4859) );
  inv_x4_sg U4572 ( .A(n4136), .X(n4975) );
  inv_x4_sg U4573 ( .A(n4132), .X(n4988) );
  inv_x4_sg U4574 ( .A(n4146), .X(n4996) );
  inv_x4_sg U4575 ( .A(n4142), .X(n4900) );
  inv_x4_sg U4576 ( .A(n4172), .X(n4876) );
  inv_x4_sg U4577 ( .A(n4134), .X(n4982) );
  inv_x4_sg U4578 ( .A(n4148), .X(n4969) );
  inv_x4_sg U4579 ( .A(n4150), .X(n4962) );
  inv_x4_sg U4580 ( .A(n4152), .X(n4956) );
  inv_x4_sg U4581 ( .A(n4154), .X(n4949) );
  inv_x4_sg U4582 ( .A(n4140), .X(n4910) );
  inv_x4_sg U4583 ( .A(n4168), .X(n4906) );
  inv_x4_sg U4584 ( .A(n4170), .X(n4856) );
  inv_x4_sg U4585 ( .A(n4158), .X(n4894) );
  inv_x4_sg U4586 ( .A(n4160), .X(n5014) );
  inv_x4_sg U4587 ( .A(n4162), .X(n4935) );
  inv_x4_sg U4588 ( .A(n4164), .X(n4916) );
  inv_x4_sg U4589 ( .A(n4166), .X(n4929) );
  inv_x4_sg U4590 ( .A(n4124), .X(n4861) );
  inv_x4_sg U4591 ( .A(n4126), .X(n4860) );
  nor_x4_sg U4592 ( .A(n2435), .B(n5020), .X(n2431) );
  nand_x4_sg U4593 ( .A(n5025), .B(mode[1]), .X(n2435) );
  inv_x4_sg U4594 ( .A(n4176), .X(n4874) );
  inv_x4_sg U4595 ( .A(n4174), .X(n4854) );
  inv_x4_sg U4596 ( .A(n4182), .X(n4870) );
  inv_x4_sg U4597 ( .A(n4180), .X(n4873) );
  inv_x4_sg U4598 ( .A(n4184), .X(n4866) );
  inv_x4_sg U4599 ( .A(n4186), .X(n4865) );
  inv_x4_sg U4600 ( .A(n4188), .X(n4864) );
  inv_x4_sg U4601 ( .A(n4190), .X(n4863) );
  inv_x4_sg U4602 ( .A(n4178), .X(n4858) );
  inv_x4_sg U4603 ( .A(n4194), .X(n4890) );
  inv_x4_sg U4604 ( .A(n4212), .X(n4872) );
  inv_x4_sg U4605 ( .A(n4222), .X(n4862) );
  inv_x4_sg U4606 ( .A(n4198), .X(n4885) );
  inv_x4_sg U4607 ( .A(n4214), .X(n4871) );
  inv_x4_sg U4608 ( .A(n4208), .X(n4879) );
  inv_x4_sg U4609 ( .A(n4202), .X(n4883) );
  inv_x4_sg U4610 ( .A(n4200), .X(n4884) );
  inv_x4_sg U4611 ( .A(n4196), .X(n4886) );
  inv_x4_sg U4612 ( .A(n4220), .X(n4867) );
  inv_x4_sg U4613 ( .A(n4216), .X(n4869) );
  inv_x4_sg U4614 ( .A(n4192), .X(n4893) );
  inv_x4_sg U4615 ( .A(n4226), .X(n4855) );
  inv_x4_sg U4616 ( .A(n4218), .X(n4868) );
  inv_x4_sg U4617 ( .A(n4224), .X(n4857) );
  inv_x4_sg U4618 ( .A(n4204), .X(n4881) );
  inv_x4_sg U4619 ( .A(n4210), .X(n4878) );
  inv_x4_sg U4620 ( .A(n4206), .X(n4880) );
  inv_x4_sg U4621 ( .A(n4234), .X(n4888) );
  inv_x4_sg U4622 ( .A(n4242), .X(n4875) );
  inv_x4_sg U4623 ( .A(n4238), .X(n4882) );
  inv_x4_sg U4624 ( .A(n4236), .X(n4887) );
  inv_x4_sg U4625 ( .A(n4232), .X(n4889) );
  inv_x4_sg U4626 ( .A(n4230), .X(n4891) );
  inv_x4_sg U4627 ( .A(n4228), .X(n4892) );
  inv_x4_sg U4628 ( .A(n4240), .X(n4877) );
  inv_x4_sg U4629 ( .A(n4333), .X(n4334) );
  inv_x4_sg U4630 ( .A(n4334), .X(n4835) );
  inv_x4_sg U4631 ( .A(n4061), .X(n4335) );
  inv_x8_sg U4632 ( .A(n4335), .X(n4336) );
  inv_x8_sg U4633 ( .A(n4336), .X(n4849) );
  nor_x8_sg U4634 ( .A(n5020), .B(mode[1]), .X(n2434) );
  inv_x8_sg U4635 ( .A(mode[0]), .X(n5020) );
  inv_x4_sg U4636 ( .A(n3989), .X(n4337) );
  inv_x8_sg U4637 ( .A(n4337), .X(n4338) );
  inv_x4_sg U4638 ( .A(n4338), .X(n4803) );
  inv_x4_sg U4639 ( .A(n4339), .X(n4340) );
  inv_x4_sg U4640 ( .A(n4017), .X(n4341) );
  inv_x8_sg U4641 ( .A(n4341), .X(n4342) );
  inv_x4_sg U4642 ( .A(n4342), .X(n4810) );
  inv_x4_sg U4643 ( .A(n4013), .X(n4343) );
  inv_x8_sg U4644 ( .A(n4343), .X(n4344) );
  inv_x4_sg U4645 ( .A(n4344), .X(n4808) );
  inv_x4_sg U4646 ( .A(n4015), .X(n4345) );
  inv_x8_sg U4647 ( .A(n4345), .X(n4346) );
  inv_x4_sg U4648 ( .A(n4346), .X(n4809) );
  inv_x4_sg U4649 ( .A(n4007), .X(n4347) );
  inv_x8_sg U4650 ( .A(n4347), .X(n4348) );
  inv_x4_sg U4651 ( .A(n4348), .X(n4806) );
  inv_x4_sg U4652 ( .A(n4011), .X(n4349) );
  inv_x8_sg U4653 ( .A(n4349), .X(n4350) );
  inv_x4_sg U4654 ( .A(n4350), .X(n4807) );
  inv_x4_sg U4655 ( .A(n4019), .X(n4351) );
  inv_x8_sg U4656 ( .A(n4351), .X(n4352) );
  inv_x4_sg U4657 ( .A(n4352), .X(n4811) );
  inv_x4_sg U4658 ( .A(n4053), .X(n4353) );
  inv_x8_sg U4659 ( .A(n4353), .X(n4354) );
  inv_x4_sg U4660 ( .A(n4354), .X(n4845) );
  inv_x4_sg U4661 ( .A(n4021), .X(n4355) );
  inv_x8_sg U4662 ( .A(n4355), .X(n4356) );
  inv_x4_sg U4663 ( .A(n4356), .X(n4812) );
  inv_x4_sg U4664 ( .A(n4057), .X(n4357) );
  inv_x8_sg U4665 ( .A(n4357), .X(n4358) );
  inv_x4_sg U4666 ( .A(n4358), .X(n4847) );
  inv_x4_sg U4667 ( .A(n4043), .X(n4359) );
  inv_x8_sg U4668 ( .A(n4359), .X(n4360) );
  inv_x4_sg U4669 ( .A(n4360), .X(n4840) );
  inv_x4_sg U4670 ( .A(n4047), .X(n4361) );
  inv_x8_sg U4671 ( .A(n4361), .X(n4362) );
  inv_x4_sg U4672 ( .A(n4362), .X(n4842) );
  inv_x4_sg U4673 ( .A(n4055), .X(n4363) );
  inv_x8_sg U4674 ( .A(n4363), .X(n4364) );
  inv_x4_sg U4675 ( .A(n4364), .X(n4846) );
  nor_x2_sg U4676 ( .A(n5031), .B(n4427), .X(n3405) );
  nor_x2_sg U4677 ( .A(n5031), .B(n1905), .X(n2026) );
  nor_x2_sg U4678 ( .A(n5031), .B(n2218), .X(n2339) );
  nor_x2_sg U4679 ( .A(n4417), .B(n5031), .X(n2744) );
  inv_x8_sg U4680 ( .A(n4244), .X(n5031) );
  nor_x2_sg U4681 ( .A(n5032), .B(n3334), .X(n3401) );
  nor_x2_sg U4682 ( .A(n5032), .B(n4421), .X(n2040) );
  nor_x2_sg U4683 ( .A(n2637), .B(n5032), .X(n2738) );
  nor_x2_sg U4684 ( .A(n5032), .B(n4411), .X(n2353) );
  inv_x8_sg U4685 ( .A(n4246), .X(n5032) );
  nor_x2_sg U4686 ( .A(n5033), .B(n4426), .X(n3397) );
  nor_x2_sg U4687 ( .A(n5033), .B(n4422), .X(n2034) );
  nor_x2_sg U4688 ( .A(n4416), .B(n5033), .X(n2732) );
  nor_x2_sg U4689 ( .A(n5033), .B(n4412), .X(n2347) );
  inv_x8_sg U4690 ( .A(n4258), .X(n5033) );
  nor_x2_sg U4691 ( .A(n5034), .B(n4427), .X(n3393) );
  nor_x2_sg U4692 ( .A(n5034), .B(n4421), .X(n1994) );
  nor_x2_sg U4693 ( .A(n4417), .B(n5034), .X(n2726) );
  nor_x2_sg U4694 ( .A(n5034), .B(n4412), .X(n2301) );
  inv_x8_sg U4695 ( .A(n4248), .X(n5034) );
  nor_x2_sg U4696 ( .A(n5035), .B(n3334), .X(n3389) );
  nor_x2_sg U4697 ( .A(n5035), .B(n4411), .X(n2307) );
  nor_x2_sg U4698 ( .A(n2637), .B(n5035), .X(n2720) );
  nor_x2_sg U4699 ( .A(n5035), .B(n4422), .X(n1988) );
  inv_x8_sg U4700 ( .A(n4250), .X(n5035) );
  nor_x2_sg U4701 ( .A(n5036), .B(n4426), .X(n3385) );
  nor_x2_sg U4702 ( .A(n5036), .B(n1905), .X(n2001) );
  nor_x2_sg U4703 ( .A(n4416), .B(n5036), .X(n2714) );
  nor_x2_sg U4704 ( .A(n5036), .B(n2218), .X(n2314) );
  inv_x8_sg U4705 ( .A(n4252), .X(n5036) );
  nor_x2_sg U4706 ( .A(n5037), .B(n4427), .X(n3381) );
  nor_x2_sg U4707 ( .A(n4417), .B(n5037), .X(n2708) );
  nor_x2_sg U4708 ( .A(n5037), .B(n4412), .X(n2320) );
  nor_x2_sg U4709 ( .A(n5037), .B(n4422), .X(n2007) );
  inv_x8_sg U4710 ( .A(n4260), .X(n5037) );
  nor_x2_sg U4711 ( .A(n5039), .B(n4426), .X(n3373) );
  nor_x2_sg U4712 ( .A(n4416), .B(n5039), .X(n2696) );
  nor_x2_sg U4713 ( .A(n5039), .B(n1905), .X(n1981) );
  nor_x2_sg U4714 ( .A(n5039), .B(n4411), .X(n2288) );
  inv_x8_sg U4715 ( .A(n4262), .X(n5039) );
  nor_x2_sg U4716 ( .A(n5044), .B(n3334), .X(n3353) );
  nor_x2_sg U4717 ( .A(n5044), .B(n4421), .X(n1933) );
  nor_x2_sg U4718 ( .A(n2637), .B(n5044), .X(n2666) );
  nor_x2_sg U4719 ( .A(n5044), .B(n4411), .X(n2246) );
  inv_x8_sg U4720 ( .A(n4264), .X(n5044) );
  nor_x2_sg U4721 ( .A(n5046), .B(n4427), .X(n3345) );
  nor_x2_sg U4722 ( .A(n4417), .B(n5046), .X(n2654) );
  nor_x2_sg U4723 ( .A(n5046), .B(n4422), .X(n1927) );
  nor_x2_sg U4724 ( .A(n5046), .B(n4412), .X(n2240) );
  inv_x8_sg U4725 ( .A(n4254), .X(n5046) );
  nor_x2_sg U4726 ( .A(n5048), .B(n4426), .X(n3337) );
  nor_x2_sg U4727 ( .A(n5048), .B(n4421), .X(n1915) );
  nor_x2_sg U4728 ( .A(n4416), .B(n5048), .X(n2642) );
  nor_x2_sg U4729 ( .A(n5048), .B(n2218), .X(n2234) );
  inv_x8_sg U4730 ( .A(n4256), .X(n5048) );
  nor_x2_sg U4731 ( .A(n5049), .B(n4427), .X(n3332) );
  nor_x2_sg U4732 ( .A(n5049), .B(n4411), .X(n2228) );
  nor_x2_sg U4733 ( .A(n4417), .B(n5049), .X(n2635) );
  nor_x2_sg U4734 ( .A(n5049), .B(n1905), .X(n1921) );
  inv_x8_sg U4735 ( .A(n4266), .X(n5049) );
  inv_x4_sg U4736 ( .A(n4035), .X(n4365) );
  inv_x8_sg U4737 ( .A(n4365), .X(n4366) );
  inv_x4_sg U4738 ( .A(n4366), .X(n4836) );
  inv_x4_sg U4739 ( .A(n4041), .X(n4367) );
  inv_x8_sg U4740 ( .A(n4367), .X(n4368) );
  inv_x4_sg U4741 ( .A(n4368), .X(n4839) );
  inv_x4_sg U4742 ( .A(n4063), .X(n4369) );
  inv_x8_sg U4743 ( .A(n4369), .X(n4370) );
  inv_x4_sg U4744 ( .A(n4370), .X(n4850) );
  inv_x4_sg U4745 ( .A(n4037), .X(n4371) );
  inv_x8_sg U4746 ( .A(n4371), .X(n4372) );
  inv_x4_sg U4747 ( .A(n4372), .X(n4837) );
  inv_x4_sg U4748 ( .A(n4003), .X(n4373) );
  inv_x4_sg U4749 ( .A(n4009), .X(n4375) );
  inv_x4_sg U4750 ( .A(n4005), .X(n4377) );
  inv_x8_sg U4751 ( .A(n4377), .X(n4378) );
  inv_x4_sg U4752 ( .A(n4049), .X(n4379) );
  inv_x8_sg U4753 ( .A(n4379), .X(n4380) );
  inv_x4_sg U4754 ( .A(n4045), .X(n4381) );
  inv_x8_sg U4755 ( .A(n4381), .X(n4382) );
  inv_x4_sg U4756 ( .A(n4065), .X(n4383) );
  inv_x8_sg U4757 ( .A(n4383), .X(n4384) );
  inv_x4_sg U4758 ( .A(n4059), .X(n4385) );
  inv_x8_sg U4759 ( .A(n4385), .X(n4386) );
  inv_x4_sg U4760 ( .A(n4039), .X(n4387) );
  inv_x8_sg U4761 ( .A(n4387), .X(n4388) );
  inv_x4_sg U4762 ( .A(n4051), .X(n4389) );
  inv_x8_sg U4763 ( .A(n4389), .X(n4390) );
  inv_x8_sg U4764 ( .A(n4110), .X(n5050) );
  inv_x8_sg U4765 ( .A(n4112), .X(n5052) );
  inv_x8_sg U4766 ( .A(n4114), .X(n5051) );
  inv_x4_sg U4767 ( .A(n4069), .X(n4391) );
  inv_x8_sg U4768 ( .A(n4391), .X(n4392) );
  inv_x4_sg U4769 ( .A(n3991), .X(n4393) );
  inv_x8_sg U4770 ( .A(n4393), .X(n4394) );
  inv_x4_sg U4771 ( .A(n3995), .X(n4395) );
  inv_x8_sg U4772 ( .A(n4395), .X(n4396) );
  inv_x4_sg U4773 ( .A(n4001), .X(n4397) );
  inv_x8_sg U4774 ( .A(n4397), .X(n4398) );
  inv_x4_sg U4775 ( .A(n3999), .X(n4399) );
  inv_x8_sg U4776 ( .A(n4399), .X(n4400) );
  inv_x4_sg U4777 ( .A(n4025), .X(n4401) );
  inv_x8_sg U4778 ( .A(n4401), .X(n4402) );
  inv_x4_sg U4779 ( .A(n4073), .X(n4403) );
  inv_x8_sg U4780 ( .A(n4403), .X(state[0]) );
  nand_x1_sg U4781 ( .A(n1709), .B(n3485), .X(n1708) );
  nand_x1_sg U4782 ( .A(n2272), .B(n2189), .X(n2184) );
  nand_x1_sg U4783 ( .A(n2197), .B(n4106), .X(n2196) );
  nand_x1_sg U4784 ( .A(n2259), .B(n2251), .X(n2200) );
  nand_x1_sg U4785 ( .A(n1880), .B(n1881), .X(n1879) );
  nand_x2_sg U4786 ( .A(n4375), .B(n1772), .X(n1867) );
  nor_x1_sg U4787 ( .A(n2738), .B(n3699), .X(n2737) );
  nor_x1_sg U4788 ( .A(n2720), .B(n3703), .X(n2719) );
  nor_x1_sg U4789 ( .A(n2702), .B(n3707), .X(n2701) );
  nor_x1_sg U4790 ( .A(n2684), .B(n3711), .X(n2683) );
  nor_x1_sg U4791 ( .A(n2726), .B(n3651), .X(n2725) );
  nor_x1_sg U4792 ( .A(n1994), .B(n3731), .X(n1993) );
  nor_x1_sg U4793 ( .A(n2001), .B(n3735), .X(n2000) );
  nor_x1_sg U4794 ( .A(n1962), .B(n3739), .X(n1961) );
  nor_x1_sg U4795 ( .A(n2744), .B(n3643), .X(n2743) );
  nor_x1_sg U4796 ( .A(n2714), .B(n3655), .X(n2713) );
  nor_x1_sg U4797 ( .A(n2708), .B(n3659), .X(n2707) );
  nor_x1_sg U4798 ( .A(n2696), .B(n3663), .X(n2695) );
  nor_x1_sg U4799 ( .A(n2690), .B(n3667), .X(n2689) );
  nor_x1_sg U4800 ( .A(n2678), .B(n3671), .X(n2677) );
  nor_x1_sg U4801 ( .A(n2672), .B(n3675), .X(n2671) );
  nor_x1_sg U4802 ( .A(n2666), .B(n3679), .X(n2665) );
  nor_x1_sg U4803 ( .A(n2660), .B(n3683), .X(n2659) );
  nor_x1_sg U4804 ( .A(n2654), .B(n3687), .X(n2653) );
  nor_x1_sg U4805 ( .A(n1927), .B(n3545), .X(n1926) );
  nor_x1_sg U4806 ( .A(n2328), .B(n3627), .X(n2327) );
  nor_x1_sg U4807 ( .A(n2026), .B(n3719), .X(n2025) );
  nor_x1_sg U4808 ( .A(n2040), .B(n3723), .X(n2039) );
  nor_x1_sg U4809 ( .A(n2034), .B(n3727), .X(n2033) );
  nor_x1_sg U4810 ( .A(n1915), .B(n3743), .X(n1914) );
  nor_x1_sg U4811 ( .A(n2307), .B(n3747), .X(n2306) );
  nor_x1_sg U4812 ( .A(n2642), .B(n3635), .X(n2641) );
  nor_x1_sg U4813 ( .A(n4120), .B(n4415), .X(\mean_pooling_0/n298 ) );
  nor_x1_sg U4814 ( .A(n4415), .B(n1723), .X(\mean_pooling_0/n242 ) );
  nand_x1_sg U4815 ( .A(n4120), .B(n3485), .X(n1720) );
  nand_x1_sg U4816 ( .A(n4108), .B(n3485), .X(n1712) );
  nand_x1_sg U4817 ( .A(n4077), .B(n3485), .X(n1696) );
  nand_x2_sg U4818 ( .A(n2633), .B(n2634), .X(n2632) );
  nor_x1_sg U4819 ( .A(n3625), .B(n3623), .X(n2633) );
  nor_x1_sg U4820 ( .A(n2635), .B(n3621), .X(n2634) );
  nor_x1_sg U4821 ( .A(n2547), .B(n4915), .X(n2622) );
  nor_x1_sg U4822 ( .A(n2540), .B(n4921), .X(n2619) );
  nor_x1_sg U4823 ( .A(n2533), .B(n4928), .X(n2616) );
  nor_x1_sg U4824 ( .A(n2526), .B(n4934), .X(n2613) );
  nor_x1_sg U4825 ( .A(n2518), .B(n4942), .X(n2610) );
  nor_x1_sg U4826 ( .A(n2512), .B(n4948), .X(n2607) );
  nor_x1_sg U4827 ( .A(n2505), .B(n4955), .X(n2604) );
  nor_x1_sg U4828 ( .A(n2497), .B(n4961), .X(n2601) );
  nor_x1_sg U4829 ( .A(n2491), .B(n4968), .X(n2598) );
  nor_x1_sg U4830 ( .A(n2484), .B(n4974), .X(n2595) );
  nor_x1_sg U4831 ( .A(n2476), .B(n4981), .X(n2592) );
  nand_x1_sg U4832 ( .A(n5006), .B(n2449), .X(n2580) );
  nand_x1_sg U4833 ( .A(n4118), .B(n3485), .X(n1718) );
  nand_x1_sg U4834 ( .A(n4116), .B(n3485), .X(n1714) );
  inv_x4_sg U4835 ( .A(n1831), .X(n4444) );
  nor_x1_sg U4836 ( .A(n3433), .B(n4424), .X(\min_pooling_0/n355 ) );
  nor_x1_sg U4837 ( .A(n3433), .B(n4423), .X(\min_pooling_0/n354 ) );
  nor_x1_sg U4838 ( .A(n4415), .B(n1717), .X(\mean_pooling_0/n222 ) );
  nor_x1_sg U4839 ( .A(n4415), .B(n1695), .X(\mean_pooling_0/n302 ) );
  nor_x1_sg U4840 ( .A(n4415), .B(n1727), .X(\mean_pooling_0/n294 ) );
  nor_x1_sg U4841 ( .A(n4415), .B(n1691), .X(\mean_pooling_0/n290 ) );
  nor_x1_sg U4842 ( .A(n4118), .B(n4415), .X(\mean_pooling_0/n286 ) );
  nor_x1_sg U4843 ( .A(n4415), .B(n1699), .X(\mean_pooling_0/n282 ) );
  nor_x1_sg U4844 ( .A(n4415), .B(n1725), .X(\mean_pooling_0/n278 ) );
  nor_x1_sg U4845 ( .A(n4108), .B(n4415), .X(\mean_pooling_0/n274 ) );
  nor_x1_sg U4846 ( .A(n4415), .B(n1711), .X(\mean_pooling_0/n270 ) );
  nor_x1_sg U4847 ( .A(n4415), .B(n1703), .X(\mean_pooling_0/n266 ) );
  nor_x1_sg U4848 ( .A(n4116), .B(n4415), .X(\mean_pooling_0/n262 ) );
  nor_x1_sg U4849 ( .A(n4415), .B(n1729), .X(\mean_pooling_0/n258 ) );
  nor_x1_sg U4850 ( .A(n4415), .B(n1701), .X(\mean_pooling_0/n254 ) );
  nor_x1_sg U4851 ( .A(n4415), .B(n1707), .X(\mean_pooling_0/n250 ) );
  nor_x1_sg U4852 ( .A(n4415), .B(n1693), .X(\mean_pooling_0/n246 ) );
  nor_x1_sg U4853 ( .A(n4415), .B(n1705), .X(\mean_pooling_0/n238 ) );
  nor_x1_sg U4854 ( .A(n4077), .B(n4415), .X(\mean_pooling_0/n234 ) );
  nand_x1_sg U4855 ( .A(n4983), .B(n1854), .X(n1853) );
  nand_x4_sg U4856 ( .A(n2551), .B(n4913), .X(n1723) );
  nor_x1_sg U4857 ( .A(n2553), .B(n2554), .X(n2552) );
  nand_x2_sg U4858 ( .A(n5027), .B(n5026), .X(n3327) );
  nor_x1_sg U4859 ( .A(n3503), .B(n2631), .X(n2630) );
  nor_x1_sg U4860 ( .A(n2568), .B(n2571), .X(n2629) );
  nor_x1_sg U4861 ( .A(n4839), .B(n2057), .X(n2250) );
  nor_x1_sg U4862 ( .A(n4850), .B(n4410), .X(n2416) );
  nor_x1_sg U4863 ( .A(n4836), .B(n4410), .X(n2360) );
  nand_x2_sg U4864 ( .A(n4957), .B(n1867), .X(n1972) );
  nand_x2_sg U4865 ( .A(n4970), .B(n1852), .X(n1851) );
  nor_x1_sg U4866 ( .A(n3062), .B(n4854), .X(n1922) );
  nor_x1_sg U4867 ( .A(n4894), .B(n4424), .X(n1924) );
  nor_x1_sg U4868 ( .A(n3071), .B(n4855), .X(n2235) );
  nor_x1_sg U4869 ( .A(n4900), .B(n4414), .X(n2237) );
  nor_x1_sg U4870 ( .A(n3062), .B(n4856), .X(n1904) );
  nor_x1_sg U4871 ( .A(n4906), .B(n4424), .X(n1907) );
  nor_x1_sg U4872 ( .A(n3071), .B(n4856), .X(n2217) );
  nor_x1_sg U4873 ( .A(n4906), .B(n4414), .X(n2220) );
  nor_x1_sg U4874 ( .A(n3062), .B(n4860), .X(n1950) );
  nor_x1_sg U4875 ( .A(n4929), .B(n4424), .X(n1952) );
  nor_x1_sg U4876 ( .A(n3071), .B(n4858), .X(n2256) );
  nor_x1_sg U4877 ( .A(n4916), .B(n4414), .X(n2258) );
  nor_x1_sg U4878 ( .A(n3071), .B(n4857), .X(n2241) );
  nor_x1_sg U4879 ( .A(n4910), .B(n4414), .X(n2243) );
  nor_x1_sg U4880 ( .A(n3071), .B(n4859), .X(n2247) );
  nor_x1_sg U4881 ( .A(n4922), .B(n4414), .X(n2249) );
  nor_x1_sg U4882 ( .A(n3062), .B(n4857), .X(n1928) );
  nor_x1_sg U4883 ( .A(n4910), .B(n4424), .X(n1930) );
  nor_x1_sg U4884 ( .A(n3062), .B(n4858), .X(n1943) );
  nor_x1_sg U4885 ( .A(n4916), .B(n4424), .X(n1945) );
  nor_x1_sg U4886 ( .A(n3071), .B(n4860), .X(n2269) );
  nor_x1_sg U4887 ( .A(n4929), .B(n4414), .X(n2271) );
  nor_x1_sg U4888 ( .A(n3071), .B(n4861), .X(n2263) );
  nor_x1_sg U4889 ( .A(n4935), .B(n4414), .X(n2265) );
  nor_x1_sg U4890 ( .A(n3071), .B(n4862), .X(n2276) );
  nor_x1_sg U4891 ( .A(n4943), .B(n4414), .X(n2278) );
  nor_x1_sg U4892 ( .A(n3071), .B(n4863), .X(n2282) );
  nor_x1_sg U4893 ( .A(n4949), .B(n4414), .X(n2284) );
  nor_x1_sg U4894 ( .A(n3071), .B(n4864), .X(n2289) );
  nor_x1_sg U4895 ( .A(n4956), .B(n4414), .X(n2291) );
  nor_x1_sg U4896 ( .A(n3062), .B(n4863), .X(n1969) );
  nor_x1_sg U4897 ( .A(n4949), .B(n4424), .X(n1971) );
  nor_x1_sg U4898 ( .A(n3062), .B(n4865), .X(n1976) );
  nor_x1_sg U4899 ( .A(n4962), .B(n4424), .X(n1978) );
  nor_x1_sg U4900 ( .A(n3062), .B(n4864), .X(n1982) );
  nor_x1_sg U4901 ( .A(n4956), .B(n4424), .X(n1984) );
  nor_x1_sg U4902 ( .A(n3062), .B(n4866), .X(n2008) );
  nor_x1_sg U4903 ( .A(n4969), .B(n4424), .X(n2010) );
  nor_x1_sg U4904 ( .A(n3062), .B(n4868), .X(n1989) );
  nor_x1_sg U4905 ( .A(n4982), .B(n4424), .X(n1991) );
  nor_x1_sg U4906 ( .A(n3071), .B(n4865), .X(n2295) );
  nor_x1_sg U4907 ( .A(n4962), .B(n4414), .X(n2297) );
  nor_x1_sg U4908 ( .A(n3071), .B(n4867), .X(n2315) );
  nor_x1_sg U4909 ( .A(n4975), .B(n4414), .X(n2317) );
  nor_x1_sg U4910 ( .A(n3071), .B(n4866), .X(n2321) );
  nor_x1_sg U4911 ( .A(n4969), .B(n4414), .X(n2323) );
  nor_x1_sg U4912 ( .A(n3071), .B(n4869), .X(n2302) );
  nor_x1_sg U4913 ( .A(n4988), .B(n4414), .X(n2304) );
  nor_x1_sg U4914 ( .A(n3071), .B(n4871), .X(n2354) );
  nor_x1_sg U4915 ( .A(n5001), .B(n4414), .X(n2356) );
  nor_x1_sg U4916 ( .A(n3071), .B(n4870), .X(n2348) );
  nor_x1_sg U4917 ( .A(n4996), .B(n4414), .X(n2350) );
  nor_x1_sg U4918 ( .A(n3062), .B(n4873), .X(n2016) );
  nor_x1_sg U4919 ( .A(n5014), .B(n4424), .X(n2018) );
  nor_x1_sg U4920 ( .A(n3163), .B(n4854), .X(n2636) );
  nor_x1_sg U4921 ( .A(n4419), .B(n4894), .X(n2639) );
  nor_x1_sg U4922 ( .A(n3162), .B(n4874), .X(n2638) );
  nor_x1_sg U4923 ( .A(n3071), .B(n4873), .X(n2329) );
  nor_x1_sg U4924 ( .A(n5014), .B(n4414), .X(n2331) );
  nor_x1_sg U4925 ( .A(n3163), .B(n4856), .X(n2649) );
  nor_x1_sg U4926 ( .A(n4419), .B(n4906), .X(n2651) );
  nor_x1_sg U4927 ( .A(n3163), .B(n4855), .X(n2643) );
  nor_x1_sg U4928 ( .A(n4419), .B(n4900), .X(n2645) );
  nor_x1_sg U4929 ( .A(n3163), .B(n4873), .X(n2754) );
  nor_x1_sg U4930 ( .A(n4419), .B(n5014), .X(n2756) );
  nor_x1_sg U4931 ( .A(n3163), .B(n4872), .X(n2745) );
  nor_x1_sg U4932 ( .A(n4419), .B(n5007), .X(n2747) );
  nor_x1_sg U4933 ( .A(n3163), .B(n4870), .X(n2733) );
  nor_x1_sg U4934 ( .A(n4419), .B(n4996), .X(n2735) );
  nor_x1_sg U4935 ( .A(n3163), .B(n4869), .X(n2727) );
  nor_x1_sg U4936 ( .A(n4419), .B(n4988), .X(n2729) );
  nor_x1_sg U4937 ( .A(n3163), .B(n4867), .X(n2715) );
  nor_x1_sg U4938 ( .A(n4419), .B(n4975), .X(n2717) );
  nor_x1_sg U4939 ( .A(n3163), .B(n4866), .X(n2709) );
  nor_x1_sg U4940 ( .A(n4419), .B(n4969), .X(n2711) );
  nor_x1_sg U4941 ( .A(n3163), .B(n4864), .X(n2697) );
  nor_x1_sg U4942 ( .A(n4419), .B(n4956), .X(n2699) );
  nor_x1_sg U4943 ( .A(n3163), .B(n4863), .X(n2691) );
  nor_x1_sg U4944 ( .A(n4419), .B(n4949), .X(n2693) );
  nor_x1_sg U4945 ( .A(n3163), .B(n4861), .X(n2679) );
  nor_x1_sg U4946 ( .A(n4419), .B(n4935), .X(n2681) );
  nor_x1_sg U4947 ( .A(n3163), .B(n4860), .X(n2673) );
  nor_x1_sg U4948 ( .A(n4419), .B(n4929), .X(n2675) );
  nor_x1_sg U4949 ( .A(n3163), .B(n4859), .X(n2667) );
  nor_x1_sg U4950 ( .A(n4419), .B(n4922), .X(n2669) );
  nor_x1_sg U4951 ( .A(n3163), .B(n4858), .X(n2661) );
  nor_x1_sg U4952 ( .A(n4419), .B(n4916), .X(n2663) );
  nor_x1_sg U4953 ( .A(n3163), .B(n4857), .X(n2655) );
  nor_x1_sg U4954 ( .A(n4419), .B(n4910), .X(n2657) );
  nor_x1_sg U4955 ( .A(n3062), .B(n4861), .X(n1956) );
  nor_x1_sg U4956 ( .A(n4935), .B(n4424), .X(n1958) );
  nor_x1_sg U4957 ( .A(n3062), .B(n4859), .X(n1934) );
  nor_x1_sg U4958 ( .A(n4922), .B(n4424), .X(n1936) );
  nor_x1_sg U4959 ( .A(n3163), .B(n4871), .X(n2739) );
  nor_x1_sg U4960 ( .A(n4419), .B(n5001), .X(n2741) );
  nor_x1_sg U4961 ( .A(n3163), .B(n4868), .X(n2721) );
  nor_x1_sg U4962 ( .A(n4419), .B(n4982), .X(n2723) );
  nor_x1_sg U4963 ( .A(n3163), .B(n4865), .X(n2703) );
  nor_x1_sg U4964 ( .A(n4419), .B(n4962), .X(n2705) );
  nor_x1_sg U4965 ( .A(n3163), .B(n4862), .X(n2685) );
  nor_x1_sg U4966 ( .A(n4419), .B(n4943), .X(n2687) );
  nor_x1_sg U4967 ( .A(n3071), .B(n4872), .X(n2340) );
  nor_x1_sg U4968 ( .A(n5007), .B(n4414), .X(n2342) );
  nor_x1_sg U4969 ( .A(n3062), .B(n4872), .X(n2027) );
  nor_x1_sg U4970 ( .A(n5007), .B(n4424), .X(n2029) );
  nor_x1_sg U4971 ( .A(n3062), .B(n4871), .X(n2041) );
  nor_x1_sg U4972 ( .A(n5001), .B(n4424), .X(n2043) );
  nor_x1_sg U4973 ( .A(n3062), .B(n4870), .X(n2035) );
  nor_x1_sg U4974 ( .A(n4996), .B(n4424), .X(n2037) );
  nor_x1_sg U4975 ( .A(n3062), .B(n4869), .X(n1995) );
  nor_x1_sg U4976 ( .A(n4988), .B(n4424), .X(n1997) );
  nor_x1_sg U4977 ( .A(n3062), .B(n4867), .X(n2002) );
  nor_x1_sg U4978 ( .A(n4975), .B(n4424), .X(n2004) );
  nor_x1_sg U4979 ( .A(n3062), .B(n4862), .X(n1963) );
  nor_x1_sg U4980 ( .A(n4943), .B(n4424), .X(n1965) );
  nor_x1_sg U4981 ( .A(n3062), .B(n4855), .X(n1916) );
  nor_x1_sg U4982 ( .A(n4900), .B(n4424), .X(n1918) );
  nor_x1_sg U4983 ( .A(n3071), .B(n4868), .X(n2308) );
  nor_x1_sg U4984 ( .A(n4982), .B(n4414), .X(n2310) );
  nor_x1_sg U4985 ( .A(n3071), .B(n4854), .X(n2229) );
  nor_x1_sg U4986 ( .A(n4894), .B(n4414), .X(n2231) );
  nor_x1_sg U4987 ( .A(n1885), .B(n1742), .X(n1884) );
  nand_x2_sg U4988 ( .A(n4810), .B(n1732), .X(n1854) );
  nand_x2_sg U4989 ( .A(n4808), .B(n1786), .X(n1852) );
  nor_x1_sg U4990 ( .A(n4094), .B(n2168), .X(n2159) );
  nor_x1_sg U4991 ( .A(n1874), .B(n1875), .X(n1872) );
  nand_x2_sg U4992 ( .A(n1886), .B(n1887), .X(n1876) );
  nand_x2_sg U4993 ( .A(n1878), .B(n1879), .X(n1877) );
  nor_x1_sg U4994 ( .A(n2455), .B(n2459), .X(n2583) );
  nand_x1_sg U4995 ( .A(n1750), .B(n4804), .X(n1898) );
  nand_x1_sg U4996 ( .A(n2557), .B(n2554), .X(n2624) );
  nor_x1_sg U4997 ( .A(n4407), .B(n2434), .X(n2433) );
  nand_x2_sg U4998 ( .A(n2080), .B(n4847), .X(n2165) );
  nand_x1_sg U4999 ( .A(n2120), .B(n4840), .X(n2195) );
  nand_x1_sg U5000 ( .A(n1764), .B(n4807), .X(n1998) );
  nor_x1_sg U5001 ( .A(n3162), .B(n4892), .X(n2746) );
  nor_x1_sg U5002 ( .A(n3162), .B(n4887), .X(n2716) );
  nor_x1_sg U5003 ( .A(n3162), .B(n4886), .X(n2710) );
  nor_x1_sg U5004 ( .A(n3162), .B(n4884), .X(n2698) );
  nor_x1_sg U5005 ( .A(n3162), .B(n4883), .X(n2692) );
  nor_x1_sg U5006 ( .A(n3162), .B(n4881), .X(n2680) );
  nor_x1_sg U5007 ( .A(n3162), .B(n4880), .X(n2674) );
  nor_x1_sg U5008 ( .A(n3162), .B(n4879), .X(n2668) );
  nor_x1_sg U5009 ( .A(n3162), .B(n4878), .X(n2662) );
  nor_x1_sg U5010 ( .A(n3162), .B(n4877), .X(n2656) );
  nor_x1_sg U5011 ( .A(n3162), .B(n4891), .X(n2740) );
  nor_x1_sg U5012 ( .A(n3162), .B(n4888), .X(n2722) );
  nor_x1_sg U5013 ( .A(n3162), .B(n4885), .X(n2704) );
  nor_x1_sg U5014 ( .A(n3162), .B(n4882), .X(n2686) );
  nand_x2_sg U5015 ( .A(n2075), .B(n4835), .X(n2225) );
  nand_x2_sg U5016 ( .A(n1893), .B(n1894), .X(n1892) );
  nand_x2_sg U5017 ( .A(n1870), .B(n1871), .X(n1869) );
  nor_x1_sg U5018 ( .A(n1818), .B(n4805), .X(n1868) );
  nor_x1_sg U5019 ( .A(n3061), .B(n4877), .X(n1929) );
  nor_x1_sg U5020 ( .A(n3070), .B(n4893), .X(n2330) );
  nor_x1_sg U5021 ( .A(n3162), .B(n4889), .X(n2728) );
  nor_x1_sg U5022 ( .A(n3061), .B(n4892), .X(n2028) );
  nor_x1_sg U5023 ( .A(n3061), .B(n4891), .X(n2042) );
  nor_x1_sg U5024 ( .A(n3061), .B(n4890), .X(n2036) );
  nor_x1_sg U5025 ( .A(n3061), .B(n4889), .X(n1996) );
  nor_x1_sg U5026 ( .A(n3061), .B(n4887), .X(n2003) );
  nor_x1_sg U5027 ( .A(n3061), .B(n4882), .X(n1964) );
  nor_x1_sg U5028 ( .A(n3061), .B(n4875), .X(n1917) );
  nor_x1_sg U5029 ( .A(n3070), .B(n4888), .X(n2309) );
  nand_x2_sg U5030 ( .A(n4992), .B(n2473), .X(n2587) );
  nand_x2_sg U5031 ( .A(n2589), .B(n3487), .X(n2588) );
  nand_x2_sg U5032 ( .A(n2125), .B(n4845), .X(n2285) );
  nor_x1_sg U5033 ( .A(n386), .B(n2431), .X(n385) );
  nor_x1_sg U5034 ( .A(n1686), .B(n2431), .X(n390) );
  nor_x1_sg U5035 ( .A(n394), .B(n2431), .X(n393) );
  nor_x1_sg U5036 ( .A(n2212), .B(n3807), .X(n2211) );
  nor_x1_sg U5037 ( .A(n4837), .B(n2070), .X(n2213) );
  nand_x2_sg U5038 ( .A(n3486), .B(n1832), .X(n1831) );
  nor_x1_sg U5039 ( .A(n3809), .B(n1846), .X(n1844) );
  nor_x1_sg U5040 ( .A(n4809), .B(n3505), .X(n1845) );
  nor_x1_sg U5041 ( .A(n2188), .B(n4952), .X(n2186) );
  nand_x2_sg U5042 ( .A(n2200), .B(n2201), .X(n2190) );
  nor_x1_sg U5043 ( .A(n3162), .B(n4875), .X(n2644) );
  nand_x4_sg U5044 ( .A(n2232), .B(n2233), .X(n2105) );
  nor_x1_sg U5045 ( .A(n3813), .B(n3519), .X(n2232) );
  nor_x1_sg U5046 ( .A(n2234), .B(n3517), .X(n2233) );
  nor_x1_sg U5047 ( .A(n3070), .B(n4875), .X(n2236) );
  nand_x4_sg U5048 ( .A(n1901), .B(n1902), .X(n1755) );
  nor_x1_sg U5049 ( .A(n3815), .B(n3523), .X(n1901) );
  nor_x1_sg U5050 ( .A(n1903), .B(n3521), .X(n1902) );
  nor_x1_sg U5051 ( .A(n3061), .B(n4876), .X(n1906) );
  nand_x4_sg U5052 ( .A(n2214), .B(n2215), .X(n2070) );
  nor_x1_sg U5053 ( .A(n3817), .B(n3527), .X(n2214) );
  nor_x1_sg U5054 ( .A(n2216), .B(n3525), .X(n2215) );
  nor_x1_sg U5055 ( .A(n3070), .B(n4876), .X(n2219) );
  nand_x4_sg U5056 ( .A(n1947), .B(n1948), .X(n1813) );
  nor_x1_sg U5057 ( .A(n3819), .B(n3531), .X(n1947) );
  nor_x1_sg U5058 ( .A(n1949), .B(n3529), .X(n1948) );
  nor_x1_sg U5059 ( .A(n3061), .B(n4880), .X(n1951) );
  nand_x4_sg U5060 ( .A(n2253), .B(n2254), .X(n2057) );
  nor_x1_sg U5061 ( .A(n3821), .B(n3535), .X(n2253) );
  nor_x1_sg U5062 ( .A(n2255), .B(n3533), .X(n2254) );
  nor_x1_sg U5063 ( .A(n3070), .B(n4878), .X(n2257) );
  nand_x4_sg U5064 ( .A(n1940), .B(n1941), .X(n1742) );
  nor_x1_sg U5065 ( .A(n3823), .B(n3551), .X(n1940) );
  nor_x1_sg U5066 ( .A(n1942), .B(n3549), .X(n1941) );
  nor_x1_sg U5067 ( .A(n3061), .B(n4878), .X(n1944) );
  nand_x4_sg U5068 ( .A(n1966), .B(n1967), .X(n1818) );
  nor_x1_sg U5069 ( .A(n3825), .B(n3575), .X(n1966) );
  nor_x1_sg U5070 ( .A(n1968), .B(n3573), .X(n1967) );
  nor_x1_sg U5071 ( .A(n3061), .B(n4883), .X(n1970) );
  nand_x4_sg U5072 ( .A(n2299), .B(n2300), .X(n2052) );
  nor_x1_sg U5073 ( .A(n3827), .B(n3607), .X(n2299) );
  nor_x1_sg U5074 ( .A(n2301), .B(n3605), .X(n2300) );
  nor_x1_sg U5075 ( .A(n3070), .B(n4889), .X(n2303) );
  nand_x4_sg U5076 ( .A(n2646), .B(n2647), .X(n2561) );
  nor_x1_sg U5077 ( .A(n3829), .B(n3633), .X(n2646) );
  nor_x1_sg U5078 ( .A(n2648), .B(n3631), .X(n2647) );
  nor_x1_sg U5079 ( .A(n3162), .B(n4876), .X(n2650) );
  nand_x2_sg U5080 ( .A(n4990), .B(n1859), .X(n1858) );
  nand_x2_sg U5081 ( .A(n1998), .B(n1852), .X(n1857) );
  nand_x4_sg U5082 ( .A(n2244), .B(n2245), .X(n2120) );
  nor_x1_sg U5083 ( .A(n3831), .B(n3543), .X(n2244) );
  nor_x1_sg U5084 ( .A(n2246), .B(n3541), .X(n2245) );
  nor_x1_sg U5085 ( .A(n3070), .B(n4879), .X(n2248) );
  nand_x4_sg U5086 ( .A(n2260), .B(n2261), .X(n2117) );
  nor_x1_sg U5087 ( .A(n3833), .B(n3559), .X(n2260) );
  nor_x1_sg U5088 ( .A(n2262), .B(n3557), .X(n2261) );
  nor_x1_sg U5089 ( .A(n3070), .B(n4881), .X(n2264) );
  nand_x4_sg U5090 ( .A(n2286), .B(n2287), .X(n2125) );
  nor_x1_sg U5091 ( .A(n3835), .B(n3571), .X(n2286) );
  nor_x1_sg U5092 ( .A(n2288), .B(n3569), .X(n2287) );
  nor_x1_sg U5093 ( .A(n3070), .B(n4884), .X(n2290) );
  nand_x4_sg U5094 ( .A(n1973), .B(n1974), .X(n1772) );
  nor_x1_sg U5095 ( .A(n3837), .B(n3579), .X(n1973) );
  nor_x1_sg U5096 ( .A(n1975), .B(n3577), .X(n1974) );
  nor_x1_sg U5097 ( .A(n3061), .B(n4885), .X(n1977) );
  nand_x4_sg U5098 ( .A(n1979), .B(n1980), .X(n1810) );
  nor_x1_sg U5099 ( .A(n3839), .B(n3583), .X(n1979) );
  nor_x1_sg U5100 ( .A(n1981), .B(n3581), .X(n1980) );
  nor_x1_sg U5101 ( .A(n3061), .B(n4884), .X(n1983) );
  nand_x4_sg U5102 ( .A(n2005), .B(n2006), .X(n1764) );
  nor_x1_sg U5103 ( .A(n3841), .B(n3587), .X(n2005) );
  nor_x1_sg U5104 ( .A(n2007), .B(n3585), .X(n2006) );
  nor_x1_sg U5105 ( .A(n3061), .B(n4886), .X(n2009) );
  nand_x4_sg U5106 ( .A(n1986), .B(n1987), .X(n1780) );
  nor_x1_sg U5107 ( .A(n3843), .B(n3591), .X(n1986) );
  nor_x1_sg U5108 ( .A(n1988), .B(n3589), .X(n1987) );
  nor_x1_sg U5109 ( .A(n3061), .B(n4888), .X(n1990) );
  nand_x4_sg U5110 ( .A(n2292), .B(n2293), .X(n2087) );
  nor_x1_sg U5111 ( .A(n3845), .B(n3595), .X(n2292) );
  nor_x1_sg U5112 ( .A(n2294), .B(n3593), .X(n2293) );
  nor_x1_sg U5113 ( .A(n3070), .B(n4885), .X(n2296) );
  nand_x4_sg U5114 ( .A(n2318), .B(n2319), .X(n2080) );
  nor_x1_sg U5115 ( .A(n3847), .B(n3603), .X(n2318) );
  nor_x1_sg U5116 ( .A(n2320), .B(n3601), .X(n2319) );
  nor_x1_sg U5117 ( .A(n3070), .B(n4886), .X(n2322) );
  nand_x4_sg U5118 ( .A(n2013), .B(n2014), .X(n1775) );
  nor_x1_sg U5119 ( .A(n3849), .B(n3619), .X(n2013) );
  nor_x1_sg U5120 ( .A(n2015), .B(n3617), .X(n2014) );
  nor_x1_sg U5121 ( .A(n3061), .B(n4893), .X(n2017) );
  nand_x4_sg U5122 ( .A(n2226), .B(n2227), .X(n2075) );
  nor_x1_sg U5123 ( .A(n3851), .B(n3753), .X(n2226) );
  nor_x1_sg U5124 ( .A(n2228), .B(n3751), .X(n2227) );
  nor_x1_sg U5125 ( .A(n3070), .B(n4874), .X(n2230) );
  nand_x4_sg U5126 ( .A(n1854), .B(n1985), .X(n1848) );
  nand_x1_sg U5127 ( .A(n1780), .B(n4809), .X(n1985) );
  nand_x4_sg U5128 ( .A(n2147), .B(n2148), .X(n2146) );
  nor_x1_sg U5129 ( .A(n2149), .B(n2150), .X(n2147) );
  nand_x1_sg U5130 ( .A(n2090), .B(n4853), .X(n2148) );
  nand_x4_sg U5131 ( .A(n2555), .B(n4909), .X(n2553) );
  nand_x1_sg U5132 ( .A(n2557), .B(n3499), .X(n2555) );
  nor_x1_sg U5133 ( .A(n3499), .B(n2557), .X(n2556) );
  nand_x4_sg U5134 ( .A(n2457), .B(n5000), .X(n2454) );
  nand_x1_sg U5135 ( .A(n2459), .B(n3500), .X(n2457) );
  nor_x1_sg U5136 ( .A(n3500), .B(n2459), .X(n2458) );
  inv_x4_sg U5137 ( .A(n4441), .X(n4440) );
  nand_x4_sg U5138 ( .A(n2022), .B(n2023), .X(n1840) );
  nand_x1_sg U5139 ( .A(n1745), .B(n4812), .X(n2022) );
  nand_x1_sg U5140 ( .A(n1826), .B(n4813), .X(n2023) );
  nor_x1_sg U5141 ( .A(n382), .B(n4406), .X(n381) );
  nor_x1_sg U5142 ( .A(n398), .B(n4406), .X(n397) );
  nor_x1_sg U5143 ( .A(n402), .B(n4406), .X(n401) );
  nor_x1_sg U5144 ( .A(n406), .B(n4406), .X(n405) );
  nor_x1_sg U5145 ( .A(n410), .B(n4406), .X(n409) );
  nor_x1_sg U5146 ( .A(n414), .B(n4406), .X(n413) );
  nor_x1_sg U5147 ( .A(n418), .B(n4406), .X(n417) );
  nor_x1_sg U5148 ( .A(n422), .B(n4406), .X(n421) );
  nor_x1_sg U5149 ( .A(n426), .B(n4406), .X(n425) );
  nor_x1_sg U5150 ( .A(n430), .B(n4406), .X(n429) );
  nor_x1_sg U5151 ( .A(n434), .B(n4406), .X(n433) );
  nor_x1_sg U5152 ( .A(n438), .B(n4406), .X(n437) );
  nor_x1_sg U5153 ( .A(n442), .B(n4406), .X(n441) );
  nor_x1_sg U5154 ( .A(n446), .B(n4406), .X(n445) );
  nor_x1_sg U5155 ( .A(n450), .B(n4406), .X(n449) );
  nor_x1_sg U5156 ( .A(n454), .B(n4406), .X(n453) );
  nor_x1_sg U5157 ( .A(n458), .B(n4406), .X(n457) );
  nor_x1_sg U5158 ( .A(n462), .B(n4406), .X(n461) );
  nor_x1_sg U5159 ( .A(n466), .B(n4406), .X(n465) );
  nor_x1_sg U5160 ( .A(n470), .B(n4406), .X(n469) );
  nor_x1_sg U5161 ( .A(n378), .B(n4406), .X(n377) );
  nor_x1_sg U5162 ( .A(n4415), .B(n1709), .X(\mean_pooling_0/n230 ) );
  nand_x4_sg U5163 ( .A(n2751), .B(n2752), .X(n2750) );
  nor_x1_sg U5164 ( .A(n3853), .B(n3641), .X(n2751) );
  nor_x1_sg U5165 ( .A(n2753), .B(n3639), .X(n2752) );
  nor_x1_sg U5166 ( .A(n3162), .B(n4893), .X(n2755) );
  nand_x2_sg U5167 ( .A(n4895), .B(n1912), .X(n1911) );
  nand_x1_sg U5168 ( .A(n1783), .B(n4803), .X(n1912) );
  nand_x4_sg U5169 ( .A(n2460), .B(n2461), .X(n1727) );
  nand_x1_sg U5170 ( .A(n2462), .B(n4999), .X(n2461) );
  nand_x4_sg U5171 ( .A(n5019), .B(n2574), .X(n1717) );
  nand_x1_sg U5172 ( .A(n4081), .B(n4086), .X(n2574) );
  nor_x1_sg U5173 ( .A(n4086), .B(n4081), .X(n2577) );
  nor_x1_sg U5174 ( .A(n1937), .B(n3879), .X(n1888) );
  nor_x1_sg U5175 ( .A(n1885), .B(n1890), .X(n1889) );
  nand_x4_sg U5176 ( .A(n1919), .B(n1920), .X(n1767) );
  nor_x1_sg U5177 ( .A(n3855), .B(n3515), .X(n1919) );
  nor_x1_sg U5178 ( .A(n1921), .B(n3513), .X(n1920) );
  nor_x1_sg U5179 ( .A(n3061), .B(n4874), .X(n1923) );
  nand_x4_sg U5180 ( .A(n2238), .B(n2239), .X(n2065) );
  nor_x1_sg U5181 ( .A(n3857), .B(n3539), .X(n2238) );
  nor_x1_sg U5182 ( .A(n2240), .B(n3537), .X(n2239) );
  nor_x1_sg U5183 ( .A(n3070), .B(n4877), .X(n2242) );
  nand_x4_sg U5184 ( .A(n2266), .B(n2267), .X(n2128) );
  nor_x1_sg U5185 ( .A(n3859), .B(n3555), .X(n2266) );
  nor_x1_sg U5186 ( .A(n2268), .B(n3553), .X(n2267) );
  nor_x1_sg U5187 ( .A(n3070), .B(n4880), .X(n2270) );
  nand_x4_sg U5188 ( .A(n2273), .B(n2274), .X(n2110) );
  nor_x1_sg U5189 ( .A(n3861), .B(n3563), .X(n2273) );
  nor_x1_sg U5190 ( .A(n2275), .B(n3561), .X(n2274) );
  nor_x1_sg U5191 ( .A(n3070), .B(n4882), .X(n2277) );
  nand_x4_sg U5192 ( .A(n2279), .B(n2280), .X(n2133) );
  nor_x1_sg U5193 ( .A(n3863), .B(n3567), .X(n2279) );
  nor_x1_sg U5194 ( .A(n2281), .B(n3565), .X(n2280) );
  nor_x1_sg U5195 ( .A(n3070), .B(n4883), .X(n2283) );
  nand_x4_sg U5196 ( .A(n2312), .B(n2313), .X(n2102) );
  nor_x1_sg U5197 ( .A(n3865), .B(n3599), .X(n2312) );
  nor_x1_sg U5198 ( .A(n2314), .B(n3597), .X(n2313) );
  nor_x1_sg U5199 ( .A(n3070), .B(n4887), .X(n2316) );
  nand_x4_sg U5200 ( .A(n2351), .B(n2352), .X(n2060) );
  nor_x1_sg U5201 ( .A(n3867), .B(n3611), .X(n2351) );
  nor_x1_sg U5202 ( .A(n2353), .B(n3609), .X(n2352) );
  nor_x1_sg U5203 ( .A(n3070), .B(n4891), .X(n2355) );
  nand_x4_sg U5204 ( .A(n2345), .B(n2346), .X(n2138) );
  nor_x1_sg U5205 ( .A(n3869), .B(n3615), .X(n2345) );
  nor_x1_sg U5206 ( .A(n2347), .B(n3613), .X(n2346) );
  nor_x1_sg U5207 ( .A(n3070), .B(n4890), .X(n2349) );
  nand_x4_sg U5208 ( .A(n2730), .B(n2731), .X(n2463) );
  nor_x1_sg U5209 ( .A(n3871), .B(n3649), .X(n2730) );
  nor_x1_sg U5210 ( .A(n2732), .B(n3647), .X(n2731) );
  nor_x1_sg U5211 ( .A(n3162), .B(n4890), .X(n2734) );
  nand_x4_sg U5212 ( .A(n1953), .B(n1954), .X(n1802) );
  nor_x1_sg U5213 ( .A(n3873), .B(n3693), .X(n1953) );
  nor_x1_sg U5214 ( .A(n1955), .B(n3691), .X(n1954) );
  nor_x1_sg U5215 ( .A(n3061), .B(n4881), .X(n1957) );
  nand_x4_sg U5216 ( .A(n1931), .B(n1932), .X(n1805) );
  nor_x1_sg U5217 ( .A(n3875), .B(n3697), .X(n1931) );
  nor_x1_sg U5218 ( .A(n1933), .B(n3695), .X(n1932) );
  nor_x1_sg U5219 ( .A(n3061), .B(n4879), .X(n1935) );
  nand_x4_sg U5220 ( .A(n2337), .B(n2338), .X(n2143) );
  nor_x1_sg U5221 ( .A(n3877), .B(n3717), .X(n2337) );
  nor_x1_sg U5222 ( .A(n2339), .B(n3715), .X(n2338) );
  nor_x1_sg U5223 ( .A(n3070), .B(n4892), .X(n2341) );
  nand_x4_sg U5224 ( .A(n2446), .B(n5012), .X(n1695) );
  nor_x1_sg U5225 ( .A(n2448), .B(n2449), .X(n2447) );
  nand_x4_sg U5226 ( .A(n2481), .B(n4979), .X(n1699) );
  nor_x1_sg U5227 ( .A(n2483), .B(n2484), .X(n2482) );
  nand_x4_sg U5228 ( .A(n2488), .B(n4972), .X(n1725) );
  nor_x1_sg U5229 ( .A(n2490), .B(n2491), .X(n2489) );
  nand_x4_sg U5230 ( .A(n2502), .B(n4959), .X(n1711) );
  nor_x1_sg U5231 ( .A(n2504), .B(n2505), .X(n2503) );
  nand_x4_sg U5232 ( .A(n2509), .B(n4953), .X(n1703) );
  nor_x1_sg U5233 ( .A(n2511), .B(n2512), .X(n2510) );
  nand_x4_sg U5234 ( .A(n2523), .B(n4940), .X(n1729) );
  nor_x1_sg U5235 ( .A(n2525), .B(n2526), .X(n2524) );
  nand_x4_sg U5236 ( .A(n2530), .B(n4932), .X(n1701) );
  nor_x1_sg U5237 ( .A(n2532), .B(n2533), .X(n2531) );
  nand_x4_sg U5238 ( .A(n2537), .B(n4926), .X(n1707) );
  nor_x1_sg U5239 ( .A(n2539), .B(n2540), .X(n2538) );
  nand_x4_sg U5240 ( .A(n2544), .B(n4919), .X(n1693) );
  nor_x1_sg U5241 ( .A(n2546), .B(n2547), .X(n2545) );
  nand_x4_sg U5242 ( .A(n2467), .B(n4993), .X(n1691) );
  nor_x1_sg U5243 ( .A(n2469), .B(n2470), .X(n2468) );
  nand_x4_sg U5244 ( .A(n4914), .B(n2623), .X(n2550) );
  nand_x1_sg U5245 ( .A(n2624), .B(n3499), .X(n2623) );
  nor_x1_sg U5246 ( .A(n2554), .B(n2557), .X(n2625) );
  nand_x4_sg U5247 ( .A(n2558), .B(n2559), .X(n1705) );
  nand_x1_sg U5248 ( .A(n2560), .B(n4079), .X(n2559) );
  nand_x2_sg U5249 ( .A(n1866), .B(n1867), .X(n1865) );
  nand_x1_sg U5250 ( .A(n1810), .B(n4806), .X(n1866) );
  nand_x2_sg U5251 ( .A(n2192), .B(n2193), .X(n2191) );
  nand_x1_sg U5252 ( .A(n2117), .B(n4842), .X(n2192) );
  nand_x2_sg U5253 ( .A(n5009), .B(n1839), .X(n1838) );
  nand_x1_sg U5254 ( .A(n4811), .B(n1821), .X(n1839) );
  nand_x4_sg U5255 ( .A(n4920), .B(n2620), .X(n2543) );
  nand_x1_sg U5256 ( .A(n4915), .B(n2547), .X(n2621) );
  nand_x4_sg U5257 ( .A(n4927), .B(n2617), .X(n2536) );
  nand_x1_sg U5258 ( .A(n4921), .B(n2540), .X(n2618) );
  nand_x4_sg U5259 ( .A(n4933), .B(n2614), .X(n2529) );
  nand_x1_sg U5260 ( .A(n4928), .B(n2533), .X(n2615) );
  nand_x4_sg U5261 ( .A(n4941), .B(n2611), .X(n2522) );
  nand_x1_sg U5262 ( .A(n4934), .B(n2526), .X(n2612) );
  nand_x4_sg U5263 ( .A(n4954), .B(n2605), .X(n2508) );
  nand_x1_sg U5264 ( .A(n4948), .B(n2512), .X(n2606) );
  nand_x4_sg U5265 ( .A(n4960), .B(n2602), .X(n2501) );
  nand_x1_sg U5266 ( .A(n4955), .B(n2505), .X(n2603) );
  nand_x4_sg U5267 ( .A(n4973), .B(n2596), .X(n2487) );
  nand_x1_sg U5268 ( .A(n4968), .B(n2491), .X(n2597) );
  nand_x4_sg U5269 ( .A(n4980), .B(n2593), .X(n2480) );
  nand_x1_sg U5270 ( .A(n4974), .B(n2484), .X(n2594) );
  nand_x2_sg U5271 ( .A(n1841), .B(n1842), .X(n1837) );
  nor_x1_sg U5272 ( .A(n1855), .B(n1856), .X(n1843) );
  nor_x1_sg U5273 ( .A(n2176), .B(n2177), .X(n2174) );
  nand_x1_sg U5274 ( .A(n2087), .B(n4846), .X(n2175) );
  nand_x1_sg U5275 ( .A(n4438), .B(n4849), .X(n2091) );
  nand_x1_sg U5276 ( .A(n4442), .B(n4911), .X(n1747) );
  nand_x1_sg U5277 ( .A(n4434), .B(n4804), .X(n1746) );
  nand_x1_sg U5278 ( .A(n4438), .B(n4853), .X(n2071) );
  nand_x1_sg U5279 ( .A(n4436), .B(n4078), .X(n2045) );
  nand_x1_sg U5280 ( .A(n4438), .B(n4850), .X(n2044) );
  nand_x1_sg U5281 ( .A(n4436), .B(n4918), .X(n2054) );
  nand_x1_sg U5282 ( .A(n4438), .B(n4839), .X(n2053) );
  nand_x1_sg U5283 ( .A(n4436), .B(n4908), .X(n2067) );
  nand_x1_sg U5284 ( .A(n4438), .B(n4837), .X(n2066) );
  nand_x1_sg U5285 ( .A(n4436), .B(n4090), .X(n2097) );
  nand_x1_sg U5286 ( .A(n4438), .B(n4836), .X(n2096) );
  nand_x1_sg U5287 ( .A(n1733), .B(n4813), .X(n1824) );
  nand_x1_sg U5288 ( .A(n4434), .B(n4812), .X(n1829) );
  nand_x1_sg U5289 ( .A(n4434), .B(n4811), .X(n1819) );
  nand_x1_sg U5290 ( .A(n4434), .B(n4810), .X(n1730) );
  nand_x1_sg U5291 ( .A(n4442), .B(n4983), .X(n1777) );
  nand_x1_sg U5292 ( .A(n4434), .B(n4809), .X(n1776) );
  nand_x1_sg U5293 ( .A(n4434), .B(n4808), .X(n1784) );
  nand_x1_sg U5294 ( .A(n4442), .B(n4970), .X(n1761) );
  nand_x1_sg U5295 ( .A(n4434), .B(n4807), .X(n1760) );
  nand_x1_sg U5296 ( .A(n4442), .B(n4957), .X(n1807) );
  nand_x1_sg U5297 ( .A(n4434), .B(n4806), .X(n1806) );
  nand_x1_sg U5298 ( .A(n4434), .B(n4803), .X(n1781) );
  nand_x1_sg U5299 ( .A(n4438), .B(n4847), .X(n2076) );
  nand_x1_sg U5300 ( .A(n4438), .B(n4846), .X(n2083) );
  nand_x1_sg U5301 ( .A(n4438), .B(n4845), .X(n2121) );
  nand_x1_sg U5302 ( .A(n4438), .B(n4842), .X(n2113) );
  nand_x1_sg U5303 ( .A(n4438), .B(n4840), .X(n2111) );
  nand_x1_sg U5304 ( .A(n4442), .B(n5015), .X(n1757) );
  nand_x1_sg U5305 ( .A(n4434), .B(n4814), .X(n1756) );
  nor_x1_sg U5306 ( .A(n4925), .B(n2204), .X(n2203) );
  nor_x1_sg U5307 ( .A(n3507), .B(n2199), .X(n2202) );
  nand_x1_sg U5308 ( .A(n4442), .B(n4950), .X(n1815) );
  nand_x1_sg U5309 ( .A(n4434), .B(n4805), .X(n1814) );
  nand_x1_sg U5310 ( .A(n4436), .B(n5003), .X(n2145) );
  nand_x1_sg U5311 ( .A(n4438), .B(n4852), .X(n2144) );
  nand_x1_sg U5312 ( .A(n4436), .B(n4998), .X(n2135) );
  nand_x1_sg U5313 ( .A(n4438), .B(n4851), .X(n2134) );
  nand_x1_sg U5314 ( .A(n4436), .B(n4977), .X(n2099) );
  nand_x1_sg U5315 ( .A(n4438), .B(n4848), .X(n2098) );
  nand_x1_sg U5316 ( .A(n4436), .B(n4951), .X(n2130) );
  nand_x1_sg U5317 ( .A(n4438), .B(n4844), .X(n2129) );
  nand_x1_sg U5318 ( .A(n4436), .B(n4945), .X(n2107) );
  nand_x1_sg U5319 ( .A(n4438), .B(n4843), .X(n2106) );
  nand_x1_sg U5320 ( .A(n4436), .B(n4931), .X(n2049) );
  nand_x1_sg U5321 ( .A(n4438), .B(n4841), .X(n2048) );
  nand_x1_sg U5322 ( .A(n4436), .B(n4912), .X(n2062) );
  nand_x1_sg U5323 ( .A(n4438), .B(n4838), .X(n2061) );
  nand_x1_sg U5324 ( .A(n4438), .B(n4835), .X(n2073) );
  nand_x1_sg U5325 ( .A(n4434), .B(n4375), .X(n1768) );
  nand_x1_sg U5326 ( .A(n4434), .B(n4373), .X(n1791) );
  nand_x1_sg U5327 ( .A(n4442), .B(n4895), .X(n1759) );
  nand_x1_sg U5328 ( .A(n4434), .B(n4088), .X(n1758) );
  nand_x2_sg U5329 ( .A(n3329), .B(output_taken), .X(n3328) );
  nor_x1_sg U5330 ( .A(state[0]), .B(n5026), .X(n3329) );
  nand_x2_sg U5331 ( .A(n5022), .B(input_ready), .X(n3326) );
  nand_x1_sg U5332 ( .A(n4449), .B(n4126), .X(n3219) );
  nand_x1_sg U5333 ( .A(n4449), .B(n4124), .X(n3221) );
  nand_x1_sg U5334 ( .A(n4449), .B(n4222), .X(n3223) );
  nand_x1_sg U5335 ( .A(n4449), .B(n4190), .X(n3225) );
  nand_x1_sg U5336 ( .A(n4449), .B(n4188), .X(n3227) );
  nand_x1_sg U5337 ( .A(n4449), .B(n4186), .X(n3229) );
  nand_x1_sg U5338 ( .A(n4449), .B(n4184), .X(n3231) );
  nand_x1_sg U5339 ( .A(n4449), .B(n4220), .X(n3233) );
  nand_x1_sg U5340 ( .A(n4449), .B(n4218), .X(n3235) );
  nand_x1_sg U5341 ( .A(n4449), .B(n4216), .X(n3237) );
  nand_x1_sg U5342 ( .A(n4449), .B(n4182), .X(n3239) );
  nand_x1_sg U5343 ( .A(n4449), .B(n4214), .X(n3241) );
  nand_x1_sg U5344 ( .A(n4449), .B(n4212), .X(n3243) );
  nand_x1_sg U5345 ( .A(n4449), .B(n4180), .X(n3245) );
  nand_x1_sg U5346 ( .A(n4449), .B(n4176), .X(n3247) );
  nand_x1_sg U5347 ( .A(n4449), .B(n4242), .X(n3249) );
  nand_x1_sg U5348 ( .A(n4449), .B(n4172), .X(n3251) );
  nand_x1_sg U5349 ( .A(n4449), .B(n4240), .X(n3253) );
  nand_x1_sg U5350 ( .A(n4449), .B(n4210), .X(n3255) );
  nand_x1_sg U5351 ( .A(n4449), .B(n4208), .X(n3257) );
  nand_x1_sg U5352 ( .A(n4449), .B(n4206), .X(n3259) );
  nand_x1_sg U5353 ( .A(n4449), .B(n4204), .X(n3261) );
  nand_x1_sg U5354 ( .A(n4449), .B(n4258), .X(n3199) );
  nand_x1_sg U5355 ( .A(n4449), .B(n4246), .X(n3201) );
  nand_x1_sg U5356 ( .A(n4449), .B(n4244), .X(n3203) );
  nand_x1_sg U5357 ( .A(n4449), .B(n4324), .X(n3205) );
  nand_x1_sg U5358 ( .A(n4449), .B(n4174), .X(n3207) );
  nand_x1_sg U5359 ( .A(n4449), .B(n4226), .X(n3209) );
  nand_x1_sg U5360 ( .A(n4449), .B(n4170), .X(n3211) );
  nand_x1_sg U5361 ( .A(n4449), .B(n4224), .X(n3213) );
  nand_x1_sg U5362 ( .A(n4449), .B(n4178), .X(n3215) );
  nand_x1_sg U5363 ( .A(n4449), .B(n4144), .X(n3217) );
  nand_x1_sg U5364 ( .A(n4449), .B(n4238), .X(n3263) );
  nand_x1_sg U5365 ( .A(n4449), .B(n4202), .X(n3265) );
  nand_x1_sg U5366 ( .A(n4449), .B(n4200), .X(n3267) );
  nand_x1_sg U5367 ( .A(n4449), .B(n4198), .X(n3269) );
  nand_x1_sg U5368 ( .A(n4449), .B(n4196), .X(n3271) );
  nand_x1_sg U5369 ( .A(n4449), .B(n4236), .X(n3273) );
  nand_x1_sg U5370 ( .A(n4449), .B(n4234), .X(n3275) );
  nand_x1_sg U5371 ( .A(n4449), .B(n4232), .X(n3277) );
  nand_x1_sg U5372 ( .A(n4449), .B(n4194), .X(n3279) );
  nand_x1_sg U5373 ( .A(n4449), .B(n4230), .X(n3281) );
  nand_x1_sg U5374 ( .A(n4449), .B(n4228), .X(n3283) );
  nand_x1_sg U5375 ( .A(n4449), .B(n4192), .X(n3285) );
  nand_x1_sg U5376 ( .A(n4449), .B(n4158), .X(n3287) );
  nand_x1_sg U5377 ( .A(n4449), .B(n4142), .X(n3289) );
  nand_x1_sg U5378 ( .A(n4449), .B(n4168), .X(n3291) );
  nand_x1_sg U5379 ( .A(n4449), .B(n4140), .X(n3293) );
  nand_x1_sg U5380 ( .A(n4449), .B(n4164), .X(n3295) );
  nand_x1_sg U5381 ( .A(n4449), .B(n4156), .X(n3297) );
  nand_x1_sg U5382 ( .A(n4449), .B(n4166), .X(n3299) );
  nand_x1_sg U5383 ( .A(n4449), .B(n4162), .X(n3301) );
  nand_x1_sg U5384 ( .A(n4449), .B(n4138), .X(n3303) );
  nand_x1_sg U5385 ( .A(n4449), .B(n4154), .X(n3305) );
  nand_x1_sg U5386 ( .A(n4449), .B(n4152), .X(n3307) );
  nand_x1_sg U5387 ( .A(n4449), .B(n4150), .X(n3309) );
  nand_x1_sg U5388 ( .A(n4449), .B(n4148), .X(n3311) );
  nand_x1_sg U5389 ( .A(n4449), .B(n4136), .X(n3313) );
  nand_x1_sg U5390 ( .A(n4449), .B(n4134), .X(n3315) );
  nand_x1_sg U5391 ( .A(n4449), .B(n4132), .X(n3317) );
  nand_x1_sg U5392 ( .A(n4449), .B(n4146), .X(n3319) );
  nand_x1_sg U5393 ( .A(n4449), .B(n4130), .X(n3321) );
  nand_x1_sg U5394 ( .A(n4449), .B(n4128), .X(n3323) );
  nand_x1_sg U5395 ( .A(n4449), .B(n4160), .X(n3325) );
  nand_x1_sg U5396 ( .A(n4449), .B(n4266), .X(n3165) );
  nand_x1_sg U5397 ( .A(n4449), .B(n4318), .X(n3183) );
  nand_x1_sg U5398 ( .A(n4449), .B(n4322), .X(n3185) );
  nand_x1_sg U5399 ( .A(n4449), .B(n4262), .X(n3187) );
  nand_x1_sg U5400 ( .A(n4451), .B(n4320), .X(n3189) );
  nand_x1_sg U5401 ( .A(n4449), .B(n4260), .X(n3191) );
  nand_x1_sg U5402 ( .A(n4449), .B(n4252), .X(n3193) );
  nand_x1_sg U5403 ( .A(n4451), .B(n4250), .X(n3195) );
  nand_x1_sg U5404 ( .A(n4449), .B(n4248), .X(n3197) );
  nand_x1_sg U5405 ( .A(n4449), .B(n4256), .X(n3169) );
  nand_x1_sg U5406 ( .A(n4449), .B(n4332), .X(n3171) );
  nand_x1_sg U5407 ( .A(n4449), .B(n4254), .X(n3173) );
  nand_x1_sg U5408 ( .A(n4449), .B(n4328), .X(n3175) );
  nand_x1_sg U5409 ( .A(n4449), .B(n4264), .X(n3177) );
  nand_x1_sg U5410 ( .A(n4449), .B(n4330), .X(n3179) );
  nand_x1_sg U5411 ( .A(n4449), .B(n4326), .X(n3181) );
  nand_x1_sg U5412 ( .A(n4316), .B(n4429), .X(n3119) );
  nand_x1_sg U5413 ( .A(n4314), .B(n4429), .X(n3147) );
  nand_x1_sg U5414 ( .A(n4312), .B(n4429), .X(n3131) );
  nand_x1_sg U5415 ( .A(n4310), .B(n4429), .X(n3145) );
  nand_x1_sg U5416 ( .A(n4308), .B(n4429), .X(n3115) );
  nand_x1_sg U5417 ( .A(n4306), .B(n4429), .X(n3135) );
  nand_x1_sg U5418 ( .A(n4304), .B(n4429), .X(n3127) );
  nand_x1_sg U5419 ( .A(n4302), .B(n4429), .X(n3143) );
  nand_x1_sg U5420 ( .A(n4300), .B(n4429), .X(n3121) );
  nand_x1_sg U5421 ( .A(n4298), .B(n4280), .X(n3133) );
  nand_x1_sg U5422 ( .A(n4296), .B(n4429), .X(n3125) );
  nand_x1_sg U5423 ( .A(n4294), .B(n4429), .X(n3141) );
  nand_x1_sg U5424 ( .A(n4292), .B(n4429), .X(n3129) );
  nand_x1_sg U5425 ( .A(n4290), .B(n4429), .X(n3149) );
  nand_x1_sg U5426 ( .A(n4288), .B(n4429), .X(n3123) );
  nand_x1_sg U5427 ( .A(n4122), .B(n4429), .X(n3151) );
  nand_x1_sg U5428 ( .A(n3117), .B(n3500), .X(n3152) );
  nand_x1_sg U5429 ( .A(n4286), .B(n4429), .X(n3139) );
  nand_x1_sg U5430 ( .A(n4284), .B(n4429), .X(n3137) );
  nand_x1_sg U5431 ( .A(n3049), .B(state[0]), .X(n3050) );
  nand_x1_sg U5432 ( .A(n3052), .B(n5022), .X(n3051) );
  nor_x1_sg U5433 ( .A(n3049), .B(n5024), .X(n3052) );
  nand_x1_sg U5434 ( .A(n3433), .B(n4102), .X(n3058) );
  nor_x1_sg U5435 ( .A(n3059), .B(n3060), .X(n3057) );
  nand_x1_sg U5436 ( .A(n3434), .B(n4100), .X(n3067) );
  nor_x1_sg U5437 ( .A(n3068), .B(n3069), .X(n3066) );
  nand_x1_sg U5438 ( .A(n4104), .B(n3435), .X(n3159) );
  nor_x1_sg U5439 ( .A(n3160), .B(n3161), .X(n3158) );
  nand_x1_sg U5440 ( .A(n3049), .B(state[1]), .X(n3047) );
  nand_x1_sg U5441 ( .A(n5022), .B(n4098), .X(n3048) );
  nand_x1_sg U5442 ( .A(n4394), .B(n3433), .X(n3340) );
  nor_x1_sg U5443 ( .A(n3341), .B(n3342), .X(n3339) );
  nand_x1_sg U5444 ( .A(n4396), .B(n3433), .X(n3348) );
  nor_x1_sg U5445 ( .A(n3349), .B(n3350), .X(n3347) );
  nand_x1_sg U5446 ( .A(n4278), .B(n3433), .X(n3352) );
  nor_x1_sg U5447 ( .A(n3353), .B(n3354), .X(n3351) );
  nand_x1_sg U5448 ( .A(n4400), .B(n3433), .X(n3356) );
  nor_x1_sg U5449 ( .A(n3357), .B(n3358), .X(n3355) );
  nand_x1_sg U5450 ( .A(n4398), .B(n3433), .X(n3360) );
  nor_x1_sg U5451 ( .A(n3361), .B(n3362), .X(n3359) );
  nand_x1_sg U5452 ( .A(n4402), .B(n3433), .X(n3408) );
  nor_x1_sg U5453 ( .A(n3409), .B(n3410), .X(n3407) );
  nand_x1_sg U5454 ( .A(n4276), .B(n3433), .X(n3344) );
  nor_x1_sg U5455 ( .A(n3345), .B(n3346), .X(n3343) );
  nand_x1_sg U5456 ( .A(n4378), .B(n3433), .X(n3368) );
  nor_x1_sg U5457 ( .A(n3369), .B(n3370), .X(n3367) );
  nand_x1_sg U5458 ( .A(n4374), .B(n3433), .X(n3364) );
  nor_x1_sg U5459 ( .A(n3365), .B(n3366), .X(n3363) );
  nand_x1_sg U5460 ( .A(n4376), .B(n3433), .X(n3376) );
  nor_x1_sg U5461 ( .A(n3377), .B(n3378), .X(n3375) );
  nand_x1_sg U5462 ( .A(n4340), .B(n3433), .X(n3331) );
  nor_x1_sg U5463 ( .A(n3332), .B(n3333), .X(n3330) );
  nand_x1_sg U5464 ( .A(n4338), .B(n3433), .X(n3336) );
  nor_x1_sg U5465 ( .A(n3337), .B(n3338), .X(n3335) );
  nand_x1_sg U5466 ( .A(n4348), .B(n3433), .X(n3372) );
  nor_x1_sg U5467 ( .A(n3373), .B(n3374), .X(n3371) );
  nand_x1_sg U5468 ( .A(n4350), .B(n3433), .X(n3380) );
  nor_x1_sg U5469 ( .A(n3381), .B(n3382), .X(n3379) );
  nand_x1_sg U5470 ( .A(n4344), .B(n3433), .X(n3384) );
  nor_x1_sg U5471 ( .A(n3385), .B(n3386), .X(n3383) );
  nand_x1_sg U5472 ( .A(n4346), .B(n3433), .X(n3388) );
  nor_x1_sg U5473 ( .A(n3389), .B(n3390), .X(n3387) );
  nand_x1_sg U5474 ( .A(n4342), .B(n3433), .X(n3392) );
  nor_x1_sg U5475 ( .A(n3393), .B(n3394), .X(n3391) );
  nand_x1_sg U5476 ( .A(n4352), .B(n3433), .X(n3396) );
  nor_x1_sg U5477 ( .A(n3397), .B(n3398), .X(n3395) );
  nand_x1_sg U5478 ( .A(n4356), .B(n3433), .X(n3400) );
  nor_x1_sg U5479 ( .A(n3401), .B(n3402), .X(n3399) );
  nand_x1_sg U5480 ( .A(n4268), .B(n3433), .X(n3404) );
  nor_x1_sg U5481 ( .A(n3405), .B(n3406), .X(n3403) );
  nand_x1_sg U5482 ( .A(n3434), .B(n4110), .X(n3093) );
  nand_x1_sg U5483 ( .A(n4431), .B(n5050), .X(n3094) );
  nand_x1_sg U5484 ( .A(n4368), .B(n3434), .X(n3079) );
  nand_x1_sg U5485 ( .A(n4362), .B(n3434), .X(n3085) );
  nand_x1_sg U5486 ( .A(n4354), .B(n3434), .X(n3091) );
  nand_x1_sg U5487 ( .A(n4336), .B(n3434), .X(n3103) );
  nand_x1_sg U5488 ( .A(n4388), .B(n3434), .X(n3073) );
  nand_x1_sg U5489 ( .A(n4390), .B(n3434), .X(n3109) );
  nand_x1_sg U5490 ( .A(n4386), .B(n3434), .X(n3097) );
  nand_x1_sg U5491 ( .A(n4334), .B(n3434), .X(n3089) );
  nand_x1_sg U5492 ( .A(n4392), .B(n3434), .X(n3111) );
  nand_x1_sg U5493 ( .A(n4382), .B(n3434), .X(n3087) );
  nand_x1_sg U5494 ( .A(n4380), .B(n3434), .X(n3095) );
  nand_x1_sg U5495 ( .A(n4384), .B(n3434), .X(n3105) );
  nand_x1_sg U5496 ( .A(n4274), .B(n3434), .X(n3101) );
  nand_x1_sg U5497 ( .A(n4272), .B(n3434), .X(n3075) );
  nand_x1_sg U5498 ( .A(n4366), .B(n3434), .X(n3081) );
  nand_x1_sg U5499 ( .A(n4372), .B(n3434), .X(n3113) );
  nand_x1_sg U5500 ( .A(n4370), .B(n3434), .X(n3099) );
  nand_x1_sg U5501 ( .A(n3433), .B(n4112), .X(n3063) );
  nand_x1_sg U5502 ( .A(n3065), .B(n5052), .X(n3064) );
  nand_x1_sg U5503 ( .A(n3435), .B(n4114), .X(n3155) );
  nand_x1_sg U5504 ( .A(n3157), .B(n5051), .X(n3156) );
  nand_x1_sg U5505 ( .A(n4360), .B(n3434), .X(n3083) );
  nand_x1_sg U5506 ( .A(n4364), .B(n3434), .X(n3107) );
  nand_x1_sg U5507 ( .A(n4358), .B(n3434), .X(n3077) );
  nor_x1_sg U5508 ( .A(n3411), .B(n3412), .X(N112) );
  nand_x1_sg U5509 ( .A(n1895), .B(n4394), .X(n1894) );
  nor_x1_sg U5510 ( .A(n1896), .B(n1755), .X(n1895) );
  nand_x1_sg U5511 ( .A(n4398), .B(n4936), .X(n1878) );
  nand_x1_sg U5512 ( .A(n1946), .B(n4400), .X(n1886) );
  nor_x1_sg U5513 ( .A(n1938), .B(n1813), .X(n1946) );
  nand_x2_sg U5514 ( .A(n4912), .B(n4388), .X(n2210) );
  nand_x1_sg U5515 ( .A(n4945), .B(n4380), .X(n2187) );
  nand_x1_sg U5516 ( .A(n1959), .B(n4374), .X(n1870) );
  nor_x1_sg U5517 ( .A(n1875), .B(n1793), .X(n1959) );
  nand_x2_sg U5518 ( .A(n4938), .B(n4362), .X(n2251) );
  nand_x1_sg U5519 ( .A(n1687), .B(n4897), .X(n2572) );
  nand_x2_sg U5520 ( .A(n2207), .B(n2208), .X(n2206) );
  nand_x2_sg U5521 ( .A(n2184), .B(n2185), .X(n2183) );
  nand_x4_sg U5522 ( .A(n1833), .B(n1834), .X(n1832) );
  nor_x1_sg U5523 ( .A(n1835), .B(n1836), .X(n1833) );
  nand_x1_sg U5524 ( .A(n4402), .B(n5015), .X(n1834) );
  nand_x4_sg U5525 ( .A(n2335), .B(n2336), .X(n2154) );
  nand_x1_sg U5526 ( .A(n5003), .B(n4274), .X(n2335) );
  nand_x1_sg U5527 ( .A(n5010), .B(n4392), .X(n2336) );
  nand_x4_sg U5528 ( .A(n2429), .B(n2430), .X(n398) );
  nand_x1_sg U5529 ( .A(n2428), .B(n4272), .X(n2430) );
  nand_x1_sg U5530 ( .A(n4407), .B(n4402), .X(n2429) );
  nand_x4_sg U5531 ( .A(n2426), .B(n2427), .X(n402) );
  nand_x1_sg U5532 ( .A(n4407), .B(n4268), .X(n2426) );
  nand_x1_sg U5533 ( .A(n2428), .B(n4392), .X(n2427) );
  nand_x4_sg U5534 ( .A(n2382), .B(n2383), .X(n446) );
  nor_x1_sg U5535 ( .A(n2384), .B(n2385), .X(n2382) );
  nand_x1_sg U5536 ( .A(n4407), .B(n4398), .X(n2383) );
  nand_x4_sg U5537 ( .A(n2378), .B(n2379), .X(n450) );
  nor_x1_sg U5538 ( .A(n2380), .B(n2381), .X(n2378) );
  nand_x1_sg U5539 ( .A(n4407), .B(n4400), .X(n2379) );
  nand_x4_sg U5540 ( .A(n2374), .B(n2375), .X(n454) );
  nor_x1_sg U5541 ( .A(n2376), .B(n2377), .X(n2374) );
  nand_x1_sg U5542 ( .A(n4407), .B(n4278), .X(n2375) );
  nand_x4_sg U5543 ( .A(n2370), .B(n2371), .X(n458) );
  nor_x1_sg U5544 ( .A(n2372), .B(n2373), .X(n2370) );
  nand_x1_sg U5545 ( .A(n4407), .B(n4396), .X(n2371) );
  nand_x4_sg U5546 ( .A(n2362), .B(n2363), .X(n466) );
  nor_x1_sg U5547 ( .A(n2364), .B(n2365), .X(n2362) );
  nand_x1_sg U5548 ( .A(n4407), .B(n4394), .X(n2363) );
  nor_x1_sg U5549 ( .A(n2169), .B(n2170), .X(n2157) );
  nand_x2_sg U5550 ( .A(n2162), .B(n2173), .X(n2172) );
  nand_x4_sg U5551 ( .A(n2251), .B(n2252), .X(n2199) );
  nand_x1_sg U5552 ( .A(n4931), .B(n4382), .X(n2252) );
  nand_x4_sg U5553 ( .A(n2390), .B(n2391), .X(n438) );
  nor_x1_sg U5554 ( .A(n2392), .B(n2393), .X(n2390) );
  nand_x1_sg U5555 ( .A(n4407), .B(n4378), .X(n2391) );
  nand_x4_sg U5556 ( .A(n2366), .B(n2367), .X(n462) );
  nor_x1_sg U5557 ( .A(n2368), .B(n2369), .X(n2366) );
  nand_x1_sg U5558 ( .A(n4407), .B(n4276), .X(n2367) );
  nand_x1_sg U5559 ( .A(n4434), .B(n4402), .X(n1773) );
  nand_x1_sg U5560 ( .A(n4434), .B(n4398), .X(n1800) );
  nand_x1_sg U5561 ( .A(n4434), .B(n4400), .X(n1811) );
  nand_x1_sg U5562 ( .A(n4434), .B(n4278), .X(n1803) );
  nand_x1_sg U5563 ( .A(n4434), .B(n4396), .X(n1740) );
  nand_x1_sg U5564 ( .A(n4434), .B(n4394), .X(n1753) );
  nand_x1_sg U5565 ( .A(n4438), .B(n4392), .X(n2141) );
  nand_x4_sg U5566 ( .A(n2398), .B(n2399), .X(n430) );
  nor_x1_sg U5567 ( .A(n2400), .B(n2401), .X(n2398) );
  nand_x1_sg U5568 ( .A(n4407), .B(n4376), .X(n2399) );
  nand_x4_sg U5569 ( .A(n2386), .B(n2387), .X(n442) );
  nor_x1_sg U5570 ( .A(n2388), .B(n2389), .X(n2386) );
  nand_x1_sg U5571 ( .A(n4407), .B(n4374), .X(n2387) );
  nand_x2_sg U5572 ( .A(n2311), .B(n2166), .X(n2171) );
  nand_x1_sg U5573 ( .A(n4971), .B(n4358), .X(n2311) );
  nor_x1_sg U5574 ( .A(n4372), .B(n4908), .X(n2209) );
  nor_x1_sg U5575 ( .A(n4380), .B(n4945), .X(n2272) );
  nand_x1_sg U5576 ( .A(n4278), .B(n4923), .X(n1882) );
  nand_x1_sg U5577 ( .A(n1884), .B(n4396), .X(n1883) );
  nand_x2_sg U5578 ( .A(n5011), .B(n2153), .X(n2152) );
  nand_x1_sg U5579 ( .A(n4998), .B(n4384), .X(n2153) );
  nand_x2_sg U5580 ( .A(n2155), .B(n2156), .X(n2151) );
  nand_x1_sg U5581 ( .A(n5016), .B(n4272), .X(n2156) );
  nor_x1_sg U5582 ( .A(n3755), .B(n2160), .X(n2158) );
  nor_x1_sg U5583 ( .A(n4382), .B(n4931), .X(n2259) );
  nor_x1_sg U5584 ( .A(n1862), .B(n1863), .X(n1860) );
  nand_x1_sg U5585 ( .A(n4376), .B(n4963), .X(n1861) );
  nand_x4_sg U5586 ( .A(n4986), .B(n2590), .X(n2473) );
  nand_x1_sg U5587 ( .A(n4981), .B(n2476), .X(n2591) );
  nand_x4_sg U5588 ( .A(n2422), .B(n2423), .X(n406) );
  nor_x1_sg U5589 ( .A(n2424), .B(n2425), .X(n2422) );
  nand_x1_sg U5590 ( .A(n4407), .B(n4356), .X(n2423) );
  nand_x4_sg U5591 ( .A(n2418), .B(n2419), .X(n410) );
  nor_x1_sg U5592 ( .A(n2420), .B(n2421), .X(n2418) );
  nand_x1_sg U5593 ( .A(n4407), .B(n4352), .X(n2419) );
  nand_x4_sg U5594 ( .A(n2414), .B(n2415), .X(n414) );
  nor_x1_sg U5595 ( .A(n3509), .B(n2417), .X(n2414) );
  nand_x1_sg U5596 ( .A(n4407), .B(n4342), .X(n2415) );
  nand_x4_sg U5597 ( .A(n2410), .B(n2411), .X(n418) );
  nor_x1_sg U5598 ( .A(n2412), .B(n2413), .X(n2410) );
  nand_x1_sg U5599 ( .A(n4407), .B(n4346), .X(n2411) );
  nand_x4_sg U5600 ( .A(n2406), .B(n2407), .X(n422) );
  nor_x1_sg U5601 ( .A(n2408), .B(n2409), .X(n2406) );
  nand_x1_sg U5602 ( .A(n4407), .B(n4344), .X(n2407) );
  nand_x4_sg U5603 ( .A(n2402), .B(n2403), .X(n426) );
  nor_x1_sg U5604 ( .A(n2404), .B(n2405), .X(n2402) );
  nand_x1_sg U5605 ( .A(n4407), .B(n4350), .X(n2403) );
  nand_x4_sg U5606 ( .A(n2394), .B(n2395), .X(n434) );
  nor_x1_sg U5607 ( .A(n2396), .B(n2397), .X(n2394) );
  nand_x1_sg U5608 ( .A(n4407), .B(n4348), .X(n2395) );
  nand_x4_sg U5609 ( .A(n2358), .B(n2359), .X(n470) );
  nor_x1_sg U5610 ( .A(n3511), .B(n2361), .X(n2358) );
  nand_x1_sg U5611 ( .A(n4407), .B(n4338), .X(n2359) );
  nand_x4_sg U5612 ( .A(n2442), .B(n2443), .X(n378) );
  nor_x1_sg U5613 ( .A(n2444), .B(n2445), .X(n2442) );
  nand_x1_sg U5614 ( .A(n4407), .B(n4340), .X(n2443) );
  nor_x1_sg U5615 ( .A(n3434), .B(n4414), .X(\max_pooling_0/n314 ) );
  nand_x1_sg U5616 ( .A(n4434), .B(n4378), .X(n1816) );
  nand_x1_sg U5617 ( .A(n4434), .B(n4276), .X(n1748) );
  nand_x1_sg U5618 ( .A(n4438), .B(n4274), .X(n2058) );
  nand_x1_sg U5619 ( .A(n4438), .B(n4384), .X(n2136) );
  nand_x1_sg U5620 ( .A(n4438), .B(n4386), .X(n2100) );
  nand_x1_sg U5621 ( .A(n4438), .B(n4390), .X(n2131) );
  nand_x1_sg U5622 ( .A(n4438), .B(n4380), .X(n2108) );
  nand_x1_sg U5623 ( .A(n4438), .B(n4382), .X(n2126) );
  nand_x1_sg U5624 ( .A(n4438), .B(n4388), .X(n2063) );
  nand_x1_sg U5625 ( .A(n4434), .B(n4376), .X(n1770) );
  nand_x1_sg U5626 ( .A(n4434), .B(n4374), .X(n1794) );
  nand_x1_sg U5627 ( .A(n4438), .B(n4272), .X(n2088) );
  nand_x2_sg U5628 ( .A(n2180), .B(n2181), .X(n2179) );
  nand_x1_sg U5629 ( .A(n4958), .B(n4354), .X(n2180) );
  nor_x1_sg U5630 ( .A(n3435), .B(n4419), .X(\mean_pooling_0/n226 ) );
  nor_x1_sg U5631 ( .A(n4368), .B(n4918), .X(n2197) );
  nand_x4_sg U5632 ( .A(n2569), .B(n2570), .X(n2567) );
  nand_x1_sg U5633 ( .A(n2571), .B(n3503), .X(n2569) );
  nand_x1_sg U5634 ( .A(n1688), .B(n4898), .X(n2570) );
  nand_x4_sg U5635 ( .A(n2541), .B(n2542), .X(n2539) );
  nand_x1_sg U5636 ( .A(n4921), .B(n3488), .X(n2541) );
  nand_x4_sg U5637 ( .A(n2485), .B(n2486), .X(n2483) );
  nand_x1_sg U5638 ( .A(n4974), .B(n3489), .X(n2485) );
  nand_x4_sg U5639 ( .A(n2492), .B(n2493), .X(n2490) );
  nand_x1_sg U5640 ( .A(n4968), .B(n3490), .X(n2492) );
  nand_x4_sg U5641 ( .A(n2506), .B(n2507), .X(n2504) );
  nand_x1_sg U5642 ( .A(n4955), .B(n3491), .X(n2506) );
  nand_x4_sg U5643 ( .A(n2513), .B(n2514), .X(n2511) );
  nand_x1_sg U5644 ( .A(n4948), .B(n3492), .X(n2513) );
  nand_x4_sg U5645 ( .A(n2527), .B(n2528), .X(n2525) );
  nand_x1_sg U5646 ( .A(n4934), .B(n3493), .X(n2527) );
  nand_x4_sg U5647 ( .A(n2534), .B(n2535), .X(n2532) );
  nand_x1_sg U5648 ( .A(n4928), .B(n3494), .X(n2534) );
  nand_x4_sg U5649 ( .A(n2478), .B(n2479), .X(n2475) );
  nand_x1_sg U5650 ( .A(n4981), .B(n3495), .X(n2478) );
  nand_x4_sg U5651 ( .A(n2499), .B(n2500), .X(n2496) );
  nand_x1_sg U5652 ( .A(n4961), .B(n3496), .X(n2499) );
  nand_x4_sg U5653 ( .A(n2520), .B(n2521), .X(n2517) );
  nand_x1_sg U5654 ( .A(n4942), .B(n3497), .X(n2520) );
  nand_x4_sg U5655 ( .A(n2450), .B(n2451), .X(n2448) );
  nand_x1_sg U5656 ( .A(n5006), .B(n3502), .X(n2450) );
  nand_x4_sg U5657 ( .A(n2548), .B(n2549), .X(n2546) );
  nand_x1_sg U5658 ( .A(n4915), .B(n3498), .X(n2548) );
  nand_x1_sg U5659 ( .A(n4438), .B(n4370), .X(n2050) );
  nand_x1_sg U5660 ( .A(n4438), .B(n4368), .X(n2055) );
  nand_x1_sg U5661 ( .A(n4438), .B(n4372), .X(n2068) );
  nand_x1_sg U5662 ( .A(n4438), .B(n4366), .X(n2103) );
  nand_x4_sg U5663 ( .A(n5005), .B(n2581), .X(n2452) );
  nand_x1_sg U5664 ( .A(n2459), .B(n2455), .X(n2582) );
  nand_x4_sg U5665 ( .A(n2471), .B(n2472), .X(n2469) );
  nand_x1_sg U5666 ( .A(n4987), .B(n3487), .X(n2471) );
  nand_x1_sg U5667 ( .A(n4434), .B(n4268), .X(n1827) );
  nand_x1_sg U5668 ( .A(n4434), .B(n4356), .X(n1743) );
  nand_x1_sg U5669 ( .A(n4434), .B(n4352), .X(n1822) );
  nand_x1_sg U5670 ( .A(n4434), .B(n4342), .X(n1736) );
  nand_x1_sg U5671 ( .A(n4434), .B(n4346), .X(n1778) );
  nand_x1_sg U5672 ( .A(n4434), .B(n4344), .X(n1787) );
  nand_x1_sg U5673 ( .A(n4434), .B(n4350), .X(n1762) );
  nand_x1_sg U5674 ( .A(n4434), .B(n4348), .X(n1808) );
  nand_x1_sg U5675 ( .A(n4434), .B(n4338), .X(n1789) );
  nand_x1_sg U5676 ( .A(n4434), .B(n4340), .X(n1765) );
  nand_x1_sg U5677 ( .A(n4438), .B(n4358), .X(n2078) );
  nand_x1_sg U5678 ( .A(n4438), .B(n4364), .X(n2085) );
  nand_x1_sg U5679 ( .A(n4438), .B(n4354), .X(n2123) );
  nand_x1_sg U5680 ( .A(n4438), .B(n4362), .X(n2115) );
  nand_x1_sg U5681 ( .A(n4438), .B(n4360), .X(n2118) );
  nand_x4_sg U5682 ( .A(n4947), .B(n2608), .X(n2515) );
  nand_x1_sg U5683 ( .A(n4942), .B(n2518), .X(n2609) );
  nand_x4_sg U5684 ( .A(n4967), .B(n2599), .X(n2494) );
  nand_x1_sg U5685 ( .A(n4961), .B(n2497), .X(n2600) );
  nand_x4_sg U5686 ( .A(n2437), .B(n2438), .X(n382) );
  nor_x1_sg U5687 ( .A(n2439), .B(n2440), .X(n2437) );
  nor_x1_sg U5688 ( .A(n3435), .B(n4418), .X(\mean_pooling_0/n225 ) );
  nor_x1_sg U5689 ( .A(n3434), .B(n4413), .X(\max_pooling_0/n313 ) );
  nand_x1_sg U5690 ( .A(n4438), .B(n4336), .X(n2094) );
  nand_x1_sg U5691 ( .A(n4438), .B(n4334), .X(n2081) );
  nand_x1_sg U5692 ( .A(n4442), .B(n4936), .X(n1799) );
  nand_x1_sg U5693 ( .A(n4442), .B(n4930), .X(n1735) );
  nand_x1_sg U5694 ( .A(n4442), .B(n4923), .X(n1797) );
  nand_x1_sg U5695 ( .A(n4442), .B(n4917), .X(n1739) );
  nand_x1_sg U5696 ( .A(n4442), .B(n4907), .X(n1752) );
  nand_x1_sg U5697 ( .A(n4436), .B(n5010), .X(n2140) );
  inv_x8_sg U5698 ( .A(n4405), .X(n4406) );
  inv_x8_sg U5699 ( .A(n2436), .X(n4407) );
  inv_x8_sg U5700 ( .A(n2434), .X(n4408) );
  inv_x8_sg U5701 ( .A(n4409), .X(n4410) );
  nand_x8_sg U5702 ( .A(n5050), .B(n4834), .X(n4411) );
  nand_x8_sg U5703 ( .A(n5050), .B(n4834), .X(n4412) );
  inv_x8_sg U5704 ( .A(n2221), .X(n4413) );
  inv_x8_sg U5705 ( .A(n4413), .X(n4414) );
  inv_x8_sg U5706 ( .A(n3157), .X(n4415) );
  nand_x8_sg U5707 ( .A(n5051), .B(n4815), .X(n4416) );
  nand_x8_sg U5708 ( .A(n5051), .B(n4815), .X(n4417) );
  inv_x8_sg U5709 ( .A(n2573), .X(n4418) );
  inv_x8_sg U5710 ( .A(n4418), .X(n4419) );
  nand_x8_sg U5711 ( .A(n4433), .B(n3485), .X(n4420) );
  nand_x8_sg U5712 ( .A(n5052), .B(n4801), .X(n4421) );
  nand_x8_sg U5713 ( .A(n5052), .B(n4801), .X(n4422) );
  inv_x8_sg U5714 ( .A(n1908), .X(n4423) );
  inv_x8_sg U5715 ( .A(n4423), .X(n4424) );
  inv_x8_sg U5716 ( .A(n3065), .X(n4425) );
  nand_x8_sg U5717 ( .A(n4433), .B(n3486), .X(n4426) );
  nand_x8_sg U5718 ( .A(n4433), .B(n3486), .X(n4427) );
  inv_x8_sg U5719 ( .A(n4428), .X(n4429) );
  nor_x8_sg U5720 ( .A(n4433), .B(n4429), .X(n3117) );
  nor_x8_sg U5721 ( .A(n4433), .B(n3434), .X(n4430) );
  nor_x8_sg U5722 ( .A(n4433), .B(n3434), .X(n4431) );
  nor_x8_sg U5723 ( .A(n4433), .B(n3434), .X(n3072) );
  inv_x8_sg U5724 ( .A(n4432), .X(n4433) );
  inv_x8_sg U5725 ( .A(n4435), .X(n4434) );
  inv_x8_sg U5726 ( .A(n4437), .X(n4436) );
  inv_x8_sg U5727 ( .A(n4439), .X(n4438) );
  inv_x8_sg U5728 ( .A(n4443), .X(n4442) );
  inv_x8_sg U5729 ( .A(n4446), .X(n4445) );
  inv_x8_sg U5730 ( .A(n4448), .X(n4447) );
  inv_x4_sg U5731 ( .A(n3167), .X(n4448) );
  inv_x8_sg U5732 ( .A(n4450), .X(n4449) );
  inv_x2_sg U6081 ( .A(n4316), .X(n4816) );
  inv_x2_sg U6082 ( .A(n4314), .X(n4817) );
  inv_x2_sg U6083 ( .A(n4312), .X(n4818) );
  inv_x2_sg U6084 ( .A(n4310), .X(n4819) );
  inv_x2_sg U6085 ( .A(n4308), .X(n4820) );
  inv_x2_sg U6086 ( .A(n4306), .X(n4821) );
  inv_x2_sg U6087 ( .A(n4304), .X(n4822) );
  inv_x2_sg U6088 ( .A(n4302), .X(n4823) );
  inv_x2_sg U6089 ( .A(n4300), .X(n4824) );
  inv_x2_sg U6090 ( .A(n4298), .X(n4825) );
  inv_x2_sg U6091 ( .A(n4296), .X(n4826) );
  inv_x2_sg U6092 ( .A(n4294), .X(n4827) );
  inv_x2_sg U6093 ( .A(n4292), .X(n4828) );
  inv_x2_sg U6094 ( .A(n4290), .X(n4829) );
  inv_x2_sg U6095 ( .A(n4288), .X(n4830) );
  inv_x2_sg U6096 ( .A(n4122), .X(n4831) );
  inv_x2_sg U6097 ( .A(n4286), .X(n4832) );
  inv_x2_sg U6098 ( .A(n4284), .X(n4833) );
  inv_x2_sg U6099 ( .A(n2090), .X(n5016) );
  inv_x2_sg U6100 ( .A(n4082), .X(n4991) );
  inv_x2_sg U6101 ( .A(n2166), .X(n4978) );
  inv_x2_sg U6102 ( .A(n2125), .X(n4958) );
  inv_x2_sg U6103 ( .A(n2189), .X(n4952) );
  inv_x2_sg U6104 ( .A(n2120), .X(n4924) );
  inv_x2_sg U6105 ( .A(n4106), .X(n4925) );
  inv_x2_sg U6106 ( .A(n2117), .X(n4938) );
  inv_x2_sg U6107 ( .A(n2181), .X(n4965) );
  inv_x2_sg U6108 ( .A(n2080), .X(n4971) );
  inv_x2_sg U6109 ( .A(n2567), .X(n4899) );
  inv_x2_sg U6110 ( .A(n2519), .X(n4946) );
  inv_x2_sg U6111 ( .A(n2498), .X(n4966) );
  inv_x2_sg U6112 ( .A(n2477), .X(n4985) );
  inv_x2_sg U6113 ( .A(n2465), .X(n4994) );
  inv_x2_sg U6114 ( .A(n2456), .X(n5004) );
  inv_x2_sg U6115 ( .A(n2580), .X(n5013) );
  inv_x2_sg U6116 ( .A(n2473), .X(n4987) );
  inv_x2_sg U6117 ( .A(n2749), .X(n5018) );
  inv_x2_sg U6118 ( .A(n4402), .X(n4814) );
  inv_x2_sg U6119 ( .A(n1764), .X(n4970) );
  inv_x2_sg U6120 ( .A(n1780), .X(n4983) );
  inv_x2_sg U6121 ( .A(n1772), .X(n4963) );
  inv_x2_sg U6122 ( .A(n1767), .X(n4895) );
  inv_x2_sg U6123 ( .A(n1810), .X(n4957) );
  inv_x2_sg U6124 ( .A(n3053), .X(n5024) );
  inv_x2_sg U6125 ( .A(state[0]), .X(n5027) );
  inv_x2_sg U6126 ( .A(n3154), .X(n5028) );
  inv_x2_sg U6127 ( .A(n3072), .X(n5029) );
endmodule

