
module transposer ( clk, reset, input_ready, output_taken, state, .in({
        \in[3][3][19] , \in[3][3][18] , \in[3][3][17] , \in[3][3][16] , 
        \in[3][3][15] , \in[3][3][14] , \in[3][3][13] , \in[3][3][12] , 
        \in[3][3][11] , \in[3][3][10] , \in[3][3][9] , \in[3][3][8] , 
        \in[3][3][7] , \in[3][3][6] , \in[3][3][5] , \in[3][3][4] , 
        \in[3][3][3] , \in[3][3][2] , \in[3][3][1] , \in[3][3][0] , 
        \in[3][2][19] , \in[3][2][18] , \in[3][2][17] , \in[3][2][16] , 
        \in[3][2][15] , \in[3][2][14] , \in[3][2][13] , \in[3][2][12] , 
        \in[3][2][11] , \in[3][2][10] , \in[3][2][9] , \in[3][2][8] , 
        \in[3][2][7] , \in[3][2][6] , \in[3][2][5] , \in[3][2][4] , 
        \in[3][2][3] , \in[3][2][2] , \in[3][2][1] , \in[3][2][0] , 
        \in[3][1][19] , \in[3][1][18] , \in[3][1][17] , \in[3][1][16] , 
        \in[3][1][15] , \in[3][1][14] , \in[3][1][13] , \in[3][1][12] , 
        \in[3][1][11] , \in[3][1][10] , \in[3][1][9] , \in[3][1][8] , 
        \in[3][1][7] , \in[3][1][6] , \in[3][1][5] , \in[3][1][4] , 
        \in[3][1][3] , \in[3][1][2] , \in[3][1][1] , \in[3][1][0] , 
        \in[3][0][19] , \in[3][0][18] , \in[3][0][17] , \in[3][0][16] , 
        \in[3][0][15] , \in[3][0][14] , \in[3][0][13] , \in[3][0][12] , 
        \in[3][0][11] , \in[3][0][10] , \in[3][0][9] , \in[3][0][8] , 
        \in[3][0][7] , \in[3][0][6] , \in[3][0][5] , \in[3][0][4] , 
        \in[3][0][3] , \in[3][0][2] , \in[3][0][1] , \in[3][0][0] , 
        \in[2][3][19] , \in[2][3][18] , \in[2][3][17] , \in[2][3][16] , 
        \in[2][3][15] , \in[2][3][14] , \in[2][3][13] , \in[2][3][12] , 
        \in[2][3][11] , \in[2][3][10] , \in[2][3][9] , \in[2][3][8] , 
        \in[2][3][7] , \in[2][3][6] , \in[2][3][5] , \in[2][3][4] , 
        \in[2][3][3] , \in[2][3][2] , \in[2][3][1] , \in[2][3][0] , 
        \in[2][2][19] , \in[2][2][18] , \in[2][2][17] , \in[2][2][16] , 
        \in[2][2][15] , \in[2][2][14] , \in[2][2][13] , \in[2][2][12] , 
        \in[2][2][11] , \in[2][2][10] , \in[2][2][9] , \in[2][2][8] , 
        \in[2][2][7] , \in[2][2][6] , \in[2][2][5] , \in[2][2][4] , 
        \in[2][2][3] , \in[2][2][2] , \in[2][2][1] , \in[2][2][0] , 
        \in[2][1][19] , \in[2][1][18] , \in[2][1][17] , \in[2][1][16] , 
        \in[2][1][15] , \in[2][1][14] , \in[2][1][13] , \in[2][1][12] , 
        \in[2][1][11] , \in[2][1][10] , \in[2][1][9] , \in[2][1][8] , 
        \in[2][1][7] , \in[2][1][6] , \in[2][1][5] , \in[2][1][4] , 
        \in[2][1][3] , \in[2][1][2] , \in[2][1][1] , \in[2][1][0] , 
        \in[2][0][19] , \in[2][0][18] , \in[2][0][17] , \in[2][0][16] , 
        \in[2][0][15] , \in[2][0][14] , \in[2][0][13] , \in[2][0][12] , 
        \in[2][0][11] , \in[2][0][10] , \in[2][0][9] , \in[2][0][8] , 
        \in[2][0][7] , \in[2][0][6] , \in[2][0][5] , \in[2][0][4] , 
        \in[2][0][3] , \in[2][0][2] , \in[2][0][1] , \in[2][0][0] , 
        \in[1][3][19] , \in[1][3][18] , \in[1][3][17] , \in[1][3][16] , 
        \in[1][3][15] , \in[1][3][14] , \in[1][3][13] , \in[1][3][12] , 
        \in[1][3][11] , \in[1][3][10] , \in[1][3][9] , \in[1][3][8] , 
        \in[1][3][7] , \in[1][3][6] , \in[1][3][5] , \in[1][3][4] , 
        \in[1][3][3] , \in[1][3][2] , \in[1][3][1] , \in[1][3][0] , 
        \in[1][2][19] , \in[1][2][18] , \in[1][2][17] , \in[1][2][16] , 
        \in[1][2][15] , \in[1][2][14] , \in[1][2][13] , \in[1][2][12] , 
        \in[1][2][11] , \in[1][2][10] , \in[1][2][9] , \in[1][2][8] , 
        \in[1][2][7] , \in[1][2][6] , \in[1][2][5] , \in[1][2][4] , 
        \in[1][2][3] , \in[1][2][2] , \in[1][2][1] , \in[1][2][0] , 
        \in[1][1][19] , \in[1][1][18] , \in[1][1][17] , \in[1][1][16] , 
        \in[1][1][15] , \in[1][1][14] , \in[1][1][13] , \in[1][1][12] , 
        \in[1][1][11] , \in[1][1][10] , \in[1][1][9] , \in[1][1][8] , 
        \in[1][1][7] , \in[1][1][6] , \in[1][1][5] , \in[1][1][4] , 
        \in[1][1][3] , \in[1][1][2] , \in[1][1][1] , \in[1][1][0] , 
        \in[1][0][19] , \in[1][0][18] , \in[1][0][17] , \in[1][0][16] , 
        \in[1][0][15] , \in[1][0][14] , \in[1][0][13] , \in[1][0][12] , 
        \in[1][0][11] , \in[1][0][10] , \in[1][0][9] , \in[1][0][8] , 
        \in[1][0][7] , \in[1][0][6] , \in[1][0][5] , \in[1][0][4] , 
        \in[1][0][3] , \in[1][0][2] , \in[1][0][1] , \in[1][0][0] , 
        \in[0][3][19] , \in[0][3][18] , \in[0][3][17] , \in[0][3][16] , 
        \in[0][3][15] , \in[0][3][14] , \in[0][3][13] , \in[0][3][12] , 
        \in[0][3][11] , \in[0][3][10] , \in[0][3][9] , \in[0][3][8] , 
        \in[0][3][7] , \in[0][3][6] , \in[0][3][5] , \in[0][3][4] , 
        \in[0][3][3] , \in[0][3][2] , \in[0][3][1] , \in[0][3][0] , 
        \in[0][2][19] , \in[0][2][18] , \in[0][2][17] , \in[0][2][16] , 
        \in[0][2][15] , \in[0][2][14] , \in[0][2][13] , \in[0][2][12] , 
        \in[0][2][11] , \in[0][2][10] , \in[0][2][9] , \in[0][2][8] , 
        \in[0][2][7] , \in[0][2][6] , \in[0][2][5] , \in[0][2][4] , 
        \in[0][2][3] , \in[0][2][2] , \in[0][2][1] , \in[0][2][0] , 
        \in[0][1][19] , \in[0][1][18] , \in[0][1][17] , \in[0][1][16] , 
        \in[0][1][15] , \in[0][1][14] , \in[0][1][13] , \in[0][1][12] , 
        \in[0][1][11] , \in[0][1][10] , \in[0][1][9] , \in[0][1][8] , 
        \in[0][1][7] , \in[0][1][6] , \in[0][1][5] , \in[0][1][4] , 
        \in[0][1][3] , \in[0][1][2] , \in[0][1][1] , \in[0][1][0] , 
        \in[0][0][19] , \in[0][0][18] , \in[0][0][17] , \in[0][0][16] , 
        \in[0][0][15] , \in[0][0][14] , \in[0][0][13] , \in[0][0][12] , 
        \in[0][0][11] , \in[0][0][10] , \in[0][0][9] , \in[0][0][8] , 
        \in[0][0][7] , \in[0][0][6] , \in[0][0][5] , \in[0][0][4] , 
        \in[0][0][3] , \in[0][0][2] , \in[0][0][1] , \in[0][0][0] }), .out({
        \out[3][3][19] , \out[3][3][18] , \out[3][3][17] , \out[3][3][16] , 
        \out[3][3][15] , \out[3][3][14] , \out[3][3][13] , \out[3][3][12] , 
        \out[3][3][11] , \out[3][3][10] , \out[3][3][9] , \out[3][3][8] , 
        \out[3][3][7] , \out[3][3][6] , \out[3][3][5] , \out[3][3][4] , 
        \out[3][3][3] , \out[3][3][2] , \out[3][3][1] , \out[3][3][0] , 
        \out[3][2][19] , \out[3][2][18] , \out[3][2][17] , \out[3][2][16] , 
        \out[3][2][15] , \out[3][2][14] , \out[3][2][13] , \out[3][2][12] , 
        \out[3][2][11] , \out[3][2][10] , \out[3][2][9] , \out[3][2][8] , 
        \out[3][2][7] , \out[3][2][6] , \out[3][2][5] , \out[3][2][4] , 
        \out[3][2][3] , \out[3][2][2] , \out[3][2][1] , \out[3][2][0] , 
        \out[3][1][19] , \out[3][1][18] , \out[3][1][17] , \out[3][1][16] , 
        \out[3][1][15] , \out[3][1][14] , \out[3][1][13] , \out[3][1][12] , 
        \out[3][1][11] , \out[3][1][10] , \out[3][1][9] , \out[3][1][8] , 
        \out[3][1][7] , \out[3][1][6] , \out[3][1][5] , \out[3][1][4] , 
        \out[3][1][3] , \out[3][1][2] , \out[3][1][1] , \out[3][1][0] , 
        \out[3][0][19] , \out[3][0][18] , \out[3][0][17] , \out[3][0][16] , 
        \out[3][0][15] , \out[3][0][14] , \out[3][0][13] , \out[3][0][12] , 
        \out[3][0][11] , \out[3][0][10] , \out[3][0][9] , \out[3][0][8] , 
        \out[3][0][7] , \out[3][0][6] , \out[3][0][5] , \out[3][0][4] , 
        \out[3][0][3] , \out[3][0][2] , \out[3][0][1] , \out[3][0][0] , 
        \out[2][3][19] , \out[2][3][18] , \out[2][3][17] , \out[2][3][16] , 
        \out[2][3][15] , \out[2][3][14] , \out[2][3][13] , \out[2][3][12] , 
        \out[2][3][11] , \out[2][3][10] , \out[2][3][9] , \out[2][3][8] , 
        \out[2][3][7] , \out[2][3][6] , \out[2][3][5] , \out[2][3][4] , 
        \out[2][3][3] , \out[2][3][2] , \out[2][3][1] , \out[2][3][0] , 
        \out[2][2][19] , \out[2][2][18] , \out[2][2][17] , \out[2][2][16] , 
        \out[2][2][15] , \out[2][2][14] , \out[2][2][13] , \out[2][2][12] , 
        \out[2][2][11] , \out[2][2][10] , \out[2][2][9] , \out[2][2][8] , 
        \out[2][2][7] , \out[2][2][6] , \out[2][2][5] , \out[2][2][4] , 
        \out[2][2][3] , \out[2][2][2] , \out[2][2][1] , \out[2][2][0] , 
        \out[2][1][19] , \out[2][1][18] , \out[2][1][17] , \out[2][1][16] , 
        \out[2][1][15] , \out[2][1][14] , \out[2][1][13] , \out[2][1][12] , 
        \out[2][1][11] , \out[2][1][10] , \out[2][1][9] , \out[2][1][8] , 
        \out[2][1][7] , \out[2][1][6] , \out[2][1][5] , \out[2][1][4] , 
        \out[2][1][3] , \out[2][1][2] , \out[2][1][1] , \out[2][1][0] , 
        \out[2][0][19] , \out[2][0][18] , \out[2][0][17] , \out[2][0][16] , 
        \out[2][0][15] , \out[2][0][14] , \out[2][0][13] , \out[2][0][12] , 
        \out[2][0][11] , \out[2][0][10] , \out[2][0][9] , \out[2][0][8] , 
        \out[2][0][7] , \out[2][0][6] , \out[2][0][5] , \out[2][0][4] , 
        \out[2][0][3] , \out[2][0][2] , \out[2][0][1] , \out[2][0][0] , 
        \out[1][3][19] , \out[1][3][18] , \out[1][3][17] , \out[1][3][16] , 
        \out[1][3][15] , \out[1][3][14] , \out[1][3][13] , \out[1][3][12] , 
        \out[1][3][11] , \out[1][3][10] , \out[1][3][9] , \out[1][3][8] , 
        \out[1][3][7] , \out[1][3][6] , \out[1][3][5] , \out[1][3][4] , 
        \out[1][3][3] , \out[1][3][2] , \out[1][3][1] , \out[1][3][0] , 
        \out[1][2][19] , \out[1][2][18] , \out[1][2][17] , \out[1][2][16] , 
        \out[1][2][15] , \out[1][2][14] , \out[1][2][13] , \out[1][2][12] , 
        \out[1][2][11] , \out[1][2][10] , \out[1][2][9] , \out[1][2][8] , 
        \out[1][2][7] , \out[1][2][6] , \out[1][2][5] , \out[1][2][4] , 
        \out[1][2][3] , \out[1][2][2] , \out[1][2][1] , \out[1][2][0] , 
        \out[1][1][19] , \out[1][1][18] , \out[1][1][17] , \out[1][1][16] , 
        \out[1][1][15] , \out[1][1][14] , \out[1][1][13] , \out[1][1][12] , 
        \out[1][1][11] , \out[1][1][10] , \out[1][1][9] , \out[1][1][8] , 
        \out[1][1][7] , \out[1][1][6] , \out[1][1][5] , \out[1][1][4] , 
        \out[1][1][3] , \out[1][1][2] , \out[1][1][1] , \out[1][1][0] , 
        \out[1][0][19] , \out[1][0][18] , \out[1][0][17] , \out[1][0][16] , 
        \out[1][0][15] , \out[1][0][14] , \out[1][0][13] , \out[1][0][12] , 
        \out[1][0][11] , \out[1][0][10] , \out[1][0][9] , \out[1][0][8] , 
        \out[1][0][7] , \out[1][0][6] , \out[1][0][5] , \out[1][0][4] , 
        \out[1][0][3] , \out[1][0][2] , \out[1][0][1] , \out[1][0][0] , 
        \out[0][3][19] , \out[0][3][18] , \out[0][3][17] , \out[0][3][16] , 
        \out[0][3][15] , \out[0][3][14] , \out[0][3][13] , \out[0][3][12] , 
        \out[0][3][11] , \out[0][3][10] , \out[0][3][9] , \out[0][3][8] , 
        \out[0][3][7] , \out[0][3][6] , \out[0][3][5] , \out[0][3][4] , 
        \out[0][3][3] , \out[0][3][2] , \out[0][3][1] , \out[0][3][0] , 
        \out[0][2][19] , \out[0][2][18] , \out[0][2][17] , \out[0][2][16] , 
        \out[0][2][15] , \out[0][2][14] , \out[0][2][13] , \out[0][2][12] , 
        \out[0][2][11] , \out[0][2][10] , \out[0][2][9] , \out[0][2][8] , 
        \out[0][2][7] , \out[0][2][6] , \out[0][2][5] , \out[0][2][4] , 
        \out[0][2][3] , \out[0][2][2] , \out[0][2][1] , \out[0][2][0] , 
        \out[0][1][19] , \out[0][1][18] , \out[0][1][17] , \out[0][1][16] , 
        \out[0][1][15] , \out[0][1][14] , \out[0][1][13] , \out[0][1][12] , 
        \out[0][1][11] , \out[0][1][10] , \out[0][1][9] , \out[0][1][8] , 
        \out[0][1][7] , \out[0][1][6] , \out[0][1][5] , \out[0][1][4] , 
        \out[0][1][3] , \out[0][1][2] , \out[0][1][1] , \out[0][1][0] , 
        \out[0][0][19] , \out[0][0][18] , \out[0][0][17] , \out[0][0][16] , 
        \out[0][0][15] , \out[0][0][14] , \out[0][0][13] , \out[0][0][12] , 
        \out[0][0][11] , \out[0][0][10] , \out[0][0][9] , \out[0][0][8] , 
        \out[0][0][7] , \out[0][0][6] , \out[0][0][5] , \out[0][0][4] , 
        \out[0][0][3] , \out[0][0][2] , \out[0][0][1] , \out[0][0][0] }) );
  output [1:0] state;
  input clk, reset, input_ready, output_taken, \in[3][3][19] , \in[3][3][18] ,
         \in[3][3][17] , \in[3][3][16] , \in[3][3][15] , \in[3][3][14] ,
         \in[3][3][13] , \in[3][3][12] , \in[3][3][11] , \in[3][3][10] ,
         \in[3][3][9] , \in[3][3][8] , \in[3][3][7] , \in[3][3][6] ,
         \in[3][3][5] , \in[3][3][4] , \in[3][3][3] , \in[3][3][2] ,
         \in[3][3][1] , \in[3][3][0] , \in[3][2][19] , \in[3][2][18] ,
         \in[3][2][17] , \in[3][2][16] , \in[3][2][15] , \in[3][2][14] ,
         \in[3][2][13] , \in[3][2][12] , \in[3][2][11] , \in[3][2][10] ,
         \in[3][2][9] , \in[3][2][8] , \in[3][2][7] , \in[3][2][6] ,
         \in[3][2][5] , \in[3][2][4] , \in[3][2][3] , \in[3][2][2] ,
         \in[3][2][1] , \in[3][2][0] , \in[3][1][19] , \in[3][1][18] ,
         \in[3][1][17] , \in[3][1][16] , \in[3][1][15] , \in[3][1][14] ,
         \in[3][1][13] , \in[3][1][12] , \in[3][1][11] , \in[3][1][10] ,
         \in[3][1][9] , \in[3][1][8] , \in[3][1][7] , \in[3][1][6] ,
         \in[3][1][5] , \in[3][1][4] , \in[3][1][3] , \in[3][1][2] ,
         \in[3][1][1] , \in[3][1][0] , \in[3][0][19] , \in[3][0][18] ,
         \in[3][0][17] , \in[3][0][16] , \in[3][0][15] , \in[3][0][14] ,
         \in[3][0][13] , \in[3][0][12] , \in[3][0][11] , \in[3][0][10] ,
         \in[3][0][9] , \in[3][0][8] , \in[3][0][7] , \in[3][0][6] ,
         \in[3][0][5] , \in[3][0][4] , \in[3][0][3] , \in[3][0][2] ,
         \in[3][0][1] , \in[3][0][0] , \in[2][3][19] , \in[2][3][18] ,
         \in[2][3][17] , \in[2][3][16] , \in[2][3][15] , \in[2][3][14] ,
         \in[2][3][13] , \in[2][3][12] , \in[2][3][11] , \in[2][3][10] ,
         \in[2][3][9] , \in[2][3][8] , \in[2][3][7] , \in[2][3][6] ,
         \in[2][3][5] , \in[2][3][4] , \in[2][3][3] , \in[2][3][2] ,
         \in[2][3][1] , \in[2][3][0] , \in[2][2][19] , \in[2][2][18] ,
         \in[2][2][17] , \in[2][2][16] , \in[2][2][15] , \in[2][2][14] ,
         \in[2][2][13] , \in[2][2][12] , \in[2][2][11] , \in[2][2][10] ,
         \in[2][2][9] , \in[2][2][8] , \in[2][2][7] , \in[2][2][6] ,
         \in[2][2][5] , \in[2][2][4] , \in[2][2][3] , \in[2][2][2] ,
         \in[2][2][1] , \in[2][2][0] , \in[2][1][19] , \in[2][1][18] ,
         \in[2][1][17] , \in[2][1][16] , \in[2][1][15] , \in[2][1][14] ,
         \in[2][1][13] , \in[2][1][12] , \in[2][1][11] , \in[2][1][10] ,
         \in[2][1][9] , \in[2][1][8] , \in[2][1][7] , \in[2][1][6] ,
         \in[2][1][5] , \in[2][1][4] , \in[2][1][3] , \in[2][1][2] ,
         \in[2][1][1] , \in[2][1][0] , \in[2][0][19] , \in[2][0][18] ,
         \in[2][0][17] , \in[2][0][16] , \in[2][0][15] , \in[2][0][14] ,
         \in[2][0][13] , \in[2][0][12] , \in[2][0][11] , \in[2][0][10] ,
         \in[2][0][9] , \in[2][0][8] , \in[2][0][7] , \in[2][0][6] ,
         \in[2][0][5] , \in[2][0][4] , \in[2][0][3] , \in[2][0][2] ,
         \in[2][0][1] , \in[2][0][0] , \in[1][3][19] , \in[1][3][18] ,
         \in[1][3][17] , \in[1][3][16] , \in[1][3][15] , \in[1][3][14] ,
         \in[1][3][13] , \in[1][3][12] , \in[1][3][11] , \in[1][3][10] ,
         \in[1][3][9] , \in[1][3][8] , \in[1][3][7] , \in[1][3][6] ,
         \in[1][3][5] , \in[1][3][4] , \in[1][3][3] , \in[1][3][2] ,
         \in[1][3][1] , \in[1][3][0] , \in[1][2][19] , \in[1][2][18] ,
         \in[1][2][17] , \in[1][2][16] , \in[1][2][15] , \in[1][2][14] ,
         \in[1][2][13] , \in[1][2][12] , \in[1][2][11] , \in[1][2][10] ,
         \in[1][2][9] , \in[1][2][8] , \in[1][2][7] , \in[1][2][6] ,
         \in[1][2][5] , \in[1][2][4] , \in[1][2][3] , \in[1][2][2] ,
         \in[1][2][1] , \in[1][2][0] , \in[1][1][19] , \in[1][1][18] ,
         \in[1][1][17] , \in[1][1][16] , \in[1][1][15] , \in[1][1][14] ,
         \in[1][1][13] , \in[1][1][12] , \in[1][1][11] , \in[1][1][10] ,
         \in[1][1][9] , \in[1][1][8] , \in[1][1][7] , \in[1][1][6] ,
         \in[1][1][5] , \in[1][1][4] , \in[1][1][3] , \in[1][1][2] ,
         \in[1][1][1] , \in[1][1][0] , \in[1][0][19] , \in[1][0][18] ,
         \in[1][0][17] , \in[1][0][16] , \in[1][0][15] , \in[1][0][14] ,
         \in[1][0][13] , \in[1][0][12] , \in[1][0][11] , \in[1][0][10] ,
         \in[1][0][9] , \in[1][0][8] , \in[1][0][7] , \in[1][0][6] ,
         \in[1][0][5] , \in[1][0][4] , \in[1][0][3] , \in[1][0][2] ,
         \in[1][0][1] , \in[1][0][0] , \in[0][3][19] , \in[0][3][18] ,
         \in[0][3][17] , \in[0][3][16] , \in[0][3][15] , \in[0][3][14] ,
         \in[0][3][13] , \in[0][3][12] , \in[0][3][11] , \in[0][3][10] ,
         \in[0][3][9] , \in[0][3][8] , \in[0][3][7] , \in[0][3][6] ,
         \in[0][3][5] , \in[0][3][4] , \in[0][3][3] , \in[0][3][2] ,
         \in[0][3][1] , \in[0][3][0] , \in[0][2][19] , \in[0][2][18] ,
         \in[0][2][17] , \in[0][2][16] , \in[0][2][15] , \in[0][2][14] ,
         \in[0][2][13] , \in[0][2][12] , \in[0][2][11] , \in[0][2][10] ,
         \in[0][2][9] , \in[0][2][8] , \in[0][2][7] , \in[0][2][6] ,
         \in[0][2][5] , \in[0][2][4] , \in[0][2][3] , \in[0][2][2] ,
         \in[0][2][1] , \in[0][2][0] , \in[0][1][19] , \in[0][1][18] ,
         \in[0][1][17] , \in[0][1][16] , \in[0][1][15] , \in[0][1][14] ,
         \in[0][1][13] , \in[0][1][12] , \in[0][1][11] , \in[0][1][10] ,
         \in[0][1][9] , \in[0][1][8] , \in[0][1][7] , \in[0][1][6] ,
         \in[0][1][5] , \in[0][1][4] , \in[0][1][3] , \in[0][1][2] ,
         \in[0][1][1] , \in[0][1][0] , \in[0][0][19] , \in[0][0][18] ,
         \in[0][0][17] , \in[0][0][16] , \in[0][0][15] , \in[0][0][14] ,
         \in[0][0][13] , \in[0][0][12] , \in[0][0][11] , \in[0][0][10] ,
         \in[0][0][9] , \in[0][0][8] , \in[0][0][7] , \in[0][0][6] ,
         \in[0][0][5] , \in[0][0][4] , \in[0][0][3] , \in[0][0][2] ,
         \in[0][0][1] , \in[0][0][0] ;
  output \out[3][3][19] , \out[3][3][18] , \out[3][3][17] , \out[3][3][16] ,
         \out[3][3][15] , \out[3][3][14] , \out[3][3][13] , \out[3][3][12] ,
         \out[3][3][11] , \out[3][3][10] , \out[3][3][9] , \out[3][3][8] ,
         \out[3][3][7] , \out[3][3][6] , \out[3][3][5] , \out[3][3][4] ,
         \out[3][3][3] , \out[3][3][2] , \out[3][3][1] , \out[3][3][0] ,
         \out[3][2][19] , \out[3][2][18] , \out[3][2][17] , \out[3][2][16] ,
         \out[3][2][15] , \out[3][2][14] , \out[3][2][13] , \out[3][2][12] ,
         \out[3][2][11] , \out[3][2][10] , \out[3][2][9] , \out[3][2][8] ,
         \out[3][2][7] , \out[3][2][6] , \out[3][2][5] , \out[3][2][4] ,
         \out[3][2][3] , \out[3][2][2] , \out[3][2][1] , \out[3][2][0] ,
         \out[3][1][19] , \out[3][1][18] , \out[3][1][17] , \out[3][1][16] ,
         \out[3][1][15] , \out[3][1][14] , \out[3][1][13] , \out[3][1][12] ,
         \out[3][1][11] , \out[3][1][10] , \out[3][1][9] , \out[3][1][8] ,
         \out[3][1][7] , \out[3][1][6] , \out[3][1][5] , \out[3][1][4] ,
         \out[3][1][3] , \out[3][1][2] , \out[3][1][1] , \out[3][1][0] ,
         \out[3][0][19] , \out[3][0][18] , \out[3][0][17] , \out[3][0][16] ,
         \out[3][0][15] , \out[3][0][14] , \out[3][0][13] , \out[3][0][12] ,
         \out[3][0][11] , \out[3][0][10] , \out[3][0][9] , \out[3][0][8] ,
         \out[3][0][7] , \out[3][0][6] , \out[3][0][5] , \out[3][0][4] ,
         \out[3][0][3] , \out[3][0][2] , \out[3][0][1] , \out[3][0][0] ,
         \out[2][3][19] , \out[2][3][18] , \out[2][3][17] , \out[2][3][16] ,
         \out[2][3][15] , \out[2][3][14] , \out[2][3][13] , \out[2][3][12] ,
         \out[2][3][11] , \out[2][3][10] , \out[2][3][9] , \out[2][3][8] ,
         \out[2][3][7] , \out[2][3][6] , \out[2][3][5] , \out[2][3][4] ,
         \out[2][3][3] , \out[2][3][2] , \out[2][3][1] , \out[2][3][0] ,
         \out[2][2][19] , \out[2][2][18] , \out[2][2][17] , \out[2][2][16] ,
         \out[2][2][15] , \out[2][2][14] , \out[2][2][13] , \out[2][2][12] ,
         \out[2][2][11] , \out[2][2][10] , \out[2][2][9] , \out[2][2][8] ,
         \out[2][2][7] , \out[2][2][6] , \out[2][2][5] , \out[2][2][4] ,
         \out[2][2][3] , \out[2][2][2] , \out[2][2][1] , \out[2][2][0] ,
         \out[2][1][19] , \out[2][1][18] , \out[2][1][17] , \out[2][1][16] ,
         \out[2][1][15] , \out[2][1][14] , \out[2][1][13] , \out[2][1][12] ,
         \out[2][1][11] , \out[2][1][10] , \out[2][1][9] , \out[2][1][8] ,
         \out[2][1][7] , \out[2][1][6] , \out[2][1][5] , \out[2][1][4] ,
         \out[2][1][3] , \out[2][1][2] , \out[2][1][1] , \out[2][1][0] ,
         \out[2][0][19] , \out[2][0][18] , \out[2][0][17] , \out[2][0][16] ,
         \out[2][0][15] , \out[2][0][14] , \out[2][0][13] , \out[2][0][12] ,
         \out[2][0][11] , \out[2][0][10] , \out[2][0][9] , \out[2][0][8] ,
         \out[2][0][7] , \out[2][0][6] , \out[2][0][5] , \out[2][0][4] ,
         \out[2][0][3] , \out[2][0][2] , \out[2][0][1] , \out[2][0][0] ,
         \out[1][3][19] , \out[1][3][18] , \out[1][3][17] , \out[1][3][16] ,
         \out[1][3][15] , \out[1][3][14] , \out[1][3][13] , \out[1][3][12] ,
         \out[1][3][11] , \out[1][3][10] , \out[1][3][9] , \out[1][3][8] ,
         \out[1][3][7] , \out[1][3][6] , \out[1][3][5] , \out[1][3][4] ,
         \out[1][3][3] , \out[1][3][2] , \out[1][3][1] , \out[1][3][0] ,
         \out[1][2][19] , \out[1][2][18] , \out[1][2][17] , \out[1][2][16] ,
         \out[1][2][15] , \out[1][2][14] , \out[1][2][13] , \out[1][2][12] ,
         \out[1][2][11] , \out[1][2][10] , \out[1][2][9] , \out[1][2][8] ,
         \out[1][2][7] , \out[1][2][6] , \out[1][2][5] , \out[1][2][4] ,
         \out[1][2][3] , \out[1][2][2] , \out[1][2][1] , \out[1][2][0] ,
         \out[1][1][19] , \out[1][1][18] , \out[1][1][17] , \out[1][1][16] ,
         \out[1][1][15] , \out[1][1][14] , \out[1][1][13] , \out[1][1][12] ,
         \out[1][1][11] , \out[1][1][10] , \out[1][1][9] , \out[1][1][8] ,
         \out[1][1][7] , \out[1][1][6] , \out[1][1][5] , \out[1][1][4] ,
         \out[1][1][3] , \out[1][1][2] , \out[1][1][1] , \out[1][1][0] ,
         \out[1][0][19] , \out[1][0][18] , \out[1][0][17] , \out[1][0][16] ,
         \out[1][0][15] , \out[1][0][14] , \out[1][0][13] , \out[1][0][12] ,
         \out[1][0][11] , \out[1][0][10] , \out[1][0][9] , \out[1][0][8] ,
         \out[1][0][7] , \out[1][0][6] , \out[1][0][5] , \out[1][0][4] ,
         \out[1][0][3] , \out[1][0][2] , \out[1][0][1] , \out[1][0][0] ,
         \out[0][3][19] , \out[0][3][18] , \out[0][3][17] , \out[0][3][16] ,
         \out[0][3][15] , \out[0][3][14] , \out[0][3][13] , \out[0][3][12] ,
         \out[0][3][11] , \out[0][3][10] , \out[0][3][9] , \out[0][3][8] ,
         \out[0][3][7] , \out[0][3][6] , \out[0][3][5] , \out[0][3][4] ,
         \out[0][3][3] , \out[0][3][2] , \out[0][3][1] , \out[0][3][0] ,
         \out[0][2][19] , \out[0][2][18] , \out[0][2][17] , \out[0][2][16] ,
         \out[0][2][15] , \out[0][2][14] , \out[0][2][13] , \out[0][2][12] ,
         \out[0][2][11] , \out[0][2][10] , \out[0][2][9] , \out[0][2][8] ,
         \out[0][2][7] , \out[0][2][6] , \out[0][2][5] , \out[0][2][4] ,
         \out[0][2][3] , \out[0][2][2] , \out[0][2][1] , \out[0][2][0] ,
         \out[0][1][19] , \out[0][1][18] , \out[0][1][17] , \out[0][1][16] ,
         \out[0][1][15] , \out[0][1][14] , \out[0][1][13] , \out[0][1][12] ,
         \out[0][1][11] , \out[0][1][10] , \out[0][1][9] , \out[0][1][8] ,
         \out[0][1][7] , \out[0][1][6] , \out[0][1][5] , \out[0][1][4] ,
         \out[0][1][3] , \out[0][1][2] , \out[0][1][1] , \out[0][1][0] ,
         \out[0][0][19] , \out[0][0][18] , \out[0][0][17] , \out[0][0][16] ,
         \out[0][0][15] , \out[0][0][14] , \out[0][0][13] , \out[0][0][12] ,
         \out[0][0][11] , \out[0][0][10] , \out[0][0][9] , \out[0][0][8] ,
         \out[0][0][7] , \out[0][0][6] , \out[0][0][5] , \out[0][0][4] ,
         \out[0][0][3] , \out[0][0][2] , \out[0][0][1] , \out[0][0][0] ;
  wire   \reg_in[3][3][19] , \reg_in[3][3][18] , \reg_in[3][3][17] ,
         \reg_in[3][3][16] , \reg_in[3][3][15] , \reg_in[3][3][14] ,
         \reg_in[3][3][13] , \reg_in[3][3][12] , \reg_in[3][3][11] ,
         \reg_in[3][3][10] , \reg_in[3][3][9] , \reg_in[3][3][8] ,
         \reg_in[3][3][7] , \reg_in[3][3][6] , \reg_in[3][3][5] ,
         \reg_in[3][3][4] , \reg_in[3][3][3] , \reg_in[3][3][2] ,
         \reg_in[3][3][1] , \reg_in[3][3][0] , \reg_in[3][2][19] ,
         \reg_in[3][2][18] , \reg_in[3][2][17] , \reg_in[3][2][16] ,
         \reg_in[3][2][15] , \reg_in[3][2][14] , \reg_in[3][2][13] ,
         \reg_in[3][2][12] , \reg_in[3][2][11] , \reg_in[3][2][10] ,
         \reg_in[3][2][9] , \reg_in[3][2][8] , \reg_in[3][2][7] ,
         \reg_in[3][2][6] , \reg_in[3][2][5] , \reg_in[3][2][4] ,
         \reg_in[3][2][3] , \reg_in[3][2][2] , \reg_in[3][2][1] ,
         \reg_in[3][2][0] , \reg_in[3][1][19] , \reg_in[3][1][18] ,
         \reg_in[3][1][17] , \reg_in[3][1][16] , \reg_in[3][1][15] ,
         \reg_in[3][1][14] , \reg_in[3][1][13] , \reg_in[3][1][12] ,
         \reg_in[3][1][11] , \reg_in[3][1][10] , \reg_in[3][1][9] ,
         \reg_in[3][1][8] , \reg_in[3][1][7] , \reg_in[3][1][6] ,
         \reg_in[3][1][5] , \reg_in[3][1][4] , \reg_in[3][1][3] ,
         \reg_in[3][1][2] , \reg_in[3][1][1] , \reg_in[3][1][0] ,
         \reg_in[3][0][19] , \reg_in[3][0][18] , \reg_in[3][0][17] ,
         \reg_in[3][0][16] , \reg_in[3][0][15] , \reg_in[3][0][14] ,
         \reg_in[3][0][13] , \reg_in[3][0][12] , \reg_in[3][0][11] ,
         \reg_in[3][0][10] , \reg_in[3][0][9] , \reg_in[3][0][8] ,
         \reg_in[3][0][7] , \reg_in[3][0][6] , \reg_in[3][0][5] ,
         \reg_in[3][0][4] , \reg_in[3][0][3] , \reg_in[3][0][2] ,
         \reg_in[3][0][1] , \reg_in[3][0][0] , \reg_in[2][3][19] ,
         \reg_in[2][3][18] , \reg_in[2][3][17] , \reg_in[2][3][16] ,
         \reg_in[2][3][15] , \reg_in[2][3][14] , \reg_in[2][3][13] ,
         \reg_in[2][3][12] , \reg_in[2][3][11] , \reg_in[2][3][10] ,
         \reg_in[2][3][9] , \reg_in[2][3][8] , \reg_in[2][3][7] ,
         \reg_in[2][3][6] , \reg_in[2][3][5] , \reg_in[2][3][4] ,
         \reg_in[2][3][3] , \reg_in[2][3][2] , \reg_in[2][3][1] ,
         \reg_in[2][3][0] , \reg_in[2][2][19] , \reg_in[2][2][18] ,
         \reg_in[2][2][17] , \reg_in[2][2][16] , \reg_in[2][2][15] ,
         \reg_in[2][2][14] , \reg_in[2][2][13] , \reg_in[2][2][12] ,
         \reg_in[2][2][11] , \reg_in[2][2][10] , \reg_in[2][2][9] ,
         \reg_in[2][2][8] , \reg_in[2][2][7] , \reg_in[2][2][6] ,
         \reg_in[2][2][5] , \reg_in[2][2][4] , \reg_in[2][2][3] ,
         \reg_in[2][2][2] , \reg_in[2][2][1] , \reg_in[2][2][0] ,
         \reg_in[2][1][19] , \reg_in[2][1][18] , \reg_in[2][1][17] ,
         \reg_in[2][1][16] , \reg_in[2][1][15] , \reg_in[2][1][14] ,
         \reg_in[2][1][13] , \reg_in[2][1][12] , \reg_in[2][1][11] ,
         \reg_in[2][1][10] , \reg_in[2][1][9] , \reg_in[2][1][8] ,
         \reg_in[2][1][7] , \reg_in[2][1][6] , \reg_in[2][1][5] ,
         \reg_in[2][1][4] , \reg_in[2][1][3] , \reg_in[2][1][2] ,
         \reg_in[2][1][1] , \reg_in[2][1][0] , \reg_in[2][0][19] ,
         \reg_in[2][0][18] , \reg_in[2][0][17] , \reg_in[2][0][16] ,
         \reg_in[2][0][15] , \reg_in[2][0][14] , \reg_in[2][0][13] ,
         \reg_in[2][0][12] , \reg_in[2][0][11] , \reg_in[2][0][10] ,
         \reg_in[2][0][9] , \reg_in[2][0][8] , \reg_in[2][0][7] ,
         \reg_in[2][0][6] , \reg_in[2][0][5] , \reg_in[2][0][4] ,
         \reg_in[2][0][3] , \reg_in[2][0][2] , \reg_in[2][0][1] ,
         \reg_in[2][0][0] , \reg_in[1][3][19] , \reg_in[1][3][18] ,
         \reg_in[1][3][17] , \reg_in[1][3][16] , \reg_in[1][3][15] ,
         \reg_in[1][3][14] , \reg_in[1][3][13] , \reg_in[1][3][12] ,
         \reg_in[1][3][11] , \reg_in[1][3][10] , \reg_in[1][3][9] ,
         \reg_in[1][3][8] , \reg_in[1][3][7] , \reg_in[1][3][6] ,
         \reg_in[1][3][5] , \reg_in[1][3][4] , \reg_in[1][3][3] ,
         \reg_in[1][3][2] , \reg_in[1][3][1] , \reg_in[1][3][0] ,
         \reg_in[1][2][19] , \reg_in[1][2][18] , \reg_in[1][2][17] ,
         \reg_in[1][2][16] , \reg_in[1][2][15] , \reg_in[1][2][14] ,
         \reg_in[1][2][13] , \reg_in[1][2][12] , \reg_in[1][2][11] ,
         \reg_in[1][2][10] , \reg_in[1][2][9] , \reg_in[1][2][8] ,
         \reg_in[1][2][7] , \reg_in[1][2][6] , \reg_in[1][2][5] ,
         \reg_in[1][2][4] , \reg_in[1][2][3] , \reg_in[1][2][2] ,
         \reg_in[1][2][1] , \reg_in[1][2][0] , \reg_in[1][1][19] ,
         \reg_in[1][1][18] , \reg_in[1][1][17] , \reg_in[1][1][16] ,
         \reg_in[1][1][15] , \reg_in[1][1][14] , \reg_in[1][1][13] ,
         \reg_in[1][1][12] , \reg_in[1][1][11] , \reg_in[1][1][10] ,
         \reg_in[1][1][9] , \reg_in[1][1][8] , \reg_in[1][1][7] ,
         \reg_in[1][1][6] , \reg_in[1][1][5] , \reg_in[1][1][4] ,
         \reg_in[1][1][3] , \reg_in[1][1][2] , \reg_in[1][1][1] ,
         \reg_in[1][1][0] , \reg_in[1][0][19] , \reg_in[1][0][18] ,
         \reg_in[1][0][17] , \reg_in[1][0][16] , \reg_in[1][0][15] ,
         \reg_in[1][0][14] , \reg_in[1][0][13] , \reg_in[1][0][12] ,
         \reg_in[1][0][11] , \reg_in[1][0][10] , \reg_in[1][0][9] ,
         \reg_in[1][0][8] , \reg_in[1][0][7] , \reg_in[1][0][6] ,
         \reg_in[1][0][5] , \reg_in[1][0][4] , \reg_in[1][0][3] ,
         \reg_in[1][0][2] , \reg_in[1][0][1] , \reg_in[1][0][0] ,
         \reg_in[0][3][19] , \reg_in[0][3][18] , \reg_in[0][3][17] ,
         \reg_in[0][3][16] , \reg_in[0][3][15] , \reg_in[0][3][14] ,
         \reg_in[0][3][13] , \reg_in[0][3][12] , \reg_in[0][3][11] ,
         \reg_in[0][3][10] , \reg_in[0][3][9] , \reg_in[0][3][8] ,
         \reg_in[0][3][7] , \reg_in[0][3][6] , \reg_in[0][3][5] ,
         \reg_in[0][3][4] , \reg_in[0][3][3] , \reg_in[0][3][2] ,
         \reg_in[0][3][1] , \reg_in[0][3][0] , \reg_in[0][2][19] ,
         \reg_in[0][2][18] , \reg_in[0][2][17] , \reg_in[0][2][16] ,
         \reg_in[0][2][15] , \reg_in[0][2][14] , \reg_in[0][2][13] ,
         \reg_in[0][2][12] , \reg_in[0][2][11] , \reg_in[0][2][10] ,
         \reg_in[0][2][9] , \reg_in[0][2][8] , \reg_in[0][2][7] ,
         \reg_in[0][2][6] , \reg_in[0][2][5] , \reg_in[0][2][4] ,
         \reg_in[0][2][3] , \reg_in[0][2][2] , \reg_in[0][2][1] ,
         \reg_in[0][2][0] , \reg_in[0][1][19] , \reg_in[0][1][18] ,
         \reg_in[0][1][17] , \reg_in[0][1][16] , \reg_in[0][1][15] ,
         \reg_in[0][1][14] , \reg_in[0][1][13] , \reg_in[0][1][12] ,
         \reg_in[0][1][11] , \reg_in[0][1][10] , \reg_in[0][1][9] ,
         \reg_in[0][1][8] , \reg_in[0][1][7] , \reg_in[0][1][6] ,
         \reg_in[0][1][5] , \reg_in[0][1][4] , \reg_in[0][1][3] ,
         \reg_in[0][1][2] , \reg_in[0][1][1] , \reg_in[0][1][0] ,
         \reg_in[0][0][19] , \reg_in[0][0][18] , \reg_in[0][0][17] ,
         \reg_in[0][0][16] , \reg_in[0][0][15] , \reg_in[0][0][14] ,
         \reg_in[0][0][13] , \reg_in[0][0][12] , \reg_in[0][0][11] ,
         \reg_in[0][0][10] , \reg_in[0][0][9] , \reg_in[0][0][8] ,
         \reg_in[0][0][7] , \reg_in[0][0][6] , \reg_in[0][0][5] ,
         \reg_in[0][0][4] , \reg_in[0][0][3] , \reg_in[0][0][2] ,
         \reg_in[0][0][1] , \reg_in[0][0][0] , n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18400, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n5145, n5141, n5137, n5133, n5129, n5125, n5121, n5117, n5113,
         n5109, n5105, n5101, n5097, n5093, n5089, n5085, n5081, n5077, n5073,
         n5069, n5065, n5061, n5057, n5053, n5049, n5045, n5041, n5037, n5033,
         n5029, n5025, n5021, n5017, n5013, n5009, n5005, n5001, n4997, n4993,
         n4989, n4985, n4981, n4977, n4973, n4969, n4965, n4961, n4957, n4953,
         n4949, n4945, n4941, n4937, n4933, n4929, n4925, n4921, n4917, n4913,
         n4909, n4905, n4901, n4897, n4893, n4889, n4885, n4881, n4877, n4873,
         n4869, n4865, n4861, n4857, n4853, n4849, n4845, n4841, n4837, n4833,
         n4829, n4825, n4821, n4817, n4813, n4809, n4805, n4801, n4797, n4793,
         n4789, n4785, n4781, n4777, n4773, n4769, n4765, n4761, n4757, n4753,
         n4749, n4745, n4741, n4737, n4733, n4729, n4725, n4721, n4717, n4713,
         n4709, n4705, n4701, n4697, n4693, n4689, n4685, n4681, n4677, n4673,
         n4669, n4665, n4661, n4657, n4653, n4649, n4645, n4641, n4637, n4633,
         n4629, n4625, n4621, n4617, n4613, n4609, n4605, n4601, n4597, n4593,
         n4589, n4585, n4581, n4577, n4573, n4569, n4565, n4561, n4557, n4553,
         n4549, n4545, n4541, n4537, n4533, n4529, n4525, n4521, n4517, n4513,
         n4509, n4505, n4501, n4497, n4493, n4489, n4485, n4481, n4477, n4473,
         n4469, n4465, n4461, n4457, n4453, n4449, n4445, n4441, n4437, n4433,
         n4429, n4425, n4421, n4417, n4413, n4409, n4405, n4401, n4397, n4393,
         n4389, n4385, n4381, n4377, n4373, n4369, n4365, n4361, n4357, n4353,
         n4349, n4345, n4341, n4337, n4333, n4329, n4325, n4321, n4317, n4313,
         n4309, n4305, n4301, n4297, n4293, n4289, n4285, n4281, n4277, n4273,
         n4269, n4265, n4261, n4257, n4253, n4249, n4245, n4241, n4237, n4233,
         n4229, n4225, n4221, n4217, n4213, n4209, n4205, n4201, n4197, n4193,
         n4189, n4185, n4181, n4177, n4173, n4169, n4165, n4161, n4157, n4153,
         n4149, n4145, n4141, n4137, n4133, n4129, n4125, n4121, n4117, n4113,
         n4109, n4105, n4101, n4097, n4093, n4089, n4085, n4081, n4077, n4073,
         n4069, n4065, n4061, n4057, n4053, n4049, n4045, n4041, n4037, n4033,
         n4029, n4025, n4021, n4017, n4013, n4009, n4005, n4001, n3997, n3993,
         n3989, n3985, n3981, n3977, n3973, n3969, n3965, n3961, n3957, n3953,
         n3949, n3945, n3941, n3937, n3933, n3929, n3925, n3921, n3917, n3913,
         n3909, n3905, n3901, n3897, n3893, n3889, n3885, n3881, n3877, n3873,
         n3869, n12859, n12858, n12857, n12856, n12855, n12854, n12853, n12852,
         n12851, n12850, n12849, n12848, n12847, n12846, n12845, n12844,
         n12843, n12842, n12841, n12840, n12839, n12838, n12837, n12836,
         n12835, n12834, n12833, n12832, n12831, n12830, n12829, n12828,
         n12827, n12826, n12825, n12824, n12823, n12822, n12821, n12820,
         n12819, n12818, n12817, n12816, n12815, n12814, n12813, n12812,
         n12811, n12810, n12809, n12808, n12807, n12806, n12805, n12804,
         n12803, n12802, n12801, n12800, n12799, n12798, n12797, n12796,
         n12795, n12794, n12793, n12792, n12791, n12790, n12789, n12788,
         n12787, n12786, n12785, n12784, n12783, n12782, n12781, n12780,
         n12779, n12778, n12777, n12776, n12775, n12774, n12773, n12772,
         n12771, n12770, n12769, n12768, n12767, n12766, n12765, n12764,
         n12763, n12762, n12761, n12760, n12759, n12758, n12757, n12756,
         n12755, n12754, n12753, n12752, n12751, n12750, n12749, n12748,
         n12747, n12746, n12745, n12744, n12743, n12742, n12741, n12740,
         n12739, n12738, n12737, n12736, n12735, n12734, n12733, n12732,
         n12731, n12730, n12729, n12728, n12727, n12726, n12725, n12724,
         n12723, n12722, n12721, n12720, n12719, n12718, n12717, n12716,
         n12715, n12714, n12713, n12712, n12711, n12710, n12709, n12708,
         n12707, n12706, n12705, n12704, n12703, n12702, n12701, n12700,
         n12699, n12698, n12697, n12696, n12695, n12694, n12693, n12692,
         n12691, n12690, n12689, n12688, n12687, n12686, n12685, n12684,
         n12683, n12682, n12681, n12680, n12679, n12678, n12677, n12676,
         n12675, n12674, n12673, n12672, n12671, n12670, n12669, n12668,
         n12667, n12666, n12665, n12664, n12663, n12662, n12661, n12660,
         n12659, n12658, n12657, n12656, n12655, n12654, n12653, n12652,
         n12651, n12650, n12649, n12648, n12647, n12646, n12645, n12644,
         n12643, n12642, n12641, n12640, n12639, n12638, n12637, n12636,
         n12635, n12634, n12633, n12632, n12631, n12630, n12629, n12628,
         n12627, n12626, n12625, n12624, n12623, n12622, n12621, n12620,
         n12619, n12618, n12617, n12616, n12615, n12614, n12613, n12612,
         n12611, n12610, n12609, n12608, n12607, n12606, n12605, n12604,
         n12603, n12602, n12601, n12600, n12599, n12598, n12597, n12596,
         n12595, n12594, n12593, n12592, n12591, n12590, n12589, n12588,
         n12587, n12586, n12585, n12584, n12583, n12582, n12581, n12580,
         n12579, n12578, n12577, n12576, n12575, n12574, n12573, n12572,
         n12571, n12570, n12569, n12568, n12567, n12566, n12565, n12564,
         n12563, n12562, n12561, n12560, n12559, n12558, n12557, n12556,
         n12555, n12554, n12553, n12552, n12551, n12550, n12549, n12548,
         n12547, n12546, n12545, n12544, n12543, n12542, n12541, n12540,
         n15445, n15446, n15447, n15448, n15449, n15451, n15453, n15455,
         n15457, n15459, n15461, n15463, n15465, n15467, n15469, n15471,
         n15473, n15475, n15477, n15479, n15481, n15483, n15485, n15487,
         n15489, n15491, n15493, n15495, n15497, n15499, n15501, n15503,
         n15505, n15507, n15509, n15511, n15513, n15515, n15517, n15519,
         n15521, n15523, n15525, n15527, n15529, n15531, n15533, n15535,
         n15537, n15539, n15541, n15543, n15545, n15547, n15549, n15551,
         n15553, n15555, n15557, n15559, n15561, n15563, n15565, n15567,
         n15569, n15571, n15573, n15575, n15577, n15579, n15581, n15583,
         n15585, n15587, n15589, n15591, n15593, n15595, n15597, n15599,
         n15601, n15603, n15605, n15607, n15609, n15611, n15613, n15615,
         n15617, n15619, n15621, n15623, n15625, n15627, n15629, n15631,
         n15633, n15635, n15637, n15639, n15641, n15643, n15645, n15647,
         n15649, n15651, n15653, n15655, n15657, n15659, n15661, n15663,
         n15665, n15667, n15669, n15671, n15673, n15675, n15677, n15679,
         n15681, n15683, n15685, n15687, n15689, n15691, n15693, n15695,
         n15697, n15699, n15701, n15703, n15705, n15707, n15709, n15711,
         n15713, n15715, n15717, n15719, n15721, n15723, n15725, n15727,
         n15729, n15731, n15733, n15735, n15737, n15739, n15741, n15743,
         n15745, n15747, n15749, n15751, n15753, n15755, n15757, n15759,
         n15761, n15763, n15765, n15767, n15769, n15771, n15773, n15775,
         n15777, n15779, n15781, n15783, n15785, n15787, n15789, n15791,
         n15793, n15795, n15797, n15799, n15801, n15803, n15805, n15807,
         n15809, n15811, n15813, n15815, n15817, n15819, n15821, n15823,
         n15825, n15827, n15829, n15831, n15833, n15835, n15837, n15839,
         n15841, n15843, n15845, n15847, n15849, n15851, n15853, n15855,
         n15857, n15859, n15861, n15863, n15865, n15867, n15869, n15871,
         n15873, n15875, n15877, n15879, n15881, n15883, n15885, n15887,
         n15889, n15891, n15893, n15895, n15897, n15899, n15901, n15903,
         n15905, n15907, n15909, n15911, n15913, n15915, n15917, n15919,
         n15921, n15923, n15925, n15927, n15929, n15931, n15933, n15935,
         n15937, n15939, n15941, n15943, n15945, n15947, n15949, n15951,
         n15953, n15955, n15957, n15959, n15961, n15963, n15965, n15967,
         n15969, n15971, n15973, n15975, n15977, n15979, n15981, n15983,
         n15985, n15987, n15989, n15991, n15993, n15995, n15997, n15999,
         n16001, n16003, n16005, n16007, n16009, n16011, n16013, n16015,
         n16017, n16019, n16021, n16023, n16025, n16027, n16029, n16031,
         n16033, n16035, n16037, n16039, n16041, n16043, n16045, n16047,
         n16049, n16051, n16053, n16055, n16057, n16059, n16061, n16063,
         n16065, n16067, n16069, n16071, n16073, n16075, n16077, n16079,
         n16081, n16083, n16085, n16087, n16089, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399;

  dff_sg \state_reg[0]  ( .D(n15444), .CP(clk), .Q(n18401) );
  dff_sg \state_reg[1]  ( .D(n15443), .CP(clk), .Q(n18400) );
  dff_sg \reg_in_reg[3][3][19]  ( .D(n15317), .CP(clk), .Q(\reg_in[3][3][19] )
         );
  dff_sg \reg_in_reg[3][3][18]  ( .D(n15321), .CP(clk), .Q(\reg_in[3][3][18] )
         );
  dff_sg \reg_in_reg[3][3][17]  ( .D(n15320), .CP(clk), .Q(\reg_in[3][3][17] )
         );
  dff_sg \reg_in_reg[3][3][16]  ( .D(n15312), .CP(clk), .Q(\reg_in[3][3][16] )
         );
  dff_sg \reg_in_reg[3][3][15]  ( .D(n15311), .CP(clk), .Q(\reg_in[3][3][15] )
         );
  dff_sg \reg_in_reg[3][3][14]  ( .D(n15315), .CP(clk), .Q(\reg_in[3][3][14] )
         );
  dff_sg \reg_in_reg[3][3][13]  ( .D(n15314), .CP(clk), .Q(\reg_in[3][3][13] )
         );
  dff_sg \reg_in_reg[3][3][12]  ( .D(n15186), .CP(clk), .Q(\reg_in[3][3][12] )
         );
  dff_sg \reg_in_reg[3][3][11]  ( .D(n15185), .CP(clk), .Q(\reg_in[3][3][11] )
         );
  dff_sg \reg_in_reg[3][3][10]  ( .D(n15189), .CP(clk), .Q(\reg_in[3][3][10] )
         );
  dff_sg \reg_in_reg[3][3][9]  ( .D(n15188), .CP(clk), .Q(\reg_in[3][3][9] )
         );
  dff_sg \reg_in_reg[3][3][8]  ( .D(n15180), .CP(clk), .Q(\reg_in[3][3][8] )
         );
  dff_sg \reg_in_reg[3][3][7]  ( .D(n15179), .CP(clk), .Q(\reg_in[3][3][7] )
         );
  dff_sg \reg_in_reg[3][3][6]  ( .D(n15183), .CP(clk), .Q(\reg_in[3][3][6] )
         );
  dff_sg \reg_in_reg[3][3][5]  ( .D(n15182), .CP(clk), .Q(\reg_in[3][3][5] )
         );
  dff_sg \reg_in_reg[3][3][4]  ( .D(n15198), .CP(clk), .Q(\reg_in[3][3][4] )
         );
  dff_sg \reg_in_reg[3][3][3]  ( .D(n15197), .CP(clk), .Q(\reg_in[3][3][3] )
         );
  dff_sg \reg_in_reg[3][3][2]  ( .D(n15201), .CP(clk), .Q(\reg_in[3][3][2] )
         );
  dff_sg \reg_in_reg[3][3][1]  ( .D(n15200), .CP(clk), .Q(\reg_in[3][3][1] )
         );
  dff_sg \reg_in_reg[3][3][0]  ( .D(n15192), .CP(clk), .Q(\reg_in[3][3][0] )
         );
  dff_sg \reg_in_reg[3][2][19]  ( .D(n15191), .CP(clk), .Q(\reg_in[3][2][19] )
         );
  dff_sg \reg_in_reg[3][2][18]  ( .D(n15195), .CP(clk), .Q(\reg_in[3][2][18] )
         );
  dff_sg \reg_in_reg[3][2][17]  ( .D(n15194), .CP(clk), .Q(\reg_in[3][2][17] )
         );
  dff_sg \reg_in_reg[3][2][16]  ( .D(n15162), .CP(clk), .Q(\reg_in[3][2][16] )
         );
  dff_sg \reg_in_reg[3][2][15]  ( .D(n15161), .CP(clk), .Q(\reg_in[3][2][15] )
         );
  dff_sg \reg_in_reg[3][2][14]  ( .D(n15165), .CP(clk), .Q(\reg_in[3][2][14] )
         );
  dff_sg \reg_in_reg[3][2][13]  ( .D(n15164), .CP(clk), .Q(\reg_in[3][2][13] )
         );
  dff_sg \reg_in_reg[3][2][12]  ( .D(n15156), .CP(clk), .Q(\reg_in[3][2][12] )
         );
  dff_sg \reg_in_reg[3][2][11]  ( .D(n15155), .CP(clk), .Q(\reg_in[3][2][11] )
         );
  dff_sg \reg_in_reg[3][2][10]  ( .D(n15159), .CP(clk), .Q(\reg_in[3][2][10] )
         );
  dff_sg \reg_in_reg[3][2][9]  ( .D(n15158), .CP(clk), .Q(\reg_in[3][2][9] )
         );
  dff_sg \reg_in_reg[3][2][8]  ( .D(n15174), .CP(clk), .Q(\reg_in[3][2][8] )
         );
  dff_sg \reg_in_reg[3][2][7]  ( .D(n15173), .CP(clk), .Q(\reg_in[3][2][7] )
         );
  dff_sg \reg_in_reg[3][2][6]  ( .D(n15177), .CP(clk), .Q(\reg_in[3][2][6] )
         );
  dff_sg \reg_in_reg[3][2][5]  ( .D(n15176), .CP(clk), .Q(\reg_in[3][2][5] )
         );
  dff_sg \reg_in_reg[3][2][4]  ( .D(n15168), .CP(clk), .Q(\reg_in[3][2][4] )
         );
  dff_sg \reg_in_reg[3][2][3]  ( .D(n15167), .CP(clk), .Q(\reg_in[3][2][3] )
         );
  dff_sg \reg_in_reg[3][2][2]  ( .D(n15171), .CP(clk), .Q(\reg_in[3][2][2] )
         );
  dff_sg \reg_in_reg[3][2][1]  ( .D(n15170), .CP(clk), .Q(\reg_in[3][2][1] )
         );
  dff_sg \reg_in_reg[3][2][0]  ( .D(n15234), .CP(clk), .Q(\reg_in[3][2][0] )
         );
  dff_sg \reg_in_reg[3][1][19]  ( .D(n15233), .CP(clk), .Q(\reg_in[3][1][19] )
         );
  dff_sg \reg_in_reg[3][1][18]  ( .D(n15237), .CP(clk), .Q(\reg_in[3][1][18] )
         );
  dff_sg \reg_in_reg[3][1][17]  ( .D(n15236), .CP(clk), .Q(\reg_in[3][1][17] )
         );
  dff_sg \reg_in_reg[3][1][16]  ( .D(n15228), .CP(clk), .Q(\reg_in[3][1][16] )
         );
  dff_sg \reg_in_reg[3][1][15]  ( .D(n15227), .CP(clk), .Q(\reg_in[3][1][15] )
         );
  dff_sg \reg_in_reg[3][1][14]  ( .D(n15231), .CP(clk), .Q(\reg_in[3][1][14] )
         );
  dff_sg \reg_in_reg[3][1][13]  ( .D(n15230), .CP(clk), .Q(\reg_in[3][1][13] )
         );
  dff_sg \reg_in_reg[3][1][12]  ( .D(n15246), .CP(clk), .Q(\reg_in[3][1][12] )
         );
  dff_sg \reg_in_reg[3][1][11]  ( .D(n15245), .CP(clk), .Q(\reg_in[3][1][11] )
         );
  dff_sg \reg_in_reg[3][1][10]  ( .D(n15249), .CP(clk), .Q(\reg_in[3][1][10] )
         );
  dff_sg \reg_in_reg[3][1][9]  ( .D(n15248), .CP(clk), .Q(\reg_in[3][1][9] )
         );
  dff_sg \reg_in_reg[3][1][8]  ( .D(n15240), .CP(clk), .Q(\reg_in[3][1][8] )
         );
  dff_sg \reg_in_reg[3][1][7]  ( .D(n15239), .CP(clk), .Q(\reg_in[3][1][7] )
         );
  dff_sg \reg_in_reg[3][1][6]  ( .D(n15243), .CP(clk), .Q(\reg_in[3][1][6] )
         );
  dff_sg \reg_in_reg[3][1][5]  ( .D(n15242), .CP(clk), .Q(\reg_in[3][1][5] )
         );
  dff_sg \reg_in_reg[3][1][4]  ( .D(n15210), .CP(clk), .Q(\reg_in[3][1][4] )
         );
  dff_sg \reg_in_reg[3][1][3]  ( .D(n15209), .CP(clk), .Q(\reg_in[3][1][3] )
         );
  dff_sg \reg_in_reg[3][1][2]  ( .D(n15213), .CP(clk), .Q(\reg_in[3][1][2] )
         );
  dff_sg \reg_in_reg[3][1][1]  ( .D(n15212), .CP(clk), .Q(\reg_in[3][1][1] )
         );
  dff_sg \reg_in_reg[3][1][0]  ( .D(n15204), .CP(clk), .Q(\reg_in[3][1][0] )
         );
  dff_sg \reg_in_reg[3][0][19]  ( .D(n15203), .CP(clk), .Q(\reg_in[3][0][19] )
         );
  dff_sg \reg_in_reg[3][0][18]  ( .D(n15207), .CP(clk), .Q(\reg_in[3][0][18] )
         );
  dff_sg \reg_in_reg[3][0][17]  ( .D(n15206), .CP(clk), .Q(\reg_in[3][0][17] )
         );
  dff_sg \reg_in_reg[3][0][16]  ( .D(n15222), .CP(clk), .Q(\reg_in[3][0][16] )
         );
  dff_sg \reg_in_reg[3][0][15]  ( .D(n15221), .CP(clk), .Q(\reg_in[3][0][15] )
         );
  dff_sg \reg_in_reg[3][0][14]  ( .D(n15225), .CP(clk), .Q(\reg_in[3][0][14] )
         );
  dff_sg \reg_in_reg[3][0][13]  ( .D(n15224), .CP(clk), .Q(\reg_in[3][0][13] )
         );
  dff_sg \reg_in_reg[3][0][12]  ( .D(n15216), .CP(clk), .Q(\reg_in[3][0][12] )
         );
  dff_sg \reg_in_reg[3][0][11]  ( .D(n15215), .CP(clk), .Q(\reg_in[3][0][11] )
         );
  dff_sg \reg_in_reg[3][0][10]  ( .D(n15219), .CP(clk), .Q(\reg_in[3][0][10] )
         );
  dff_sg \reg_in_reg[3][0][9]  ( .D(n15218), .CP(clk), .Q(\reg_in[3][0][9] )
         );
  dff_sg \reg_in_reg[3][0][8]  ( .D(n15379), .CP(clk), .Q(\reg_in[3][0][8] )
         );
  dff_sg \reg_in_reg[3][0][7]  ( .D(n15378), .CP(clk), .Q(\reg_in[3][0][7] )
         );
  dff_sg \reg_in_reg[3][0][6]  ( .D(n15382), .CP(clk), .Q(\reg_in[3][0][6] )
         );
  dff_sg \reg_in_reg[3][0][5]  ( .D(n15381), .CP(clk), .Q(\reg_in[3][0][5] )
         );
  dff_sg \reg_in_reg[3][0][4]  ( .D(n15373), .CP(clk), .Q(\reg_in[3][0][4] )
         );
  dff_sg \reg_in_reg[3][0][3]  ( .D(n15372), .CP(clk), .Q(\reg_in[3][0][3] )
         );
  dff_sg \reg_in_reg[3][0][2]  ( .D(n15376), .CP(clk), .Q(\reg_in[3][0][2] )
         );
  dff_sg \reg_in_reg[3][0][1]  ( .D(n15375), .CP(clk), .Q(\reg_in[3][0][1] )
         );
  dff_sg \reg_in_reg[3][0][0]  ( .D(n15391), .CP(clk), .Q(\reg_in[3][0][0] )
         );
  dff_sg \reg_in_reg[2][3][19]  ( .D(n15390), .CP(clk), .Q(\reg_in[2][3][19] )
         );
  dff_sg \reg_in_reg[2][3][18]  ( .D(n15394), .CP(clk), .Q(\reg_in[2][3][18] )
         );
  dff_sg \reg_in_reg[2][3][17]  ( .D(n15393), .CP(clk), .Q(\reg_in[2][3][17] )
         );
  dff_sg \reg_in_reg[2][3][16]  ( .D(n15385), .CP(clk), .Q(\reg_in[2][3][16] )
         );
  dff_sg \reg_in_reg[2][3][15]  ( .D(n15384), .CP(clk), .Q(\reg_in[2][3][15] )
         );
  dff_sg \reg_in_reg[2][3][14]  ( .D(n15388), .CP(clk), .Q(\reg_in[2][3][14] )
         );
  dff_sg \reg_in_reg[2][3][13]  ( .D(n15387), .CP(clk), .Q(\reg_in[2][3][13] )
         );
  dff_sg \reg_in_reg[2][3][12]  ( .D(n15355), .CP(clk), .Q(\reg_in[2][3][12] )
         );
  dff_sg \reg_in_reg[2][3][11]  ( .D(n15354), .CP(clk), .Q(\reg_in[2][3][11] )
         );
  dff_sg \reg_in_reg[2][3][10]  ( .D(n15358), .CP(clk), .Q(\reg_in[2][3][10] )
         );
  dff_sg \reg_in_reg[2][3][9]  ( .D(n15357), .CP(clk), .Q(\reg_in[2][3][9] )
         );
  dff_sg \reg_in_reg[2][3][8]  ( .D(n15349), .CP(clk), .Q(\reg_in[2][3][8] )
         );
  dff_sg \reg_in_reg[2][3][7]  ( .D(n15348), .CP(clk), .Q(\reg_in[2][3][7] )
         );
  dff_sg \reg_in_reg[2][3][6]  ( .D(n15352), .CP(clk), .Q(\reg_in[2][3][6] )
         );
  dff_sg \reg_in_reg[2][3][5]  ( .D(n15351), .CP(clk), .Q(\reg_in[2][3][5] )
         );
  dff_sg \reg_in_reg[2][3][4]  ( .D(n15367), .CP(clk), .Q(\reg_in[2][3][4] )
         );
  dff_sg \reg_in_reg[2][3][3]  ( .D(n15366), .CP(clk), .Q(\reg_in[2][3][3] )
         );
  dff_sg \reg_in_reg[2][3][2]  ( .D(n15370), .CP(clk), .Q(\reg_in[2][3][2] )
         );
  dff_sg \reg_in_reg[2][3][1]  ( .D(n15369), .CP(clk), .Q(\reg_in[2][3][1] )
         );
  dff_sg \reg_in_reg[2][3][0]  ( .D(n15361), .CP(clk), .Q(\reg_in[2][3][0] )
         );
  dff_sg \reg_in_reg[2][2][19]  ( .D(n15360), .CP(clk), .Q(\reg_in[2][2][19] )
         );
  dff_sg \reg_in_reg[2][2][18]  ( .D(n15364), .CP(clk), .Q(\reg_in[2][2][18] )
         );
  dff_sg \reg_in_reg[2][2][17]  ( .D(n15363), .CP(clk), .Q(\reg_in[2][2][17] )
         );
  dff_sg \reg_in_reg[2][2][16]  ( .D(n15427), .CP(clk), .Q(\reg_in[2][2][16] )
         );
  dff_sg \reg_in_reg[2][2][15]  ( .D(n15426), .CP(clk), .Q(\reg_in[2][2][15] )
         );
  dff_sg \reg_in_reg[2][2][14]  ( .D(n15430), .CP(clk), .Q(\reg_in[2][2][14] )
         );
  dff_sg \reg_in_reg[2][2][13]  ( .D(n15429), .CP(clk), .Q(\reg_in[2][2][13] )
         );
  dff_sg \reg_in_reg[2][2][12]  ( .D(n15421), .CP(clk), .Q(\reg_in[2][2][12] )
         );
  dff_sg \reg_in_reg[2][2][11]  ( .D(n15420), .CP(clk), .Q(\reg_in[2][2][11] )
         );
  dff_sg \reg_in_reg[2][2][10]  ( .D(n15424), .CP(clk), .Q(\reg_in[2][2][10] )
         );
  dff_sg \reg_in_reg[2][2][9]  ( .D(n15423), .CP(clk), .Q(\reg_in[2][2][9] )
         );
  dff_sg \reg_in_reg[2][2][8]  ( .D(n15439), .CP(clk), .Q(\reg_in[2][2][8] )
         );
  dff_sg \reg_in_reg[2][2][7]  ( .D(n15438), .CP(clk), .Q(\reg_in[2][2][7] )
         );
  dff_sg \reg_in_reg[2][2][6]  ( .D(n15442), .CP(clk), .Q(\reg_in[2][2][6] )
         );
  dff_sg \reg_in_reg[2][2][5]  ( .D(n15441), .CP(clk), .Q(\reg_in[2][2][5] )
         );
  dff_sg \reg_in_reg[2][2][4]  ( .D(n15433), .CP(clk), .Q(\reg_in[2][2][4] )
         );
  dff_sg \reg_in_reg[2][2][3]  ( .D(n15432), .CP(clk), .Q(\reg_in[2][2][3] )
         );
  dff_sg \reg_in_reg[2][2][2]  ( .D(n15436), .CP(clk), .Q(\reg_in[2][2][2] )
         );
  dff_sg \reg_in_reg[2][2][1]  ( .D(n15435), .CP(clk), .Q(\reg_in[2][2][1] )
         );
  dff_sg \reg_in_reg[2][2][0]  ( .D(n15403), .CP(clk), .Q(\reg_in[2][2][0] )
         );
  dff_sg \reg_in_reg[2][1][19]  ( .D(n15402), .CP(clk), .Q(\reg_in[2][1][19] )
         );
  dff_sg \reg_in_reg[2][1][18]  ( .D(n15406), .CP(clk), .Q(\reg_in[2][1][18] )
         );
  dff_sg \reg_in_reg[2][1][17]  ( .D(n15405), .CP(clk), .Q(\reg_in[2][1][17] )
         );
  dff_sg \reg_in_reg[2][1][16]  ( .D(n15397), .CP(clk), .Q(\reg_in[2][1][16] )
         );
  dff_sg \reg_in_reg[2][1][15]  ( .D(n15396), .CP(clk), .Q(\reg_in[2][1][15] )
         );
  dff_sg \reg_in_reg[2][1][14]  ( .D(n15400), .CP(clk), .Q(\reg_in[2][1][14] )
         );
  dff_sg \reg_in_reg[2][1][13]  ( .D(n15399), .CP(clk), .Q(\reg_in[2][1][13] )
         );
  dff_sg \reg_in_reg[2][1][12]  ( .D(n15415), .CP(clk), .Q(\reg_in[2][1][12] )
         );
  dff_sg \reg_in_reg[2][1][11]  ( .D(n15414), .CP(clk), .Q(\reg_in[2][1][11] )
         );
  dff_sg \reg_in_reg[2][1][10]  ( .D(n15418), .CP(clk), .Q(\reg_in[2][1][10] )
         );
  dff_sg \reg_in_reg[2][1][9]  ( .D(n15417), .CP(clk), .Q(\reg_in[2][1][9] )
         );
  dff_sg \reg_in_reg[2][1][8]  ( .D(n15409), .CP(clk), .Q(\reg_in[2][1][8] )
         );
  dff_sg \reg_in_reg[2][1][7]  ( .D(n15408), .CP(clk), .Q(\reg_in[2][1][7] )
         );
  dff_sg \reg_in_reg[2][1][6]  ( .D(n15412), .CP(clk), .Q(\reg_in[2][1][6] )
         );
  dff_sg \reg_in_reg[2][1][5]  ( .D(n15411), .CP(clk), .Q(\reg_in[2][1][5] )
         );
  dff_sg \reg_in_reg[2][1][4]  ( .D(n15250), .CP(clk), .Q(\reg_in[2][1][4] )
         );
  dff_sg \reg_in_reg[2][1][3]  ( .D(n15141), .CP(clk), .Q(\reg_in[2][1][3] )
         );
  dff_sg \reg_in_reg[2][1][2]  ( .D(n15199), .CP(clk), .Q(\reg_in[2][1][2] )
         );
  dff_sg \reg_in_reg[2][1][1]  ( .D(n15241), .CP(clk), .Q(\reg_in[2][1][1] )
         );
  dff_sg \reg_in_reg[2][1][0]  ( .D(n15190), .CP(clk), .Q(\reg_in[2][1][0] )
         );
  dff_sg \reg_in_reg[2][0][19]  ( .D(n15142), .CP(clk), .Q(\reg_in[2][0][19] )
         );
  dff_sg \reg_in_reg[2][0][18]  ( .D(n15184), .CP(clk), .Q(\reg_in[2][0][18] )
         );
  dff_sg \reg_in_reg[2][0][17]  ( .D(n15181), .CP(clk), .Q(\reg_in[2][0][17] )
         );
  dff_sg \reg_in_reg[2][0][16]  ( .D(n15226), .CP(clk), .Q(\reg_in[2][0][16] )
         );
  dff_sg \reg_in_reg[2][0][15]  ( .D(n15223), .CP(clk), .Q(\reg_in[2][0][15] )
         );
  dff_sg \reg_in_reg[2][0][14]  ( .D(n15211), .CP(clk), .Q(\reg_in[2][0][14] )
         );
  dff_sg \reg_in_reg[2][0][13]  ( .D(n15208), .CP(clk), .Q(\reg_in[2][0][13] )
         );
  dff_sg \reg_in_reg[2][0][12]  ( .D(n15247), .CP(clk), .Q(\reg_in[2][0][12] )
         );
  dff_sg \reg_in_reg[2][0][11]  ( .D(n15244), .CP(clk), .Q(\reg_in[2][0][11] )
         );
  dff_sg \reg_in_reg[2][0][10]  ( .D(n15232), .CP(clk), .Q(\reg_in[2][0][10] )
         );
  dff_sg \reg_in_reg[2][0][9]  ( .D(n15229), .CP(clk), .Q(\reg_in[2][0][9] )
         );
  dff_sg \reg_in_reg[2][0][8]  ( .D(n15437), .CP(clk), .Q(\reg_in[2][0][8] )
         );
  dff_sg \reg_in_reg[2][0][7]  ( .D(n15163), .CP(clk), .Q(\reg_in[2][0][7] )
         );
  dff_sg \reg_in_reg[2][0][6]  ( .D(n15428), .CP(clk), .Q(\reg_in[2][0][6] )
         );
  dff_sg \reg_in_reg[2][0][5]  ( .D(n15425), .CP(clk), .Q(\reg_in[2][0][5] )
         );
  dff_sg \reg_in_reg[2][0][4]  ( .D(n15365), .CP(clk), .Q(\reg_in[2][0][4] )
         );
  dff_sg \reg_in_reg[2][0][3]  ( .D(n15160), .CP(clk), .Q(\reg_in[2][0][3] )
         );
  dff_sg \reg_in_reg[2][0][2]  ( .D(n15356), .CP(clk), .Q(\reg_in[2][0][2] )
         );
  dff_sg \reg_in_reg[2][0][1]  ( .D(n15350), .CP(clk), .Q(\reg_in[2][0][1] )
         );
  dff_sg \reg_in_reg[2][0][0]  ( .D(n15175), .CP(clk), .Q(\reg_in[2][0][0] )
         );
  dff_sg \reg_in_reg[1][3][19]  ( .D(n15172), .CP(clk), .Q(\reg_in[1][3][19] )
         );
  dff_sg \reg_in_reg[1][3][18]  ( .D(n15166), .CP(clk), .Q(\reg_in[1][3][18] )
         );
  dff_sg \reg_in_reg[1][3][17]  ( .D(n15152), .CP(clk), .Q(\reg_in[1][3][17] )
         );
  dff_sg \reg_in_reg[1][3][16]  ( .D(n15410), .CP(clk), .Q(\reg_in[1][3][16] )
         );
  dff_sg \reg_in_reg[1][3][15]  ( .D(n15407), .CP(clk), .Q(\reg_in[1][3][15] )
         );
  dff_sg \reg_in_reg[1][3][14]  ( .D(n15129), .CP(clk), .Q(\reg_in[1][3][14] )
         );
  dff_sg \reg_in_reg[1][3][13]  ( .D(n15151), .CP(clk), .Q(\reg_in[1][3][13] )
         );
  dff_sg \reg_in_reg[1][3][12]  ( .D(n15147), .CP(clk), .Q(\reg_in[1][3][12] )
         );
  dff_sg \reg_in_reg[1][3][11]  ( .D(n15146), .CP(clk), .Q(\reg_in[1][3][11] )
         );
  dff_sg \reg_in_reg[1][3][10]  ( .D(n15150), .CP(clk), .Q(\reg_in[1][3][10] )
         );
  dff_sg \reg_in_reg[1][3][9]  ( .D(n15149), .CP(clk), .Q(\reg_in[1][3][9] )
         );
  dff_sg \reg_in_reg[1][3][8]  ( .D(n15295), .CP(clk), .Q(\reg_in[1][3][8] )
         );
  dff_sg \reg_in_reg[1][3][7]  ( .D(n15292), .CP(clk), .Q(\reg_in[1][3][7] )
         );
  dff_sg \reg_in_reg[1][3][6]  ( .D(n15289), .CP(clk), .Q(\reg_in[1][3][6] )
         );
  dff_sg \reg_in_reg[1][3][5]  ( .D(n15286), .CP(clk), .Q(\reg_in[1][3][5] )
         );
  dff_sg \reg_in_reg[1][3][4]  ( .D(n15340), .CP(clk), .Q(\reg_in[1][3][4] )
         );
  dff_sg \reg_in_reg[1][3][3]  ( .D(n15337), .CP(clk), .Q(\reg_in[1][3][3] )
         );
  dff_sg \reg_in_reg[1][3][2]  ( .D(n15331), .CP(clk), .Q(\reg_in[1][3][2] )
         );
  dff_sg \reg_in_reg[1][3][1]  ( .D(n15328), .CP(clk), .Q(\reg_in[1][3][1] )
         );
  dff_sg \reg_in_reg[1][3][0]  ( .D(n15139), .CP(clk), .Q(\reg_in[1][3][0] )
         );
  dff_sg \reg_in_reg[1][2][19]  ( .D(n15138), .CP(clk), .Q(\reg_in[1][2][19] )
         );
  dff_sg \reg_in_reg[1][2][18]  ( .D(n15202), .CP(clk), .Q(\reg_in[1][2][18] )
         );
  dff_sg \reg_in_reg[1][2][17]  ( .D(n15214), .CP(clk), .Q(\reg_in[1][2][17] )
         );
  dff_sg \reg_in_reg[1][2][16]  ( .D(n15265), .CP(clk), .Q(\reg_in[1][2][16] )
         );
  dff_sg \reg_in_reg[1][2][15]  ( .D(n15262), .CP(clk), .Q(\reg_in[1][2][15] )
         );
  dff_sg \reg_in_reg[1][2][14]  ( .D(n15259), .CP(clk), .Q(\reg_in[1][2][14] )
         );
  dff_sg \reg_in_reg[1][2][13]  ( .D(n15256), .CP(clk), .Q(\reg_in[1][2][13] )
         );
  dff_sg \reg_in_reg[1][2][12]  ( .D(n15280), .CP(clk), .Q(\reg_in[1][2][12] )
         );
  dff_sg \reg_in_reg[1][2][11]  ( .D(n15125), .CP(clk), .Q(\reg_in[1][2][11] )
         );
  dff_sg \reg_in_reg[1][2][10]  ( .D(n15271), .CP(clk), .Q(\reg_in[1][2][10] )
         );
  dff_sg \reg_in_reg[1][2][9]  ( .D(n15268), .CP(clk), .Q(\reg_in[1][2][9] )
         );
  dff_sg \reg_in_reg[1][2][8]  ( .D(n15124), .CP(clk), .Q(\reg_in[1][2][8] )
         );
  dff_sg \reg_in_reg[1][2][7]  ( .D(n15123), .CP(clk), .Q(\reg_in[1][2][7] )
         );
  dff_sg \reg_in_reg[1][2][6]  ( .D(n15313), .CP(clk), .Q(\reg_in[1][2][6] )
         );
  dff_sg \reg_in_reg[1][2][5]  ( .D(n15310), .CP(clk), .Q(\reg_in[1][2][5] )
         );
  dff_sg \reg_in_reg[1][2][4]  ( .D(n15322), .CP(clk), .Q(\reg_in[1][2][4] )
         );
  dff_sg \reg_in_reg[1][2][3]  ( .D(n15319), .CP(clk), .Q(\reg_in[1][2][3] )
         );
  dff_sg \reg_in_reg[1][2][2]  ( .D(n15304), .CP(clk), .Q(\reg_in[1][2][2] )
         );
  dff_sg \reg_in_reg[1][2][1]  ( .D(n15301), .CP(clk), .Q(\reg_in[1][2][1] )
         );
  dff_sg \reg_in_reg[1][2][0]  ( .D(n15153), .CP(clk), .Q(\reg_in[1][2][0] )
         );
  dff_sg \reg_in_reg[1][1][19]  ( .D(n15343), .CP(clk), .Q(\reg_in[1][1][19] )
         );
  dff_sg \reg_in_reg[1][1][18]  ( .D(n15137), .CP(clk), .Q(\reg_in[1][1][18] )
         );
  dff_sg \reg_in_reg[1][1][17]  ( .D(n15148), .CP(clk), .Q(\reg_in[1][1][17] )
         );
  dff_sg \reg_in_reg[1][1][16]  ( .D(n15422), .CP(clk), .Q(\reg_in[1][1][16] )
         );
  dff_sg \reg_in_reg[1][1][15]  ( .D(n15220), .CP(clk), .Q(\reg_in[1][1][15] )
         );
  dff_sg \reg_in_reg[1][1][14]  ( .D(n15392), .CP(clk), .Q(\reg_in[1][1][14] )
         );
  dff_sg \reg_in_reg[1][1][13]  ( .D(n15413), .CP(clk), .Q(\reg_in[1][1][13] )
         );
  dff_sg \reg_in_reg[1][1][12]  ( .D(n15386), .CP(clk), .Q(\reg_in[1][1][12] )
         );
  dff_sg \reg_in_reg[1][1][11]  ( .D(n15383), .CP(clk), .Q(\reg_in[1][1][11] )
         );
  dff_sg \reg_in_reg[1][1][10]  ( .D(n15362), .CP(clk), .Q(\reg_in[1][1][10] )
         );
  dff_sg \reg_in_reg[1][1][9]  ( .D(n15416), .CP(clk), .Q(\reg_in[1][1][9] )
         );
  dff_sg \reg_in_reg[1][1][8]  ( .D(n15401), .CP(clk), .Q(\reg_in[1][1][8] )
         );
  dff_sg \reg_in_reg[1][1][7]  ( .D(n15419), .CP(clk), .Q(\reg_in[1][1][7] )
         );
  dff_sg \reg_in_reg[1][1][6]  ( .D(n15398), .CP(clk), .Q(\reg_in[1][1][6] )
         );
  dff_sg \reg_in_reg[1][1][5]  ( .D(n15395), .CP(clk), .Q(\reg_in[1][1][5] )
         );
  dff_sg \reg_in_reg[1][1][4]  ( .D(n15298), .CP(clk), .Q(\reg_in[1][1][4] )
         );
  dff_sg \reg_in_reg[1][1][3]  ( .D(n15132), .CP(clk), .Q(\reg_in[1][1][3] )
         );
  dff_sg \reg_in_reg[1][1][2]  ( .D(n15253), .CP(clk), .Q(\reg_in[1][1][2] )
         );
  dff_sg \reg_in_reg[1][1][1]  ( .D(n15283), .CP(clk), .Q(\reg_in[1][1][1] )
         );
  dff_sg \reg_in_reg[1][1][0]  ( .D(n15145), .CP(clk), .Q(\reg_in[1][1][0] )
         );
  dff_sg \reg_in_reg[1][0][19]  ( .D(n15131), .CP(clk), .Q(\reg_in[1][0][19] )
         );
  dff_sg \reg_in_reg[1][0][18]  ( .D(n15135), .CP(clk), .Q(\reg_in[1][0][18] )
         );
  dff_sg \reg_in_reg[1][0][17]  ( .D(n15307), .CP(clk), .Q(\reg_in[1][0][17] )
         );
  dff_sg \reg_in_reg[1][0][16]  ( .D(n15440), .CP(clk), .Q(\reg_in[1][0][16] )
         );
  dff_sg \reg_in_reg[1][0][15]  ( .D(n15134), .CP(clk), .Q(\reg_in[1][0][15] )
         );
  dff_sg \reg_in_reg[1][0][14]  ( .D(n15187), .CP(clk), .Q(\reg_in[1][0][14] )
         );
  dff_sg \reg_in_reg[1][0][13]  ( .D(n15334), .CP(clk), .Q(\reg_in[1][0][13] )
         );
  dff_sg \reg_in_reg[1][0][12]  ( .D(n15136), .CP(clk), .Q(\reg_in[1][0][12] )
         );
  dff_sg \reg_in_reg[1][0][11]  ( .D(n15133), .CP(clk), .Q(\reg_in[1][0][11] )
         );
  dff_sg \reg_in_reg[1][0][10]  ( .D(n15143), .CP(clk), .Q(\reg_in[1][0][10] )
         );
  dff_sg \reg_in_reg[1][0][9]  ( .D(n15144), .CP(clk), .Q(\reg_in[1][0][9] )
         );
  dff_sg \reg_in_reg[1][0][8]  ( .D(n15389), .CP(clk), .Q(\reg_in[1][0][8] )
         );
  dff_sg \reg_in_reg[1][0][7]  ( .D(n15380), .CP(clk), .Q(\reg_in[1][0][7] )
         );
  dff_sg \reg_in_reg[1][0][6]  ( .D(n15377), .CP(clk), .Q(\reg_in[1][0][6] )
         );
  dff_sg \reg_in_reg[1][0][5]  ( .D(n15374), .CP(clk), .Q(\reg_in[1][0][5] )
         );
  dff_sg \reg_in_reg[1][0][4]  ( .D(n15434), .CP(clk), .Q(\reg_in[1][0][4] )
         );
  dff_sg \reg_in_reg[1][0][3]  ( .D(n15325), .CP(clk), .Q(\reg_in[1][0][3] )
         );
  dff_sg \reg_in_reg[1][0][2]  ( .D(n15368), .CP(clk), .Q(\reg_in[1][0][2] )
         );
  dff_sg \reg_in_reg[1][0][1]  ( .D(n15359), .CP(clk), .Q(\reg_in[1][0][1] )
         );
  dff_sg \reg_in_reg[1][0][0]  ( .D(n15205), .CP(clk), .Q(\reg_in[1][0][0] )
         );
  dff_sg \reg_in_reg[0][3][19]  ( .D(n15193), .CP(clk), .Q(\reg_in[0][3][19] )
         );
  dff_sg \reg_in_reg[0][3][18]  ( .D(n15169), .CP(clk), .Q(\reg_in[0][3][18] )
         );
  dff_sg \reg_in_reg[0][3][17]  ( .D(n15178), .CP(clk), .Q(\reg_in[0][3][17] )
         );
  dff_sg \reg_in_reg[0][3][16]  ( .D(n15277), .CP(clk), .Q(\reg_in[0][3][16] )
         );
  dff_sg \reg_in_reg[0][3][15]  ( .D(n15127), .CP(clk), .Q(\reg_in[0][3][15] )
         );
  dff_sg \reg_in_reg[0][3][14]  ( .D(n15217), .CP(clk), .Q(\reg_in[0][3][14] )
         );
  dff_sg \reg_in_reg[0][3][13]  ( .D(n15235), .CP(clk), .Q(\reg_in[0][3][13] )
         );
  dff_sg \reg_in_reg[0][3][12]  ( .D(n15128), .CP(clk), .Q(\reg_in[0][3][12] )
         );
  dff_sg \reg_in_reg[0][3][11]  ( .D(n15238), .CP(clk), .Q(\reg_in[0][3][11] )
         );
  dff_sg \reg_in_reg[0][3][10]  ( .D(n15126), .CP(clk), .Q(\reg_in[0][3][10] )
         );
  dff_sg \reg_in_reg[0][3][9]  ( .D(n15371), .CP(clk), .Q(\reg_in[0][3][9] )
         );
  dff_sg \reg_in_reg[0][3][8]  ( .D(n15274), .CP(clk), .Q(\reg_in[0][3][8] )
         );
  dff_sg \reg_in_reg[0][3][7]  ( .D(n15196), .CP(clk), .Q(\reg_in[0][3][7] )
         );
  dff_sg \reg_in_reg[0][3][6]  ( .D(n15353), .CP(clk), .Q(\reg_in[0][3][6] )
         );
  dff_sg \reg_in_reg[0][3][5]  ( .D(n15316), .CP(clk), .Q(\reg_in[0][3][5] )
         );
  dff_sg \reg_in_reg[0][3][4]  ( .D(n15154), .CP(clk), .Q(\reg_in[0][3][4] )
         );
  dff_sg \reg_in_reg[0][3][3]  ( .D(n15431), .CP(clk), .Q(\reg_in[0][3][3] )
         );
  dff_sg \reg_in_reg[0][3][2]  ( .D(n15130), .CP(clk), .Q(\reg_in[0][3][2] )
         );
  dff_sg \reg_in_reg[0][3][1]  ( .D(n15140), .CP(clk), .Q(\reg_in[0][3][1] )
         );
  dff_sg \reg_in_reg[0][3][0]  ( .D(n15346), .CP(clk), .Q(\reg_in[0][3][0] )
         );
  dff_sg \reg_in_reg[0][2][19]  ( .D(n15404), .CP(clk), .Q(\reg_in[0][2][19] )
         );
  dff_sg \reg_in_reg[0][2][18]  ( .D(n15347), .CP(clk), .Q(\reg_in[0][2][18] )
         );
  dff_sg \reg_in_reg[0][2][17]  ( .D(n15157), .CP(clk), .Q(\reg_in[0][2][17] )
         );
  dff_sg \reg_in_reg[0][2][16]  ( .D(n15282), .CP(clk), .Q(\reg_in[0][2][16] )
         );
  dff_sg \reg_in_reg[0][2][15]  ( .D(n15281), .CP(clk), .Q(\reg_in[0][2][15] )
         );
  dff_sg \reg_in_reg[0][2][14]  ( .D(n15285), .CP(clk), .Q(\reg_in[0][2][14] )
         );
  dff_sg \reg_in_reg[0][2][13]  ( .D(n15284), .CP(clk), .Q(\reg_in[0][2][13] )
         );
  dff_sg \reg_in_reg[0][2][12]  ( .D(n15276), .CP(clk), .Q(\reg_in[0][2][12] )
         );
  dff_sg \reg_in_reg[0][2][11]  ( .D(n15275), .CP(clk), .Q(\reg_in[0][2][11] )
         );
  dff_sg \reg_in_reg[0][2][10]  ( .D(n15279), .CP(clk), .Q(\reg_in[0][2][10] )
         );
  dff_sg \reg_in_reg[0][2][9]  ( .D(n15278), .CP(clk), .Q(\reg_in[0][2][9] )
         );
  dff_sg \reg_in_reg[0][2][8]  ( .D(n15294), .CP(clk), .Q(\reg_in[0][2][8] )
         );
  dff_sg \reg_in_reg[0][2][7]  ( .D(n15293), .CP(clk), .Q(\reg_in[0][2][7] )
         );
  dff_sg \reg_in_reg[0][2][6]  ( .D(n15297), .CP(clk), .Q(\reg_in[0][2][6] )
         );
  dff_sg \reg_in_reg[0][2][5]  ( .D(n15296), .CP(clk), .Q(\reg_in[0][2][5] )
         );
  dff_sg \reg_in_reg[0][2][4]  ( .D(n15288), .CP(clk), .Q(\reg_in[0][2][4] )
         );
  dff_sg \reg_in_reg[0][2][3]  ( .D(n15287), .CP(clk), .Q(\reg_in[0][2][3] )
         );
  dff_sg \reg_in_reg[0][2][2]  ( .D(n15291), .CP(clk), .Q(\reg_in[0][2][2] )
         );
  dff_sg \reg_in_reg[0][2][1]  ( .D(n15290), .CP(clk), .Q(\reg_in[0][2][1] )
         );
  dff_sg \reg_in_reg[0][2][0]  ( .D(n15258), .CP(clk), .Q(\reg_in[0][2][0] )
         );
  dff_sg \reg_in_reg[0][1][19]  ( .D(n15257), .CP(clk), .Q(\reg_in[0][1][19] )
         );
  dff_sg \reg_in_reg[0][1][18]  ( .D(n15261), .CP(clk), .Q(\reg_in[0][1][18] )
         );
  dff_sg \reg_in_reg[0][1][17]  ( .D(n15260), .CP(clk), .Q(\reg_in[0][1][17] )
         );
  dff_sg \reg_in_reg[0][1][16]  ( .D(n15252), .CP(clk), .Q(\reg_in[0][1][16] )
         );
  dff_sg \reg_in_reg[0][1][15]  ( .D(n15251), .CP(clk), .Q(\reg_in[0][1][15] )
         );
  dff_sg \reg_in_reg[0][1][14]  ( .D(n15255), .CP(clk), .Q(\reg_in[0][1][14] )
         );
  dff_sg \reg_in_reg[0][1][13]  ( .D(n15254), .CP(clk), .Q(\reg_in[0][1][13] )
         );
  dff_sg \reg_in_reg[0][1][12]  ( .D(n15270), .CP(clk), .Q(\reg_in[0][1][12] )
         );
  dff_sg \reg_in_reg[0][1][11]  ( .D(n15269), .CP(clk), .Q(\reg_in[0][1][11] )
         );
  dff_sg \reg_in_reg[0][1][10]  ( .D(n15273), .CP(clk), .Q(\reg_in[0][1][10] )
         );
  dff_sg \reg_in_reg[0][1][9]  ( .D(n15272), .CP(clk), .Q(\reg_in[0][1][9] )
         );
  dff_sg \reg_in_reg[0][1][8]  ( .D(n15264), .CP(clk), .Q(\reg_in[0][1][8] )
         );
  dff_sg \reg_in_reg[0][1][7]  ( .D(n15263), .CP(clk), .Q(\reg_in[0][1][7] )
         );
  dff_sg \reg_in_reg[0][1][6]  ( .D(n15267), .CP(clk), .Q(\reg_in[0][1][6] )
         );
  dff_sg \reg_in_reg[0][1][5]  ( .D(n15266), .CP(clk), .Q(\reg_in[0][1][5] )
         );
  dff_sg \reg_in_reg[0][1][4]  ( .D(n15330), .CP(clk), .Q(\reg_in[0][1][4] )
         );
  dff_sg \reg_in_reg[0][1][3]  ( .D(n15329), .CP(clk), .Q(\reg_in[0][1][3] )
         );
  dff_sg \reg_in_reg[0][1][2]  ( .D(n15333), .CP(clk), .Q(\reg_in[0][1][2] )
         );
  dff_sg \reg_in_reg[0][1][1]  ( .D(n15332), .CP(clk), .Q(\reg_in[0][1][1] )
         );
  dff_sg \reg_in_reg[0][1][0]  ( .D(n15324), .CP(clk), .Q(\reg_in[0][1][0] )
         );
  dff_sg \reg_in_reg[0][0][19]  ( .D(n15323), .CP(clk), .Q(\reg_in[0][0][19] )
         );
  dff_sg \reg_in_reg[0][0][18]  ( .D(n15327), .CP(clk), .Q(\reg_in[0][0][18] )
         );
  dff_sg \reg_in_reg[0][0][17]  ( .D(n15326), .CP(clk), .Q(\reg_in[0][0][17] )
         );
  dff_sg \reg_in_reg[0][0][16]  ( .D(n15342), .CP(clk), .Q(\reg_in[0][0][16] )
         );
  dff_sg \reg_in_reg[0][0][15]  ( .D(n15341), .CP(clk), .Q(\reg_in[0][0][15] )
         );
  dff_sg \reg_in_reg[0][0][14]  ( .D(n15345), .CP(clk), .Q(\reg_in[0][0][14] )
         );
  dff_sg \reg_in_reg[0][0][13]  ( .D(n15344), .CP(clk), .Q(\reg_in[0][0][13] )
         );
  dff_sg \reg_in_reg[0][0][12]  ( .D(n15336), .CP(clk), .Q(\reg_in[0][0][12] )
         );
  dff_sg \reg_in_reg[0][0][11]  ( .D(n15335), .CP(clk), .Q(\reg_in[0][0][11] )
         );
  dff_sg \reg_in_reg[0][0][10]  ( .D(n15339), .CP(clk), .Q(\reg_in[0][0][10] )
         );
  dff_sg \reg_in_reg[0][0][9]  ( .D(n15338), .CP(clk), .Q(\reg_in[0][0][9] )
         );
  dff_sg \reg_in_reg[0][0][8]  ( .D(n15306), .CP(clk), .Q(\reg_in[0][0][8] )
         );
  dff_sg \reg_in_reg[0][0][7]  ( .D(n15305), .CP(clk), .Q(\reg_in[0][0][7] )
         );
  dff_sg \reg_in_reg[0][0][6]  ( .D(n15309), .CP(clk), .Q(\reg_in[0][0][6] )
         );
  dff_sg \reg_in_reg[0][0][5]  ( .D(n15308), .CP(clk), .Q(\reg_in[0][0][5] )
         );
  dff_sg \reg_in_reg[0][0][4]  ( .D(n15300), .CP(clk), .Q(\reg_in[0][0][4] )
         );
  dff_sg \reg_in_reg[0][0][3]  ( .D(n15299), .CP(clk), .Q(\reg_in[0][0][3] )
         );
  dff_sg \reg_in_reg[0][0][2]  ( .D(n15303), .CP(clk), .Q(\reg_in[0][0][2] )
         );
  dff_sg \reg_in_reg[0][0][1]  ( .D(n15302), .CP(clk), .Q(\reg_in[0][0][1] )
         );
  dff_sg \reg_in_reg[0][0][0]  ( .D(n15318), .CP(clk), .Q(\reg_in[0][0][0] )
         );
  dff_sg \out_reg[3][3][19]  ( .D(n14921), .CP(clk), .Q(n18402) );
  dff_sg \out_reg[3][3][18]  ( .D(n14821), .CP(clk), .Q(n18403) );
  dff_sg \out_reg[3][3][17]  ( .D(n14879), .CP(clk), .Q(n18404) );
  dff_sg \out_reg[3][3][16]  ( .D(n14876), .CP(clk), .Q(n18405) );
  dff_sg \out_reg[3][3][15]  ( .D(n14867), .CP(clk), .Q(n18406) );
  dff_sg \out_reg[3][3][14]  ( .D(n14822), .CP(clk), .Q(n18407) );
  dff_sg \out_reg[3][3][13]  ( .D(n14864), .CP(clk), .Q(n18408) );
  dff_sg \out_reg[3][3][12]  ( .D(n14861), .CP(clk), .Q(n18409) );
  dff_sg \out_reg[3][3][11]  ( .D(n14894), .CP(clk), .Q(n18410) );
  dff_sg \out_reg[3][3][10]  ( .D(n14918), .CP(clk), .Q(n18411) );
  dff_sg \out_reg[3][3][9]  ( .D(n14888), .CP(clk), .Q(n18412) );
  dff_sg \out_reg[3][3][8]  ( .D(n14885), .CP(clk), .Q(n18413) );
  dff_sg \out_reg[3][3][7]  ( .D(n14915), .CP(clk), .Q(n18414) );
  dff_sg \out_reg[3][3][6]  ( .D(n14912), .CP(clk), .Q(n18415) );
  dff_sg \out_reg[3][3][5]  ( .D(n14903), .CP(clk), .Q(n18416) );
  dff_sg \out_reg[3][3][4]  ( .D(n14900), .CP(clk), .Q(n18417) );
  dff_sg \out_reg[3][3][3]  ( .D(n15093), .CP(clk), .Q(n18418) );
  dff_sg \out_reg[3][3][2]  ( .D(n14809), .CP(clk), .Q(n18419) );
  dff_sg \out_reg[3][3][1]  ( .D(n15078), .CP(clk), .Q(n18420) );
  dff_sg \out_reg[3][3][0]  ( .D(n15075), .CP(clk), .Q(n18421) );
  dff_sg \out_reg[3][2][19]  ( .D(n15117), .CP(clk), .Q(n18422) );
  dff_sg \out_reg[3][2][18]  ( .D(n14840), .CP(clk), .Q(n18423) );
  dff_sg \out_reg[3][2][17]  ( .D(n15111), .CP(clk), .Q(n18424) );
  dff_sg \out_reg[3][2][16]  ( .D(n15108), .CP(clk), .Q(n18425) );
  dff_sg \out_reg[3][2][15]  ( .D(n14852), .CP(clk), .Q(n18426) );
  dff_sg \out_reg[3][2][14]  ( .D(n14805), .CP(clk), .Q(n18427) );
  dff_sg \out_reg[3][2][13]  ( .D(n14846), .CP(clk), .Q(n18428) );
  dff_sg \out_reg[3][2][12]  ( .D(n14843), .CP(clk), .Q(n18429) );
  dff_sg \out_reg[3][2][11]  ( .D(n15084), .CP(clk), .Q(n18430) );
  dff_sg \out_reg[3][2][10]  ( .D(n15087), .CP(clk), .Q(n18431) );
  dff_sg \out_reg[3][2][9]  ( .D(n14804), .CP(clk), .Q(n18432) );
  dff_sg \out_reg[3][2][8]  ( .D(n14803), .CP(clk), .Q(n18433) );
  dff_sg \out_reg[3][2][7]  ( .D(n14827), .CP(clk), .Q(n18434) );
  dff_sg \out_reg[3][2][6]  ( .D(n14826), .CP(clk), .Q(n18435) );
  dff_sg \out_reg[3][2][5]  ( .D(n14830), .CP(clk), .Q(n18436) );
  dff_sg \out_reg[3][2][4]  ( .D(n14829), .CP(clk), .Q(n18437) );
  dff_sg \out_reg[3][2][3]  ( .D(n14993), .CP(clk), .Q(n18438) );
  dff_sg \out_reg[3][2][2]  ( .D(n14990), .CP(clk), .Q(n18439) );
  dff_sg \out_reg[3][2][1]  ( .D(n14984), .CP(clk), .Q(n18440) );
  dff_sg \out_reg[3][2][0]  ( .D(n14981), .CP(clk), .Q(n18441) );
  dff_sg \out_reg[3][1][19]  ( .D(n15008), .CP(clk), .Q(n18442) );
  dff_sg \out_reg[3][1][18]  ( .D(n14833), .CP(clk), .Q(n18443) );
  dff_sg \out_reg[3][1][17]  ( .D(n15005), .CP(clk), .Q(n18444) );
  dff_sg \out_reg[3][1][16]  ( .D(n15002), .CP(clk), .Q(n18445) );
  dff_sg \out_reg[3][1][15]  ( .D(n15023), .CP(clk), .Q(n18446) );
  dff_sg \out_reg[3][1][14]  ( .D(n14832), .CP(clk), .Q(n18447) );
  dff_sg \out_reg[3][1][13]  ( .D(n15020), .CP(clk), .Q(n18448) );
  dff_sg \out_reg[3][1][12]  ( .D(n15017), .CP(clk), .Q(n18449) );
  dff_sg \out_reg[3][1][11]  ( .D(n14936), .CP(clk), .Q(n18450) );
  dff_sg \out_reg[3][1][10]  ( .D(n14933), .CP(clk), .Q(n18451) );
  dff_sg \out_reg[3][1][9]  ( .D(n14930), .CP(clk), .Q(n18452) );
  dff_sg \out_reg[3][1][8]  ( .D(n14927), .CP(clk), .Q(n18453) );
  dff_sg \out_reg[3][1][7]  ( .D(n14954), .CP(clk), .Q(n18454) );
  dff_sg \out_reg[3][1][6]  ( .D(n14951), .CP(clk), .Q(n18455) );
  dff_sg \out_reg[3][1][5]  ( .D(n14945), .CP(clk), .Q(n18456) );
  dff_sg \out_reg[3][1][4]  ( .D(n14942), .CP(clk), .Q(n18457) );
  dff_sg \out_reg[3][1][3]  ( .D(n14978), .CP(clk), .Q(n18458) );
  dff_sg \out_reg[3][1][2]  ( .D(n14975), .CP(clk), .Q(n18459) );
  dff_sg \out_reg[3][1][1]  ( .D(n14972), .CP(clk), .Q(n18460) );
  dff_sg \out_reg[3][1][0]  ( .D(n14969), .CP(clk), .Q(n18461) );
  dff_sg \out_reg[3][0][19]  ( .D(n14818), .CP(clk), .Q(n18462) );
  dff_sg \out_reg[3][0][18]  ( .D(n14817), .CP(clk), .Q(n18463) );
  dff_sg \out_reg[3][0][17]  ( .D(n14963), .CP(clk), .Q(n18464) );
  dff_sg \out_reg[3][0][16]  ( .D(n14960), .CP(clk), .Q(n18465) );
  dff_sg \out_reg[3][0][15]  ( .D(n15014), .CP(clk), .Q(n18466) );
  dff_sg \out_reg[3][0][14]  ( .D(n14831), .CP(clk), .Q(n18467) );
  dff_sg \out_reg[3][0][13]  ( .D(n14828), .CP(clk), .Q(n18468) );
  dff_sg \out_reg[3][0][12]  ( .D(n14825), .CP(clk), .Q(n18469) );
  dff_sg \out_reg[3][0][11]  ( .D(n15033), .CP(clk), .Q(n18470) );
  dff_sg \out_reg[3][0][10]  ( .D(n14823), .CP(clk), .Q(n18471) );
  dff_sg \out_reg[3][0][9]  ( .D(n15066), .CP(clk), .Q(n18472) );
  dff_sg \out_reg[3][0][8]  ( .D(n14999), .CP(clk), .Q(n18473) );
  dff_sg \out_reg[3][0][7]  ( .D(n15105), .CP(clk), .Q(n18474) );
  dff_sg \out_reg[3][0][6]  ( .D(n15048), .CP(clk), .Q(n18475) );
  dff_sg \out_reg[3][0][5]  ( .D(n15042), .CP(clk), .Q(n18476) );
  dff_sg \out_reg[3][0][4]  ( .D(n15060), .CP(clk), .Q(n18477) );
  dff_sg \out_reg[3][0][3]  ( .D(n15045), .CP(clk), .Q(n18478) );
  dff_sg \out_reg[3][0][2]  ( .D(n15072), .CP(clk), .Q(n18479) );
  dff_sg \out_reg[3][0][1]  ( .D(n15039), .CP(clk), .Q(n18480) );
  dff_sg \out_reg[3][0][0]  ( .D(n15036), .CP(clk), .Q(n18481) );
  dff_sg \out_reg[2][3][19]  ( .D(n14924), .CP(clk), .Q(n18482) );
  dff_sg \out_reg[2][3][18]  ( .D(n14812), .CP(clk), .Q(n18483) );
  dff_sg \out_reg[2][3][17]  ( .D(n14957), .CP(clk), .Q(n18484) );
  dff_sg \out_reg[2][3][16]  ( .D(n14939), .CP(clk), .Q(n18485) );
  dff_sg \out_reg[2][3][15]  ( .D(n14811), .CP(clk), .Q(n18486) );
  dff_sg \out_reg[2][3][14]  ( .D(n14810), .CP(clk), .Q(n18487) );
  dff_sg \out_reg[2][3][13]  ( .D(n14815), .CP(clk), .Q(n18488) );
  dff_sg \out_reg[2][3][12]  ( .D(n14819), .CP(clk), .Q(n18489) );
  dff_sg \out_reg[2][3][11]  ( .D(n15120), .CP(clk), .Q(n18490) );
  dff_sg \out_reg[2][3][10]  ( .D(n14814), .CP(clk), .Q(n18491) );
  dff_sg \out_reg[2][3][9]  ( .D(n14816), .CP(clk), .Q(n18492) );
  dff_sg \out_reg[2][3][8]  ( .D(n15011), .CP(clk), .Q(n18493) );
  dff_sg \out_reg[2][3][7]  ( .D(n15063), .CP(clk), .Q(n18494) );
  dff_sg \out_reg[2][3][6]  ( .D(n14813), .CP(clk), .Q(n18495) );
  dff_sg \out_reg[2][3][5]  ( .D(n14824), .CP(clk), .Q(n18496) );
  dff_sg \out_reg[2][3][4]  ( .D(n14966), .CP(clk), .Q(n18497) );
  dff_sg \out_reg[2][3][3]  ( .D(n15096), .CP(clk), .Q(n18498) );
  dff_sg \out_reg[2][3][2]  ( .D(n15069), .CP(clk), .Q(n18499) );
  dff_sg \out_reg[2][3][1]  ( .D(n15057), .CP(clk), .Q(n18500) );
  dff_sg \out_reg[2][3][0]  ( .D(n15054), .CP(clk), .Q(n18501) );
  dff_sg \out_reg[2][2][19]  ( .D(n15114), .CP(clk), .Q(n18502) );
  dff_sg \out_reg[2][2][18]  ( .D(n14996), .CP(clk), .Q(n18503) );
  dff_sg \out_reg[2][2][17]  ( .D(n15030), .CP(clk), .Q(n18504) );
  dff_sg \out_reg[2][2][16]  ( .D(n15027), .CP(clk), .Q(n18505) );
  dff_sg \out_reg[2][2][15]  ( .D(n14855), .CP(clk), .Q(n18506) );
  dff_sg \out_reg[2][2][14]  ( .D(n14873), .CP(clk), .Q(n18507) );
  dff_sg \out_reg[2][2][13]  ( .D(n14834), .CP(clk), .Q(n18508) );
  dff_sg \out_reg[2][2][12]  ( .D(n15081), .CP(clk), .Q(n18509) );
  dff_sg \out_reg[2][2][11]  ( .D(n14891), .CP(clk), .Q(n18510) );
  dff_sg \out_reg[2][2][10]  ( .D(n14807), .CP(clk), .Q(n18511) );
  dff_sg \out_reg[2][2][9]  ( .D(n14906), .CP(clk), .Q(n18512) );
  dff_sg \out_reg[2][2][8]  ( .D(n14909), .CP(clk), .Q(n18513) );
  dff_sg \out_reg[2][2][7]  ( .D(n14808), .CP(clk), .Q(n18514) );
  dff_sg \out_reg[2][2][6]  ( .D(n14849), .CP(clk), .Q(n18515) );
  dff_sg \out_reg[2][2][5]  ( .D(n14806), .CP(clk), .Q(n18516) );
  dff_sg \out_reg[2][2][4]  ( .D(n15051), .CP(clk), .Q(n18517) );
  dff_sg \out_reg[2][2][3]  ( .D(n14987), .CP(clk), .Q(n18518) );
  dff_sg \out_reg[2][2][2]  ( .D(n15099), .CP(clk), .Q(n18519) );
  dff_sg \out_reg[2][2][1]  ( .D(n15090), .CP(clk), .Q(n18520) );
  dff_sg \out_reg[2][2][0]  ( .D(n14948), .CP(clk), .Q(n18521) );
  dff_sg \out_reg[2][1][19]  ( .D(n14897), .CP(clk), .Q(n18522) );
  dff_sg \out_reg[2][1][18]  ( .D(n14882), .CP(clk), .Q(n18523) );
  dff_sg \out_reg[2][1][17]  ( .D(n14858), .CP(clk), .Q(n18524) );
  dff_sg \out_reg[2][1][16]  ( .D(n14820), .CP(clk), .Q(n18525) );
  dff_sg \out_reg[2][1][15]  ( .D(n15026), .CP(clk), .Q(n18526) );
  dff_sg \out_reg[2][1][14]  ( .D(n14870), .CP(clk), .Q(n18527) );
  dff_sg \out_reg[2][1][13]  ( .D(n15102), .CP(clk), .Q(n18528) );
  dff_sg \out_reg[2][1][12]  ( .D(n14837), .CP(clk), .Q(n18529) );
  dff_sg \out_reg[2][1][11]  ( .D(n14962), .CP(clk), .Q(n18530) );
  dff_sg \out_reg[2][1][10]  ( .D(n14961), .CP(clk), .Q(n18531) );
  dff_sg \out_reg[2][1][9]  ( .D(n14965), .CP(clk), .Q(n18532) );
  dff_sg \out_reg[2][1][8]  ( .D(n14964), .CP(clk), .Q(n18533) );
  dff_sg \out_reg[2][1][7]  ( .D(n14956), .CP(clk), .Q(n18534) );
  dff_sg \out_reg[2][1][6]  ( .D(n14955), .CP(clk), .Q(n18535) );
  dff_sg \out_reg[2][1][5]  ( .D(n14959), .CP(clk), .Q(n18536) );
  dff_sg \out_reg[2][1][4]  ( .D(n14958), .CP(clk), .Q(n18537) );
  dff_sg \out_reg[2][1][3]  ( .D(n14974), .CP(clk), .Q(n18538) );
  dff_sg \out_reg[2][1][2]  ( .D(n14973), .CP(clk), .Q(n18539) );
  dff_sg \out_reg[2][1][1]  ( .D(n14977), .CP(clk), .Q(n18540) );
  dff_sg \out_reg[2][1][0]  ( .D(n14976), .CP(clk), .Q(n18541) );
  dff_sg \out_reg[2][0][19]  ( .D(n14968), .CP(clk), .Q(n18542) );
  dff_sg \out_reg[2][0][18]  ( .D(n14967), .CP(clk), .Q(n18543) );
  dff_sg \out_reg[2][0][17]  ( .D(n14971), .CP(clk), .Q(n18544) );
  dff_sg \out_reg[2][0][16]  ( .D(n14970), .CP(clk), .Q(n18545) );
  dff_sg \out_reg[2][0][15]  ( .D(n14938), .CP(clk), .Q(n18546) );
  dff_sg \out_reg[2][0][14]  ( .D(n14937), .CP(clk), .Q(n18547) );
  dff_sg \out_reg[2][0][13]  ( .D(n14941), .CP(clk), .Q(n18548) );
  dff_sg \out_reg[2][0][12]  ( .D(n14940), .CP(clk), .Q(n18549) );
  dff_sg \out_reg[2][0][11]  ( .D(n14932), .CP(clk), .Q(n18550) );
  dff_sg \out_reg[2][0][10]  ( .D(n14931), .CP(clk), .Q(n18551) );
  dff_sg \out_reg[2][0][9]  ( .D(n14935), .CP(clk), .Q(n18552) );
  dff_sg \out_reg[2][0][8]  ( .D(n14934), .CP(clk), .Q(n18553) );
  dff_sg \out_reg[2][0][7]  ( .D(n14950), .CP(clk), .Q(n18554) );
  dff_sg \out_reg[2][0][6]  ( .D(n14949), .CP(clk), .Q(n18555) );
  dff_sg \out_reg[2][0][5]  ( .D(n14953), .CP(clk), .Q(n18556) );
  dff_sg \out_reg[2][0][4]  ( .D(n14952), .CP(clk), .Q(n18557) );
  dff_sg \out_reg[2][0][3]  ( .D(n14944), .CP(clk), .Q(n18558) );
  dff_sg \out_reg[2][0][2]  ( .D(n14943), .CP(clk), .Q(n18559) );
  dff_sg \out_reg[2][0][1]  ( .D(n14947), .CP(clk), .Q(n18560) );
  dff_sg \out_reg[2][0][0]  ( .D(n14946), .CP(clk), .Q(n18561) );
  dff_sg \out_reg[1][3][19]  ( .D(n15010), .CP(clk), .Q(n18562) );
  dff_sg \out_reg[1][3][18]  ( .D(n15009), .CP(clk), .Q(n18563) );
  dff_sg \out_reg[1][3][17]  ( .D(n15013), .CP(clk), .Q(n18564) );
  dff_sg \out_reg[1][3][16]  ( .D(n15012), .CP(clk), .Q(n18565) );
  dff_sg \out_reg[1][3][15]  ( .D(n15004), .CP(clk), .Q(n18566) );
  dff_sg \out_reg[1][3][14]  ( .D(n15003), .CP(clk), .Q(n18567) );
  dff_sg \out_reg[1][3][13]  ( .D(n15007), .CP(clk), .Q(n18568) );
  dff_sg \out_reg[1][3][12]  ( .D(n15006), .CP(clk), .Q(n18569) );
  dff_sg \out_reg[1][3][11]  ( .D(n15022), .CP(clk), .Q(n18570) );
  dff_sg \out_reg[1][3][10]  ( .D(n15021), .CP(clk), .Q(n18571) );
  dff_sg \out_reg[1][3][9]  ( .D(n15025), .CP(clk), .Q(n18572) );
  dff_sg \out_reg[1][3][8]  ( .D(n15024), .CP(clk), .Q(n18573) );
  dff_sg \out_reg[1][3][7]  ( .D(n15016), .CP(clk), .Q(n18574) );
  dff_sg \out_reg[1][3][6]  ( .D(n15015), .CP(clk), .Q(n18575) );
  dff_sg \out_reg[1][3][5]  ( .D(n15019), .CP(clk), .Q(n18576) );
  dff_sg \out_reg[1][3][4]  ( .D(n15018), .CP(clk), .Q(n18577) );
  dff_sg \out_reg[1][3][3]  ( .D(n14986), .CP(clk), .Q(n18578) );
  dff_sg \out_reg[1][3][2]  ( .D(n14985), .CP(clk), .Q(n18579) );
  dff_sg \out_reg[1][3][1]  ( .D(n14989), .CP(clk), .Q(n18580) );
  dff_sg \out_reg[1][3][0]  ( .D(n14988), .CP(clk), .Q(n18581) );
  dff_sg \out_reg[1][2][19]  ( .D(n14980), .CP(clk), .Q(n18582) );
  dff_sg \out_reg[1][2][18]  ( .D(n14979), .CP(clk), .Q(n18583) );
  dff_sg \out_reg[1][2][17]  ( .D(n14983), .CP(clk), .Q(n18584) );
  dff_sg \out_reg[1][2][16]  ( .D(n14982), .CP(clk), .Q(n18585) );
  dff_sg \out_reg[1][2][15]  ( .D(n14998), .CP(clk), .Q(n18586) );
  dff_sg \out_reg[1][2][14]  ( .D(n14997), .CP(clk), .Q(n18587) );
  dff_sg \out_reg[1][2][13]  ( .D(n15001), .CP(clk), .Q(n18588) );
  dff_sg \out_reg[1][2][12]  ( .D(n15000), .CP(clk), .Q(n18589) );
  dff_sg \out_reg[1][2][11]  ( .D(n14992), .CP(clk), .Q(n18590) );
  dff_sg \out_reg[1][2][10]  ( .D(n14991), .CP(clk), .Q(n18591) );
  dff_sg \out_reg[1][2][9]  ( .D(n14995), .CP(clk), .Q(n18592) );
  dff_sg \out_reg[1][2][8]  ( .D(n14994), .CP(clk), .Q(n18593) );
  dff_sg \out_reg[1][2][7]  ( .D(n14866), .CP(clk), .Q(n18594) );
  dff_sg \out_reg[1][2][6]  ( .D(n14865), .CP(clk), .Q(n18595) );
  dff_sg \out_reg[1][2][5]  ( .D(n14869), .CP(clk), .Q(n18596) );
  dff_sg \out_reg[1][2][4]  ( .D(n14868), .CP(clk), .Q(n18597) );
  dff_sg \out_reg[1][2][3]  ( .D(n14860), .CP(clk), .Q(n18598) );
  dff_sg \out_reg[1][2][2]  ( .D(n14859), .CP(clk), .Q(n18599) );
  dff_sg \out_reg[1][2][1]  ( .D(n14863), .CP(clk), .Q(n18600) );
  dff_sg \out_reg[1][2][0]  ( .D(n14862), .CP(clk), .Q(n18601) );
  dff_sg \out_reg[1][1][19]  ( .D(n14878), .CP(clk), .Q(n18602) );
  dff_sg \out_reg[1][1][18]  ( .D(n14877), .CP(clk), .Q(n18603) );
  dff_sg \out_reg[1][1][17]  ( .D(n14881), .CP(clk), .Q(n18604) );
  dff_sg \out_reg[1][1][16]  ( .D(n14880), .CP(clk), .Q(n18605) );
  dff_sg \out_reg[1][1][15]  ( .D(n14872), .CP(clk), .Q(n18606) );
  dff_sg \out_reg[1][1][14]  ( .D(n14871), .CP(clk), .Q(n18607) );
  dff_sg \out_reg[1][1][13]  ( .D(n14875), .CP(clk), .Q(n18608) );
  dff_sg \out_reg[1][1][12]  ( .D(n14874), .CP(clk), .Q(n18609) );
  dff_sg \out_reg[1][1][11]  ( .D(n14842), .CP(clk), .Q(n18610) );
  dff_sg \out_reg[1][1][10]  ( .D(n14841), .CP(clk), .Q(n18611) );
  dff_sg \out_reg[1][1][9]  ( .D(n14845), .CP(clk), .Q(n18612) );
  dff_sg \out_reg[1][1][8]  ( .D(n14844), .CP(clk), .Q(n18613) );
  dff_sg \out_reg[1][1][7]  ( .D(n14836), .CP(clk), .Q(n18614) );
  dff_sg \out_reg[1][1][6]  ( .D(n14835), .CP(clk), .Q(n18615) );
  dff_sg \out_reg[1][1][5]  ( .D(n14839), .CP(clk), .Q(n18616) );
  dff_sg \out_reg[1][1][4]  ( .D(n14838), .CP(clk), .Q(n18617) );
  dff_sg \out_reg[1][1][3]  ( .D(n14854), .CP(clk), .Q(n18618) );
  dff_sg \out_reg[1][1][2]  ( .D(n14853), .CP(clk), .Q(n18619) );
  dff_sg \out_reg[1][1][1]  ( .D(n14857), .CP(clk), .Q(n18620) );
  dff_sg \out_reg[1][1][0]  ( .D(n14856), .CP(clk), .Q(n18621) );
  dff_sg \out_reg[1][0][19]  ( .D(n14848), .CP(clk), .Q(n18622) );
  dff_sg \out_reg[1][0][18]  ( .D(n14847), .CP(clk), .Q(n18623) );
  dff_sg \out_reg[1][0][17]  ( .D(n14851), .CP(clk), .Q(n18624) );
  dff_sg \out_reg[1][0][16]  ( .D(n14850), .CP(clk), .Q(n18625) );
  dff_sg \out_reg[1][0][15]  ( .D(n14914), .CP(clk), .Q(n18626) );
  dff_sg \out_reg[1][0][14]  ( .D(n14913), .CP(clk), .Q(n18627) );
  dff_sg \out_reg[1][0][13]  ( .D(n14917), .CP(clk), .Q(n18628) );
  dff_sg \out_reg[1][0][12]  ( .D(n14916), .CP(clk), .Q(n18629) );
  dff_sg \out_reg[1][0][11]  ( .D(n14908), .CP(clk), .Q(n18630) );
  dff_sg \out_reg[1][0][10]  ( .D(n14907), .CP(clk), .Q(n18631) );
  dff_sg \out_reg[1][0][9]  ( .D(n14911), .CP(clk), .Q(n18632) );
  dff_sg \out_reg[1][0][8]  ( .D(n14910), .CP(clk), .Q(n18633) );
  dff_sg \out_reg[1][0][7]  ( .D(n14926), .CP(clk), .Q(n18634) );
  dff_sg \out_reg[1][0][6]  ( .D(n14925), .CP(clk), .Q(n18635) );
  dff_sg \out_reg[1][0][5]  ( .D(n14929), .CP(clk), .Q(n18636) );
  dff_sg \out_reg[1][0][4]  ( .D(n14928), .CP(clk), .Q(n18637) );
  dff_sg \out_reg[1][0][3]  ( .D(n14920), .CP(clk), .Q(n18638) );
  dff_sg \out_reg[1][0][2]  ( .D(n14919), .CP(clk), .Q(n18639) );
  dff_sg \out_reg[1][0][1]  ( .D(n14923), .CP(clk), .Q(n18640) );
  dff_sg \out_reg[1][0][0]  ( .D(n14922), .CP(clk), .Q(n18641) );
  dff_sg \out_reg[0][3][19]  ( .D(n14890), .CP(clk), .Q(n18642) );
  dff_sg \out_reg[0][3][18]  ( .D(n14889), .CP(clk), .Q(n18643) );
  dff_sg \out_reg[0][3][17]  ( .D(n14893), .CP(clk), .Q(n18644) );
  dff_sg \out_reg[0][3][16]  ( .D(n14892), .CP(clk), .Q(n18645) );
  dff_sg \out_reg[0][3][15]  ( .D(n14884), .CP(clk), .Q(n18646) );
  dff_sg \out_reg[0][3][14]  ( .D(n14883), .CP(clk), .Q(n18647) );
  dff_sg \out_reg[0][3][13]  ( .D(n14887), .CP(clk), .Q(n18648) );
  dff_sg \out_reg[0][3][12]  ( .D(n14886), .CP(clk), .Q(n18649) );
  dff_sg \out_reg[0][3][11]  ( .D(n14902), .CP(clk), .Q(n18650) );
  dff_sg \out_reg[0][3][10]  ( .D(n14901), .CP(clk), .Q(n18651) );
  dff_sg \out_reg[0][3][9]  ( .D(n14905), .CP(clk), .Q(n18652) );
  dff_sg \out_reg[0][3][8]  ( .D(n14904), .CP(clk), .Q(n18653) );
  dff_sg \out_reg[0][3][7]  ( .D(n14896), .CP(clk), .Q(n18654) );
  dff_sg \out_reg[0][3][6]  ( .D(n14895), .CP(clk), .Q(n18655) );
  dff_sg \out_reg[0][3][5]  ( .D(n14899), .CP(clk), .Q(n18656) );
  dff_sg \out_reg[0][3][4]  ( .D(n14898), .CP(clk), .Q(n18657) );
  dff_sg \out_reg[0][3][3]  ( .D(n15059), .CP(clk), .Q(n18658) );
  dff_sg \out_reg[0][3][2]  ( .D(n15058), .CP(clk), .Q(n18659) );
  dff_sg \out_reg[0][3][1]  ( .D(n15062), .CP(clk), .Q(n18660) );
  dff_sg \out_reg[0][3][0]  ( .D(n15061), .CP(clk), .Q(n18661) );
  dff_sg \out_reg[0][2][19]  ( .D(n15053), .CP(clk), .Q(n18662) );
  dff_sg \out_reg[0][2][18]  ( .D(n15052), .CP(clk), .Q(n18663) );
  dff_sg \out_reg[0][2][17]  ( .D(n15056), .CP(clk), .Q(n18664) );
  dff_sg \out_reg[0][2][16]  ( .D(n15055), .CP(clk), .Q(n18665) );
  dff_sg \out_reg[0][2][15]  ( .D(n15071), .CP(clk), .Q(n18666) );
  dff_sg \out_reg[0][2][14]  ( .D(n15070), .CP(clk), .Q(n18667) );
  dff_sg \out_reg[0][2][13]  ( .D(n15074), .CP(clk), .Q(n18668) );
  dff_sg \out_reg[0][2][12]  ( .D(n15073), .CP(clk), .Q(n18669) );
  dff_sg \out_reg[0][2][11]  ( .D(n15065), .CP(clk), .Q(n18670) );
  dff_sg \out_reg[0][2][10]  ( .D(n15064), .CP(clk), .Q(n18671) );
  dff_sg \out_reg[0][2][9]  ( .D(n15068), .CP(clk), .Q(n18672) );
  dff_sg \out_reg[0][2][8]  ( .D(n15067), .CP(clk), .Q(n18673) );
  dff_sg \out_reg[0][2][7]  ( .D(n15035), .CP(clk), .Q(n18674) );
  dff_sg \out_reg[0][2][6]  ( .D(n15034), .CP(clk), .Q(n18675) );
  dff_sg \out_reg[0][2][5]  ( .D(n15038), .CP(clk), .Q(n18676) );
  dff_sg \out_reg[0][2][4]  ( .D(n15037), .CP(clk), .Q(n18677) );
  dff_sg \out_reg[0][2][3]  ( .D(n15029), .CP(clk), .Q(n18678) );
  dff_sg \out_reg[0][2][2]  ( .D(n15028), .CP(clk), .Q(n18679) );
  dff_sg \out_reg[0][2][1]  ( .D(n15032), .CP(clk), .Q(n18680) );
  dff_sg \out_reg[0][2][0]  ( .D(n15031), .CP(clk), .Q(n18681) );
  dff_sg \out_reg[0][1][19]  ( .D(n15047), .CP(clk), .Q(n18682) );
  dff_sg \out_reg[0][1][18]  ( .D(n15046), .CP(clk), .Q(n18683) );
  dff_sg \out_reg[0][1][17]  ( .D(n15050), .CP(clk), .Q(n18684) );
  dff_sg \out_reg[0][1][16]  ( .D(n15049), .CP(clk), .Q(n18685) );
  dff_sg \out_reg[0][1][15]  ( .D(n15041), .CP(clk), .Q(n18686) );
  dff_sg \out_reg[0][1][14]  ( .D(n15040), .CP(clk), .Q(n18687) );
  dff_sg \out_reg[0][1][13]  ( .D(n15044), .CP(clk), .Q(n18688) );
  dff_sg \out_reg[0][1][12]  ( .D(n15043), .CP(clk), .Q(n18689) );
  dff_sg \out_reg[0][1][11]  ( .D(n15107), .CP(clk), .Q(n18690) );
  dff_sg \out_reg[0][1][10]  ( .D(n15106), .CP(clk), .Q(n18691) );
  dff_sg \out_reg[0][1][9]  ( .D(n15110), .CP(clk), .Q(n18692) );
  dff_sg \out_reg[0][1][8]  ( .D(n15109), .CP(clk), .Q(n18693) );
  dff_sg \out_reg[0][1][7]  ( .D(n15101), .CP(clk), .Q(n18694) );
  dff_sg \out_reg[0][1][6]  ( .D(n15100), .CP(clk), .Q(n18695) );
  dff_sg \out_reg[0][1][5]  ( .D(n15104), .CP(clk), .Q(n18696) );
  dff_sg \out_reg[0][1][4]  ( .D(n15103), .CP(clk), .Q(n18697) );
  dff_sg \out_reg[0][1][3]  ( .D(n15119), .CP(clk), .Q(n18698) );
  dff_sg \out_reg[0][1][2]  ( .D(n15118), .CP(clk), .Q(n18699) );
  dff_sg \out_reg[0][1][1]  ( .D(n15122), .CP(clk), .Q(n18700) );
  dff_sg \out_reg[0][1][0]  ( .D(n15121), .CP(clk), .Q(n18701) );
  dff_sg \out_reg[0][0][19]  ( .D(n15113), .CP(clk), .Q(n18702) );
  dff_sg \out_reg[0][0][18]  ( .D(n15112), .CP(clk), .Q(n18703) );
  dff_sg \out_reg[0][0][17]  ( .D(n15116), .CP(clk), .Q(n18704) );
  dff_sg \out_reg[0][0][16]  ( .D(n15115), .CP(clk), .Q(n18705) );
  dff_sg \out_reg[0][0][15]  ( .D(n15083), .CP(clk), .Q(n18706) );
  dff_sg \out_reg[0][0][14]  ( .D(n15082), .CP(clk), .Q(n18707) );
  dff_sg \out_reg[0][0][13]  ( .D(n15086), .CP(clk), .Q(n18708) );
  dff_sg \out_reg[0][0][12]  ( .D(n15085), .CP(clk), .Q(n18709) );
  dff_sg \out_reg[0][0][11]  ( .D(n15077), .CP(clk), .Q(n18710) );
  dff_sg \out_reg[0][0][10]  ( .D(n15076), .CP(clk), .Q(n18711) );
  dff_sg \out_reg[0][0][9]  ( .D(n15080), .CP(clk), .Q(n18712) );
  dff_sg \out_reg[0][0][8]  ( .D(n15079), .CP(clk), .Q(n18713) );
  dff_sg \out_reg[0][0][7]  ( .D(n15095), .CP(clk), .Q(n18714) );
  dff_sg \out_reg[0][0][6]  ( .D(n15094), .CP(clk), .Q(n18715) );
  dff_sg \out_reg[0][0][5]  ( .D(n15098), .CP(clk), .Q(n18716) );
  dff_sg \out_reg[0][0][4]  ( .D(n15097), .CP(clk), .Q(n18717) );
  dff_sg \out_reg[0][0][3]  ( .D(n15089), .CP(clk), .Q(n18718) );
  dff_sg \out_reg[0][0][2]  ( .D(n15088), .CP(clk), .Q(n18719) );
  dff_sg \out_reg[0][0][1]  ( .D(n15092), .CP(clk), .Q(n18720) );
  dff_sg \out_reg[0][0][0]  ( .D(n15091), .CP(clk), .Q(n18721) );
  \**FFGEN**  \reg_out_reg[3][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3873), .force_10(n18078), .force_11(1'b0), 
        .Q(n14802) );
  \**FFGEN**  \reg_out_reg[3][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3877), .force_10(n18079), .force_11(1'b0), 
        .Q(n14801) );
  \**FFGEN**  \reg_out_reg[3][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3881), .force_10(n18080), .force_11(1'b0), 
        .Q(n14800) );
  \**FFGEN**  \reg_out_reg[3][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3885), .force_10(n18081), .force_11(1'b0), 
        .Q(n14799) );
  \**FFGEN**  \reg_out_reg[3][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3889), .force_10(n18082), .force_11(1'b0), 
        .Q(n14798) );
  \**FFGEN**  \reg_out_reg[3][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3893), .force_10(n18083), .force_11(1'b0), 
        .Q(n14797) );
  \**FFGEN**  \reg_out_reg[3][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3897), .force_10(n18084), .force_11(1'b0), 
        .Q(n14796) );
  \**FFGEN**  \reg_out_reg[3][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3901), .force_10(n18085), .force_11(1'b0), 
        .Q(n14795) );
  \**FFGEN**  \reg_out_reg[3][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3905), .force_10(n18086), .force_11(1'b0), 
        .Q(n14794) );
  \**FFGEN**  \reg_out_reg[3][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3909), .force_10(n18087), .force_11(1'b0), 
        .Q(n14793) );
  \**FFGEN**  \reg_out_reg[3][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3913), .force_10(n18088), .force_11(1'b0), 
        .Q(n14792) );
  \**FFGEN**  \reg_out_reg[3][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3917), .force_10(n18089), .force_11(1'b0), 
        .Q(n14791) );
  \**FFGEN**  \reg_out_reg[3][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3921), .force_10(n18090), .force_11(1'b0), 
        .Q(n14790) );
  \**FFGEN**  \reg_out_reg[3][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3925), .force_10(n18091), .force_11(1'b0), 
        .Q(n14789) );
  \**FFGEN**  \reg_out_reg[3][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3929), .force_10(n18092), .force_11(1'b0), 
        .Q(n14788) );
  \**FFGEN**  \reg_out_reg[3][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3933), .force_10(n18093), .force_11(1'b0), 
        .Q(n14787) );
  \**FFGEN**  \reg_out_reg[3][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3937), .force_10(n18094), .force_11(1'b0), 
        .Q(n14786) );
  \**FFGEN**  \reg_out_reg[3][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3941), .force_10(n18095), .force_11(1'b0), 
        .Q(n14785) );
  \**FFGEN**  \reg_out_reg[3][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3945), .force_10(n18096), .force_11(1'b0), 
        .Q(n14784) );
  \**FFGEN**  \reg_out_reg[3][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3949), .force_10(n18097), .force_11(1'b0), 
        .Q(n14783) );
  \**FFGEN**  \reg_out_reg[3][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3953), .force_10(n18098), .force_11(1'b0), 
        .Q(n14782) );
  \**FFGEN**  \reg_out_reg[3][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3957), .force_10(n18099), .force_11(1'b0), 
        .Q(n14781) );
  \**FFGEN**  \reg_out_reg[3][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3961), .force_10(n18100), .force_11(1'b0), 
        .Q(n14780) );
  \**FFGEN**  \reg_out_reg[3][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3965), .force_10(n18101), .force_11(1'b0), 
        .Q(n14779) );
  \**FFGEN**  \reg_out_reg[3][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3969), .force_10(n18102), .force_11(1'b0), 
        .Q(n14778) );
  \**FFGEN**  \reg_out_reg[3][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3973), .force_10(n18103), .force_11(1'b0), 
        .Q(n14777) );
  \**FFGEN**  \reg_out_reg[3][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3977), .force_10(n18104), .force_11(1'b0), 
        .Q(n14776) );
  \**FFGEN**  \reg_out_reg[3][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3981), .force_10(n18105), .force_11(1'b0), 
        .Q(n14775) );
  \**FFGEN**  \reg_out_reg[3][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3985), .force_10(n18106), .force_11(1'b0), 
        .Q(n14774) );
  \**FFGEN**  \reg_out_reg[3][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3989), .force_10(n18107), .force_11(1'b0), 
        .Q(n14773) );
  \**FFGEN**  \reg_out_reg[3][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3993), .force_10(n18108), .force_11(1'b0), 
        .Q(n14772) );
  \**FFGEN**  \reg_out_reg[3][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3997), .force_10(n18109), .force_11(1'b0), 
        .Q(n14771) );
  \**FFGEN**  \reg_out_reg[3][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4001), .force_10(n18110), .force_11(1'b0), 
        .Q(n14770) );
  \**FFGEN**  \reg_out_reg[3][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4005), .force_10(n18111), .force_11(1'b0), 
        .Q(n14769) );
  \**FFGEN**  \reg_out_reg[3][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4009), .force_10(n18112), .force_11(1'b0), 
        .Q(n14768) );
  \**FFGEN**  \reg_out_reg[3][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4013), .force_10(n18113), .force_11(1'b0), 
        .Q(n14767) );
  \**FFGEN**  \reg_out_reg[3][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4017), .force_10(n18114), .force_11(1'b0), 
        .Q(n14766) );
  \**FFGEN**  \reg_out_reg[3][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4021), .force_10(n18115), .force_11(1'b0), 
        .Q(n14765) );
  \**FFGEN**  \reg_out_reg[3][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4025), .force_10(n18116), .force_11(1'b0), 
        .Q(n14764) );
  \**FFGEN**  \reg_out_reg[3][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4029), .force_10(n18117), .force_11(1'b0), 
        .Q(n14763) );
  \**FFGEN**  \reg_out_reg[3][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4033), .force_10(n18118), .force_11(1'b0), 
        .Q(n14762) );
  \**FFGEN**  \reg_out_reg[3][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4037), .force_10(n18119), .force_11(1'b0), 
        .Q(n14761) );
  \**FFGEN**  \reg_out_reg[3][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4041), .force_10(n18120), .force_11(1'b0), 
        .Q(n14760) );
  \**FFGEN**  \reg_out_reg[3][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4045), .force_10(n18121), .force_11(1'b0), 
        .Q(n14759) );
  \**FFGEN**  \reg_out_reg[3][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4049), .force_10(n18122), .force_11(1'b0), 
        .Q(n14758) );
  \**FFGEN**  \reg_out_reg[3][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4053), .force_10(n18123), .force_11(1'b0), 
        .Q(n14757) );
  \**FFGEN**  \reg_out_reg[3][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4057), .force_10(n18124), .force_11(1'b0), 
        .Q(n14756) );
  \**FFGEN**  \reg_out_reg[3][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4061), .force_10(n18125), .force_11(1'b0), 
        .Q(n14755) );
  \**FFGEN**  \reg_out_reg[3][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4065), .force_10(n18126), .force_11(1'b0), 
        .Q(n14754) );
  \**FFGEN**  \reg_out_reg[3][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4069), .force_10(n18127), .force_11(1'b0), 
        .Q(n14753) );
  \**FFGEN**  \reg_out_reg[3][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4073), .force_10(n18128), .force_11(1'b0), 
        .Q(n14752) );
  \**FFGEN**  \reg_out_reg[3][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4077), .force_10(n18129), .force_11(1'b0), 
        .Q(n14751) );
  \**FFGEN**  \reg_out_reg[3][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4081), .force_10(n18130), .force_11(1'b0), 
        .Q(n14750) );
  \**FFGEN**  \reg_out_reg[3][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4085), .force_10(n18131), .force_11(1'b0), 
        .Q(n14749) );
  \**FFGEN**  \reg_out_reg[3][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4089), .force_10(n18132), .force_11(1'b0), 
        .Q(n14748) );
  \**FFGEN**  \reg_out_reg[3][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4093), .force_10(n18133), .force_11(1'b0), 
        .Q(n14747) );
  \**FFGEN**  \reg_out_reg[3][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4097), .force_10(n18134), .force_11(1'b0), 
        .Q(n14746) );
  \**FFGEN**  \reg_out_reg[3][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4101), .force_10(n18135), .force_11(1'b0), 
        .Q(n14745) );
  \**FFGEN**  \reg_out_reg[3][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4105), .force_10(n18136), .force_11(1'b0), 
        .Q(n14744) );
  \**FFGEN**  \reg_out_reg[3][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4109), .force_10(n18137), .force_11(1'b0), 
        .Q(n14743) );
  \**FFGEN**  \reg_out_reg[3][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4113), .force_10(n18138), .force_11(1'b0), 
        .Q(n14742) );
  \**FFGEN**  \reg_out_reg[3][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4117), .force_10(n18139), .force_11(1'b0), 
        .Q(n14741) );
  \**FFGEN**  \reg_out_reg[3][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4121), .force_10(n18140), .force_11(1'b0), 
        .Q(n14740) );
  \**FFGEN**  \reg_out_reg[3][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4125), .force_10(n18141), .force_11(1'b0), 
        .Q(n14739) );
  \**FFGEN**  \reg_out_reg[3][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4129), .force_10(n18142), .force_11(1'b0), 
        .Q(n14738) );
  \**FFGEN**  \reg_out_reg[3][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4133), .force_10(n18143), .force_11(1'b0), 
        .Q(n14737) );
  \**FFGEN**  \reg_out_reg[3][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4137), .force_10(n18144), .force_11(1'b0), 
        .Q(n14736) );
  \**FFGEN**  \reg_out_reg[3][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4141), .force_10(n18145), .force_11(1'b0), 
        .Q(n14735) );
  \**FFGEN**  \reg_out_reg[3][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4145), .force_10(n18146), .force_11(1'b0), 
        .Q(n14734) );
  \**FFGEN**  \reg_out_reg[3][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4149), .force_10(n18147), .force_11(1'b0), 
        .Q(n14733) );
  \**FFGEN**  \reg_out_reg[3][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4153), .force_10(n18148), .force_11(1'b0), 
        .Q(n14732) );
  \**FFGEN**  \reg_out_reg[3][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4157), .force_10(n18149), .force_11(1'b0), 
        .Q(n14731) );
  \**FFGEN**  \reg_out_reg[3][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4161), .force_10(n18150), .force_11(1'b0), 
        .Q(n14730) );
  \**FFGEN**  \reg_out_reg[3][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4165), .force_10(n18151), .force_11(1'b0), 
        .Q(n14729) );
  \**FFGEN**  \reg_out_reg[3][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4169), .force_10(n18152), .force_11(1'b0), 
        .Q(n14728) );
  \**FFGEN**  \reg_out_reg[3][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4173), .force_10(n18153), .force_11(1'b0), 
        .Q(n14727) );
  \**FFGEN**  \reg_out_reg[3][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4177), .force_10(n18154), .force_11(1'b0), 
        .Q(n14726) );
  \**FFGEN**  \reg_out_reg[3][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4181), .force_10(n18155), .force_11(1'b0), 
        .Q(n14725) );
  \**FFGEN**  \reg_out_reg[3][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4185), .force_10(n18156), .force_11(1'b0), 
        .Q(n14724) );
  \**FFGEN**  \reg_out_reg[3][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4189), .force_10(n18157), .force_11(1'b0), 
        .Q(n14723) );
  \**FFGEN**  \reg_out_reg[2][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4193), .force_10(n18158), .force_11(1'b0), 
        .Q(n14722) );
  \**FFGEN**  \reg_out_reg[2][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4197), .force_10(n18159), .force_11(1'b0), 
        .Q(n14721) );
  \**FFGEN**  \reg_out_reg[2][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4201), .force_10(n18160), .force_11(1'b0), 
        .Q(n14720) );
  \**FFGEN**  \reg_out_reg[2][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4205), .force_10(n18161), .force_11(1'b0), 
        .Q(n14719) );
  \**FFGEN**  \reg_out_reg[2][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4209), .force_10(n18162), .force_11(1'b0), 
        .Q(n14718) );
  \**FFGEN**  \reg_out_reg[2][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4213), .force_10(n18163), .force_11(1'b0), 
        .Q(n14717) );
  \**FFGEN**  \reg_out_reg[2][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4217), .force_10(n18164), .force_11(1'b0), 
        .Q(n14716) );
  \**FFGEN**  \reg_out_reg[2][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4221), .force_10(n18165), .force_11(1'b0), 
        .Q(n14715) );
  \**FFGEN**  \reg_out_reg[2][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4225), .force_10(n18166), .force_11(1'b0), 
        .Q(n14714) );
  \**FFGEN**  \reg_out_reg[2][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4229), .force_10(n18167), .force_11(1'b0), 
        .Q(n14713) );
  \**FFGEN**  \reg_out_reg[2][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4233), .force_10(n18168), .force_11(1'b0), 
        .Q(n14712) );
  \**FFGEN**  \reg_out_reg[2][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4237), .force_10(n18169), .force_11(1'b0), 
        .Q(n14711) );
  \**FFGEN**  \reg_out_reg[2][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4241), .force_10(n18170), .force_11(1'b0), 
        .Q(n14710) );
  \**FFGEN**  \reg_out_reg[2][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4245), .force_10(n18171), .force_11(1'b0), 
        .Q(n14709) );
  \**FFGEN**  \reg_out_reg[2][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4249), .force_10(n18172), .force_11(1'b0), 
        .Q(n14708) );
  \**FFGEN**  \reg_out_reg[2][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4253), .force_10(n18173), .force_11(1'b0), 
        .Q(n14707) );
  \**FFGEN**  \reg_out_reg[2][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4257), .force_10(n18174), .force_11(1'b0), 
        .Q(n14706) );
  \**FFGEN**  \reg_out_reg[2][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4261), .force_10(n18175), .force_11(1'b0), 
        .Q(n14705) );
  \**FFGEN**  \reg_out_reg[2][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4265), .force_10(n18176), .force_11(1'b0), 
        .Q(n14704) );
  \**FFGEN**  \reg_out_reg[2][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4269), .force_10(n18177), .force_11(1'b0), 
        .Q(n14703) );
  \**FFGEN**  \reg_out_reg[2][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4273), .force_10(n18178), .force_11(1'b0), 
        .Q(n14702) );
  \**FFGEN**  \reg_out_reg[2][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4277), .force_10(n18179), .force_11(1'b0), 
        .Q(n14701) );
  \**FFGEN**  \reg_out_reg[2][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4281), .force_10(n18180), .force_11(1'b0), 
        .Q(n14700) );
  \**FFGEN**  \reg_out_reg[2][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4285), .force_10(n18181), .force_11(1'b0), 
        .Q(n14699) );
  \**FFGEN**  \reg_out_reg[2][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4289), .force_10(n18182), .force_11(1'b0), 
        .Q(n14698) );
  \**FFGEN**  \reg_out_reg[2][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4293), .force_10(n18183), .force_11(1'b0), 
        .Q(n14697) );
  \**FFGEN**  \reg_out_reg[2][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4297), .force_10(n18184), .force_11(1'b0), 
        .Q(n14696) );
  \**FFGEN**  \reg_out_reg[2][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4301), .force_10(n18185), .force_11(1'b0), 
        .Q(n14695) );
  \**FFGEN**  \reg_out_reg[2][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4305), .force_10(n18186), .force_11(1'b0), 
        .Q(n14694) );
  \**FFGEN**  \reg_out_reg[2][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4309), .force_10(n18187), .force_11(1'b0), 
        .Q(n14693) );
  \**FFGEN**  \reg_out_reg[2][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4313), .force_10(n18188), .force_11(1'b0), 
        .Q(n14692) );
  \**FFGEN**  \reg_out_reg[2][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4317), .force_10(n18189), .force_11(1'b0), 
        .Q(n14691) );
  \**FFGEN**  \reg_out_reg[2][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4321), .force_10(n18190), .force_11(1'b0), 
        .Q(n14690) );
  \**FFGEN**  \reg_out_reg[2][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4325), .force_10(n18191), .force_11(1'b0), 
        .Q(n14689) );
  \**FFGEN**  \reg_out_reg[2][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4329), .force_10(n18192), .force_11(1'b0), 
        .Q(n14688) );
  \**FFGEN**  \reg_out_reg[2][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4333), .force_10(n18193), .force_11(1'b0), 
        .Q(n14687) );
  \**FFGEN**  \reg_out_reg[2][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4337), .force_10(n18194), .force_11(1'b0), 
        .Q(n14686) );
  \**FFGEN**  \reg_out_reg[2][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4341), .force_10(n18195), .force_11(1'b0), 
        .Q(n14685) );
  \**FFGEN**  \reg_out_reg[2][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4345), .force_10(n18196), .force_11(1'b0), 
        .Q(n14684) );
  \**FFGEN**  \reg_out_reg[2][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4349), .force_10(n18197), .force_11(1'b0), 
        .Q(n14683) );
  \**FFGEN**  \reg_out_reg[2][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4353), .force_10(n18198), .force_11(1'b0), 
        .Q(n14682) );
  \**FFGEN**  \reg_out_reg[2][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4357), .force_10(n18199), .force_11(1'b0), 
        .Q(n14681) );
  \**FFGEN**  \reg_out_reg[2][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4361), .force_10(n18200), .force_11(1'b0), 
        .Q(n14680) );
  \**FFGEN**  \reg_out_reg[2][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4365), .force_10(n18201), .force_11(1'b0), 
        .Q(n14679) );
  \**FFGEN**  \reg_out_reg[2][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4369), .force_10(n18202), .force_11(1'b0), 
        .Q(n14678) );
  \**FFGEN**  \reg_out_reg[2][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4373), .force_10(n18203), .force_11(1'b0), 
        .Q(n14677) );
  \**FFGEN**  \reg_out_reg[2][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4377), .force_10(n18204), .force_11(1'b0), 
        .Q(n14676) );
  \**FFGEN**  \reg_out_reg[2][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4381), .force_10(n18205), .force_11(1'b0), 
        .Q(n14675) );
  \**FFGEN**  \reg_out_reg[2][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4385), .force_10(n18206), .force_11(1'b0), 
        .Q(n14674) );
  \**FFGEN**  \reg_out_reg[2][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4389), .force_10(n18207), .force_11(1'b0), 
        .Q(n14673) );
  \**FFGEN**  \reg_out_reg[2][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4393), .force_10(n18208), .force_11(1'b0), 
        .Q(n14672) );
  \**FFGEN**  \reg_out_reg[2][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4397), .force_10(n18209), .force_11(1'b0), 
        .Q(n14671) );
  \**FFGEN**  \reg_out_reg[2][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4401), .force_10(n18210), .force_11(1'b0), 
        .Q(n14670) );
  \**FFGEN**  \reg_out_reg[2][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4405), .force_10(n18211), .force_11(1'b0), 
        .Q(n14669) );
  \**FFGEN**  \reg_out_reg[2][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4409), .force_10(n18212), .force_11(1'b0), 
        .Q(n14668) );
  \**FFGEN**  \reg_out_reg[2][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4413), .force_10(n18213), .force_11(1'b0), 
        .Q(n14667) );
  \**FFGEN**  \reg_out_reg[2][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4417), .force_10(n18214), .force_11(1'b0), 
        .Q(n14666) );
  \**FFGEN**  \reg_out_reg[2][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4421), .force_10(n18215), .force_11(1'b0), 
        .Q(n14665) );
  \**FFGEN**  \reg_out_reg[2][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4425), .force_10(n18216), .force_11(1'b0), 
        .Q(n14664) );
  \**FFGEN**  \reg_out_reg[2][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4429), .force_10(n18217), .force_11(1'b0), 
        .Q(n14663) );
  \**FFGEN**  \reg_out_reg[2][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4433), .force_10(n18218), .force_11(1'b0), 
        .Q(n14662) );
  \**FFGEN**  \reg_out_reg[2][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4437), .force_10(n18219), .force_11(1'b0), 
        .Q(n14661) );
  \**FFGEN**  \reg_out_reg[2][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4441), .force_10(n18220), .force_11(1'b0), 
        .Q(n14660) );
  \**FFGEN**  \reg_out_reg[2][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4445), .force_10(n18221), .force_11(1'b0), 
        .Q(n14659) );
  \**FFGEN**  \reg_out_reg[2][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4449), .force_10(n18222), .force_11(1'b0), 
        .Q(n14658) );
  \**FFGEN**  \reg_out_reg[2][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4453), .force_10(n18223), .force_11(1'b0), 
        .Q(n14657) );
  \**FFGEN**  \reg_out_reg[2][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4457), .force_10(n18224), .force_11(1'b0), 
        .Q(n14656) );
  \**FFGEN**  \reg_out_reg[2][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4461), .force_10(n18225), .force_11(1'b0), 
        .Q(n14655) );
  \**FFGEN**  \reg_out_reg[2][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4465), .force_10(n18226), .force_11(1'b0), 
        .Q(n14654) );
  \**FFGEN**  \reg_out_reg[2][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4469), .force_10(n18227), .force_11(1'b0), 
        .Q(n14653) );
  \**FFGEN**  \reg_out_reg[2][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4473), .force_10(n18228), .force_11(1'b0), 
        .Q(n14652) );
  \**FFGEN**  \reg_out_reg[2][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4477), .force_10(n18229), .force_11(1'b0), 
        .Q(n14651) );
  \**FFGEN**  \reg_out_reg[2][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4481), .force_10(n18230), .force_11(1'b0), 
        .Q(n14650) );
  \**FFGEN**  \reg_out_reg[2][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4485), .force_10(n18231), .force_11(1'b0), 
        .Q(n14649) );
  \**FFGEN**  \reg_out_reg[2][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4489), .force_10(n18232), .force_11(1'b0), 
        .Q(n14648) );
  \**FFGEN**  \reg_out_reg[2][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4493), .force_10(n18233), .force_11(1'b0), 
        .Q(n14647) );
  \**FFGEN**  \reg_out_reg[2][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4497), .force_10(n18234), .force_11(1'b0), 
        .Q(n14646) );
  \**FFGEN**  \reg_out_reg[2][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4501), .force_10(n18235), .force_11(1'b0), 
        .Q(n14645) );
  \**FFGEN**  \reg_out_reg[2][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4505), .force_10(n18236), .force_11(1'b0), 
        .Q(n14644) );
  \**FFGEN**  \reg_out_reg[2][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4509), .force_10(n18237), .force_11(1'b0), 
        .Q(n14643) );
  \**FFGEN**  \reg_out_reg[1][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4513), .force_10(n18238), .force_11(1'b0), 
        .Q(n14642) );
  \**FFGEN**  \reg_out_reg[1][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4517), .force_10(n18239), .force_11(1'b0), 
        .Q(n14641) );
  \**FFGEN**  \reg_out_reg[1][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4521), .force_10(n18240), .force_11(1'b0), 
        .Q(n14640) );
  \**FFGEN**  \reg_out_reg[1][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4525), .force_10(n18241), .force_11(1'b0), 
        .Q(n14639) );
  \**FFGEN**  \reg_out_reg[1][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4529), .force_10(n18242), .force_11(1'b0), 
        .Q(n14638) );
  \**FFGEN**  \reg_out_reg[1][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4533), .force_10(n18243), .force_11(1'b0), 
        .Q(n14637) );
  \**FFGEN**  \reg_out_reg[1][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4537), .force_10(n18244), .force_11(1'b0), 
        .Q(n14636) );
  \**FFGEN**  \reg_out_reg[1][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4541), .force_10(n18245), .force_11(1'b0), 
        .Q(n14635) );
  \**FFGEN**  \reg_out_reg[1][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4545), .force_10(n18246), .force_11(1'b0), 
        .Q(n14634) );
  \**FFGEN**  \reg_out_reg[1][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4549), .force_10(n18247), .force_11(1'b0), 
        .Q(n14633) );
  \**FFGEN**  \reg_out_reg[1][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4553), .force_10(n18248), .force_11(1'b0), 
        .Q(n14632) );
  \**FFGEN**  \reg_out_reg[1][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4557), .force_10(n18249), .force_11(1'b0), 
        .Q(n14631) );
  \**FFGEN**  \reg_out_reg[1][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4561), .force_10(n18250), .force_11(1'b0), 
        .Q(n14630) );
  \**FFGEN**  \reg_out_reg[1][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4565), .force_10(n18251), .force_11(1'b0), 
        .Q(n14629) );
  \**FFGEN**  \reg_out_reg[1][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4569), .force_10(n18252), .force_11(1'b0), 
        .Q(n14628) );
  \**FFGEN**  \reg_out_reg[1][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4573), .force_10(n18253), .force_11(1'b0), 
        .Q(n14627) );
  \**FFGEN**  \reg_out_reg[1][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4577), .force_10(n18254), .force_11(1'b0), 
        .Q(n14626) );
  \**FFGEN**  \reg_out_reg[1][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4581), .force_10(n18255), .force_11(1'b0), 
        .Q(n14625) );
  \**FFGEN**  \reg_out_reg[1][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4585), .force_10(n18256), .force_11(1'b0), 
        .Q(n14624) );
  \**FFGEN**  \reg_out_reg[1][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4589), .force_10(n18257), .force_11(1'b0), 
        .Q(n14623) );
  \**FFGEN**  \reg_out_reg[1][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4593), .force_10(n18258), .force_11(1'b0), 
        .Q(n14622) );
  \**FFGEN**  \reg_out_reg[1][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4597), .force_10(n18259), .force_11(1'b0), 
        .Q(n14621) );
  \**FFGEN**  \reg_out_reg[1][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4601), .force_10(n18260), .force_11(1'b0), 
        .Q(n14620) );
  \**FFGEN**  \reg_out_reg[1][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4605), .force_10(n18261), .force_11(1'b0), 
        .Q(n14619) );
  \**FFGEN**  \reg_out_reg[1][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4609), .force_10(n18262), .force_11(1'b0), 
        .Q(n14618) );
  \**FFGEN**  \reg_out_reg[1][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4613), .force_10(n18263), .force_11(1'b0), 
        .Q(n14617) );
  \**FFGEN**  \reg_out_reg[1][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4617), .force_10(n18264), .force_11(1'b0), 
        .Q(n14616) );
  \**FFGEN**  \reg_out_reg[1][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4621), .force_10(n18265), .force_11(1'b0), 
        .Q(n14615) );
  \**FFGEN**  \reg_out_reg[1][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4625), .force_10(n18266), .force_11(1'b0), 
        .Q(n14614) );
  \**FFGEN**  \reg_out_reg[1][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4629), .force_10(n18267), .force_11(1'b0), 
        .Q(n14613) );
  \**FFGEN**  \reg_out_reg[1][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4633), .force_10(n18268), .force_11(1'b0), 
        .Q(n14612) );
  \**FFGEN**  \reg_out_reg[1][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4637), .force_10(n18269), .force_11(1'b0), 
        .Q(n14611) );
  \**FFGEN**  \reg_out_reg[1][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4641), .force_10(n18270), .force_11(1'b0), 
        .Q(n14610) );
  \**FFGEN**  \reg_out_reg[1][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4645), .force_10(n18271), .force_11(1'b0), 
        .Q(n14609) );
  \**FFGEN**  \reg_out_reg[1][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4649), .force_10(n18272), .force_11(1'b0), 
        .Q(n14608) );
  \**FFGEN**  \reg_out_reg[1][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4653), .force_10(n18273), .force_11(1'b0), 
        .Q(n14607) );
  \**FFGEN**  \reg_out_reg[1][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4657), .force_10(n18274), .force_11(1'b0), 
        .Q(n14606) );
  \**FFGEN**  \reg_out_reg[1][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4661), .force_10(n18275), .force_11(1'b0), 
        .Q(n14605) );
  \**FFGEN**  \reg_out_reg[1][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4665), .force_10(n18276), .force_11(1'b0), 
        .Q(n14604) );
  \**FFGEN**  \reg_out_reg[1][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4669), .force_10(n18277), .force_11(1'b0), 
        .Q(n14603) );
  \**FFGEN**  \reg_out_reg[1][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4673), .force_10(n18278), .force_11(1'b0), 
        .Q(n14602) );
  \**FFGEN**  \reg_out_reg[1][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4677), .force_10(n18279), .force_11(1'b0), 
        .Q(n14601) );
  \**FFGEN**  \reg_out_reg[1][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4681), .force_10(n18280), .force_11(1'b0), 
        .Q(n14600) );
  \**FFGEN**  \reg_out_reg[1][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4685), .force_10(n18281), .force_11(1'b0), 
        .Q(n14599) );
  \**FFGEN**  \reg_out_reg[1][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4689), .force_10(n18282), .force_11(1'b0), 
        .Q(n14598) );
  \**FFGEN**  \reg_out_reg[1][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4693), .force_10(n18283), .force_11(1'b0), 
        .Q(n14597) );
  \**FFGEN**  \reg_out_reg[1][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4697), .force_10(n18284), .force_11(1'b0), 
        .Q(n14596) );
  \**FFGEN**  \reg_out_reg[1][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4701), .force_10(n18285), .force_11(1'b0), 
        .Q(n14595) );
  \**FFGEN**  \reg_out_reg[1][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4705), .force_10(n18286), .force_11(1'b0), 
        .Q(n14594) );
  \**FFGEN**  \reg_out_reg[1][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4709), .force_10(n18287), .force_11(1'b0), 
        .Q(n14593) );
  \**FFGEN**  \reg_out_reg[1][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4713), .force_10(n18288), .force_11(1'b0), 
        .Q(n14592) );
  \**FFGEN**  \reg_out_reg[1][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4717), .force_10(n18289), .force_11(1'b0), 
        .Q(n14591) );
  \**FFGEN**  \reg_out_reg[1][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4721), .force_10(n18290), .force_11(1'b0), 
        .Q(n14590) );
  \**FFGEN**  \reg_out_reg[1][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4725), .force_10(n18291), .force_11(1'b0), 
        .Q(n14589) );
  \**FFGEN**  \reg_out_reg[1][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4729), .force_10(n18292), .force_11(1'b0), 
        .Q(n14588) );
  \**FFGEN**  \reg_out_reg[1][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4733), .force_10(n18293), .force_11(1'b0), 
        .Q(n14587) );
  \**FFGEN**  \reg_out_reg[1][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4737), .force_10(n18294), .force_11(1'b0), 
        .Q(n14586) );
  \**FFGEN**  \reg_out_reg[1][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4741), .force_10(n18295), .force_11(1'b0), 
        .Q(n14585) );
  \**FFGEN**  \reg_out_reg[1][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4745), .force_10(n18296), .force_11(1'b0), 
        .Q(n14584) );
  \**FFGEN**  \reg_out_reg[1][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4749), .force_10(n18297), .force_11(1'b0), 
        .Q(n14583) );
  \**FFGEN**  \reg_out_reg[1][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4753), .force_10(n18298), .force_11(1'b0), 
        .Q(n14582) );
  \**FFGEN**  \reg_out_reg[1][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4757), .force_10(n18299), .force_11(1'b0), 
        .Q(n14581) );
  \**FFGEN**  \reg_out_reg[1][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4761), .force_10(n18300), .force_11(1'b0), 
        .Q(n14580) );
  \**FFGEN**  \reg_out_reg[1][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4765), .force_10(n18301), .force_11(1'b0), 
        .Q(n14579) );
  \**FFGEN**  \reg_out_reg[1][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4769), .force_10(n18302), .force_11(1'b0), 
        .Q(n14578) );
  \**FFGEN**  \reg_out_reg[1][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4773), .force_10(n18303), .force_11(1'b0), 
        .Q(n14577) );
  \**FFGEN**  \reg_out_reg[1][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4777), .force_10(n18304), .force_11(1'b0), 
        .Q(n14576) );
  \**FFGEN**  \reg_out_reg[1][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4781), .force_10(n18305), .force_11(1'b0), 
        .Q(n14575) );
  \**FFGEN**  \reg_out_reg[1][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4785), .force_10(n18306), .force_11(1'b0), 
        .Q(n14574) );
  \**FFGEN**  \reg_out_reg[1][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4789), .force_10(n18307), .force_11(1'b0), 
        .Q(n14573) );
  \**FFGEN**  \reg_out_reg[1][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4793), .force_10(n18308), .force_11(1'b0), 
        .Q(n14572) );
  \**FFGEN**  \reg_out_reg[1][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4797), .force_10(n18309), .force_11(1'b0), 
        .Q(n14571) );
  \**FFGEN**  \reg_out_reg[1][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4801), .force_10(n18310), .force_11(1'b0), 
        .Q(n14570) );
  \**FFGEN**  \reg_out_reg[1][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4805), .force_10(n18311), .force_11(1'b0), 
        .Q(n14569) );
  \**FFGEN**  \reg_out_reg[1][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4809), .force_10(n18312), .force_11(1'b0), 
        .Q(n14568) );
  \**FFGEN**  \reg_out_reg[1][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4813), .force_10(n18313), .force_11(1'b0), 
        .Q(n14567) );
  \**FFGEN**  \reg_out_reg[1][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4817), .force_10(n18314), .force_11(1'b0), 
        .Q(n14566) );
  \**FFGEN**  \reg_out_reg[1][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4821), .force_10(n18315), .force_11(1'b0), 
        .Q(n14565) );
  \**FFGEN**  \reg_out_reg[1][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4825), .force_10(n18316), .force_11(1'b0), 
        .Q(n14564) );
  \**FFGEN**  \reg_out_reg[1][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4829), .force_10(n18317), .force_11(1'b0), 
        .Q(n14563) );
  \**FFGEN**  \reg_out_reg[0][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4833), .force_10(n18318), .force_11(1'b0), 
        .Q(n14562) );
  \**FFGEN**  \reg_out_reg[0][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4837), .force_10(n18319), .force_11(1'b0), 
        .Q(n14561) );
  \**FFGEN**  \reg_out_reg[0][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4841), .force_10(n18320), .force_11(1'b0), 
        .Q(n14560) );
  \**FFGEN**  \reg_out_reg[0][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4845), .force_10(n18321), .force_11(1'b0), 
        .Q(n14559) );
  \**FFGEN**  \reg_out_reg[0][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4849), .force_10(n18322), .force_11(1'b0), 
        .Q(n14558) );
  \**FFGEN**  \reg_out_reg[0][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4853), .force_10(n18323), .force_11(1'b0), 
        .Q(n14557) );
  \**FFGEN**  \reg_out_reg[0][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4857), .force_10(n18324), .force_11(1'b0), 
        .Q(n14556) );
  \**FFGEN**  \reg_out_reg[0][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4861), .force_10(n18325), .force_11(1'b0), 
        .Q(n14555) );
  \**FFGEN**  \reg_out_reg[0][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4865), .force_10(n18326), .force_11(1'b0), 
        .Q(n14554) );
  \**FFGEN**  \reg_out_reg[0][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4869), .force_10(n18327), .force_11(1'b0), 
        .Q(n14553) );
  \**FFGEN**  \reg_out_reg[0][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4873), .force_10(n18328), .force_11(1'b0), 
        .Q(n14552) );
  \**FFGEN**  \reg_out_reg[0][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4877), .force_10(n18329), .force_11(1'b0), 
        .Q(n14551) );
  \**FFGEN**  \reg_out_reg[0][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4881), .force_10(n18330), .force_11(1'b0), 
        .Q(n14550) );
  \**FFGEN**  \reg_out_reg[0][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4885), .force_10(n18331), .force_11(1'b0), 
        .Q(n14549) );
  \**FFGEN**  \reg_out_reg[0][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4889), .force_10(n18332), .force_11(1'b0), 
        .Q(n14548) );
  \**FFGEN**  \reg_out_reg[0][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4893), .force_10(n18333), .force_11(1'b0), 
        .Q(n14547) );
  \**FFGEN**  \reg_out_reg[0][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4897), .force_10(n18334), .force_11(1'b0), 
        .Q(n14546) );
  \**FFGEN**  \reg_out_reg[0][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4901), .force_10(n18335), .force_11(1'b0), 
        .Q(n14545) );
  \**FFGEN**  \reg_out_reg[0][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4905), .force_10(n18336), .force_11(1'b0), 
        .Q(n14544) );
  \**FFGEN**  \reg_out_reg[0][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4909), .force_10(n18337), .force_11(1'b0), 
        .Q(n14543) );
  \**FFGEN**  \reg_out_reg[0][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4913), .force_10(n18338), .force_11(1'b0), 
        .Q(n14542) );
  \**FFGEN**  \reg_out_reg[0][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4917), .force_10(n18339), .force_11(1'b0), 
        .Q(n14541) );
  \**FFGEN**  \reg_out_reg[0][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4921), .force_10(n18340), .force_11(1'b0), 
        .Q(n14540) );
  \**FFGEN**  \reg_out_reg[0][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4925), .force_10(n18341), .force_11(1'b0), 
        .Q(n14539) );
  \**FFGEN**  \reg_out_reg[0][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4929), .force_10(n18342), .force_11(1'b0), 
        .Q(n14538) );
  \**FFGEN**  \reg_out_reg[0][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4933), .force_10(n18343), .force_11(1'b0), 
        .Q(n14537) );
  \**FFGEN**  \reg_out_reg[0][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4937), .force_10(n18344), .force_11(1'b0), 
        .Q(n14536) );
  \**FFGEN**  \reg_out_reg[0][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4941), .force_10(n18345), .force_11(1'b0), 
        .Q(n14535) );
  \**FFGEN**  \reg_out_reg[0][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4945), .force_10(n18346), .force_11(1'b0), 
        .Q(n14534) );
  \**FFGEN**  \reg_out_reg[0][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4949), .force_10(n18347), .force_11(1'b0), 
        .Q(n14533) );
  \**FFGEN**  \reg_out_reg[0][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4953), .force_10(n18348), .force_11(1'b0), 
        .Q(n14532) );
  \**FFGEN**  \reg_out_reg[0][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4957), .force_10(n18349), .force_11(1'b0), 
        .Q(n14531) );
  \**FFGEN**  \reg_out_reg[0][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4961), .force_10(n18350), .force_11(1'b0), 
        .Q(n14530) );
  \**FFGEN**  \reg_out_reg[0][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4965), .force_10(n18351), .force_11(1'b0), 
        .Q(n14529) );
  \**FFGEN**  \reg_out_reg[0][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4969), .force_10(n18352), .force_11(1'b0), 
        .Q(n14528) );
  \**FFGEN**  \reg_out_reg[0][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4973), .force_10(n18353), .force_11(1'b0), 
        .Q(n14527) );
  \**FFGEN**  \reg_out_reg[0][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4977), .force_10(n18354), .force_11(1'b0), 
        .Q(n14526) );
  \**FFGEN**  \reg_out_reg[0][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4981), .force_10(n18355), .force_11(1'b0), 
        .Q(n14525) );
  \**FFGEN**  \reg_out_reg[0][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4985), .force_10(n18356), .force_11(1'b0), 
        .Q(n14524) );
  \**FFGEN**  \reg_out_reg[0][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4989), .force_10(n18357), .force_11(1'b0), 
        .Q(n14523) );
  \**FFGEN**  \reg_out_reg[0][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4993), .force_10(n18358), .force_11(1'b0), 
        .Q(n14522) );
  \**FFGEN**  \reg_out_reg[0][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n4997), .force_10(n18359), .force_11(1'b0), 
        .Q(n14521) );
  \**FFGEN**  \reg_out_reg[0][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5001), .force_10(n18360), .force_11(1'b0), 
        .Q(n14520) );
  \**FFGEN**  \reg_out_reg[0][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5005), .force_10(n18361), .force_11(1'b0), 
        .Q(n14519) );
  \**FFGEN**  \reg_out_reg[0][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5009), .force_10(n18362), .force_11(1'b0), 
        .Q(n14518) );
  \**FFGEN**  \reg_out_reg[0][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5013), .force_10(n18363), .force_11(1'b0), 
        .Q(n14517) );
  \**FFGEN**  \reg_out_reg[0][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5017), .force_10(n18364), .force_11(1'b0), 
        .Q(n14516) );
  \**FFGEN**  \reg_out_reg[0][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5021), .force_10(n18365), .force_11(1'b0), 
        .Q(n14515) );
  \**FFGEN**  \reg_out_reg[0][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5025), .force_10(n18366), .force_11(1'b0), 
        .Q(n14514) );
  \**FFGEN**  \reg_out_reg[0][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5029), .force_10(n18367), .force_11(1'b0), 
        .Q(n14513) );
  \**FFGEN**  \reg_out_reg[0][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5033), .force_10(n18368), .force_11(1'b0), 
        .Q(n14512) );
  \**FFGEN**  \reg_out_reg[0][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5037), .force_10(n18369), .force_11(1'b0), 
        .Q(n14511) );
  \**FFGEN**  \reg_out_reg[0][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5041), .force_10(n18370), .force_11(1'b0), 
        .Q(n14510) );
  \**FFGEN**  \reg_out_reg[0][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5045), .force_10(n18371), .force_11(1'b0), 
        .Q(n14509) );
  \**FFGEN**  \reg_out_reg[0][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5049), .force_10(n18372), .force_11(1'b0), 
        .Q(n14508) );
  \**FFGEN**  \reg_out_reg[0][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5053), .force_10(n18373), .force_11(1'b0), 
        .Q(n14507) );
  \**FFGEN**  \reg_out_reg[0][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5057), .force_10(n18374), .force_11(1'b0), 
        .Q(n14506) );
  \**FFGEN**  \reg_out_reg[0][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5061), .force_10(n18375), .force_11(1'b0), 
        .Q(n14505) );
  \**FFGEN**  \reg_out_reg[0][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5065), .force_10(n18376), .force_11(1'b0), 
        .Q(n14504) );
  \**FFGEN**  \reg_out_reg[0][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5069), .force_10(n18377), .force_11(1'b0), 
        .Q(n14503) );
  \**FFGEN**  \reg_out_reg[0][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5073), .force_10(n18378), .force_11(1'b0), 
        .Q(n14502) );
  \**FFGEN**  \reg_out_reg[0][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5077), .force_10(n18379), .force_11(1'b0), 
        .Q(n14501) );
  \**FFGEN**  \reg_out_reg[0][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5081), .force_10(n18380), .force_11(1'b0), 
        .Q(n14500) );
  \**FFGEN**  \reg_out_reg[0][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5085), .force_10(n18381), .force_11(1'b0), 
        .Q(n14499) );
  \**FFGEN**  \reg_out_reg[0][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5089), .force_10(n18382), .force_11(1'b0), 
        .Q(n14498) );
  \**FFGEN**  \reg_out_reg[0][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5093), .force_10(n18383), .force_11(1'b0), 
        .Q(n14497) );
  \**FFGEN**  \reg_out_reg[0][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5097), .force_10(n18384), .force_11(1'b0), 
        .Q(n14496) );
  \**FFGEN**  \reg_out_reg[0][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5101), .force_10(n18385), .force_11(1'b0), 
        .Q(n14495) );
  \**FFGEN**  \reg_out_reg[0][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5105), .force_10(n18386), .force_11(1'b0), 
        .Q(n14494) );
  \**FFGEN**  \reg_out_reg[0][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5109), .force_10(n18387), .force_11(1'b0), 
        .Q(n14493) );
  \**FFGEN**  \reg_out_reg[0][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5113), .force_10(n18388), .force_11(1'b0), 
        .Q(n14492) );
  \**FFGEN**  \reg_out_reg[0][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5117), .force_10(n18389), .force_11(1'b0), 
        .Q(n14491) );
  \**FFGEN**  \reg_out_reg[0][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5121), .force_10(n18390), .force_11(1'b0), 
        .Q(n14490) );
  \**FFGEN**  \reg_out_reg[0][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5125), .force_10(n18391), .force_11(1'b0), 
        .Q(n14489) );
  \**FFGEN**  \reg_out_reg[0][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5129), .force_10(n18392), .force_11(1'b0), 
        .Q(n14488) );
  \**FFGEN**  \reg_out_reg[0][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5133), .force_10(n18393), .force_11(1'b0), 
        .Q(n14487) );
  \**FFGEN**  \reg_out_reg[0][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5137), .force_10(n18394), .force_11(1'b0), 
        .Q(n14486) );
  \**FFGEN**  \reg_out_reg[0][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5141), .force_10(n18395), .force_11(1'b0), 
        .Q(n14485) );
  \**FFGEN**  \reg_out_reg[0][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5145), .force_10(n18396), .force_11(1'b0), 
        .Q(n14484) );
  \**FFGEN**  \reg_out_reg[0][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3869), .force_10(n18077), .force_11(1'b0), 
        .Q(n14483) );
  nand_x8_sg U7711 ( .A(state[0]), .B(n18399), .X(n14475) );
  inv_x4_sg U9655 ( .A(n16776), .X(n16775) );
  inv_x4_sg U9656 ( .A(n16743), .X(n16742) );
  inv_x4_sg U9657 ( .A(n16777), .X(n16776) );
  inv_x2_sg U9658 ( .A(n13189), .X(n16777) );
  nor_x1_sg U9659 ( .A(n14475), .B(n18397), .X(n13189) );
  inv_x4_sg U9660 ( .A(n16744), .X(n16743) );
  inv_x2_sg U9661 ( .A(n13831), .X(n16744) );
  nor_x1_sg U9662 ( .A(n14470), .B(n14471), .X(n13831) );
  inv_x2_sg U9663 ( .A(n13188), .X(n16796) );
  nor_x1_sg U9664 ( .A(n18397), .B(n16774), .X(n13188) );
  inv_x2_sg U9665 ( .A(n13830), .X(n16760) );
  nor_x1_sg U9666 ( .A(n18397), .B(n16741), .X(n13830) );
  inv_x4_sg U9667 ( .A(n16795), .X(n16794) );
  inv_x4_sg U9668 ( .A(n16759), .X(n16758) );
  inv_x4_sg U9669 ( .A(n16796), .X(n16795) );
  inv_x4_sg U9670 ( .A(n16760), .X(n16759) );
  inv_x1_sg U9671 ( .A(n18400), .X(n15445) );
  inv_x2_sg U9672 ( .A(n15445), .X(n15446) );
  inv_x1_sg U9673 ( .A(n18401), .X(n15447) );
  inv_x2_sg U9674 ( .A(n15447), .X(n15448) );
  nor_x4_sg U9675 ( .A(n14479), .B(n18397), .X(n14474) );
  nand_x4_sg U9676 ( .A(n14475), .B(n14482), .X(n14479) );
  inv_x8_sg U9677 ( .A(n14480), .X(n18398) );
  nand_x4_sg U9678 ( .A(n14481), .B(output_taken), .X(n14480) );
  inv_x8_sg U9679 ( .A(n14472), .X(n18397) );
  nor_x8_sg U9680 ( .A(n18398), .B(reset), .X(n14472) );
  inv_x1_sg U9681 ( .A(n18721), .X(n16089) );
  inv_x1_sg U9682 ( .A(n18720), .X(n16087) );
  inv_x1_sg U9683 ( .A(n18719), .X(n16085) );
  inv_x1_sg U9684 ( .A(n18718), .X(n16083) );
  inv_x1_sg U9685 ( .A(n18717), .X(n16081) );
  inv_x1_sg U9686 ( .A(n18716), .X(n16079) );
  inv_x1_sg U9687 ( .A(n18715), .X(n16077) );
  inv_x1_sg U9688 ( .A(n18714), .X(n16075) );
  inv_x1_sg U9689 ( .A(n18713), .X(n16073) );
  inv_x1_sg U9690 ( .A(n18712), .X(n16071) );
  inv_x1_sg U9691 ( .A(n18711), .X(n16069) );
  inv_x1_sg U9692 ( .A(n18710), .X(n16067) );
  inv_x1_sg U9693 ( .A(n18709), .X(n16065) );
  inv_x1_sg U9694 ( .A(n18708), .X(n16063) );
  inv_x1_sg U9695 ( .A(n18707), .X(n16061) );
  inv_x1_sg U9696 ( .A(n18706), .X(n16059) );
  inv_x1_sg U9697 ( .A(n18705), .X(n16057) );
  inv_x1_sg U9698 ( .A(n18704), .X(n16055) );
  inv_x1_sg U9699 ( .A(n18703), .X(n16053) );
  inv_x1_sg U9700 ( .A(n18702), .X(n16051) );
  inv_x1_sg U9701 ( .A(n18701), .X(n16049) );
  inv_x1_sg U9702 ( .A(n18700), .X(n16047) );
  inv_x1_sg U9703 ( .A(n18699), .X(n16045) );
  inv_x1_sg U9704 ( .A(n18698), .X(n16043) );
  inv_x1_sg U9705 ( .A(n18697), .X(n16041) );
  inv_x1_sg U9706 ( .A(n18696), .X(n16039) );
  inv_x1_sg U9707 ( .A(n18695), .X(n16037) );
  inv_x1_sg U9708 ( .A(n18694), .X(n16035) );
  inv_x1_sg U9709 ( .A(n18693), .X(n16033) );
  inv_x1_sg U9710 ( .A(n18692), .X(n16031) );
  inv_x1_sg U9711 ( .A(n18691), .X(n16029) );
  inv_x1_sg U9712 ( .A(n18690), .X(n16027) );
  inv_x1_sg U9713 ( .A(n18689), .X(n16025) );
  inv_x1_sg U9714 ( .A(n18688), .X(n16023) );
  inv_x1_sg U9715 ( .A(n18687), .X(n16021) );
  inv_x1_sg U9716 ( .A(n18686), .X(n16019) );
  inv_x1_sg U9717 ( .A(n18685), .X(n16017) );
  inv_x1_sg U9718 ( .A(n18684), .X(n16015) );
  inv_x1_sg U9719 ( .A(n18683), .X(n16013) );
  inv_x1_sg U9720 ( .A(n18682), .X(n16011) );
  inv_x1_sg U9721 ( .A(n18681), .X(n16009) );
  inv_x1_sg U9722 ( .A(n18680), .X(n16007) );
  inv_x1_sg U9723 ( .A(n18679), .X(n16005) );
  inv_x1_sg U9724 ( .A(n18678), .X(n16003) );
  inv_x1_sg U9725 ( .A(n18677), .X(n16001) );
  inv_x1_sg U9726 ( .A(n18676), .X(n15999) );
  inv_x1_sg U9727 ( .A(n18675), .X(n15997) );
  inv_x1_sg U9728 ( .A(n18674), .X(n15995) );
  inv_x1_sg U9729 ( .A(n18673), .X(n15993) );
  inv_x1_sg U9730 ( .A(n18672), .X(n15991) );
  inv_x1_sg U9731 ( .A(n18671), .X(n15989) );
  inv_x1_sg U9732 ( .A(n18670), .X(n15987) );
  inv_x1_sg U9733 ( .A(n18669), .X(n15985) );
  inv_x1_sg U9734 ( .A(n18668), .X(n15983) );
  inv_x1_sg U9735 ( .A(n18667), .X(n15981) );
  inv_x1_sg U9736 ( .A(n18666), .X(n15979) );
  inv_x1_sg U9737 ( .A(n18665), .X(n15977) );
  inv_x1_sg U9738 ( .A(n18664), .X(n15975) );
  inv_x1_sg U9739 ( .A(n18663), .X(n15973) );
  inv_x1_sg U9740 ( .A(n18662), .X(n15971) );
  inv_x1_sg U9741 ( .A(n18661), .X(n15969) );
  inv_x1_sg U9742 ( .A(n18660), .X(n15967) );
  inv_x1_sg U9743 ( .A(n18659), .X(n15965) );
  inv_x1_sg U9744 ( .A(n18658), .X(n15963) );
  inv_x1_sg U9745 ( .A(n18657), .X(n15961) );
  inv_x1_sg U9746 ( .A(n18656), .X(n15959) );
  inv_x1_sg U9747 ( .A(n18655), .X(n15957) );
  inv_x1_sg U9748 ( .A(n18654), .X(n15955) );
  inv_x1_sg U9749 ( .A(n18653), .X(n15953) );
  inv_x1_sg U9750 ( .A(n18652), .X(n15951) );
  inv_x1_sg U9751 ( .A(n18651), .X(n15949) );
  inv_x1_sg U9752 ( .A(n18650), .X(n15947) );
  inv_x1_sg U9753 ( .A(n18649), .X(n15945) );
  inv_x1_sg U9754 ( .A(n18648), .X(n15943) );
  inv_x1_sg U9755 ( .A(n18647), .X(n15941) );
  inv_x1_sg U9756 ( .A(n18646), .X(n15939) );
  inv_x1_sg U9757 ( .A(n18645), .X(n15937) );
  inv_x1_sg U9758 ( .A(n18644), .X(n15935) );
  inv_x1_sg U9759 ( .A(n18643), .X(n15933) );
  inv_x1_sg U9760 ( .A(n18642), .X(n15931) );
  inv_x1_sg U9761 ( .A(n18641), .X(n15929) );
  inv_x1_sg U9762 ( .A(n18640), .X(n15927) );
  inv_x1_sg U9763 ( .A(n18639), .X(n15925) );
  inv_x1_sg U9764 ( .A(n18638), .X(n15923) );
  inv_x1_sg U9765 ( .A(n18637), .X(n15921) );
  inv_x1_sg U9766 ( .A(n18636), .X(n15919) );
  inv_x1_sg U9767 ( .A(n18635), .X(n15917) );
  inv_x1_sg U9768 ( .A(n18634), .X(n15915) );
  inv_x1_sg U9769 ( .A(n18633), .X(n15913) );
  inv_x1_sg U9770 ( .A(n18632), .X(n15911) );
  inv_x1_sg U9771 ( .A(n18631), .X(n15909) );
  inv_x1_sg U9772 ( .A(n18630), .X(n15907) );
  inv_x1_sg U9773 ( .A(n18629), .X(n15905) );
  inv_x1_sg U9774 ( .A(n18628), .X(n15903) );
  inv_x1_sg U9775 ( .A(n18627), .X(n15901) );
  inv_x1_sg U9776 ( .A(n18626), .X(n15899) );
  inv_x1_sg U9777 ( .A(n18625), .X(n15897) );
  inv_x1_sg U9778 ( .A(n18624), .X(n15895) );
  inv_x1_sg U9779 ( .A(n18623), .X(n15893) );
  inv_x1_sg U9780 ( .A(n18622), .X(n15891) );
  inv_x1_sg U9781 ( .A(n18621), .X(n15889) );
  inv_x1_sg U9782 ( .A(n18620), .X(n15887) );
  inv_x1_sg U9783 ( .A(n18619), .X(n15885) );
  inv_x1_sg U9784 ( .A(n18618), .X(n15883) );
  inv_x1_sg U9785 ( .A(n18617), .X(n15881) );
  inv_x1_sg U9786 ( .A(n18616), .X(n15879) );
  inv_x1_sg U9787 ( .A(n18615), .X(n15877) );
  inv_x1_sg U9788 ( .A(n18614), .X(n15875) );
  inv_x1_sg U9789 ( .A(n18613), .X(n15873) );
  inv_x1_sg U9790 ( .A(n18612), .X(n15871) );
  inv_x1_sg U9791 ( .A(n18611), .X(n15869) );
  inv_x1_sg U9792 ( .A(n18610), .X(n15867) );
  inv_x1_sg U9793 ( .A(n18609), .X(n15865) );
  inv_x1_sg U9794 ( .A(n18608), .X(n15863) );
  inv_x1_sg U9795 ( .A(n18607), .X(n15861) );
  inv_x1_sg U9796 ( .A(n18606), .X(n15859) );
  inv_x1_sg U9797 ( .A(n18605), .X(n15857) );
  inv_x1_sg U9798 ( .A(n18604), .X(n15855) );
  inv_x1_sg U9799 ( .A(n18603), .X(n15853) );
  inv_x1_sg U9800 ( .A(n18602), .X(n15851) );
  inv_x1_sg U9801 ( .A(n18601), .X(n15849) );
  inv_x1_sg U9802 ( .A(n18600), .X(n15847) );
  inv_x1_sg U9803 ( .A(n18599), .X(n15845) );
  inv_x1_sg U9804 ( .A(n18598), .X(n15843) );
  inv_x1_sg U9805 ( .A(n18597), .X(n15841) );
  inv_x1_sg U9806 ( .A(n18596), .X(n15839) );
  inv_x1_sg U9807 ( .A(n18595), .X(n15837) );
  inv_x1_sg U9808 ( .A(n18594), .X(n15835) );
  inv_x1_sg U9809 ( .A(n18593), .X(n15833) );
  inv_x1_sg U9810 ( .A(n18592), .X(n15831) );
  inv_x1_sg U9811 ( .A(n18591), .X(n15829) );
  inv_x1_sg U9812 ( .A(n18590), .X(n15827) );
  inv_x1_sg U9813 ( .A(n18589), .X(n15825) );
  inv_x1_sg U9814 ( .A(n18588), .X(n15823) );
  inv_x1_sg U9815 ( .A(n18587), .X(n15821) );
  inv_x1_sg U9816 ( .A(n18586), .X(n15819) );
  inv_x1_sg U9817 ( .A(n18585), .X(n15817) );
  inv_x1_sg U9818 ( .A(n18584), .X(n15815) );
  inv_x1_sg U9819 ( .A(n18583), .X(n15813) );
  inv_x1_sg U9820 ( .A(n18582), .X(n15811) );
  inv_x1_sg U9821 ( .A(n18581), .X(n15809) );
  inv_x1_sg U9822 ( .A(n18580), .X(n15807) );
  inv_x1_sg U9823 ( .A(n18579), .X(n15805) );
  inv_x1_sg U9824 ( .A(n18578), .X(n15803) );
  inv_x1_sg U9825 ( .A(n18577), .X(n15801) );
  inv_x1_sg U9826 ( .A(n18576), .X(n15799) );
  inv_x1_sg U9827 ( .A(n18575), .X(n15797) );
  inv_x1_sg U9828 ( .A(n18574), .X(n15795) );
  inv_x1_sg U9829 ( .A(n18573), .X(n15793) );
  inv_x1_sg U9830 ( .A(n18572), .X(n15791) );
  inv_x1_sg U9831 ( .A(n18571), .X(n15789) );
  inv_x1_sg U9832 ( .A(n18570), .X(n15787) );
  inv_x1_sg U9833 ( .A(n18569), .X(n15785) );
  inv_x1_sg U9834 ( .A(n18568), .X(n15783) );
  inv_x1_sg U9835 ( .A(n18567), .X(n15781) );
  inv_x1_sg U9836 ( .A(n18566), .X(n15779) );
  inv_x1_sg U9837 ( .A(n18565), .X(n15777) );
  inv_x1_sg U9838 ( .A(n18564), .X(n15775) );
  inv_x1_sg U9839 ( .A(n18563), .X(n15773) );
  inv_x1_sg U9840 ( .A(n18562), .X(n15771) );
  inv_x1_sg U9841 ( .A(n18561), .X(n15769) );
  inv_x1_sg U9842 ( .A(n18560), .X(n15767) );
  inv_x1_sg U9843 ( .A(n18559), .X(n15765) );
  inv_x1_sg U9844 ( .A(n18558), .X(n15763) );
  inv_x1_sg U9845 ( .A(n18557), .X(n15761) );
  inv_x1_sg U9846 ( .A(n18556), .X(n15759) );
  inv_x1_sg U9847 ( .A(n18555), .X(n15757) );
  inv_x1_sg U9848 ( .A(n18554), .X(n15755) );
  inv_x1_sg U9849 ( .A(n18553), .X(n15753) );
  inv_x1_sg U9850 ( .A(n18552), .X(n15751) );
  inv_x1_sg U9851 ( .A(n18551), .X(n15749) );
  inv_x1_sg U9852 ( .A(n18550), .X(n15747) );
  inv_x1_sg U9853 ( .A(n18549), .X(n15745) );
  inv_x1_sg U9854 ( .A(n18548), .X(n15743) );
  inv_x1_sg U9855 ( .A(n18547), .X(n15741) );
  inv_x1_sg U9856 ( .A(n18546), .X(n15739) );
  inv_x1_sg U9857 ( .A(n18545), .X(n15737) );
  inv_x1_sg U9858 ( .A(n18544), .X(n15735) );
  inv_x1_sg U9859 ( .A(n18543), .X(n15733) );
  inv_x1_sg U9860 ( .A(n18542), .X(n15731) );
  inv_x1_sg U9861 ( .A(n18541), .X(n15729) );
  inv_x1_sg U9862 ( .A(n18540), .X(n15727) );
  inv_x1_sg U9863 ( .A(n18539), .X(n15725) );
  inv_x1_sg U9864 ( .A(n18538), .X(n15723) );
  inv_x1_sg U9865 ( .A(n18537), .X(n15721) );
  inv_x1_sg U9866 ( .A(n18536), .X(n15719) );
  inv_x1_sg U9867 ( .A(n18535), .X(n15717) );
  inv_x1_sg U9868 ( .A(n18534), .X(n15715) );
  inv_x1_sg U9869 ( .A(n18533), .X(n15713) );
  inv_x1_sg U9870 ( .A(n18532), .X(n15711) );
  inv_x1_sg U9871 ( .A(n18531), .X(n15709) );
  inv_x1_sg U9872 ( .A(n18530), .X(n15707) );
  inv_x1_sg U9873 ( .A(n18529), .X(n15705) );
  inv_x1_sg U9874 ( .A(n18528), .X(n15703) );
  inv_x1_sg U9875 ( .A(n18527), .X(n15701) );
  inv_x1_sg U9876 ( .A(n18526), .X(n15699) );
  inv_x1_sg U9877 ( .A(n18525), .X(n15697) );
  inv_x1_sg U9878 ( .A(n18524), .X(n15695) );
  inv_x1_sg U9879 ( .A(n18523), .X(n15693) );
  inv_x1_sg U9880 ( .A(n18522), .X(n15691) );
  inv_x1_sg U9881 ( .A(n18521), .X(n15689) );
  inv_x1_sg U9882 ( .A(n18520), .X(n15687) );
  inv_x1_sg U9883 ( .A(n18519), .X(n15685) );
  inv_x1_sg U9884 ( .A(n18518), .X(n15683) );
  inv_x1_sg U9885 ( .A(n18517), .X(n15681) );
  inv_x1_sg U9886 ( .A(n18516), .X(n15679) );
  inv_x1_sg U9887 ( .A(n18515), .X(n15677) );
  inv_x1_sg U9888 ( .A(n18514), .X(n15675) );
  inv_x1_sg U9889 ( .A(n18513), .X(n15673) );
  inv_x1_sg U9890 ( .A(n18512), .X(n15671) );
  inv_x1_sg U9891 ( .A(n18511), .X(n15669) );
  inv_x1_sg U9892 ( .A(n18510), .X(n15667) );
  inv_x1_sg U9893 ( .A(n18509), .X(n15665) );
  inv_x1_sg U9894 ( .A(n18508), .X(n15663) );
  inv_x1_sg U9895 ( .A(n18507), .X(n15661) );
  inv_x1_sg U9896 ( .A(n18506), .X(n15659) );
  inv_x1_sg U9897 ( .A(n18505), .X(n15657) );
  inv_x1_sg U9898 ( .A(n18504), .X(n15655) );
  inv_x1_sg U9899 ( .A(n18503), .X(n15653) );
  inv_x1_sg U9900 ( .A(n18502), .X(n15651) );
  inv_x1_sg U9901 ( .A(n18501), .X(n15649) );
  inv_x1_sg U9902 ( .A(n18500), .X(n15647) );
  inv_x1_sg U9903 ( .A(n18499), .X(n15645) );
  inv_x1_sg U9904 ( .A(n18498), .X(n15643) );
  inv_x1_sg U9905 ( .A(n18497), .X(n15641) );
  inv_x1_sg U9906 ( .A(n18496), .X(n15639) );
  inv_x1_sg U9907 ( .A(n18495), .X(n15637) );
  inv_x1_sg U9908 ( .A(n18494), .X(n15635) );
  inv_x1_sg U9909 ( .A(n18493), .X(n15633) );
  inv_x1_sg U9910 ( .A(n18492), .X(n15631) );
  inv_x1_sg U9911 ( .A(n18491), .X(n15629) );
  inv_x1_sg U9912 ( .A(n18490), .X(n15627) );
  inv_x1_sg U9913 ( .A(n18489), .X(n15625) );
  inv_x1_sg U9914 ( .A(n18488), .X(n15623) );
  inv_x1_sg U9915 ( .A(n18487), .X(n15621) );
  inv_x1_sg U9916 ( .A(n18486), .X(n15619) );
  inv_x1_sg U9917 ( .A(n18485), .X(n15617) );
  inv_x1_sg U9918 ( .A(n18484), .X(n15615) );
  inv_x1_sg U9919 ( .A(n18483), .X(n15613) );
  inv_x1_sg U9920 ( .A(n18482), .X(n15611) );
  inv_x1_sg U9921 ( .A(n18481), .X(n15609) );
  inv_x1_sg U9922 ( .A(n18480), .X(n15607) );
  inv_x1_sg U9923 ( .A(n18479), .X(n15605) );
  inv_x1_sg U9924 ( .A(n18478), .X(n15603) );
  inv_x1_sg U9925 ( .A(n18477), .X(n15601) );
  inv_x1_sg U9926 ( .A(n18476), .X(n15599) );
  inv_x1_sg U9927 ( .A(n18475), .X(n15597) );
  inv_x1_sg U9928 ( .A(n18474), .X(n15595) );
  inv_x1_sg U9929 ( .A(n18473), .X(n15593) );
  inv_x1_sg U9930 ( .A(n18472), .X(n15591) );
  inv_x1_sg U9931 ( .A(n18471), .X(n15589) );
  inv_x1_sg U9932 ( .A(n18470), .X(n15587) );
  inv_x1_sg U9933 ( .A(n18469), .X(n15585) );
  inv_x1_sg U9934 ( .A(n18468), .X(n15583) );
  inv_x1_sg U9935 ( .A(n18467), .X(n15581) );
  inv_x1_sg U9936 ( .A(n18466), .X(n15579) );
  inv_x1_sg U9937 ( .A(n18465), .X(n15577) );
  inv_x1_sg U9938 ( .A(n18464), .X(n15575) );
  inv_x1_sg U9939 ( .A(n18463), .X(n15573) );
  inv_x1_sg U9940 ( .A(n18462), .X(n15571) );
  inv_x1_sg U9941 ( .A(n18461), .X(n15569) );
  inv_x1_sg U9942 ( .A(n18460), .X(n15567) );
  inv_x1_sg U9943 ( .A(n18459), .X(n15565) );
  inv_x1_sg U9944 ( .A(n18458), .X(n15563) );
  inv_x1_sg U9945 ( .A(n18457), .X(n15561) );
  inv_x1_sg U9946 ( .A(n18456), .X(n15559) );
  inv_x1_sg U9947 ( .A(n18455), .X(n15557) );
  inv_x1_sg U9948 ( .A(n18454), .X(n15555) );
  inv_x1_sg U9949 ( .A(n18453), .X(n15553) );
  inv_x1_sg U9950 ( .A(n18452), .X(n15551) );
  inv_x1_sg U9951 ( .A(n18451), .X(n15549) );
  inv_x1_sg U9952 ( .A(n18450), .X(n15547) );
  inv_x1_sg U9953 ( .A(n18449), .X(n15545) );
  inv_x1_sg U9954 ( .A(n18448), .X(n15543) );
  inv_x1_sg U9955 ( .A(n18447), .X(n15541) );
  inv_x1_sg U9956 ( .A(n18446), .X(n15539) );
  inv_x1_sg U9957 ( .A(n18445), .X(n15537) );
  inv_x1_sg U9958 ( .A(n18444), .X(n15535) );
  inv_x1_sg U9959 ( .A(n18443), .X(n15533) );
  inv_x1_sg U9960 ( .A(n18442), .X(n15531) );
  inv_x1_sg U9961 ( .A(n18441), .X(n15529) );
  inv_x1_sg U9962 ( .A(n18440), .X(n15527) );
  inv_x1_sg U9963 ( .A(n18439), .X(n15525) );
  inv_x1_sg U9964 ( .A(n18438), .X(n15523) );
  inv_x1_sg U9965 ( .A(n18437), .X(n15521) );
  inv_x1_sg U9966 ( .A(n18436), .X(n15519) );
  inv_x1_sg U9967 ( .A(n18435), .X(n15517) );
  inv_x1_sg U9968 ( .A(n18434), .X(n15515) );
  inv_x1_sg U9969 ( .A(n18433), .X(n15513) );
  inv_x1_sg U9970 ( .A(n18432), .X(n15511) );
  inv_x1_sg U9971 ( .A(n18431), .X(n15509) );
  inv_x1_sg U9972 ( .A(n18430), .X(n15507) );
  inv_x1_sg U9973 ( .A(n18429), .X(n15505) );
  inv_x1_sg U9974 ( .A(n18428), .X(n15503) );
  inv_x1_sg U9975 ( .A(n18427), .X(n15501) );
  inv_x1_sg U9976 ( .A(n18426), .X(n15499) );
  inv_x1_sg U9977 ( .A(n18425), .X(n15497) );
  inv_x1_sg U9978 ( .A(n18424), .X(n15495) );
  inv_x1_sg U9979 ( .A(n18423), .X(n15493) );
  inv_x1_sg U9980 ( .A(n18422), .X(n15491) );
  inv_x1_sg U9981 ( .A(n18421), .X(n15489) );
  inv_x1_sg U9982 ( .A(n18420), .X(n15487) );
  inv_x1_sg U9983 ( .A(n18419), .X(n15485) );
  inv_x1_sg U9984 ( .A(n18418), .X(n15483) );
  inv_x1_sg U9985 ( .A(n18417), .X(n15481) );
  inv_x1_sg U9986 ( .A(n18416), .X(n15479) );
  inv_x1_sg U9987 ( .A(n18415), .X(n15477) );
  inv_x1_sg U9988 ( .A(n18414), .X(n15475) );
  inv_x1_sg U9989 ( .A(n18413), .X(n15473) );
  inv_x1_sg U9990 ( .A(n18412), .X(n15471) );
  inv_x1_sg U9991 ( .A(n18411), .X(n15469) );
  inv_x1_sg U9992 ( .A(n18410), .X(n15467) );
  inv_x1_sg U9993 ( .A(n18409), .X(n15465) );
  inv_x1_sg U9994 ( .A(n18408), .X(n15463) );
  inv_x1_sg U9995 ( .A(n18407), .X(n15461) );
  inv_x1_sg U9996 ( .A(n18406), .X(n15459) );
  inv_x1_sg U9997 ( .A(n18405), .X(n15457) );
  inv_x1_sg U9998 ( .A(n18404), .X(n15455) );
  inv_x1_sg U9999 ( .A(n18403), .X(n15453) );
  inv_x1_sg U10000 ( .A(n18402), .X(n15451) );
  inv_x1_sg U10001 ( .A(n12859), .X(n18077) );
  inv_x1_sg U10002 ( .A(n12540), .X(n18396) );
  inv_x1_sg U10003 ( .A(n12541), .X(n18395) );
  inv_x1_sg U10004 ( .A(n12542), .X(n18394) );
  inv_x1_sg U10005 ( .A(n12543), .X(n18393) );
  inv_x1_sg U10006 ( .A(n12544), .X(n18392) );
  inv_x1_sg U10007 ( .A(n12545), .X(n18391) );
  inv_x1_sg U10008 ( .A(n12546), .X(n18390) );
  inv_x1_sg U10009 ( .A(n12547), .X(n18389) );
  inv_x1_sg U10010 ( .A(n12548), .X(n18388) );
  inv_x1_sg U10011 ( .A(n12549), .X(n18387) );
  inv_x1_sg U10012 ( .A(n12550), .X(n18386) );
  inv_x1_sg U10013 ( .A(n12551), .X(n18385) );
  inv_x1_sg U10014 ( .A(n12552), .X(n18384) );
  inv_x1_sg U10015 ( .A(n12553), .X(n18383) );
  inv_x1_sg U10016 ( .A(n12554), .X(n18382) );
  inv_x1_sg U10017 ( .A(n12555), .X(n18381) );
  inv_x1_sg U10018 ( .A(n12556), .X(n18380) );
  inv_x1_sg U10019 ( .A(n12557), .X(n18379) );
  inv_x1_sg U10020 ( .A(n12558), .X(n18378) );
  inv_x1_sg U10021 ( .A(n12559), .X(n18377) );
  inv_x1_sg U10022 ( .A(n12560), .X(n18376) );
  inv_x1_sg U10023 ( .A(n12561), .X(n18375) );
  inv_x1_sg U10024 ( .A(n12562), .X(n18374) );
  inv_x1_sg U10025 ( .A(n12563), .X(n18373) );
  inv_x1_sg U10026 ( .A(n12564), .X(n18372) );
  inv_x1_sg U10027 ( .A(n12565), .X(n18371) );
  inv_x1_sg U10028 ( .A(n12566), .X(n18370) );
  inv_x1_sg U10029 ( .A(n12567), .X(n18369) );
  inv_x1_sg U10030 ( .A(n12568), .X(n18368) );
  inv_x1_sg U10031 ( .A(n12569), .X(n18367) );
  inv_x1_sg U10032 ( .A(n12570), .X(n18366) );
  inv_x1_sg U10033 ( .A(n12571), .X(n18365) );
  inv_x1_sg U10034 ( .A(n12572), .X(n18364) );
  inv_x1_sg U10035 ( .A(n12573), .X(n18363) );
  inv_x1_sg U10036 ( .A(n12574), .X(n18362) );
  inv_x1_sg U10037 ( .A(n12575), .X(n18361) );
  inv_x1_sg U10038 ( .A(n12576), .X(n18360) );
  inv_x1_sg U10039 ( .A(n12577), .X(n18359) );
  inv_x1_sg U10040 ( .A(n12578), .X(n18358) );
  inv_x1_sg U10041 ( .A(n12579), .X(n18357) );
  inv_x1_sg U10042 ( .A(n12580), .X(n18356) );
  inv_x1_sg U10043 ( .A(n12581), .X(n18355) );
  inv_x1_sg U10044 ( .A(n12582), .X(n18354) );
  inv_x1_sg U10045 ( .A(n12583), .X(n18353) );
  inv_x1_sg U10046 ( .A(n12584), .X(n18352) );
  inv_x1_sg U10047 ( .A(n12585), .X(n18351) );
  inv_x1_sg U10048 ( .A(n12586), .X(n18350) );
  inv_x1_sg U10049 ( .A(n12587), .X(n18349) );
  inv_x1_sg U10050 ( .A(n12588), .X(n18348) );
  inv_x1_sg U10051 ( .A(n12589), .X(n18347) );
  inv_x1_sg U10052 ( .A(n12590), .X(n18346) );
  inv_x1_sg U10053 ( .A(n12591), .X(n18345) );
  inv_x1_sg U10054 ( .A(n12592), .X(n18344) );
  inv_x1_sg U10055 ( .A(n12593), .X(n18343) );
  inv_x1_sg U10056 ( .A(n12594), .X(n18342) );
  inv_x1_sg U10057 ( .A(n12595), .X(n18341) );
  inv_x1_sg U10058 ( .A(n12596), .X(n18340) );
  inv_x1_sg U10059 ( .A(n12597), .X(n18339) );
  inv_x1_sg U10060 ( .A(n12598), .X(n18338) );
  inv_x1_sg U10061 ( .A(n12599), .X(n18337) );
  inv_x1_sg U10062 ( .A(n12600), .X(n18336) );
  inv_x1_sg U10063 ( .A(n12601), .X(n18335) );
  inv_x1_sg U10064 ( .A(n12602), .X(n18334) );
  inv_x1_sg U10065 ( .A(n12603), .X(n18333) );
  inv_x1_sg U10066 ( .A(n12604), .X(n18332) );
  inv_x1_sg U10067 ( .A(n12605), .X(n18331) );
  inv_x1_sg U10068 ( .A(n12606), .X(n18330) );
  inv_x1_sg U10069 ( .A(n12607), .X(n18329) );
  inv_x1_sg U10070 ( .A(n12608), .X(n18328) );
  inv_x1_sg U10071 ( .A(n12609), .X(n18327) );
  inv_x1_sg U10072 ( .A(n12610), .X(n18326) );
  inv_x1_sg U10073 ( .A(n12611), .X(n18325) );
  inv_x1_sg U10074 ( .A(n12612), .X(n18324) );
  inv_x1_sg U10075 ( .A(n12613), .X(n18323) );
  inv_x1_sg U10076 ( .A(n12614), .X(n18322) );
  inv_x1_sg U10077 ( .A(n12615), .X(n18321) );
  inv_x1_sg U10078 ( .A(n12616), .X(n18320) );
  inv_x1_sg U10079 ( .A(n12617), .X(n18319) );
  inv_x1_sg U10080 ( .A(n12618), .X(n18318) );
  inv_x1_sg U10081 ( .A(n12619), .X(n18317) );
  inv_x1_sg U10082 ( .A(n12620), .X(n18316) );
  inv_x1_sg U10083 ( .A(n12621), .X(n18315) );
  inv_x1_sg U10084 ( .A(n12622), .X(n18314) );
  inv_x1_sg U10085 ( .A(n12623), .X(n18313) );
  inv_x1_sg U10086 ( .A(n12624), .X(n18312) );
  inv_x1_sg U10087 ( .A(n12625), .X(n18311) );
  inv_x1_sg U10088 ( .A(n12626), .X(n18310) );
  inv_x1_sg U10089 ( .A(n12627), .X(n18309) );
  inv_x1_sg U10090 ( .A(n12628), .X(n18308) );
  inv_x1_sg U10091 ( .A(n12629), .X(n18307) );
  inv_x1_sg U10092 ( .A(n12630), .X(n18306) );
  inv_x1_sg U10093 ( .A(n12631), .X(n18305) );
  inv_x1_sg U10094 ( .A(n12632), .X(n18304) );
  inv_x1_sg U10095 ( .A(n12633), .X(n18303) );
  inv_x1_sg U10096 ( .A(n12634), .X(n18302) );
  inv_x1_sg U10097 ( .A(n12635), .X(n18301) );
  inv_x1_sg U10098 ( .A(n12636), .X(n18300) );
  inv_x1_sg U10099 ( .A(n12637), .X(n18299) );
  inv_x1_sg U10100 ( .A(n12638), .X(n18298) );
  inv_x1_sg U10101 ( .A(n12639), .X(n18297) );
  inv_x1_sg U10102 ( .A(n12640), .X(n18296) );
  inv_x1_sg U10103 ( .A(n12641), .X(n18295) );
  inv_x1_sg U10104 ( .A(n12642), .X(n18294) );
  inv_x1_sg U10105 ( .A(n12643), .X(n18293) );
  inv_x1_sg U10106 ( .A(n12644), .X(n18292) );
  inv_x1_sg U10107 ( .A(n12645), .X(n18291) );
  inv_x1_sg U10108 ( .A(n12646), .X(n18290) );
  inv_x1_sg U10109 ( .A(n12647), .X(n18289) );
  inv_x1_sg U10110 ( .A(n12648), .X(n18288) );
  inv_x1_sg U10111 ( .A(n12649), .X(n18287) );
  inv_x1_sg U10112 ( .A(n12650), .X(n18286) );
  inv_x1_sg U10113 ( .A(n12651), .X(n18285) );
  inv_x1_sg U10114 ( .A(n12652), .X(n18284) );
  inv_x1_sg U10115 ( .A(n12653), .X(n18283) );
  inv_x1_sg U10116 ( .A(n12654), .X(n18282) );
  inv_x1_sg U10117 ( .A(n12655), .X(n18281) );
  inv_x1_sg U10118 ( .A(n12656), .X(n18280) );
  inv_x1_sg U10119 ( .A(n12657), .X(n18279) );
  inv_x1_sg U10120 ( .A(n12658), .X(n18278) );
  inv_x1_sg U10121 ( .A(n12659), .X(n18277) );
  inv_x1_sg U10122 ( .A(n12660), .X(n18276) );
  inv_x1_sg U10123 ( .A(n12661), .X(n18275) );
  inv_x1_sg U10124 ( .A(n12662), .X(n18274) );
  inv_x1_sg U10125 ( .A(n12663), .X(n18273) );
  inv_x1_sg U10126 ( .A(n12664), .X(n18272) );
  inv_x1_sg U10127 ( .A(n12665), .X(n18271) );
  inv_x1_sg U10128 ( .A(n12666), .X(n18270) );
  inv_x1_sg U10129 ( .A(n12667), .X(n18269) );
  inv_x1_sg U10130 ( .A(n12668), .X(n18268) );
  inv_x1_sg U10131 ( .A(n12669), .X(n18267) );
  inv_x1_sg U10132 ( .A(n12670), .X(n18266) );
  inv_x1_sg U10133 ( .A(n12671), .X(n18265) );
  inv_x1_sg U10134 ( .A(n12672), .X(n18264) );
  inv_x1_sg U10135 ( .A(n12673), .X(n18263) );
  inv_x1_sg U10136 ( .A(n12674), .X(n18262) );
  inv_x1_sg U10137 ( .A(n12675), .X(n18261) );
  inv_x1_sg U10138 ( .A(n12676), .X(n18260) );
  inv_x1_sg U10139 ( .A(n12677), .X(n18259) );
  inv_x1_sg U10140 ( .A(n12678), .X(n18258) );
  inv_x1_sg U10141 ( .A(n12679), .X(n18257) );
  inv_x1_sg U10142 ( .A(n12680), .X(n18256) );
  inv_x1_sg U10143 ( .A(n12681), .X(n18255) );
  inv_x1_sg U10144 ( .A(n12682), .X(n18254) );
  inv_x1_sg U10145 ( .A(n12683), .X(n18253) );
  inv_x1_sg U10146 ( .A(n12684), .X(n18252) );
  inv_x1_sg U10147 ( .A(n12685), .X(n18251) );
  inv_x1_sg U10148 ( .A(n12686), .X(n18250) );
  inv_x1_sg U10149 ( .A(n12687), .X(n18249) );
  inv_x1_sg U10150 ( .A(n12688), .X(n18248) );
  inv_x1_sg U10151 ( .A(n12689), .X(n18247) );
  inv_x1_sg U10152 ( .A(n12690), .X(n18246) );
  inv_x1_sg U10153 ( .A(n12691), .X(n18245) );
  inv_x1_sg U10154 ( .A(n12692), .X(n18244) );
  inv_x1_sg U10155 ( .A(n12693), .X(n18243) );
  inv_x1_sg U10156 ( .A(n12694), .X(n18242) );
  inv_x1_sg U10157 ( .A(n12695), .X(n18241) );
  inv_x1_sg U10158 ( .A(n12696), .X(n18240) );
  inv_x1_sg U10159 ( .A(n12697), .X(n18239) );
  inv_x1_sg U10160 ( .A(n12698), .X(n18238) );
  inv_x1_sg U10161 ( .A(n12699), .X(n18237) );
  inv_x1_sg U10162 ( .A(n12700), .X(n18236) );
  inv_x1_sg U10163 ( .A(n12701), .X(n18235) );
  inv_x1_sg U10164 ( .A(n12702), .X(n18234) );
  inv_x1_sg U10165 ( .A(n12703), .X(n18233) );
  inv_x1_sg U10166 ( .A(n12704), .X(n18232) );
  inv_x1_sg U10167 ( .A(n12705), .X(n18231) );
  inv_x1_sg U10168 ( .A(n12706), .X(n18230) );
  inv_x1_sg U10169 ( .A(n12707), .X(n18229) );
  inv_x1_sg U10170 ( .A(n12708), .X(n18228) );
  inv_x1_sg U10171 ( .A(n12709), .X(n18227) );
  inv_x1_sg U10172 ( .A(n12710), .X(n18226) );
  inv_x1_sg U10173 ( .A(n12711), .X(n18225) );
  inv_x1_sg U10174 ( .A(n12712), .X(n18224) );
  inv_x1_sg U10175 ( .A(n12713), .X(n18223) );
  inv_x1_sg U10176 ( .A(n12714), .X(n18222) );
  inv_x1_sg U10177 ( .A(n12715), .X(n18221) );
  inv_x1_sg U10178 ( .A(n12716), .X(n18220) );
  inv_x1_sg U10179 ( .A(n12717), .X(n18219) );
  inv_x1_sg U10180 ( .A(n12718), .X(n18218) );
  inv_x1_sg U10181 ( .A(n12719), .X(n18217) );
  inv_x1_sg U10182 ( .A(n12720), .X(n18216) );
  inv_x1_sg U10183 ( .A(n12721), .X(n18215) );
  inv_x1_sg U10184 ( .A(n12722), .X(n18214) );
  inv_x1_sg U10185 ( .A(n12723), .X(n18213) );
  inv_x1_sg U10186 ( .A(n12724), .X(n18212) );
  inv_x1_sg U10187 ( .A(n12725), .X(n18211) );
  inv_x1_sg U10188 ( .A(n12726), .X(n18210) );
  inv_x1_sg U10189 ( .A(n12727), .X(n18209) );
  inv_x1_sg U10190 ( .A(n12728), .X(n18208) );
  inv_x1_sg U10191 ( .A(n12729), .X(n18207) );
  inv_x1_sg U10192 ( .A(n12730), .X(n18206) );
  inv_x1_sg U10193 ( .A(n12731), .X(n18205) );
  inv_x1_sg U10194 ( .A(n12732), .X(n18204) );
  inv_x1_sg U10195 ( .A(n12733), .X(n18203) );
  inv_x1_sg U10196 ( .A(n12734), .X(n18202) );
  inv_x1_sg U10197 ( .A(n12735), .X(n18201) );
  inv_x1_sg U10198 ( .A(n12736), .X(n18200) );
  inv_x1_sg U10199 ( .A(n12737), .X(n18199) );
  inv_x1_sg U10200 ( .A(n12738), .X(n18198) );
  inv_x1_sg U10201 ( .A(n12739), .X(n18197) );
  inv_x1_sg U10202 ( .A(n12740), .X(n18196) );
  inv_x1_sg U10203 ( .A(n12741), .X(n18195) );
  inv_x1_sg U10204 ( .A(n12742), .X(n18194) );
  inv_x1_sg U10205 ( .A(n12743), .X(n18193) );
  inv_x1_sg U10206 ( .A(n12744), .X(n18192) );
  inv_x1_sg U10207 ( .A(n12745), .X(n18191) );
  inv_x1_sg U10208 ( .A(n12746), .X(n18190) );
  inv_x1_sg U10209 ( .A(n12747), .X(n18189) );
  inv_x1_sg U10210 ( .A(n12748), .X(n18188) );
  inv_x1_sg U10211 ( .A(n12749), .X(n18187) );
  inv_x1_sg U10212 ( .A(n12750), .X(n18186) );
  inv_x1_sg U10213 ( .A(n12751), .X(n18185) );
  inv_x1_sg U10214 ( .A(n12752), .X(n18184) );
  inv_x1_sg U10215 ( .A(n12753), .X(n18183) );
  inv_x1_sg U10216 ( .A(n12754), .X(n18182) );
  inv_x1_sg U10217 ( .A(n12755), .X(n18181) );
  inv_x1_sg U10218 ( .A(n12756), .X(n18180) );
  inv_x1_sg U10219 ( .A(n12757), .X(n18179) );
  inv_x1_sg U10220 ( .A(n12758), .X(n18178) );
  inv_x1_sg U10221 ( .A(n12759), .X(n18177) );
  inv_x1_sg U10222 ( .A(n12760), .X(n18176) );
  inv_x1_sg U10223 ( .A(n12761), .X(n18175) );
  inv_x1_sg U10224 ( .A(n12762), .X(n18174) );
  inv_x1_sg U10225 ( .A(n12763), .X(n18173) );
  inv_x1_sg U10226 ( .A(n12764), .X(n18172) );
  inv_x1_sg U10227 ( .A(n12765), .X(n18171) );
  inv_x1_sg U10228 ( .A(n12766), .X(n18170) );
  inv_x1_sg U10229 ( .A(n12767), .X(n18169) );
  inv_x1_sg U10230 ( .A(n12768), .X(n18168) );
  inv_x1_sg U10231 ( .A(n12769), .X(n18167) );
  inv_x1_sg U10232 ( .A(n12770), .X(n18166) );
  inv_x1_sg U10233 ( .A(n12771), .X(n18165) );
  inv_x1_sg U10234 ( .A(n12772), .X(n18164) );
  inv_x1_sg U10235 ( .A(n12773), .X(n18163) );
  inv_x1_sg U10236 ( .A(n12774), .X(n18162) );
  inv_x1_sg U10237 ( .A(n12775), .X(n18161) );
  inv_x1_sg U10238 ( .A(n12776), .X(n18160) );
  inv_x1_sg U10239 ( .A(n12777), .X(n18159) );
  inv_x1_sg U10240 ( .A(n12778), .X(n18158) );
  inv_x1_sg U10241 ( .A(n12779), .X(n18157) );
  inv_x1_sg U10242 ( .A(n12780), .X(n18156) );
  inv_x1_sg U10243 ( .A(n12781), .X(n18155) );
  inv_x1_sg U10244 ( .A(n12782), .X(n18154) );
  inv_x1_sg U10245 ( .A(n12783), .X(n18153) );
  inv_x1_sg U10246 ( .A(n12784), .X(n18152) );
  inv_x1_sg U10247 ( .A(n12785), .X(n18151) );
  inv_x1_sg U10248 ( .A(n12786), .X(n18150) );
  inv_x1_sg U10249 ( .A(n12787), .X(n18149) );
  inv_x1_sg U10250 ( .A(n12788), .X(n18148) );
  inv_x1_sg U10251 ( .A(n12789), .X(n18147) );
  inv_x1_sg U10252 ( .A(n12790), .X(n18146) );
  inv_x1_sg U10253 ( .A(n12791), .X(n18145) );
  inv_x1_sg U10254 ( .A(n12792), .X(n18144) );
  inv_x1_sg U10255 ( .A(n12793), .X(n18143) );
  inv_x1_sg U10256 ( .A(n12794), .X(n18142) );
  inv_x1_sg U10257 ( .A(n12795), .X(n18141) );
  inv_x1_sg U10258 ( .A(n12796), .X(n18140) );
  inv_x1_sg U10259 ( .A(n12797), .X(n18139) );
  inv_x1_sg U10260 ( .A(n12798), .X(n18138) );
  inv_x1_sg U10261 ( .A(n12799), .X(n18137) );
  inv_x1_sg U10262 ( .A(n12800), .X(n18136) );
  inv_x1_sg U10263 ( .A(n12801), .X(n18135) );
  inv_x1_sg U10264 ( .A(n12802), .X(n18134) );
  inv_x1_sg U10265 ( .A(n12803), .X(n18133) );
  inv_x1_sg U10266 ( .A(n12804), .X(n18132) );
  inv_x1_sg U10267 ( .A(n12805), .X(n18131) );
  inv_x1_sg U10268 ( .A(n12806), .X(n18130) );
  inv_x1_sg U10269 ( .A(n12807), .X(n18129) );
  inv_x1_sg U10270 ( .A(n12808), .X(n18128) );
  inv_x1_sg U10271 ( .A(n12809), .X(n18127) );
  inv_x1_sg U10272 ( .A(n12810), .X(n18126) );
  inv_x1_sg U10273 ( .A(n12811), .X(n18125) );
  inv_x1_sg U10274 ( .A(n12812), .X(n18124) );
  inv_x1_sg U10275 ( .A(n12813), .X(n18123) );
  inv_x1_sg U10276 ( .A(n12814), .X(n18122) );
  inv_x1_sg U10277 ( .A(n12815), .X(n18121) );
  inv_x1_sg U10278 ( .A(n12816), .X(n18120) );
  inv_x1_sg U10279 ( .A(n12817), .X(n18119) );
  inv_x1_sg U10280 ( .A(n12818), .X(n18118) );
  inv_x1_sg U10281 ( .A(n12819), .X(n18117) );
  inv_x1_sg U10282 ( .A(n12820), .X(n18116) );
  inv_x1_sg U10283 ( .A(n12821), .X(n18115) );
  inv_x1_sg U10284 ( .A(n12822), .X(n18114) );
  inv_x1_sg U10285 ( .A(n12823), .X(n18113) );
  inv_x1_sg U10286 ( .A(n12824), .X(n18112) );
  inv_x1_sg U10287 ( .A(n12825), .X(n18111) );
  inv_x1_sg U10288 ( .A(n12826), .X(n18110) );
  inv_x1_sg U10289 ( .A(n12827), .X(n18109) );
  inv_x1_sg U10290 ( .A(n12828), .X(n18108) );
  inv_x1_sg U10291 ( .A(n12829), .X(n18107) );
  inv_x1_sg U10292 ( .A(n12830), .X(n18106) );
  inv_x1_sg U10293 ( .A(n12831), .X(n18105) );
  inv_x1_sg U10294 ( .A(n12832), .X(n18104) );
  inv_x1_sg U10295 ( .A(n12833), .X(n18103) );
  inv_x1_sg U10296 ( .A(n12834), .X(n18102) );
  inv_x1_sg U10297 ( .A(n12835), .X(n18101) );
  inv_x1_sg U10298 ( .A(n12836), .X(n18100) );
  inv_x1_sg U10299 ( .A(n12837), .X(n18099) );
  inv_x1_sg U10300 ( .A(n12838), .X(n18098) );
  inv_x1_sg U10301 ( .A(n12839), .X(n18097) );
  inv_x1_sg U10302 ( .A(n12840), .X(n18096) );
  inv_x1_sg U10303 ( .A(n12841), .X(n18095) );
  inv_x1_sg U10304 ( .A(n12842), .X(n18094) );
  inv_x1_sg U10305 ( .A(n12843), .X(n18093) );
  inv_x1_sg U10306 ( .A(n12844), .X(n18092) );
  inv_x1_sg U10307 ( .A(n12845), .X(n18091) );
  inv_x1_sg U10308 ( .A(n12846), .X(n18090) );
  inv_x1_sg U10309 ( .A(n12847), .X(n18089) );
  inv_x1_sg U10310 ( .A(n12848), .X(n18088) );
  inv_x1_sg U10311 ( .A(n12849), .X(n18087) );
  inv_x1_sg U10312 ( .A(n12850), .X(n18086) );
  inv_x1_sg U10313 ( .A(n12851), .X(n18085) );
  inv_x1_sg U10314 ( .A(n12852), .X(n18084) );
  inv_x1_sg U10315 ( .A(n12853), .X(n18083) );
  inv_x1_sg U10316 ( .A(n12854), .X(n18082) );
  inv_x1_sg U10317 ( .A(n12855), .X(n18081) );
  inv_x1_sg U10318 ( .A(n12856), .X(n18080) );
  inv_x1_sg U10319 ( .A(n12857), .X(n18079) );
  inv_x1_sg U10320 ( .A(n12858), .X(n18078) );
  nand_x1_sg U10321 ( .A(n13764), .B(n13765), .X(n15091) );
  nand_x1_sg U10322 ( .A(n14483), .B(n16763), .X(n13764) );
  nand_x1_sg U10323 ( .A(n13766), .B(n13767), .X(n15092) );
  nand_x1_sg U10324 ( .A(n14484), .B(n16763), .X(n13766) );
  nand_x1_sg U10325 ( .A(n13758), .B(n13759), .X(n15088) );
  nand_x1_sg U10326 ( .A(n14485), .B(n16763), .X(n13758) );
  nand_x1_sg U10327 ( .A(n13760), .B(n13761), .X(n15089) );
  nand_x1_sg U10328 ( .A(n14486), .B(n16763), .X(n13760) );
  nand_x1_sg U10329 ( .A(n13776), .B(n13777), .X(n15097) );
  nand_x1_sg U10330 ( .A(n14487), .B(n16762), .X(n13776) );
  nand_x1_sg U10331 ( .A(n13778), .B(n13779), .X(n15098) );
  nand_x1_sg U10332 ( .A(n14488), .B(n16762), .X(n13778) );
  nand_x1_sg U10333 ( .A(n13770), .B(n13771), .X(n15094) );
  nand_x1_sg U10334 ( .A(n14489), .B(n16762), .X(n13770) );
  nand_x1_sg U10335 ( .A(n13772), .B(n13773), .X(n15095) );
  nand_x1_sg U10336 ( .A(n14490), .B(n16762), .X(n13772) );
  nand_x1_sg U10337 ( .A(n13740), .B(n13741), .X(n15079) );
  nand_x1_sg U10338 ( .A(n14491), .B(n16764), .X(n13740) );
  nand_x1_sg U10339 ( .A(n13742), .B(n13743), .X(n15080) );
  nand_x1_sg U10340 ( .A(n14492), .B(n16764), .X(n13742) );
  nand_x1_sg U10341 ( .A(n13734), .B(n13735), .X(n15076) );
  nand_x1_sg U10342 ( .A(n14493), .B(n16764), .X(n13734) );
  nand_x1_sg U10343 ( .A(n13736), .B(n13737), .X(n15077) );
  nand_x1_sg U10344 ( .A(n14494), .B(n16764), .X(n13736) );
  nand_x1_sg U10345 ( .A(n13752), .B(n13753), .X(n15085) );
  nand_x1_sg U10346 ( .A(n14495), .B(n16763), .X(n13752) );
  nand_x1_sg U10347 ( .A(n13754), .B(n13755), .X(n15086) );
  nand_x1_sg U10348 ( .A(n14496), .B(n16763), .X(n13754) );
  nand_x1_sg U10349 ( .A(n13746), .B(n13747), .X(n15082) );
  nand_x1_sg U10350 ( .A(n14497), .B(n16764), .X(n13746) );
  nand_x1_sg U10351 ( .A(n13748), .B(n13749), .X(n15083) );
  nand_x1_sg U10352 ( .A(n14498), .B(n16764), .X(n13748) );
  nand_x1_sg U10353 ( .A(n13812), .B(n13813), .X(n15115) );
  nand_x1_sg U10354 ( .A(n14499), .B(n16772), .X(n13812) );
  nand_x1_sg U10355 ( .A(n13814), .B(n13815), .X(n15116) );
  nand_x1_sg U10356 ( .A(n14500), .B(n16771), .X(n13814) );
  nand_x1_sg U10357 ( .A(n13806), .B(n13807), .X(n15112) );
  nand_x1_sg U10358 ( .A(n14501), .B(n16772), .X(n13806) );
  nand_x1_sg U10359 ( .A(n13808), .B(n13809), .X(n15113) );
  nand_x1_sg U10360 ( .A(n14502), .B(n16771), .X(n13808) );
  nand_x1_sg U10361 ( .A(n13824), .B(n13825), .X(n15121) );
  nand_x1_sg U10362 ( .A(n14503), .B(n16768), .X(n13824) );
  nand_x1_sg U10363 ( .A(n13826), .B(n13827), .X(n15122) );
  nand_x1_sg U10364 ( .A(n14504), .B(n16771), .X(n13826) );
  nand_x1_sg U10365 ( .A(n13818), .B(n13819), .X(n15118) );
  nand_x1_sg U10366 ( .A(n14505), .B(n16771), .X(n13818) );
  nand_x1_sg U10367 ( .A(n13820), .B(n13821), .X(n15119) );
  nand_x1_sg U10368 ( .A(n14506), .B(n16771), .X(n13820) );
  nand_x1_sg U10369 ( .A(n13788), .B(n13789), .X(n15103) );
  nand_x1_sg U10370 ( .A(n14507), .B(n16771), .X(n13788) );
  nand_x1_sg U10371 ( .A(n13790), .B(n13791), .X(n15104) );
  nand_x1_sg U10372 ( .A(n14508), .B(n16761), .X(n13790) );
  nand_x1_sg U10373 ( .A(n13782), .B(n13783), .X(n15100) );
  nand_x1_sg U10374 ( .A(n14509), .B(n16762), .X(n13782) );
  nand_x1_sg U10375 ( .A(n13784), .B(n13785), .X(n15101) );
  nand_x1_sg U10376 ( .A(n14510), .B(n16762), .X(n13784) );
  nand_x1_sg U10377 ( .A(n13800), .B(n13801), .X(n15109) );
  nand_x1_sg U10378 ( .A(n14511), .B(n16772), .X(n13800) );
  nand_x1_sg U10379 ( .A(n13802), .B(n13803), .X(n15110) );
  nand_x1_sg U10380 ( .A(n14512), .B(n16771), .X(n13802) );
  nand_x1_sg U10381 ( .A(n13794), .B(n13795), .X(n15106) );
  nand_x1_sg U10382 ( .A(n14513), .B(n16771), .X(n13794) );
  nand_x1_sg U10383 ( .A(n13796), .B(n13797), .X(n15107) );
  nand_x1_sg U10384 ( .A(n14514), .B(n16761), .X(n13796) );
  nand_x1_sg U10385 ( .A(n13668), .B(n13669), .X(n15043) );
  nand_x1_sg U10386 ( .A(n14515), .B(n16768), .X(n13668) );
  nand_x1_sg U10387 ( .A(n13670), .B(n13671), .X(n15044) );
  nand_x1_sg U10388 ( .A(n14516), .B(n16768), .X(n13670) );
  nand_x1_sg U10389 ( .A(n13662), .B(n13663), .X(n15040) );
  nand_x1_sg U10390 ( .A(n14517), .B(n16769), .X(n13662) );
  nand_x1_sg U10391 ( .A(n13664), .B(n13665), .X(n15041) );
  nand_x1_sg U10392 ( .A(n14518), .B(n16768), .X(n13664) );
  nand_x1_sg U10393 ( .A(n13680), .B(n13681), .X(n15049) );
  nand_x1_sg U10394 ( .A(n14519), .B(n16767), .X(n13680) );
  nand_x1_sg U10395 ( .A(n13682), .B(n13683), .X(n15050) );
  nand_x1_sg U10396 ( .A(n14520), .B(n16767), .X(n13682) );
  nand_x1_sg U10397 ( .A(n13674), .B(n13675), .X(n15046) );
  nand_x1_sg U10398 ( .A(n14521), .B(n16768), .X(n13674) );
  nand_x1_sg U10399 ( .A(n13676), .B(n13677), .X(n15047) );
  nand_x1_sg U10400 ( .A(n14522), .B(n16768), .X(n13676) );
  nand_x1_sg U10401 ( .A(n13644), .B(n13645), .X(n15031) );
  nand_x1_sg U10402 ( .A(n14523), .B(n16771), .X(n13644) );
  nand_x1_sg U10403 ( .A(n13646), .B(n13647), .X(n15032) );
  nand_x1_sg U10404 ( .A(n14524), .B(n16769), .X(n13646) );
  nand_x1_sg U10405 ( .A(n13638), .B(n13639), .X(n15028) );
  nand_x1_sg U10406 ( .A(n14525), .B(n16761), .X(n13638) );
  nand_x1_sg U10407 ( .A(n13640), .B(n13641), .X(n15029) );
  nand_x1_sg U10408 ( .A(n14526), .B(n16761), .X(n13640) );
  nand_x1_sg U10409 ( .A(n13656), .B(n13657), .X(n15037) );
  nand_x1_sg U10410 ( .A(n14527), .B(n16769), .X(n13656) );
  nand_x1_sg U10411 ( .A(n13658), .B(n13659), .X(n15038) );
  nand_x1_sg U10412 ( .A(n14528), .B(n16769), .X(n13658) );
  nand_x1_sg U10413 ( .A(n13650), .B(n13651), .X(n15034) );
  nand_x1_sg U10414 ( .A(n14529), .B(n16769), .X(n13650) );
  nand_x1_sg U10415 ( .A(n13652), .B(n13653), .X(n15035) );
  nand_x1_sg U10416 ( .A(n14530), .B(n16769), .X(n13652) );
  nand_x1_sg U10417 ( .A(n13716), .B(n13717), .X(n15067) );
  nand_x1_sg U10418 ( .A(n14531), .B(n16765), .X(n13716) );
  nand_x1_sg U10419 ( .A(n13718), .B(n13719), .X(n15068) );
  nand_x1_sg U10420 ( .A(n14532), .B(n16765), .X(n13718) );
  nand_x1_sg U10421 ( .A(n13710), .B(n13711), .X(n15064) );
  nand_x1_sg U10422 ( .A(n14533), .B(n16766), .X(n13710) );
  nand_x1_sg U10423 ( .A(n13712), .B(n13713), .X(n15065) );
  nand_x1_sg U10424 ( .A(n14534), .B(n16766), .X(n13712) );
  nand_x1_sg U10425 ( .A(n13728), .B(n13729), .X(n15073) );
  nand_x1_sg U10426 ( .A(n14535), .B(n16765), .X(n13728) );
  nand_x1_sg U10427 ( .A(n13730), .B(n13731), .X(n15074) );
  nand_x1_sg U10428 ( .A(n14536), .B(n16765), .X(n13730) );
  nand_x1_sg U10429 ( .A(n13722), .B(n13723), .X(n15070) );
  nand_x1_sg U10430 ( .A(n14537), .B(n16765), .X(n13722) );
  nand_x1_sg U10431 ( .A(n13724), .B(n13725), .X(n15071) );
  nand_x1_sg U10432 ( .A(n14538), .B(n16765), .X(n13724) );
  nand_x1_sg U10433 ( .A(n13692), .B(n13693), .X(n15055) );
  nand_x1_sg U10434 ( .A(n14539), .B(n16767), .X(n13692) );
  nand_x1_sg U10435 ( .A(n13694), .B(n13695), .X(n15056) );
  nand_x1_sg U10436 ( .A(n14540), .B(n16767), .X(n13694) );
  nand_x1_sg U10437 ( .A(n13686), .B(n13687), .X(n15052) );
  nand_x1_sg U10438 ( .A(n14541), .B(n16767), .X(n13686) );
  nand_x1_sg U10439 ( .A(n13688), .B(n13689), .X(n15053) );
  nand_x1_sg U10440 ( .A(n14542), .B(n16767), .X(n13688) );
  nand_x1_sg U10441 ( .A(n13704), .B(n13705), .X(n15061) );
  nand_x1_sg U10442 ( .A(n14543), .B(n16766), .X(n13704) );
  nand_x1_sg U10443 ( .A(n13706), .B(n13707), .X(n15062) );
  nand_x1_sg U10444 ( .A(n14544), .B(n16766), .X(n13706) );
  nand_x1_sg U10445 ( .A(n13698), .B(n13699), .X(n15058) );
  nand_x1_sg U10446 ( .A(n14545), .B(n16766), .X(n13698) );
  nand_x1_sg U10447 ( .A(n13700), .B(n13701), .X(n15059) );
  nand_x1_sg U10448 ( .A(n14546), .B(n16766), .X(n13700) );
  nand_x1_sg U10449 ( .A(n13378), .B(n13379), .X(n14898) );
  nand_x1_sg U10450 ( .A(n14547), .B(n16772), .X(n13378) );
  nand_x1_sg U10451 ( .A(n13380), .B(n13381), .X(n14899) );
  nand_x1_sg U10452 ( .A(n14548), .B(n16772), .X(n13380) );
  nand_x1_sg U10453 ( .A(n13372), .B(n13373), .X(n14895) );
  nand_x1_sg U10454 ( .A(n14549), .B(n16761), .X(n13372) );
  nand_x1_sg U10455 ( .A(n13374), .B(n13375), .X(n14896) );
  nand_x1_sg U10456 ( .A(n14550), .B(n16771), .X(n13374) );
  nand_x1_sg U10457 ( .A(n13390), .B(n13391), .X(n14904) );
  nand_x1_sg U10458 ( .A(n14551), .B(n16761), .X(n13390) );
  nand_x1_sg U10459 ( .A(n13392), .B(n13393), .X(n14905) );
  nand_x1_sg U10460 ( .A(n14552), .B(n16772), .X(n13392) );
  nand_x1_sg U10461 ( .A(n13384), .B(n13385), .X(n14901) );
  nand_x1_sg U10462 ( .A(n14553), .B(n16771), .X(n13384) );
  nand_x1_sg U10463 ( .A(n13386), .B(n13387), .X(n14902) );
  nand_x1_sg U10464 ( .A(n14554), .B(n16772), .X(n13386) );
  nand_x1_sg U10465 ( .A(n13354), .B(n13355), .X(n14886) );
  nand_x1_sg U10466 ( .A(n14555), .B(n16771), .X(n13354) );
  nand_x1_sg U10467 ( .A(n13356), .B(n13357), .X(n14887) );
  nand_x1_sg U10468 ( .A(n14556), .B(n16771), .X(n13356) );
  nand_x1_sg U10469 ( .A(n13348), .B(n13349), .X(n14883) );
  nand_x1_sg U10470 ( .A(n14557), .B(n16771), .X(n13348) );
  nand_x1_sg U10471 ( .A(n13350), .B(n13351), .X(n14884) );
  nand_x1_sg U10472 ( .A(n14558), .B(n16772), .X(n13350) );
  nand_x1_sg U10473 ( .A(n13366), .B(n13367), .X(n14892) );
  nand_x1_sg U10474 ( .A(n14559), .B(n16772), .X(n13366) );
  nand_x1_sg U10475 ( .A(n13368), .B(n13369), .X(n14893) );
  nand_x1_sg U10476 ( .A(n14560), .B(n16761), .X(n13368) );
  nand_x1_sg U10477 ( .A(n13360), .B(n13361), .X(n14889) );
  nand_x1_sg U10478 ( .A(n14561), .B(n16772), .X(n13360) );
  nand_x1_sg U10479 ( .A(n13362), .B(n13363), .X(n14890) );
  nand_x1_sg U10480 ( .A(n14562), .B(n16761), .X(n13362) );
  nand_x1_sg U10481 ( .A(n13426), .B(n13427), .X(n14922) );
  nand_x1_sg U10482 ( .A(n14563), .B(n16761), .X(n13426) );
  nand_x1_sg U10483 ( .A(n13428), .B(n13429), .X(n14923) );
  nand_x1_sg U10484 ( .A(n14564), .B(n16761), .X(n13428) );
  nand_x1_sg U10485 ( .A(n13420), .B(n13421), .X(n14919) );
  nand_x1_sg U10486 ( .A(n14565), .B(n16771), .X(n13420) );
  nand_x1_sg U10487 ( .A(n13422), .B(n13423), .X(n14920) );
  nand_x1_sg U10488 ( .A(n14566), .B(n16771), .X(n13422) );
  nand_x1_sg U10489 ( .A(n13438), .B(n13439), .X(n14928) );
  nand_x1_sg U10490 ( .A(n14567), .B(n16772), .X(n13438) );
  nand_x1_sg U10491 ( .A(n13440), .B(n13441), .X(n14929) );
  nand_x1_sg U10492 ( .A(n14568), .B(n16761), .X(n13440) );
  nand_x1_sg U10493 ( .A(n13432), .B(n13433), .X(n14925) );
  nand_x1_sg U10494 ( .A(n14569), .B(n16771), .X(n13432) );
  nand_x1_sg U10495 ( .A(n13434), .B(n13435), .X(n14926) );
  nand_x1_sg U10496 ( .A(n14570), .B(n16771), .X(n13434) );
  nand_x1_sg U10497 ( .A(n13402), .B(n13403), .X(n14910) );
  nand_x1_sg U10498 ( .A(n14571), .B(n16772), .X(n13402) );
  nand_x1_sg U10499 ( .A(n13404), .B(n13405), .X(n14911) );
  nand_x1_sg U10500 ( .A(n14572), .B(n16761), .X(n13404) );
  nand_x1_sg U10501 ( .A(n13396), .B(n13397), .X(n14907) );
  nand_x1_sg U10502 ( .A(n14573), .B(n16761), .X(n13396) );
  nand_x1_sg U10503 ( .A(n13398), .B(n13399), .X(n14908) );
  nand_x1_sg U10504 ( .A(n14574), .B(n16761), .X(n13398) );
  nand_x1_sg U10505 ( .A(n13414), .B(n13415), .X(n14916) );
  nand_x1_sg U10506 ( .A(n14575), .B(n16771), .X(n13414) );
  nand_x1_sg U10507 ( .A(n13416), .B(n13417), .X(n14917) );
  nand_x1_sg U10508 ( .A(n14576), .B(n16771), .X(n13416) );
  nand_x1_sg U10509 ( .A(n13408), .B(n13409), .X(n14913) );
  nand_x1_sg U10510 ( .A(n14577), .B(n16772), .X(n13408) );
  nand_x1_sg U10511 ( .A(n13410), .B(n13411), .X(n14914) );
  nand_x1_sg U10512 ( .A(n14578), .B(n16761), .X(n13410) );
  nand_x1_sg U10513 ( .A(n13282), .B(n13283), .X(n14850) );
  nand_x1_sg U10514 ( .A(n14579), .B(n16772), .X(n13282) );
  nand_x1_sg U10515 ( .A(n13284), .B(n13285), .X(n14851) );
  nand_x1_sg U10516 ( .A(n14580), .B(n16771), .X(n13284) );
  nand_x1_sg U10517 ( .A(n13276), .B(n13277), .X(n14847) );
  nand_x1_sg U10518 ( .A(n14581), .B(n16771), .X(n13276) );
  nand_x1_sg U10519 ( .A(n13278), .B(n13279), .X(n14848) );
  nand_x1_sg U10520 ( .A(n14582), .B(n16772), .X(n13278) );
  nand_x1_sg U10521 ( .A(n13294), .B(n13295), .X(n14856) );
  nand_x1_sg U10522 ( .A(n14583), .B(n16761), .X(n13294) );
  nand_x1_sg U10523 ( .A(n13296), .B(n13297), .X(n14857) );
  nand_x1_sg U10524 ( .A(n14584), .B(n16771), .X(n13296) );
  nand_x1_sg U10525 ( .A(n13288), .B(n13289), .X(n14853) );
  nand_x1_sg U10526 ( .A(n14585), .B(n16761), .X(n13288) );
  nand_x1_sg U10527 ( .A(n13290), .B(n13291), .X(n14854) );
  nand_x1_sg U10528 ( .A(n14586), .B(n16771), .X(n13290) );
  nand_x1_sg U10529 ( .A(n13258), .B(n13259), .X(n14838) );
  nand_x1_sg U10530 ( .A(n14587), .B(n16761), .X(n13258) );
  nand_x1_sg U10531 ( .A(n13260), .B(n13261), .X(n14839) );
  nand_x1_sg U10532 ( .A(n14588), .B(n16771), .X(n13260) );
  nand_x1_sg U10533 ( .A(n13252), .B(n13253), .X(n14835) );
  nand_x1_sg U10534 ( .A(n14589), .B(n16761), .X(n13252) );
  nand_x1_sg U10535 ( .A(n13254), .B(n13255), .X(n14836) );
  nand_x1_sg U10536 ( .A(n14590), .B(n16761), .X(n13254) );
  nand_x1_sg U10537 ( .A(n13270), .B(n13271), .X(n14844) );
  nand_x1_sg U10538 ( .A(n14591), .B(n16771), .X(n13270) );
  nand_x1_sg U10539 ( .A(n13272), .B(n13273), .X(n14845) );
  nand_x1_sg U10540 ( .A(n14592), .B(n16761), .X(n13272) );
  nand_x1_sg U10541 ( .A(n13264), .B(n13265), .X(n14841) );
  nand_x1_sg U10542 ( .A(n14593), .B(n16771), .X(n13264) );
  nand_x1_sg U10543 ( .A(n13266), .B(n13267), .X(n14842) );
  nand_x1_sg U10544 ( .A(n14594), .B(n16771), .X(n13266) );
  nand_x1_sg U10545 ( .A(n13330), .B(n13331), .X(n14874) );
  nand_x1_sg U10546 ( .A(n14595), .B(n16761), .X(n13330) );
  nand_x1_sg U10547 ( .A(n13332), .B(n13333), .X(n14875) );
  nand_x1_sg U10548 ( .A(n14596), .B(n16772), .X(n13332) );
  nand_x1_sg U10549 ( .A(n13324), .B(n13325), .X(n14871) );
  nand_x1_sg U10550 ( .A(n14597), .B(n16771), .X(n13324) );
  nand_x1_sg U10551 ( .A(n13326), .B(n13327), .X(n14872) );
  nand_x1_sg U10552 ( .A(n14598), .B(n16761), .X(n13326) );
  nand_x1_sg U10553 ( .A(n13342), .B(n13343), .X(n14880) );
  nand_x1_sg U10554 ( .A(n14599), .B(n16771), .X(n13342) );
  nand_x1_sg U10555 ( .A(n13344), .B(n13345), .X(n14881) );
  nand_x1_sg U10556 ( .A(n14600), .B(n16761), .X(n13344) );
  nand_x1_sg U10557 ( .A(n13336), .B(n13337), .X(n14877) );
  nand_x1_sg U10558 ( .A(n14601), .B(n16761), .X(n13336) );
  nand_x1_sg U10559 ( .A(n13338), .B(n13339), .X(n14878) );
  nand_x1_sg U10560 ( .A(n14602), .B(n16771), .X(n13338) );
  nand_x1_sg U10561 ( .A(n13306), .B(n13307), .X(n14862) );
  nand_x1_sg U10562 ( .A(n14603), .B(n16772), .X(n13306) );
  nand_x1_sg U10563 ( .A(n13308), .B(n13309), .X(n14863) );
  nand_x1_sg U10564 ( .A(n14604), .B(n16761), .X(n13308) );
  nand_x1_sg U10565 ( .A(n13300), .B(n13301), .X(n14859) );
  nand_x1_sg U10566 ( .A(n14605), .B(n16761), .X(n13300) );
  nand_x1_sg U10567 ( .A(n13302), .B(n13303), .X(n14860) );
  nand_x1_sg U10568 ( .A(n14606), .B(n16761), .X(n13302) );
  nand_x1_sg U10569 ( .A(n13318), .B(n13319), .X(n14868) );
  nand_x1_sg U10570 ( .A(n14607), .B(n16761), .X(n13318) );
  nand_x1_sg U10571 ( .A(n13320), .B(n13321), .X(n14869) );
  nand_x1_sg U10572 ( .A(n14608), .B(n16771), .X(n13320) );
  nand_x1_sg U10573 ( .A(n13312), .B(n13313), .X(n14865) );
  nand_x1_sg U10574 ( .A(n14609), .B(n16772), .X(n13312) );
  nand_x1_sg U10575 ( .A(n13314), .B(n13315), .X(n14866) );
  nand_x1_sg U10576 ( .A(n14610), .B(n16772), .X(n13314) );
  nand_x1_sg U10577 ( .A(n13570), .B(n13571), .X(n14994) );
  nand_x1_sg U10578 ( .A(n14611), .B(n16761), .X(n13570) );
  nand_x1_sg U10579 ( .A(n13572), .B(n13573), .X(n14995) );
  nand_x1_sg U10580 ( .A(n14612), .B(n16772), .X(n13572) );
  nand_x1_sg U10581 ( .A(n13564), .B(n13565), .X(n14991) );
  nand_x1_sg U10582 ( .A(n14613), .B(n16761), .X(n13564) );
  nand_x1_sg U10583 ( .A(n13566), .B(n13567), .X(n14992) );
  nand_x1_sg U10584 ( .A(n14614), .B(n16772), .X(n13566) );
  nand_x1_sg U10585 ( .A(n13582), .B(n13583), .X(n15000) );
  nand_x1_sg U10586 ( .A(n14615), .B(n16772), .X(n13582) );
  nand_x1_sg U10587 ( .A(n13584), .B(n13585), .X(n15001) );
  nand_x1_sg U10588 ( .A(n14616), .B(n16761), .X(n13584) );
  nand_x1_sg U10589 ( .A(n13576), .B(n13577), .X(n14997) );
  nand_x1_sg U10590 ( .A(n14617), .B(n16761), .X(n13576) );
  nand_x1_sg U10591 ( .A(n13578), .B(n13579), .X(n14998) );
  nand_x1_sg U10592 ( .A(n14618), .B(n16772), .X(n13578) );
  nand_x1_sg U10593 ( .A(n13546), .B(n13547), .X(n14982) );
  nand_x1_sg U10594 ( .A(n14619), .B(n16772), .X(n13546) );
  nand_x1_sg U10595 ( .A(n13548), .B(n13549), .X(n14983) );
  nand_x1_sg U10596 ( .A(n14620), .B(n16772), .X(n13548) );
  nand_x1_sg U10597 ( .A(n13540), .B(n13541), .X(n14979) );
  nand_x1_sg U10598 ( .A(n14621), .B(n16772), .X(n13540) );
  nand_x1_sg U10599 ( .A(n13542), .B(n13543), .X(n14980) );
  nand_x1_sg U10600 ( .A(n14622), .B(n16771), .X(n13542) );
  nand_x1_sg U10601 ( .A(n13558), .B(n13559), .X(n14988) );
  nand_x1_sg U10602 ( .A(n14623), .B(n16771), .X(n13558) );
  nand_x1_sg U10603 ( .A(n13560), .B(n13561), .X(n14989) );
  nand_x1_sg U10604 ( .A(n14624), .B(n16771), .X(n13560) );
  nand_x1_sg U10605 ( .A(n13552), .B(n13553), .X(n14985) );
  nand_x1_sg U10606 ( .A(n14625), .B(n16771), .X(n13552) );
  nand_x1_sg U10607 ( .A(n13554), .B(n13555), .X(n14986) );
  nand_x1_sg U10608 ( .A(n14626), .B(n16774), .X(n13554) );
  nand_x1_sg U10609 ( .A(n13618), .B(n13619), .X(n15018) );
  nand_x1_sg U10610 ( .A(n14627), .B(n16761), .X(n13618) );
  nand_x1_sg U10611 ( .A(n13620), .B(n13621), .X(n15019) );
  nand_x1_sg U10612 ( .A(n14628), .B(n16761), .X(n13620) );
  nand_x1_sg U10613 ( .A(n13612), .B(n13613), .X(n15015) );
  nand_x1_sg U10614 ( .A(n14629), .B(n16771), .X(n13612) );
  nand_x1_sg U10615 ( .A(n13614), .B(n13615), .X(n15016) );
  nand_x1_sg U10616 ( .A(n14630), .B(n16772), .X(n13614) );
  nand_x1_sg U10617 ( .A(n13630), .B(n13631), .X(n15024) );
  nand_x1_sg U10618 ( .A(n14631), .B(n16772), .X(n13630) );
  nand_x1_sg U10619 ( .A(n13632), .B(n13633), .X(n15025) );
  nand_x1_sg U10620 ( .A(n14632), .B(n16761), .X(n13632) );
  nand_x1_sg U10621 ( .A(n13624), .B(n13625), .X(n15021) );
  nand_x1_sg U10622 ( .A(n14633), .B(n16771), .X(n13624) );
  nand_x1_sg U10623 ( .A(n13626), .B(n13627), .X(n15022) );
  nand_x1_sg U10624 ( .A(n14634), .B(n16771), .X(n13626) );
  nand_x1_sg U10625 ( .A(n13594), .B(n13595), .X(n15006) );
  nand_x1_sg U10626 ( .A(n14635), .B(n16771), .X(n13594) );
  nand_x1_sg U10627 ( .A(n13596), .B(n13597), .X(n15007) );
  nand_x1_sg U10628 ( .A(n14636), .B(n16772), .X(n13596) );
  nand_x1_sg U10629 ( .A(n13588), .B(n13589), .X(n15003) );
  nand_x1_sg U10630 ( .A(n14637), .B(n16772), .X(n13588) );
  nand_x1_sg U10631 ( .A(n13590), .B(n13591), .X(n15004) );
  nand_x1_sg U10632 ( .A(n14638), .B(n16761), .X(n13590) );
  nand_x1_sg U10633 ( .A(n13606), .B(n13607), .X(n15012) );
  nand_x1_sg U10634 ( .A(n14639), .B(n16774), .X(n13606) );
  nand_x1_sg U10635 ( .A(n13608), .B(n13609), .X(n15013) );
  nand_x1_sg U10636 ( .A(n14640), .B(n16774), .X(n13608) );
  nand_x1_sg U10637 ( .A(n13600), .B(n13601), .X(n15009) );
  nand_x1_sg U10638 ( .A(n14641), .B(n16761), .X(n13600) );
  nand_x1_sg U10639 ( .A(n13602), .B(n13603), .X(n15010) );
  nand_x1_sg U10640 ( .A(n14642), .B(n16771), .X(n13602) );
  nand_x1_sg U10641 ( .A(n13474), .B(n13475), .X(n14946) );
  nand_x1_sg U10642 ( .A(n14643), .B(n16772), .X(n13474) );
  nand_x1_sg U10643 ( .A(n13476), .B(n13477), .X(n14947) );
  nand_x1_sg U10644 ( .A(n14644), .B(n16771), .X(n13476) );
  nand_x1_sg U10645 ( .A(n13468), .B(n13469), .X(n14943) );
  nand_x1_sg U10646 ( .A(n14645), .B(n16761), .X(n13468) );
  nand_x1_sg U10647 ( .A(n13470), .B(n13471), .X(n14944) );
  nand_x1_sg U10648 ( .A(n14646), .B(n16771), .X(n13470) );
  nand_x1_sg U10649 ( .A(n13486), .B(n13487), .X(n14952) );
  nand_x1_sg U10650 ( .A(n14647), .B(n16772), .X(n13486) );
  nand_x1_sg U10651 ( .A(n13488), .B(n13489), .X(n14953) );
  nand_x1_sg U10652 ( .A(n14648), .B(n16771), .X(n13488) );
  nand_x1_sg U10653 ( .A(n13480), .B(n13481), .X(n14949) );
  nand_x1_sg U10654 ( .A(n14649), .B(n16772), .X(n13480) );
  nand_x1_sg U10655 ( .A(n13482), .B(n13483), .X(n14950) );
  nand_x1_sg U10656 ( .A(n14650), .B(n16771), .X(n13482) );
  nand_x1_sg U10657 ( .A(n13450), .B(n13451), .X(n14934) );
  nand_x1_sg U10658 ( .A(n14651), .B(n16771), .X(n13450) );
  nand_x1_sg U10659 ( .A(n13452), .B(n13453), .X(n14935) );
  nand_x1_sg U10660 ( .A(n14652), .B(n16774), .X(n13452) );
  nand_x1_sg U10661 ( .A(n13444), .B(n13445), .X(n14931) );
  nand_x1_sg U10662 ( .A(n14653), .B(n16772), .X(n13444) );
  nand_x1_sg U10663 ( .A(n13446), .B(n13447), .X(n14932) );
  nand_x1_sg U10664 ( .A(n14654), .B(n16771), .X(n13446) );
  nand_x1_sg U10665 ( .A(n13462), .B(n13463), .X(n14940) );
  nand_x1_sg U10666 ( .A(n14655), .B(n16761), .X(n13462) );
  nand_x1_sg U10667 ( .A(n13464), .B(n13465), .X(n14941) );
  nand_x1_sg U10668 ( .A(n14656), .B(n16771), .X(n13464) );
  nand_x1_sg U10669 ( .A(n13456), .B(n13457), .X(n14937) );
  nand_x1_sg U10670 ( .A(n14657), .B(n16771), .X(n13456) );
  nand_x1_sg U10671 ( .A(n13458), .B(n13459), .X(n14938) );
  nand_x1_sg U10672 ( .A(n14658), .B(n16772), .X(n13458) );
  nand_x1_sg U10673 ( .A(n13522), .B(n13523), .X(n14970) );
  nand_x1_sg U10674 ( .A(n14659), .B(n16772), .X(n13522) );
  nand_x1_sg U10675 ( .A(n13524), .B(n13525), .X(n14971) );
  nand_x1_sg U10676 ( .A(n14660), .B(n16761), .X(n13524) );
  nand_x1_sg U10677 ( .A(n13516), .B(n13517), .X(n14967) );
  nand_x1_sg U10678 ( .A(n14661), .B(n16761), .X(n13516) );
  nand_x1_sg U10679 ( .A(n13518), .B(n13519), .X(n14968) );
  nand_x1_sg U10680 ( .A(n14662), .B(n16772), .X(n13518) );
  nand_x1_sg U10681 ( .A(n13534), .B(n13535), .X(n14976) );
  nand_x1_sg U10682 ( .A(n14663), .B(n16772), .X(n13534) );
  nand_x1_sg U10683 ( .A(n13536), .B(n13537), .X(n14977) );
  nand_x1_sg U10684 ( .A(n14664), .B(n16761), .X(n13536) );
  nand_x1_sg U10685 ( .A(n13528), .B(n13529), .X(n14973) );
  nand_x1_sg U10686 ( .A(n14665), .B(n16772), .X(n13528) );
  nand_x1_sg U10687 ( .A(n13530), .B(n13531), .X(n14974) );
  nand_x1_sg U10688 ( .A(n14666), .B(n16771), .X(n13530) );
  nand_x1_sg U10689 ( .A(n13498), .B(n13499), .X(n14958) );
  nand_x1_sg U10690 ( .A(n14667), .B(n16772), .X(n13498) );
  nand_x1_sg U10691 ( .A(n13500), .B(n13501), .X(n14959) );
  nand_x1_sg U10692 ( .A(n14668), .B(n16761), .X(n13500) );
  nand_x1_sg U10693 ( .A(n13492), .B(n13493), .X(n14955) );
  nand_x1_sg U10694 ( .A(n14669), .B(n16771), .X(n13492) );
  nand_x1_sg U10695 ( .A(n13494), .B(n13495), .X(n14956) );
  nand_x1_sg U10696 ( .A(n14670), .B(n16771), .X(n13494) );
  nand_x1_sg U10697 ( .A(n13510), .B(n13511), .X(n14964) );
  nand_x1_sg U10698 ( .A(n14671), .B(n16772), .X(n13510) );
  nand_x1_sg U10699 ( .A(n13512), .B(n13513), .X(n14965) );
  nand_x1_sg U10700 ( .A(n14672), .B(n16771), .X(n13512) );
  nand_x1_sg U10701 ( .A(n13504), .B(n13505), .X(n14961) );
  nand_x1_sg U10702 ( .A(n14673), .B(n16776), .X(n13504) );
  nand_x1_sg U10703 ( .A(n13506), .B(n13507), .X(n14962) );
  nand_x1_sg U10704 ( .A(n14674), .B(n16772), .X(n13506) );
  nand_x1_sg U10705 ( .A(n13256), .B(n13257), .X(n14837) );
  nand_x1_sg U10706 ( .A(n14675), .B(n16761), .X(n13256) );
  nand_x1_sg U10707 ( .A(n13786), .B(n13787), .X(n15102) );
  nand_x1_sg U10708 ( .A(n14676), .B(n16762), .X(n13786) );
  nand_x1_sg U10709 ( .A(n13322), .B(n13323), .X(n14870) );
  nand_x1_sg U10710 ( .A(n14677), .B(n16761), .X(n13322) );
  nand_x1_sg U10711 ( .A(n13634), .B(n13635), .X(n15026) );
  nand_x1_sg U10712 ( .A(n14678), .B(n16771), .X(n13634) );
  nand_x1_sg U10713 ( .A(n13222), .B(n13223), .X(n14820) );
  nand_x1_sg U10714 ( .A(n14679), .B(n16772), .X(n13222) );
  nand_x1_sg U10715 ( .A(n13298), .B(n13299), .X(n14858) );
  nand_x1_sg U10716 ( .A(n14680), .B(n16771), .X(n13298) );
  nand_x1_sg U10717 ( .A(n13346), .B(n13347), .X(n14882) );
  nand_x1_sg U10718 ( .A(n14681), .B(n16771), .X(n13346) );
  nand_x1_sg U10719 ( .A(n13376), .B(n13377), .X(n14897) );
  nand_x1_sg U10720 ( .A(n14682), .B(n16761), .X(n13376) );
  nand_x1_sg U10721 ( .A(n13478), .B(n13479), .X(n14948) );
  nand_x1_sg U10722 ( .A(n14683), .B(n16772), .X(n13478) );
  nand_x1_sg U10723 ( .A(n13762), .B(n13763), .X(n15090) );
  nand_x1_sg U10724 ( .A(n14684), .B(n16763), .X(n13762) );
  nand_x1_sg U10725 ( .A(n13780), .B(n13781), .X(n15099) );
  nand_x1_sg U10726 ( .A(n14685), .B(n16762), .X(n13780) );
  nand_x1_sg U10727 ( .A(n13556), .B(n13557), .X(n14987) );
  nand_x1_sg U10728 ( .A(n14686), .B(n16761), .X(n13556) );
  nand_x1_sg U10729 ( .A(n13684), .B(n13685), .X(n15051) );
  nand_x1_sg U10730 ( .A(n14687), .B(n16767), .X(n13684) );
  nand_x1_sg U10731 ( .A(n13194), .B(n13195), .X(n14806) );
  nand_x1_sg U10732 ( .A(n14688), .B(n16771), .X(n13194) );
  nand_x1_sg U10733 ( .A(n13280), .B(n13281), .X(n14849) );
  nand_x1_sg U10734 ( .A(n14689), .B(n16772), .X(n13280) );
  nand_x1_sg U10735 ( .A(n13198), .B(n13199), .X(n14808) );
  nand_x1_sg U10736 ( .A(n14690), .B(n16761), .X(n13198) );
  nand_x1_sg U10737 ( .A(n13400), .B(n13401), .X(n14909) );
  nand_x1_sg U10738 ( .A(n14691), .B(n16772), .X(n13400) );
  nand_x1_sg U10739 ( .A(n13394), .B(n13395), .X(n14906) );
  nand_x1_sg U10740 ( .A(n14692), .B(n16772), .X(n13394) );
  nand_x1_sg U10741 ( .A(n13196), .B(n13197), .X(n14807) );
  nand_x1_sg U10742 ( .A(n14693), .B(n16761), .X(n13196) );
  nand_x1_sg U10743 ( .A(n13364), .B(n13365), .X(n14891) );
  nand_x1_sg U10744 ( .A(n14694), .B(n16761), .X(n13364) );
  nand_x1_sg U10745 ( .A(n13744), .B(n13745), .X(n15081) );
  nand_x1_sg U10746 ( .A(n14695), .B(n16764), .X(n13744) );
  nand_x1_sg U10747 ( .A(n13250), .B(n13251), .X(n14834) );
  nand_x1_sg U10748 ( .A(n14696), .B(n16761), .X(n13250) );
  nand_x1_sg U10749 ( .A(n13328), .B(n13329), .X(n14873) );
  nand_x1_sg U10750 ( .A(n14697), .B(n16772), .X(n13328) );
  nand_x1_sg U10751 ( .A(n13292), .B(n13293), .X(n14855) );
  nand_x1_sg U10752 ( .A(n14698), .B(n16761), .X(n13292) );
  nand_x1_sg U10753 ( .A(n13636), .B(n13637), .X(n15027) );
  nand_x1_sg U10754 ( .A(n14699), .B(n16761), .X(n13636) );
  nand_x1_sg U10755 ( .A(n13642), .B(n13643), .X(n15030) );
  nand_x1_sg U10756 ( .A(n14700), .B(n16772), .X(n13642) );
  nand_x1_sg U10757 ( .A(n13574), .B(n13575), .X(n14996) );
  nand_x1_sg U10758 ( .A(n14701), .B(n16761), .X(n13574) );
  nand_x1_sg U10759 ( .A(n13810), .B(n13811), .X(n15114) );
  nand_x1_sg U10760 ( .A(n14702), .B(n16761), .X(n13810) );
  nand_x1_sg U10761 ( .A(n13690), .B(n13691), .X(n15054) );
  nand_x1_sg U10762 ( .A(n14703), .B(n16767), .X(n13690) );
  nand_x1_sg U10763 ( .A(n13696), .B(n13697), .X(n15057) );
  nand_x1_sg U10764 ( .A(n14704), .B(n16767), .X(n13696) );
  nand_x1_sg U10765 ( .A(n13720), .B(n13721), .X(n15069) );
  nand_x1_sg U10766 ( .A(n14705), .B(n16765), .X(n13720) );
  nand_x1_sg U10767 ( .A(n13774), .B(n13775), .X(n15096) );
  nand_x1_sg U10768 ( .A(n14706), .B(n16762), .X(n13774) );
  nand_x1_sg U10769 ( .A(n13514), .B(n13515), .X(n14966) );
  nand_x1_sg U10770 ( .A(n14707), .B(n16761), .X(n13514) );
  nand_x1_sg U10771 ( .A(n13230), .B(n13231), .X(n14824) );
  nand_x1_sg U10772 ( .A(n14708), .B(n16771), .X(n13230) );
  nand_x1_sg U10773 ( .A(n13208), .B(n13209), .X(n14813) );
  nand_x1_sg U10774 ( .A(n14709), .B(n16771), .X(n13208) );
  nand_x1_sg U10775 ( .A(n13708), .B(n13709), .X(n15063) );
  nand_x1_sg U10776 ( .A(n14710), .B(n16766), .X(n13708) );
  nand_x1_sg U10777 ( .A(n13604), .B(n13605), .X(n15011) );
  nand_x1_sg U10778 ( .A(n14711), .B(n16771), .X(n13604) );
  nand_x1_sg U10779 ( .A(n13214), .B(n13215), .X(n14816) );
  nand_x1_sg U10780 ( .A(n14712), .B(n16761), .X(n13214) );
  nand_x1_sg U10781 ( .A(n13210), .B(n13211), .X(n14814) );
  nand_x1_sg U10782 ( .A(n14713), .B(n16771), .X(n13210) );
  nand_x1_sg U10783 ( .A(n13822), .B(n13823), .X(n15120) );
  nand_x1_sg U10784 ( .A(n14714), .B(n16771), .X(n13822) );
  nand_x1_sg U10785 ( .A(n13220), .B(n13221), .X(n14819) );
  nand_x1_sg U10786 ( .A(n14715), .B(n16772), .X(n13220) );
  nand_x1_sg U10787 ( .A(n13212), .B(n13213), .X(n14815) );
  nand_x1_sg U10788 ( .A(n14716), .B(n16761), .X(n13212) );
  nand_x1_sg U10789 ( .A(n13202), .B(n13203), .X(n14810) );
  nand_x1_sg U10790 ( .A(n14717), .B(n16761), .X(n13202) );
  nand_x1_sg U10791 ( .A(n13204), .B(n13205), .X(n14811) );
  nand_x1_sg U10792 ( .A(n14718), .B(n16761), .X(n13204) );
  nand_x1_sg U10793 ( .A(n13460), .B(n13461), .X(n14939) );
  nand_x1_sg U10794 ( .A(n14719), .B(n16761), .X(n13460) );
  nand_x1_sg U10795 ( .A(n13496), .B(n13497), .X(n14957) );
  nand_x1_sg U10796 ( .A(n14720), .B(n16771), .X(n13496) );
  nand_x1_sg U10797 ( .A(n13206), .B(n13207), .X(n14812) );
  nand_x1_sg U10798 ( .A(n14721), .B(n16772), .X(n13206) );
  nand_x1_sg U10799 ( .A(n13430), .B(n13431), .X(n14924) );
  nand_x1_sg U10800 ( .A(n14722), .B(n16772), .X(n13430) );
  nand_x1_sg U10801 ( .A(n13654), .B(n13655), .X(n15036) );
  nand_x1_sg U10802 ( .A(n14723), .B(n16769), .X(n13654) );
  nand_x1_sg U10803 ( .A(n13660), .B(n13661), .X(n15039) );
  nand_x1_sg U10804 ( .A(n14724), .B(n16769), .X(n13660) );
  nand_x1_sg U10805 ( .A(n13726), .B(n13727), .X(n15072) );
  nand_x1_sg U10806 ( .A(n14725), .B(n16765), .X(n13726) );
  nand_x1_sg U10807 ( .A(n13672), .B(n13673), .X(n15045) );
  nand_x1_sg U10808 ( .A(n14726), .B(n16768), .X(n13672) );
  nand_x1_sg U10809 ( .A(n13702), .B(n13703), .X(n15060) );
  nand_x1_sg U10810 ( .A(n14727), .B(n16766), .X(n13702) );
  nand_x1_sg U10811 ( .A(n13666), .B(n13667), .X(n15042) );
  nand_x1_sg U10812 ( .A(n14728), .B(n16768), .X(n13666) );
  nand_x1_sg U10813 ( .A(n13678), .B(n13679), .X(n15048) );
  nand_x1_sg U10814 ( .A(n14729), .B(n16768), .X(n13678) );
  nand_x1_sg U10815 ( .A(n13792), .B(n13793), .X(n15105) );
  nand_x1_sg U10816 ( .A(n14730), .B(n16771), .X(n13792) );
  nand_x1_sg U10817 ( .A(n13580), .B(n13581), .X(n14999) );
  nand_x1_sg U10818 ( .A(n14731), .B(n16771), .X(n13580) );
  nand_x1_sg U10819 ( .A(n13714), .B(n13715), .X(n15066) );
  nand_x1_sg U10820 ( .A(n14732), .B(n16766), .X(n13714) );
  nand_x1_sg U10821 ( .A(n13228), .B(n13229), .X(n14823) );
  nand_x1_sg U10822 ( .A(n14733), .B(n16772), .X(n13228) );
  nand_x1_sg U10823 ( .A(n13648), .B(n13649), .X(n15033) );
  nand_x1_sg U10824 ( .A(n14734), .B(n16769), .X(n13648) );
  nand_x1_sg U10825 ( .A(n13232), .B(n13233), .X(n14825) );
  nand_x1_sg U10826 ( .A(n14735), .B(n16761), .X(n13232) );
  nand_x1_sg U10827 ( .A(n13238), .B(n13239), .X(n14828) );
  nand_x1_sg U10828 ( .A(n14736), .B(n16761), .X(n13238) );
  nand_x1_sg U10829 ( .A(n13244), .B(n13245), .X(n14831) );
  nand_x1_sg U10830 ( .A(n14737), .B(n16761), .X(n13244) );
  nand_x1_sg U10831 ( .A(n13610), .B(n13611), .X(n15014) );
  nand_x1_sg U10832 ( .A(n14738), .B(n16772), .X(n13610) );
  nand_x1_sg U10833 ( .A(n13502), .B(n13503), .X(n14960) );
  nand_x1_sg U10834 ( .A(n14739), .B(n16772), .X(n13502) );
  nand_x1_sg U10835 ( .A(n13508), .B(n13509), .X(n14963) );
  nand_x1_sg U10836 ( .A(n14740), .B(n16771), .X(n13508) );
  nand_x1_sg U10837 ( .A(n13216), .B(n13217), .X(n14817) );
  nand_x1_sg U10838 ( .A(n14741), .B(n16771), .X(n13216) );
  nand_x1_sg U10839 ( .A(n13218), .B(n13219), .X(n14818) );
  nand_x1_sg U10840 ( .A(n14742), .B(n16761), .X(n13218) );
  nand_x1_sg U10841 ( .A(n13520), .B(n13521), .X(n14969) );
  nand_x1_sg U10842 ( .A(n14743), .B(n16771), .X(n13520) );
  nand_x1_sg U10843 ( .A(n13526), .B(n13527), .X(n14972) );
  nand_x1_sg U10844 ( .A(n14744), .B(n16771), .X(n13526) );
  nand_x1_sg U10845 ( .A(n13532), .B(n13533), .X(n14975) );
  nand_x1_sg U10846 ( .A(n14745), .B(n16761), .X(n13532) );
  nand_x1_sg U10847 ( .A(n13538), .B(n13539), .X(n14978) );
  nand_x1_sg U10848 ( .A(n14746), .B(n16771), .X(n13538) );
  nand_x1_sg U10849 ( .A(n13466), .B(n13467), .X(n14942) );
  nand_x1_sg U10850 ( .A(n14747), .B(n16761), .X(n13466) );
  nand_x1_sg U10851 ( .A(n13472), .B(n13473), .X(n14945) );
  nand_x1_sg U10852 ( .A(n14748), .B(n16772), .X(n13472) );
  nand_x1_sg U10853 ( .A(n13484), .B(n13485), .X(n14951) );
  nand_x1_sg U10854 ( .A(n14749), .B(n16774), .X(n13484) );
  nand_x1_sg U10855 ( .A(n13490), .B(n13491), .X(n14954) );
  nand_x1_sg U10856 ( .A(n14750), .B(n16771), .X(n13490) );
  nand_x1_sg U10857 ( .A(n13436), .B(n13437), .X(n14927) );
  nand_x1_sg U10858 ( .A(n14751), .B(n16761), .X(n13436) );
  nand_x1_sg U10859 ( .A(n13442), .B(n13443), .X(n14930) );
  nand_x1_sg U10860 ( .A(n14752), .B(n16774), .X(n13442) );
  nand_x1_sg U10861 ( .A(n13448), .B(n13449), .X(n14933) );
  nand_x1_sg U10862 ( .A(n14753), .B(n16771), .X(n13448) );
  nand_x1_sg U10863 ( .A(n13454), .B(n13455), .X(n14936) );
  nand_x1_sg U10864 ( .A(n14754), .B(n16772), .X(n13454) );
  nand_x1_sg U10865 ( .A(n13616), .B(n13617), .X(n15017) );
  nand_x1_sg U10866 ( .A(n14755), .B(n16772), .X(n13616) );
  nand_x1_sg U10867 ( .A(n13622), .B(n13623), .X(n15020) );
  nand_x1_sg U10868 ( .A(n14756), .B(n16761), .X(n13622) );
  nand_x1_sg U10869 ( .A(n13246), .B(n13247), .X(n14832) );
  nand_x1_sg U10870 ( .A(n14757), .B(n16761), .X(n13246) );
  nand_x1_sg U10871 ( .A(n13628), .B(n13629), .X(n15023) );
  nand_x1_sg U10872 ( .A(n14758), .B(n16761), .X(n13628) );
  nand_x1_sg U10873 ( .A(n13586), .B(n13587), .X(n15002) );
  nand_x1_sg U10874 ( .A(n14759), .B(n16771), .X(n13586) );
  nand_x1_sg U10875 ( .A(n13592), .B(n13593), .X(n15005) );
  nand_x1_sg U10876 ( .A(n14760), .B(n16772), .X(n13592) );
  nand_x1_sg U10877 ( .A(n13248), .B(n13249), .X(n14833) );
  nand_x1_sg U10878 ( .A(n14761), .B(n16761), .X(n13248) );
  nand_x1_sg U10879 ( .A(n13598), .B(n13599), .X(n15008) );
  nand_x1_sg U10880 ( .A(n14762), .B(n16772), .X(n13598) );
  nand_x1_sg U10881 ( .A(n13544), .B(n13545), .X(n14981) );
  nand_x1_sg U10882 ( .A(n14763), .B(n16771), .X(n13544) );
  nand_x1_sg U10883 ( .A(n13550), .B(n13551), .X(n14984) );
  nand_x1_sg U10884 ( .A(n14764), .B(n16774), .X(n13550) );
  nand_x1_sg U10885 ( .A(n13562), .B(n13563), .X(n14990) );
  nand_x1_sg U10886 ( .A(n14765), .B(n16761), .X(n13562) );
  nand_x1_sg U10887 ( .A(n13568), .B(n13569), .X(n14993) );
  nand_x1_sg U10888 ( .A(n14766), .B(n16771), .X(n13568) );
  nand_x1_sg U10889 ( .A(n13240), .B(n13241), .X(n14829) );
  nand_x1_sg U10890 ( .A(n14767), .B(n16771), .X(n13240) );
  nand_x1_sg U10891 ( .A(n13242), .B(n13243), .X(n14830) );
  nand_x1_sg U10892 ( .A(n14768), .B(n16761), .X(n13242) );
  nand_x1_sg U10893 ( .A(n13234), .B(n13235), .X(n14826) );
  nand_x1_sg U10894 ( .A(n14769), .B(n16771), .X(n13234) );
  nand_x1_sg U10895 ( .A(n13236), .B(n13237), .X(n14827) );
  nand_x1_sg U10896 ( .A(n14770), .B(n16772), .X(n13236) );
  nand_x1_sg U10897 ( .A(n13186), .B(n13187), .X(n14803) );
  nand_x1_sg U10898 ( .A(n14771), .B(n16771), .X(n13186) );
  nand_x1_sg U10899 ( .A(n13190), .B(n13191), .X(n14804) );
  nand_x1_sg U10900 ( .A(n14772), .B(n16771), .X(n13190) );
  nand_x1_sg U10901 ( .A(n13756), .B(n13757), .X(n15087) );
  nand_x1_sg U10902 ( .A(n14773), .B(n16763), .X(n13756) );
  nand_x1_sg U10903 ( .A(n13750), .B(n13751), .X(n15084) );
  nand_x1_sg U10904 ( .A(n14774), .B(n16764), .X(n13750) );
  nand_x1_sg U10905 ( .A(n13268), .B(n13269), .X(n14843) );
  nand_x1_sg U10906 ( .A(n14775), .B(n16771), .X(n13268) );
  nand_x1_sg U10907 ( .A(n13274), .B(n13275), .X(n14846) );
  nand_x1_sg U10908 ( .A(n14776), .B(n16771), .X(n13274) );
  nand_x1_sg U10909 ( .A(n13192), .B(n13193), .X(n14805) );
  nand_x1_sg U10910 ( .A(n14777), .B(n16761), .X(n13192) );
  nand_x1_sg U10911 ( .A(n13286), .B(n13287), .X(n14852) );
  nand_x1_sg U10912 ( .A(n14778), .B(n16771), .X(n13286) );
  nand_x1_sg U10913 ( .A(n13798), .B(n13799), .X(n15108) );
  nand_x1_sg U10914 ( .A(n14779), .B(n16761), .X(n13798) );
  nand_x1_sg U10915 ( .A(n13804), .B(n13805), .X(n15111) );
  nand_x1_sg U10916 ( .A(n14780), .B(n16761), .X(n13804) );
  nand_x1_sg U10917 ( .A(n13262), .B(n13263), .X(n14840) );
  nand_x1_sg U10918 ( .A(n14781), .B(n16761), .X(n13262) );
  nand_x1_sg U10919 ( .A(n13816), .B(n13817), .X(n15117) );
  nand_x1_sg U10920 ( .A(n14782), .B(n16772), .X(n13816) );
  nand_x1_sg U10921 ( .A(n13732), .B(n13733), .X(n15075) );
  nand_x1_sg U10922 ( .A(n14783), .B(n16765), .X(n13732) );
  nand_x1_sg U10923 ( .A(n13738), .B(n13739), .X(n15078) );
  nand_x1_sg U10924 ( .A(n14784), .B(n16764), .X(n13738) );
  nand_x1_sg U10925 ( .A(n13200), .B(n13201), .X(n14809) );
  nand_x1_sg U10926 ( .A(n14785), .B(n16772), .X(n13200) );
  nand_x1_sg U10927 ( .A(n13768), .B(n13769), .X(n15093) );
  nand_x1_sg U10928 ( .A(n14786), .B(n16763), .X(n13768) );
  nand_x1_sg U10929 ( .A(n13382), .B(n13383), .X(n14900) );
  nand_x1_sg U10930 ( .A(n14787), .B(n16772), .X(n13382) );
  nand_x1_sg U10931 ( .A(n13388), .B(n13389), .X(n14903) );
  nand_x1_sg U10932 ( .A(n14788), .B(n16771), .X(n13388) );
  nand_x1_sg U10933 ( .A(n13406), .B(n13407), .X(n14912) );
  nand_x1_sg U10934 ( .A(n14789), .B(n16771), .X(n13406) );
  nand_x1_sg U10935 ( .A(n13412), .B(n13413), .X(n14915) );
  nand_x1_sg U10936 ( .A(n14790), .B(n16771), .X(n13412) );
  nand_x1_sg U10937 ( .A(n13352), .B(n13353), .X(n14885) );
  nand_x1_sg U10938 ( .A(n14791), .B(n16772), .X(n13352) );
  nand_x1_sg U10939 ( .A(n13358), .B(n13359), .X(n14888) );
  nand_x1_sg U10940 ( .A(n14792), .B(n16772), .X(n13358) );
  nand_x1_sg U10941 ( .A(n13418), .B(n13419), .X(n14918) );
  nand_x1_sg U10942 ( .A(n14793), .B(n16761), .X(n13418) );
  nand_x1_sg U10943 ( .A(n13370), .B(n13371), .X(n14894) );
  nand_x1_sg U10944 ( .A(n14794), .B(n16761), .X(n13370) );
  nand_x1_sg U10945 ( .A(n13304), .B(n13305), .X(n14861) );
  nand_x1_sg U10946 ( .A(n14795), .B(n16772), .X(n13304) );
  nand_x1_sg U10947 ( .A(n13310), .B(n13311), .X(n14864) );
  nand_x1_sg U10948 ( .A(n14796), .B(n16761), .X(n13310) );
  nand_x1_sg U10949 ( .A(n13226), .B(n13227), .X(n14822) );
  nand_x1_sg U10950 ( .A(n14797), .B(n16771), .X(n13226) );
  nand_x1_sg U10951 ( .A(n13316), .B(n13317), .X(n14867) );
  nand_x1_sg U10952 ( .A(n14798), .B(n16761), .X(n13316) );
  nand_x1_sg U10953 ( .A(n13334), .B(n13335), .X(n14876) );
  nand_x1_sg U10954 ( .A(n14799), .B(n16771), .X(n13334) );
  nand_x1_sg U10955 ( .A(n13340), .B(n13341), .X(n14879) );
  nand_x1_sg U10956 ( .A(n14800), .B(n16772), .X(n13340) );
  nand_x1_sg U10957 ( .A(n13224), .B(n13225), .X(n14821) );
  nand_x1_sg U10958 ( .A(n14801), .B(n16772), .X(n13224) );
  nand_x1_sg U10959 ( .A(n13424), .B(n13425), .X(n14921) );
  nand_x1_sg U10960 ( .A(n14802), .B(n16772), .X(n13424) );
  nand_x1_sg U10961 ( .A(n14220), .B(n14221), .X(n15318) );
  nand_x1_sg U10962 ( .A(\in[0][0][0] ), .B(n16737), .X(n14220) );
  nand_x1_sg U10963 ( .A(n14188), .B(n14189), .X(n15302) );
  nand_x1_sg U10964 ( .A(\in[0][0][1] ), .B(n16738), .X(n14188) );
  nand_x1_sg U10965 ( .A(n14190), .B(n14191), .X(n15303) );
  nand_x1_sg U10966 ( .A(\in[0][0][2] ), .B(n16739), .X(n14190) );
  nand_x1_sg U10967 ( .A(n14182), .B(n14183), .X(n15299) );
  nand_x1_sg U10968 ( .A(\in[0][0][3] ), .B(n16738), .X(n14182) );
  nand_x1_sg U10969 ( .A(n14184), .B(n14185), .X(n15300) );
  nand_x1_sg U10970 ( .A(\in[0][0][4] ), .B(n16739), .X(n14184) );
  nand_x1_sg U10971 ( .A(n14200), .B(n14201), .X(n15308) );
  nand_x1_sg U10972 ( .A(\in[0][0][5] ), .B(n16737), .X(n14200) );
  nand_x1_sg U10973 ( .A(n14202), .B(n14203), .X(n15309) );
  nand_x1_sg U10974 ( .A(\in[0][0][6] ), .B(n16739), .X(n14202) );
  nand_x1_sg U10975 ( .A(n14194), .B(n14195), .X(n15305) );
  nand_x1_sg U10976 ( .A(\in[0][0][7] ), .B(n16738), .X(n14194) );
  nand_x1_sg U10977 ( .A(n14196), .B(n14197), .X(n15306) );
  nand_x1_sg U10978 ( .A(\in[0][0][8] ), .B(n16739), .X(n14196) );
  nand_x1_sg U10979 ( .A(n14260), .B(n14261), .X(n15338) );
  nand_x1_sg U10980 ( .A(\in[0][0][9] ), .B(n16739), .X(n14260) );
  nand_x1_sg U10981 ( .A(n14262), .B(n14263), .X(n15339) );
  nand_x1_sg U10982 ( .A(\in[0][0][10] ), .B(n16739), .X(n14262) );
  nand_x1_sg U10983 ( .A(n14254), .B(n14255), .X(n15335) );
  nand_x1_sg U10984 ( .A(\in[0][0][11] ), .B(n16739), .X(n14254) );
  nand_x1_sg U10985 ( .A(n14256), .B(n14257), .X(n15336) );
  nand_x1_sg U10986 ( .A(\in[0][0][12] ), .B(n16739), .X(n14256) );
  nand_x1_sg U10987 ( .A(n14272), .B(n14273), .X(n15344) );
  nand_x1_sg U10988 ( .A(\in[0][0][13] ), .B(n16738), .X(n14272) );
  nand_x1_sg U10989 ( .A(n14274), .B(n14275), .X(n15345) );
  nand_x1_sg U10990 ( .A(\in[0][0][14] ), .B(n16738), .X(n14274) );
  nand_x1_sg U10991 ( .A(n14266), .B(n14267), .X(n15341) );
  nand_x1_sg U10992 ( .A(\in[0][0][15] ), .B(n16739), .X(n14266) );
  nand_x1_sg U10993 ( .A(n14268), .B(n14269), .X(n15342) );
  nand_x1_sg U10994 ( .A(\in[0][0][16] ), .B(n16739), .X(n14268) );
  nand_x1_sg U10995 ( .A(n14236), .B(n14237), .X(n15326) );
  nand_x1_sg U10996 ( .A(\in[0][0][17] ), .B(n16736), .X(n14236) );
  nand_x1_sg U10997 ( .A(n14238), .B(n14239), .X(n15327) );
  nand_x1_sg U10998 ( .A(\in[0][0][18] ), .B(n16736), .X(n14238) );
  nand_x1_sg U10999 ( .A(n14230), .B(n14231), .X(n15323) );
  nand_x1_sg U11000 ( .A(\in[0][0][19] ), .B(n16736), .X(n14230) );
  nand_x1_sg U11001 ( .A(n14232), .B(n14233), .X(n15324) );
  nand_x1_sg U11002 ( .A(\in[0][1][0] ), .B(n16738), .X(n14232) );
  nand_x1_sg U11003 ( .A(n14248), .B(n14249), .X(n15332) );
  nand_x1_sg U11004 ( .A(\in[0][1][1] ), .B(n16737), .X(n14248) );
  nand_x1_sg U11005 ( .A(n14250), .B(n14251), .X(n15333) );
  nand_x1_sg U11006 ( .A(\in[0][1][2] ), .B(n16738), .X(n14250) );
  nand_x1_sg U11007 ( .A(n14242), .B(n14243), .X(n15329) );
  nand_x1_sg U11008 ( .A(\in[0][1][3] ), .B(n16736), .X(n14242) );
  nand_x1_sg U11009 ( .A(n14244), .B(n14245), .X(n15330) );
  nand_x1_sg U11010 ( .A(\in[0][1][4] ), .B(n16737), .X(n14244) );
  nand_x1_sg U11011 ( .A(n14116), .B(n14117), .X(n15266) );
  nand_x1_sg U11012 ( .A(\in[0][1][5] ), .B(n16741), .X(n14116) );
  nand_x1_sg U11013 ( .A(n14118), .B(n14119), .X(n15267) );
  nand_x1_sg U11014 ( .A(\in[0][1][6] ), .B(n16741), .X(n14118) );
  nand_x1_sg U11015 ( .A(n14110), .B(n14111), .X(n15263) );
  nand_x1_sg U11016 ( .A(\in[0][1][7] ), .B(n16736), .X(n14110) );
  nand_x1_sg U11017 ( .A(n14112), .B(n14113), .X(n15264) );
  nand_x1_sg U11018 ( .A(\in[0][1][8] ), .B(n16736), .X(n14112) );
  nand_x1_sg U11019 ( .A(n14128), .B(n14129), .X(n15272) );
  nand_x1_sg U11020 ( .A(\in[0][1][9] ), .B(n16736), .X(n14128) );
  nand_x1_sg U11021 ( .A(n14130), .B(n14131), .X(n15273) );
  nand_x1_sg U11022 ( .A(\in[0][1][10] ), .B(n16736), .X(n14130) );
  nand_x1_sg U11023 ( .A(n14122), .B(n14123), .X(n15269) );
  nand_x1_sg U11024 ( .A(\in[0][1][11] ), .B(n16741), .X(n14122) );
  nand_x1_sg U11025 ( .A(n14124), .B(n14125), .X(n15270) );
  nand_x1_sg U11026 ( .A(\in[0][1][12] ), .B(n16737), .X(n14124) );
  nand_x1_sg U11027 ( .A(n14092), .B(n14093), .X(n15254) );
  nand_x1_sg U11028 ( .A(\in[0][1][13] ), .B(n16736), .X(n14092) );
  nand_x1_sg U11029 ( .A(n14094), .B(n14095), .X(n15255) );
  nand_x1_sg U11030 ( .A(\in[0][1][14] ), .B(n16738), .X(n14094) );
  nand_x1_sg U11031 ( .A(n14086), .B(n14087), .X(n15251) );
  nand_x1_sg U11032 ( .A(\in[0][1][15] ), .B(n16739), .X(n14086) );
  nand_x1_sg U11033 ( .A(n14088), .B(n14089), .X(n15252) );
  nand_x1_sg U11034 ( .A(\in[0][1][16] ), .B(n16736), .X(n14088) );
  nand_x1_sg U11035 ( .A(n14104), .B(n14105), .X(n15260) );
  nand_x1_sg U11036 ( .A(\in[0][1][17] ), .B(n16736), .X(n14104) );
  nand_x1_sg U11037 ( .A(n14106), .B(n14107), .X(n15261) );
  nand_x1_sg U11038 ( .A(\in[0][1][18] ), .B(n16736), .X(n14106) );
  nand_x1_sg U11039 ( .A(n14098), .B(n14099), .X(n15257) );
  nand_x1_sg U11040 ( .A(\in[0][1][19] ), .B(n16736), .X(n14098) );
  nand_x1_sg U11041 ( .A(n14100), .B(n14101), .X(n15258) );
  nand_x1_sg U11042 ( .A(\in[0][2][0] ), .B(n16736), .X(n14100) );
  nand_x1_sg U11043 ( .A(n14164), .B(n14165), .X(n15290) );
  nand_x1_sg U11044 ( .A(\in[0][2][1] ), .B(n16738), .X(n14164) );
  nand_x1_sg U11045 ( .A(n14166), .B(n14167), .X(n15291) );
  nand_x1_sg U11046 ( .A(\in[0][2][2] ), .B(n16736), .X(n14166) );
  nand_x1_sg U11047 ( .A(n14158), .B(n14159), .X(n15287) );
  nand_x1_sg U11048 ( .A(\in[0][2][3] ), .B(n16736), .X(n14158) );
  nand_x1_sg U11049 ( .A(n14160), .B(n14161), .X(n15288) );
  nand_x1_sg U11050 ( .A(\in[0][2][4] ), .B(n16738), .X(n14160) );
  nand_x1_sg U11051 ( .A(n14176), .B(n14177), .X(n15296) );
  nand_x1_sg U11052 ( .A(\in[0][2][5] ), .B(n16738), .X(n14176) );
  nand_x1_sg U11053 ( .A(n14178), .B(n14179), .X(n15297) );
  nand_x1_sg U11054 ( .A(\in[0][2][6] ), .B(n16739), .X(n14178) );
  nand_x1_sg U11055 ( .A(n14170), .B(n14171), .X(n15293) );
  nand_x1_sg U11056 ( .A(\in[0][2][7] ), .B(n16737), .X(n14170) );
  nand_x1_sg U11057 ( .A(n14172), .B(n14173), .X(n15294) );
  nand_x1_sg U11058 ( .A(\in[0][2][8] ), .B(n16736), .X(n14172) );
  nand_x1_sg U11059 ( .A(n14140), .B(n14141), .X(n15278) );
  nand_x1_sg U11060 ( .A(\in[0][2][9] ), .B(n16736), .X(n14140) );
  nand_x1_sg U11061 ( .A(n14142), .B(n14143), .X(n15279) );
  nand_x1_sg U11062 ( .A(\in[0][2][10] ), .B(n16738), .X(n14142) );
  nand_x1_sg U11063 ( .A(n14134), .B(n14135), .X(n15275) );
  nand_x1_sg U11064 ( .A(\in[0][2][11] ), .B(n16743), .X(n14134) );
  nand_x1_sg U11065 ( .A(n14136), .B(n14137), .X(n15276) );
  nand_x1_sg U11066 ( .A(\in[0][2][12] ), .B(n16737), .X(n14136) );
  nand_x1_sg U11067 ( .A(n14152), .B(n14153), .X(n15284) );
  nand_x1_sg U11068 ( .A(\in[0][2][13] ), .B(n16739), .X(n14152) );
  nand_x1_sg U11069 ( .A(n14154), .B(n14155), .X(n15285) );
  nand_x1_sg U11070 ( .A(\in[0][2][14] ), .B(n16737), .X(n14154) );
  nand_x1_sg U11071 ( .A(n14146), .B(n14147), .X(n15281) );
  nand_x1_sg U11072 ( .A(\in[0][2][15] ), .B(n16736), .X(n14146) );
  nand_x1_sg U11073 ( .A(n14148), .B(n14149), .X(n15282) );
  nand_x1_sg U11074 ( .A(\in[0][2][16] ), .B(n16738), .X(n14148) );
  nand_x1_sg U11075 ( .A(n13898), .B(n13899), .X(n15157) );
  nand_x1_sg U11076 ( .A(\in[0][2][17] ), .B(n16739), .X(n13898) );
  nand_x1_sg U11077 ( .A(n14278), .B(n14279), .X(n15347) );
  nand_x1_sg U11078 ( .A(\in[0][2][18] ), .B(n16738), .X(n14278) );
  nand_x1_sg U11079 ( .A(n14392), .B(n14393), .X(n15404) );
  nand_x1_sg U11080 ( .A(\in[0][2][19] ), .B(n16736), .X(n14392) );
  nand_x1_sg U11081 ( .A(n14276), .B(n14277), .X(n15346) );
  nand_x1_sg U11082 ( .A(\in[0][3][0] ), .B(n16738), .X(n14276) );
  nand_x1_sg U11083 ( .A(n13864), .B(n13865), .X(n15140) );
  nand_x1_sg U11084 ( .A(\in[0][3][1] ), .B(n16737), .X(n13864) );
  nand_x1_sg U11085 ( .A(n13844), .B(n13845), .X(n15130) );
  nand_x1_sg U11086 ( .A(\in[0][3][2] ), .B(n16737), .X(n13844) );
  nand_x1_sg U11087 ( .A(n14446), .B(n14447), .X(n15431) );
  nand_x1_sg U11088 ( .A(\in[0][3][3] ), .B(n16736), .X(n14446) );
  nand_x1_sg U11089 ( .A(n13892), .B(n13893), .X(n15154) );
  nand_x1_sg U11090 ( .A(\in[0][3][4] ), .B(n16738), .X(n13892) );
  nand_x1_sg U11091 ( .A(n14216), .B(n14217), .X(n15316) );
  nand_x1_sg U11092 ( .A(\in[0][3][5] ), .B(n16737), .X(n14216) );
  nand_x1_sg U11093 ( .A(n14290), .B(n14291), .X(n15353) );
  nand_x1_sg U11094 ( .A(\in[0][3][6] ), .B(n16736), .X(n14290) );
  nand_x1_sg U11095 ( .A(n13976), .B(n13977), .X(n15196) );
  nand_x1_sg U11096 ( .A(\in[0][3][7] ), .B(n16737), .X(n13976) );
  nand_x1_sg U11097 ( .A(n14132), .B(n14133), .X(n15274) );
  nand_x1_sg U11098 ( .A(\in[0][3][8] ), .B(n16737), .X(n14132) );
  nand_x1_sg U11099 ( .A(n14326), .B(n14327), .X(n15371) );
  nand_x1_sg U11100 ( .A(\in[0][3][9] ), .B(n16737), .X(n14326) );
  nand_x1_sg U11101 ( .A(n13836), .B(n13837), .X(n15126) );
  nand_x1_sg U11102 ( .A(\in[0][3][10] ), .B(n16739), .X(n13836) );
  nand_x1_sg U11103 ( .A(n14060), .B(n14061), .X(n15238) );
  nand_x1_sg U11104 ( .A(\in[0][3][11] ), .B(n16736), .X(n14060) );
  nand_x1_sg U11105 ( .A(n13840), .B(n13841), .X(n15128) );
  nand_x1_sg U11106 ( .A(\in[0][3][12] ), .B(n16739), .X(n13840) );
  nand_x1_sg U11107 ( .A(n14054), .B(n14055), .X(n15235) );
  nand_x1_sg U11108 ( .A(\in[0][3][13] ), .B(n16736), .X(n14054) );
  nand_x1_sg U11109 ( .A(n14018), .B(n14019), .X(n15217) );
  nand_x1_sg U11110 ( .A(\in[0][3][14] ), .B(n16737), .X(n14018) );
  nand_x1_sg U11111 ( .A(n13838), .B(n13839), .X(n15127) );
  nand_x1_sg U11112 ( .A(\in[0][3][15] ), .B(n16737), .X(n13838) );
  nand_x1_sg U11113 ( .A(n14138), .B(n14139), .X(n15277) );
  nand_x1_sg U11114 ( .A(\in[0][3][16] ), .B(n16736), .X(n14138) );
  nand_x1_sg U11115 ( .A(n13940), .B(n13941), .X(n15178) );
  nand_x1_sg U11116 ( .A(\in[0][3][17] ), .B(n16737), .X(n13940) );
  nand_x1_sg U11117 ( .A(n13922), .B(n13923), .X(n15169) );
  nand_x1_sg U11118 ( .A(\in[0][3][18] ), .B(n16736), .X(n13922) );
  nand_x1_sg U11119 ( .A(n13970), .B(n13971), .X(n15193) );
  nand_x1_sg U11120 ( .A(\in[0][3][19] ), .B(n16737), .X(n13970) );
  nand_x1_sg U11121 ( .A(n13994), .B(n13995), .X(n15205) );
  nand_x1_sg U11122 ( .A(\in[1][0][0] ), .B(n16737), .X(n13994) );
  nand_x1_sg U11123 ( .A(n14302), .B(n14303), .X(n15359) );
  nand_x1_sg U11124 ( .A(\in[1][0][1] ), .B(n16736), .X(n14302) );
  nand_x1_sg U11125 ( .A(n14320), .B(n14321), .X(n15368) );
  nand_x1_sg U11126 ( .A(\in[1][0][2] ), .B(n16738), .X(n14320) );
  nand_x1_sg U11127 ( .A(n14234), .B(n14235), .X(n15325) );
  nand_x1_sg U11128 ( .A(\in[1][0][3] ), .B(n16739), .X(n14234) );
  nand_x1_sg U11129 ( .A(n14452), .B(n14453), .X(n15434) );
  nand_x1_sg U11130 ( .A(\in[1][0][4] ), .B(n16738), .X(n14452) );
  nand_x1_sg U11131 ( .A(n14332), .B(n14333), .X(n15374) );
  nand_x1_sg U11132 ( .A(\in[1][0][5] ), .B(n16737), .X(n14332) );
  nand_x1_sg U11133 ( .A(n14338), .B(n14339), .X(n15377) );
  nand_x1_sg U11134 ( .A(\in[1][0][6] ), .B(n16739), .X(n14338) );
  nand_x1_sg U11135 ( .A(n14344), .B(n14345), .X(n15380) );
  nand_x1_sg U11136 ( .A(\in[1][0][7] ), .B(n16738), .X(n14344) );
  nand_x1_sg U11137 ( .A(n14362), .B(n14363), .X(n15389) );
  nand_x1_sg U11138 ( .A(\in[1][0][8] ), .B(n16739), .X(n14362) );
  nand_x1_sg U11139 ( .A(n13872), .B(n13873), .X(n15144) );
  nand_x1_sg U11140 ( .A(\in[1][0][9] ), .B(n16739), .X(n13872) );
  nand_x1_sg U11141 ( .A(n13870), .B(n13871), .X(n15143) );
  nand_x1_sg U11142 ( .A(\in[1][0][10] ), .B(n16738), .X(n13870) );
  nand_x1_sg U11143 ( .A(n13850), .B(n13851), .X(n15133) );
  nand_x1_sg U11144 ( .A(\in[1][0][11] ), .B(n16738), .X(n13850) );
  nand_x1_sg U11145 ( .A(n13856), .B(n13857), .X(n15136) );
  nand_x1_sg U11146 ( .A(\in[1][0][12] ), .B(n16738), .X(n13856) );
  nand_x1_sg U11147 ( .A(n14252), .B(n14253), .X(n15334) );
  nand_x1_sg U11148 ( .A(\in[1][0][13] ), .B(n16739), .X(n14252) );
  nand_x1_sg U11149 ( .A(n13958), .B(n13959), .X(n15187) );
  nand_x1_sg U11150 ( .A(\in[1][0][14] ), .B(n16738), .X(n13958) );
  nand_x1_sg U11151 ( .A(n13852), .B(n13853), .X(n15134) );
  nand_x1_sg U11152 ( .A(\in[1][0][15] ), .B(n16736), .X(n13852) );
  nand_x1_sg U11153 ( .A(n14464), .B(n14465), .X(n15440) );
  nand_x1_sg U11154 ( .A(\in[1][0][16] ), .B(n16739), .X(n14464) );
  nand_x1_sg U11155 ( .A(n14198), .B(n14199), .X(n15307) );
  nand_x1_sg U11156 ( .A(\in[1][0][17] ), .B(n16737), .X(n14198) );
  nand_x1_sg U11157 ( .A(n13854), .B(n13855), .X(n15135) );
  nand_x1_sg U11158 ( .A(\in[1][0][18] ), .B(n16737), .X(n13854) );
  nand_x1_sg U11159 ( .A(n13846), .B(n13847), .X(n15131) );
  nand_x1_sg U11160 ( .A(\in[1][0][19] ), .B(n16739), .X(n13846) );
  nand_x1_sg U11161 ( .A(n13874), .B(n13875), .X(n15145) );
  nand_x1_sg U11162 ( .A(\in[1][1][0] ), .B(n16739), .X(n13874) );
  nand_x1_sg U11163 ( .A(n14150), .B(n14151), .X(n15283) );
  nand_x1_sg U11164 ( .A(\in[1][1][1] ), .B(n16738), .X(n14150) );
  nand_x1_sg U11165 ( .A(n14090), .B(n14091), .X(n15253) );
  nand_x1_sg U11166 ( .A(\in[1][1][2] ), .B(n16739), .X(n14090) );
  nand_x1_sg U11167 ( .A(n13848), .B(n13849), .X(n15132) );
  nand_x1_sg U11168 ( .A(\in[1][1][3] ), .B(n16737), .X(n13848) );
  nand_x1_sg U11169 ( .A(n14180), .B(n14181), .X(n15298) );
  nand_x1_sg U11170 ( .A(\in[1][1][4] ), .B(n16738), .X(n14180) );
  nand_x1_sg U11171 ( .A(n14374), .B(n14375), .X(n15395) );
  nand_x1_sg U11172 ( .A(\in[1][1][5] ), .B(n16739), .X(n14374) );
  nand_x1_sg U11173 ( .A(n14380), .B(n14381), .X(n15398) );
  nand_x1_sg U11174 ( .A(\in[1][1][6] ), .B(n16738), .X(n14380) );
  nand_x1_sg U11175 ( .A(n14422), .B(n14423), .X(n15419) );
  nand_x1_sg U11176 ( .A(\in[1][1][7] ), .B(n16738), .X(n14422) );
  nand_x1_sg U11177 ( .A(n14386), .B(n14387), .X(n15401) );
  nand_x1_sg U11178 ( .A(\in[1][1][8] ), .B(n16739), .X(n14386) );
  nand_x1_sg U11179 ( .A(n14416), .B(n14417), .X(n15416) );
  nand_x1_sg U11180 ( .A(\in[1][1][9] ), .B(n16737), .X(n14416) );
  nand_x1_sg U11181 ( .A(n14308), .B(n14309), .X(n15362) );
  nand_x1_sg U11182 ( .A(\in[1][1][10] ), .B(n16736), .X(n14308) );
  nand_x1_sg U11183 ( .A(n14350), .B(n14351), .X(n15383) );
  nand_x1_sg U11184 ( .A(\in[1][1][11] ), .B(n16738), .X(n14350) );
  nand_x1_sg U11185 ( .A(n14356), .B(n14357), .X(n15386) );
  nand_x1_sg U11186 ( .A(\in[1][1][12] ), .B(n16739), .X(n14356) );
  nand_x1_sg U11187 ( .A(n14410), .B(n14411), .X(n15413) );
  nand_x1_sg U11188 ( .A(\in[1][1][13] ), .B(n16737), .X(n14410) );
  nand_x1_sg U11189 ( .A(n14368), .B(n14369), .X(n15392) );
  nand_x1_sg U11190 ( .A(\in[1][1][14] ), .B(n16738), .X(n14368) );
  nand_x1_sg U11191 ( .A(n14024), .B(n14025), .X(n15220) );
  nand_x1_sg U11192 ( .A(\in[1][1][15] ), .B(n16739), .X(n14024) );
  nand_x1_sg U11193 ( .A(n14428), .B(n14429), .X(n15422) );
  nand_x1_sg U11194 ( .A(\in[1][1][16] ), .B(n16738), .X(n14428) );
  nand_x1_sg U11195 ( .A(n13880), .B(n13881), .X(n15148) );
  nand_x1_sg U11196 ( .A(\in[1][1][17] ), .B(n16738), .X(n13880) );
  nand_x1_sg U11197 ( .A(n13858), .B(n13859), .X(n15137) );
  nand_x1_sg U11198 ( .A(\in[1][1][18] ), .B(n16739), .X(n13858) );
  nand_x1_sg U11199 ( .A(n14270), .B(n14271), .X(n15343) );
  nand_x1_sg U11200 ( .A(\in[1][1][19] ), .B(n16738), .X(n14270) );
  nand_x1_sg U11201 ( .A(n13890), .B(n13891), .X(n15153) );
  nand_x1_sg U11202 ( .A(\in[1][2][0] ), .B(n16739), .X(n13890) );
  nand_x1_sg U11203 ( .A(n14186), .B(n14187), .X(n15301) );
  nand_x1_sg U11204 ( .A(\in[1][2][1] ), .B(n16739), .X(n14186) );
  nand_x1_sg U11205 ( .A(n14192), .B(n14193), .X(n15304) );
  nand_x1_sg U11206 ( .A(\in[1][2][2] ), .B(n16738), .X(n14192) );
  nand_x1_sg U11207 ( .A(n14222), .B(n14223), .X(n15319) );
  nand_x1_sg U11208 ( .A(\in[1][2][3] ), .B(n16736), .X(n14222) );
  nand_x1_sg U11209 ( .A(n14228), .B(n14229), .X(n15322) );
  nand_x1_sg U11210 ( .A(\in[1][2][4] ), .B(n16738), .X(n14228) );
  nand_x1_sg U11211 ( .A(n14204), .B(n14205), .X(n15310) );
  nand_x1_sg U11212 ( .A(\in[1][2][5] ), .B(n16738), .X(n14204) );
  nand_x1_sg U11213 ( .A(n14210), .B(n14211), .X(n15313) );
  nand_x1_sg U11214 ( .A(\in[1][2][6] ), .B(n16738), .X(n14210) );
  nand_x1_sg U11215 ( .A(n13828), .B(n13829), .X(n15123) );
  nand_x1_sg U11216 ( .A(\in[1][2][7] ), .B(n16737), .X(n13828) );
  nand_x1_sg U11217 ( .A(n13832), .B(n13833), .X(n15124) );
  nand_x1_sg U11218 ( .A(\in[1][2][8] ), .B(n16739), .X(n13832) );
  nand_x1_sg U11219 ( .A(n14120), .B(n14121), .X(n15268) );
  nand_x1_sg U11220 ( .A(\in[1][2][9] ), .B(n16741), .X(n14120) );
  nand_x1_sg U11221 ( .A(n14126), .B(n14127), .X(n15271) );
  nand_x1_sg U11222 ( .A(\in[1][2][10] ), .B(n16736), .X(n14126) );
  nand_x1_sg U11223 ( .A(n13834), .B(n13835), .X(n15125) );
  nand_x1_sg U11224 ( .A(\in[1][2][11] ), .B(n16737), .X(n13834) );
  nand_x1_sg U11225 ( .A(n14144), .B(n14145), .X(n15280) );
  nand_x1_sg U11226 ( .A(\in[1][2][12] ), .B(n16738), .X(n14144) );
  nand_x1_sg U11227 ( .A(n14096), .B(n14097), .X(n15256) );
  nand_x1_sg U11228 ( .A(\in[1][2][13] ), .B(n16738), .X(n14096) );
  nand_x1_sg U11229 ( .A(n14102), .B(n14103), .X(n15259) );
  nand_x1_sg U11230 ( .A(\in[1][2][14] ), .B(n16736), .X(n14102) );
  nand_x1_sg U11231 ( .A(n14108), .B(n14109), .X(n15262) );
  nand_x1_sg U11232 ( .A(\in[1][2][15] ), .B(n16736), .X(n14108) );
  nand_x1_sg U11233 ( .A(n14114), .B(n14115), .X(n15265) );
  nand_x1_sg U11234 ( .A(\in[1][2][16] ), .B(n16736), .X(n14114) );
  nand_x1_sg U11235 ( .A(n14012), .B(n14013), .X(n15214) );
  nand_x1_sg U11236 ( .A(\in[1][2][17] ), .B(n16739), .X(n14012) );
  nand_x1_sg U11237 ( .A(n13988), .B(n13989), .X(n15202) );
  nand_x1_sg U11238 ( .A(\in[1][2][18] ), .B(n16739), .X(n13988) );
  nand_x1_sg U11239 ( .A(n13860), .B(n13861), .X(n15138) );
  nand_x1_sg U11240 ( .A(\in[1][2][19] ), .B(n16737), .X(n13860) );
  nand_x1_sg U11241 ( .A(n13862), .B(n13863), .X(n15139) );
  nand_x1_sg U11242 ( .A(\in[1][3][0] ), .B(n16736), .X(n13862) );
  nand_x1_sg U11243 ( .A(n14240), .B(n14241), .X(n15328) );
  nand_x1_sg U11244 ( .A(\in[1][3][1] ), .B(n16739), .X(n14240) );
  nand_x1_sg U11245 ( .A(n14246), .B(n14247), .X(n15331) );
  nand_x1_sg U11246 ( .A(\in[1][3][2] ), .B(n16736), .X(n14246) );
  nand_x1_sg U11247 ( .A(n14258), .B(n14259), .X(n15337) );
  nand_x1_sg U11248 ( .A(\in[1][3][3] ), .B(n16739), .X(n14258) );
  nand_x1_sg U11249 ( .A(n14264), .B(n14265), .X(n15340) );
  nand_x1_sg U11250 ( .A(\in[1][3][4] ), .B(n16739), .X(n14264) );
  nand_x1_sg U11251 ( .A(n14156), .B(n14157), .X(n15286) );
  nand_x1_sg U11252 ( .A(\in[1][3][5] ), .B(n16739), .X(n14156) );
  nand_x1_sg U11253 ( .A(n14162), .B(n14163), .X(n15289) );
  nand_x1_sg U11254 ( .A(\in[1][3][6] ), .B(n16737), .X(n14162) );
  nand_x1_sg U11255 ( .A(n14168), .B(n14169), .X(n15292) );
  nand_x1_sg U11256 ( .A(\in[1][3][7] ), .B(n16739), .X(n14168) );
  nand_x1_sg U11257 ( .A(n14174), .B(n14175), .X(n15295) );
  nand_x1_sg U11258 ( .A(\in[1][3][8] ), .B(n16738), .X(n14174) );
  nand_x1_sg U11259 ( .A(n13882), .B(n13883), .X(n15149) );
  nand_x1_sg U11260 ( .A(\in[1][3][9] ), .B(n16739), .X(n13882) );
  nand_x1_sg U11261 ( .A(n13884), .B(n13885), .X(n15150) );
  nand_x1_sg U11262 ( .A(\in[1][3][10] ), .B(n16738), .X(n13884) );
  nand_x1_sg U11263 ( .A(n13876), .B(n13877), .X(n15146) );
  nand_x1_sg U11264 ( .A(\in[1][3][11] ), .B(n16738), .X(n13876) );
  nand_x1_sg U11265 ( .A(n13878), .B(n13879), .X(n15147) );
  nand_x1_sg U11266 ( .A(\in[1][3][12] ), .B(n16739), .X(n13878) );
  nand_x1_sg U11267 ( .A(n13886), .B(n13887), .X(n15151) );
  nand_x1_sg U11268 ( .A(\in[1][3][13] ), .B(n16739), .X(n13886) );
  nand_x1_sg U11269 ( .A(n13842), .B(n13843), .X(n15129) );
  nand_x1_sg U11270 ( .A(\in[1][3][14] ), .B(n16736), .X(n13842) );
  nand_x1_sg U11271 ( .A(n14398), .B(n14399), .X(n15407) );
  nand_x1_sg U11272 ( .A(\in[1][3][15] ), .B(n16738), .X(n14398) );
  nand_x1_sg U11273 ( .A(n14404), .B(n14405), .X(n15410) );
  nand_x1_sg U11274 ( .A(\in[1][3][16] ), .B(n16736), .X(n14404) );
  nand_x1_sg U11275 ( .A(n13888), .B(n13889), .X(n15152) );
  nand_x1_sg U11276 ( .A(\in[1][3][17] ), .B(n16738), .X(n13888) );
  nand_x1_sg U11277 ( .A(n13916), .B(n13917), .X(n15166) );
  nand_x1_sg U11278 ( .A(\in[1][3][18] ), .B(n16737), .X(n13916) );
  nand_x1_sg U11279 ( .A(n13928), .B(n13929), .X(n15172) );
  nand_x1_sg U11280 ( .A(\in[1][3][19] ), .B(n16736), .X(n13928) );
  nand_x1_sg U11281 ( .A(n13934), .B(n13935), .X(n15175) );
  nand_x1_sg U11282 ( .A(\in[2][0][0] ), .B(n16736), .X(n13934) );
  nand_x1_sg U11283 ( .A(n14284), .B(n14285), .X(n15350) );
  nand_x1_sg U11284 ( .A(\in[2][0][1] ), .B(n16738), .X(n14284) );
  nand_x1_sg U11285 ( .A(n14296), .B(n14297), .X(n15356) );
  nand_x1_sg U11286 ( .A(\in[2][0][2] ), .B(n16738), .X(n14296) );
  nand_x1_sg U11287 ( .A(n13904), .B(n13905), .X(n15160) );
  nand_x1_sg U11288 ( .A(\in[2][0][3] ), .B(n16737), .X(n13904) );
  nand_x1_sg U11289 ( .A(n14314), .B(n14315), .X(n15365) );
  nand_x1_sg U11290 ( .A(\in[2][0][4] ), .B(n16739), .X(n14314) );
  nand_x1_sg U11291 ( .A(n14434), .B(n14435), .X(n15425) );
  nand_x1_sg U11292 ( .A(\in[2][0][5] ), .B(n16736), .X(n14434) );
  nand_x1_sg U11293 ( .A(n14440), .B(n14441), .X(n15428) );
  nand_x1_sg U11294 ( .A(\in[2][0][6] ), .B(n16739), .X(n14440) );
  nand_x1_sg U11295 ( .A(n13910), .B(n13911), .X(n15163) );
  nand_x1_sg U11296 ( .A(\in[2][0][7] ), .B(n16737), .X(n13910) );
  nand_x1_sg U11297 ( .A(n14458), .B(n14459), .X(n15437) );
  nand_x1_sg U11298 ( .A(\in[2][0][8] ), .B(n16737), .X(n14458) );
  nand_x1_sg U11299 ( .A(n14042), .B(n14043), .X(n15229) );
  nand_x1_sg U11300 ( .A(\in[2][0][9] ), .B(n16737), .X(n14042) );
  nand_x1_sg U11301 ( .A(n14048), .B(n14049), .X(n15232) );
  nand_x1_sg U11302 ( .A(\in[2][0][10] ), .B(n16738), .X(n14048) );
  nand_x1_sg U11303 ( .A(n14072), .B(n14073), .X(n15244) );
  nand_x1_sg U11304 ( .A(\in[2][0][11] ), .B(n16738), .X(n14072) );
  nand_x1_sg U11305 ( .A(n14078), .B(n14079), .X(n15247) );
  nand_x1_sg U11306 ( .A(\in[2][0][12] ), .B(n16736), .X(n14078) );
  nand_x1_sg U11307 ( .A(n14000), .B(n14001), .X(n15208) );
  nand_x1_sg U11308 ( .A(\in[2][0][13] ), .B(n16737), .X(n14000) );
  nand_x1_sg U11309 ( .A(n14006), .B(n14007), .X(n15211) );
  nand_x1_sg U11310 ( .A(\in[2][0][14] ), .B(n16737), .X(n14006) );
  nand_x1_sg U11311 ( .A(n14030), .B(n14031), .X(n15223) );
  nand_x1_sg U11312 ( .A(\in[2][0][15] ), .B(n16738), .X(n14030) );
  nand_x1_sg U11313 ( .A(n14036), .B(n14037), .X(n15226) );
  nand_x1_sg U11314 ( .A(\in[2][0][16] ), .B(n16738), .X(n14036) );
  nand_x1_sg U11315 ( .A(n13946), .B(n13947), .X(n15181) );
  nand_x1_sg U11316 ( .A(\in[2][0][17] ), .B(n16736), .X(n13946) );
  nand_x1_sg U11317 ( .A(n13952), .B(n13953), .X(n15184) );
  nand_x1_sg U11318 ( .A(\in[2][0][18] ), .B(n16736), .X(n13952) );
  nand_x1_sg U11319 ( .A(n13868), .B(n13869), .X(n15142) );
  nand_x1_sg U11320 ( .A(\in[2][0][19] ), .B(n16738), .X(n13868) );
  nand_x1_sg U11321 ( .A(n13964), .B(n13965), .X(n15190) );
  nand_x1_sg U11322 ( .A(\in[2][1][0] ), .B(n16739), .X(n13964) );
  nand_x1_sg U11323 ( .A(n14066), .B(n14067), .X(n15241) );
  nand_x1_sg U11324 ( .A(\in[2][1][1] ), .B(n16737), .X(n14066) );
  nand_x1_sg U11325 ( .A(n13982), .B(n13983), .X(n15199) );
  nand_x1_sg U11326 ( .A(\in[2][1][2] ), .B(n16736), .X(n13982) );
  nand_x1_sg U11327 ( .A(n13866), .B(n13867), .X(n15141) );
  nand_x1_sg U11328 ( .A(\in[2][1][3] ), .B(n16739), .X(n13866) );
  nand_x1_sg U11329 ( .A(n14084), .B(n14085), .X(n15250) );
  nand_x1_sg U11330 ( .A(\in[2][1][4] ), .B(n16739), .X(n14084) );
  nand_x1_sg U11331 ( .A(n14406), .B(n14407), .X(n15411) );
  nand_x1_sg U11332 ( .A(\in[2][1][5] ), .B(n16738), .X(n14406) );
  nand_x1_sg U11333 ( .A(n14408), .B(n14409), .X(n15412) );
  nand_x1_sg U11334 ( .A(\in[2][1][6] ), .B(n16739), .X(n14408) );
  nand_x1_sg U11335 ( .A(n14400), .B(n14401), .X(n15408) );
  nand_x1_sg U11336 ( .A(\in[2][1][7] ), .B(n16739), .X(n14400) );
  nand_x1_sg U11337 ( .A(n14402), .B(n14403), .X(n15409) );
  nand_x1_sg U11338 ( .A(\in[2][1][8] ), .B(n16739), .X(n14402) );
  nand_x1_sg U11339 ( .A(n14418), .B(n14419), .X(n15417) );
  nand_x1_sg U11340 ( .A(\in[2][1][9] ), .B(n16736), .X(n14418) );
  nand_x1_sg U11341 ( .A(n14420), .B(n14421), .X(n15418) );
  nand_x1_sg U11342 ( .A(\in[2][1][10] ), .B(n16739), .X(n14420) );
  nand_x1_sg U11343 ( .A(n14412), .B(n14413), .X(n15414) );
  nand_x1_sg U11344 ( .A(\in[2][1][11] ), .B(n16737), .X(n14412) );
  nand_x1_sg U11345 ( .A(n14414), .B(n14415), .X(n15415) );
  nand_x1_sg U11346 ( .A(\in[2][1][12] ), .B(n16738), .X(n14414) );
  nand_x1_sg U11347 ( .A(n14382), .B(n14383), .X(n15399) );
  nand_x1_sg U11348 ( .A(\in[2][1][13] ), .B(n16738), .X(n14382) );
  nand_x1_sg U11349 ( .A(n14384), .B(n14385), .X(n15400) );
  nand_x1_sg U11350 ( .A(\in[2][1][14] ), .B(n16736), .X(n14384) );
  nand_x1_sg U11351 ( .A(n14376), .B(n14377), .X(n15396) );
  nand_x1_sg U11352 ( .A(\in[2][1][15] ), .B(n16738), .X(n14376) );
  nand_x1_sg U11353 ( .A(n14378), .B(n14379), .X(n15397) );
  nand_x1_sg U11354 ( .A(\in[2][1][16] ), .B(n16738), .X(n14378) );
  nand_x1_sg U11355 ( .A(n14394), .B(n14395), .X(n15405) );
  nand_x1_sg U11356 ( .A(\in[2][1][17] ), .B(n16737), .X(n14394) );
  nand_x1_sg U11357 ( .A(n14396), .B(n14397), .X(n15406) );
  nand_x1_sg U11358 ( .A(\in[2][1][18] ), .B(n16737), .X(n14396) );
  nand_x1_sg U11359 ( .A(n14388), .B(n14389), .X(n15402) );
  nand_x1_sg U11360 ( .A(\in[2][1][19] ), .B(n16738), .X(n14388) );
  nand_x1_sg U11361 ( .A(n14390), .B(n14391), .X(n15403) );
  nand_x1_sg U11362 ( .A(\in[2][2][0] ), .B(n16738), .X(n14390) );
  nand_x1_sg U11363 ( .A(n14454), .B(n14455), .X(n15435) );
  nand_x1_sg U11364 ( .A(\in[2][2][1] ), .B(n16739), .X(n14454) );
  nand_x1_sg U11365 ( .A(n14456), .B(n14457), .X(n15436) );
  nand_x1_sg U11366 ( .A(\in[2][2][2] ), .B(n16738), .X(n14456) );
  nand_x1_sg U11367 ( .A(n14448), .B(n14449), .X(n15432) );
  nand_x1_sg U11368 ( .A(\in[2][2][3] ), .B(n16736), .X(n14448) );
  nand_x1_sg U11369 ( .A(n14450), .B(n14451), .X(n15433) );
  nand_x1_sg U11370 ( .A(\in[2][2][4] ), .B(n16739), .X(n14450) );
  nand_x1_sg U11371 ( .A(n14466), .B(n14467), .X(n15441) );
  nand_x1_sg U11372 ( .A(\in[2][2][5] ), .B(n16737), .X(n14466) );
  nand_x1_sg U11373 ( .A(n14468), .B(n14469), .X(n15442) );
  nand_x1_sg U11374 ( .A(\in[2][2][6] ), .B(n16737), .X(n14468) );
  nand_x1_sg U11375 ( .A(n14460), .B(n14461), .X(n15438) );
  nand_x1_sg U11376 ( .A(\in[2][2][7] ), .B(n16737), .X(n14460) );
  nand_x1_sg U11377 ( .A(n14462), .B(n14463), .X(n15439) );
  nand_x1_sg U11378 ( .A(\in[2][2][8] ), .B(n16738), .X(n14462) );
  nand_x1_sg U11379 ( .A(n14430), .B(n14431), .X(n15423) );
  nand_x1_sg U11380 ( .A(\in[2][2][9] ), .B(n16738), .X(n14430) );
  nand_x1_sg U11381 ( .A(n14432), .B(n14433), .X(n15424) );
  nand_x1_sg U11382 ( .A(\in[2][2][10] ), .B(n16737), .X(n14432) );
  nand_x1_sg U11383 ( .A(n14424), .B(n14425), .X(n15420) );
  nand_x1_sg U11384 ( .A(\in[2][2][11] ), .B(n16736), .X(n14424) );
  nand_x1_sg U11385 ( .A(n14426), .B(n14427), .X(n15421) );
  nand_x1_sg U11386 ( .A(\in[2][2][12] ), .B(n16737), .X(n14426) );
  nand_x1_sg U11387 ( .A(n14442), .B(n14443), .X(n15429) );
  nand_x1_sg U11388 ( .A(\in[2][2][13] ), .B(n16738), .X(n14442) );
  nand_x1_sg U11389 ( .A(n14444), .B(n14445), .X(n15430) );
  nand_x1_sg U11390 ( .A(\in[2][2][14] ), .B(n16737), .X(n14444) );
  nand_x1_sg U11391 ( .A(n14436), .B(n14437), .X(n15426) );
  nand_x1_sg U11392 ( .A(\in[2][2][15] ), .B(n16736), .X(n14436) );
  nand_x1_sg U11393 ( .A(n14438), .B(n14439), .X(n15427) );
  nand_x1_sg U11394 ( .A(\in[2][2][16] ), .B(n16738), .X(n14438) );
  nand_x1_sg U11395 ( .A(n14310), .B(n14311), .X(n15363) );
  nand_x1_sg U11396 ( .A(\in[2][2][17] ), .B(n16736), .X(n14310) );
  nand_x1_sg U11397 ( .A(n14312), .B(n14313), .X(n15364) );
  nand_x1_sg U11398 ( .A(\in[2][2][18] ), .B(n16739), .X(n14312) );
  nand_x1_sg U11399 ( .A(n14304), .B(n14305), .X(n15360) );
  nand_x1_sg U11400 ( .A(\in[2][2][19] ), .B(n16739), .X(n14304) );
  nand_x1_sg U11401 ( .A(n14306), .B(n14307), .X(n15361) );
  nand_x1_sg U11402 ( .A(\in[2][3][0] ), .B(n16737), .X(n14306) );
  nand_x1_sg U11403 ( .A(n14322), .B(n14323), .X(n15369) );
  nand_x1_sg U11404 ( .A(\in[2][3][1] ), .B(n16736), .X(n14322) );
  nand_x1_sg U11405 ( .A(n14324), .B(n14325), .X(n15370) );
  nand_x1_sg U11406 ( .A(\in[2][3][2] ), .B(n16737), .X(n14324) );
  nand_x1_sg U11407 ( .A(n14316), .B(n14317), .X(n15366) );
  nand_x1_sg U11408 ( .A(\in[2][3][3] ), .B(n16738), .X(n14316) );
  nand_x1_sg U11409 ( .A(n14318), .B(n14319), .X(n15367) );
  nand_x1_sg U11410 ( .A(\in[2][3][4] ), .B(n16739), .X(n14318) );
  nand_x1_sg U11411 ( .A(n14286), .B(n14287), .X(n15351) );
  nand_x1_sg U11412 ( .A(\in[2][3][5] ), .B(n16738), .X(n14286) );
  nand_x1_sg U11413 ( .A(n14288), .B(n14289), .X(n15352) );
  nand_x1_sg U11414 ( .A(\in[2][3][6] ), .B(n16737), .X(n14288) );
  nand_x1_sg U11415 ( .A(n14280), .B(n14281), .X(n15348) );
  nand_x1_sg U11416 ( .A(\in[2][3][7] ), .B(n16738), .X(n14280) );
  nand_x1_sg U11417 ( .A(n14282), .B(n14283), .X(n15349) );
  nand_x1_sg U11418 ( .A(\in[2][3][8] ), .B(n16738), .X(n14282) );
  nand_x1_sg U11419 ( .A(n14298), .B(n14299), .X(n15357) );
  nand_x1_sg U11420 ( .A(\in[2][3][9] ), .B(n16738), .X(n14298) );
  nand_x1_sg U11421 ( .A(n14300), .B(n14301), .X(n15358) );
  nand_x1_sg U11422 ( .A(\in[2][3][10] ), .B(n16736), .X(n14300) );
  nand_x1_sg U11423 ( .A(n14292), .B(n14293), .X(n15354) );
  nand_x1_sg U11424 ( .A(\in[2][3][11] ), .B(n16736), .X(n14292) );
  nand_x1_sg U11425 ( .A(n14294), .B(n14295), .X(n15355) );
  nand_x1_sg U11426 ( .A(\in[2][3][12] ), .B(n16737), .X(n14294) );
  nand_x1_sg U11427 ( .A(n14358), .B(n14359), .X(n15387) );
  nand_x1_sg U11428 ( .A(\in[2][3][13] ), .B(n16738), .X(n14358) );
  nand_x1_sg U11429 ( .A(n14360), .B(n14361), .X(n15388) );
  nand_x1_sg U11430 ( .A(\in[2][3][14] ), .B(n16736), .X(n14360) );
  nand_x1_sg U11431 ( .A(n14352), .B(n14353), .X(n15384) );
  nand_x1_sg U11432 ( .A(\in[2][3][15] ), .B(n16737), .X(n14352) );
  nand_x1_sg U11433 ( .A(n14354), .B(n14355), .X(n15385) );
  nand_x1_sg U11434 ( .A(\in[2][3][16] ), .B(n16736), .X(n14354) );
  nand_x1_sg U11435 ( .A(n14370), .B(n14371), .X(n15393) );
  nand_x1_sg U11436 ( .A(\in[2][3][17] ), .B(n16737), .X(n14370) );
  nand_x1_sg U11437 ( .A(n14372), .B(n14373), .X(n15394) );
  nand_x1_sg U11438 ( .A(\in[2][3][18] ), .B(n16739), .X(n14372) );
  nand_x1_sg U11439 ( .A(n14364), .B(n14365), .X(n15390) );
  nand_x1_sg U11440 ( .A(\in[2][3][19] ), .B(n16739), .X(n14364) );
  nand_x1_sg U11441 ( .A(n14366), .B(n14367), .X(n15391) );
  nand_x1_sg U11442 ( .A(\in[3][0][0] ), .B(n16736), .X(n14366) );
  nand_x1_sg U11443 ( .A(n14334), .B(n14335), .X(n15375) );
  nand_x1_sg U11444 ( .A(\in[3][0][1] ), .B(n16739), .X(n14334) );
  nand_x1_sg U11445 ( .A(n14336), .B(n14337), .X(n15376) );
  nand_x1_sg U11446 ( .A(\in[3][0][2] ), .B(n16739), .X(n14336) );
  nand_x1_sg U11447 ( .A(n14328), .B(n14329), .X(n15372) );
  nand_x1_sg U11448 ( .A(\in[3][0][3] ), .B(n16736), .X(n14328) );
  nand_x1_sg U11449 ( .A(n14330), .B(n14331), .X(n15373) );
  nand_x1_sg U11450 ( .A(\in[3][0][4] ), .B(n16736), .X(n14330) );
  nand_x1_sg U11451 ( .A(n14346), .B(n14347), .X(n15381) );
  nand_x1_sg U11452 ( .A(\in[3][0][5] ), .B(n16739), .X(n14346) );
  nand_x1_sg U11453 ( .A(n14348), .B(n14349), .X(n15382) );
  nand_x1_sg U11454 ( .A(\in[3][0][6] ), .B(n16738), .X(n14348) );
  nand_x1_sg U11455 ( .A(n14340), .B(n14341), .X(n15378) );
  nand_x1_sg U11456 ( .A(\in[3][0][7] ), .B(n16737), .X(n14340) );
  nand_x1_sg U11457 ( .A(n14342), .B(n14343), .X(n15379) );
  nand_x1_sg U11458 ( .A(\in[3][0][8] ), .B(n16741), .X(n14342) );
  nand_x1_sg U11459 ( .A(n14020), .B(n14021), .X(n15218) );
  nand_x1_sg U11460 ( .A(\in[3][0][9] ), .B(n16736), .X(n14020) );
  nand_x1_sg U11461 ( .A(n14022), .B(n14023), .X(n15219) );
  nand_x1_sg U11462 ( .A(\in[3][0][10] ), .B(n16737), .X(n14022) );
  nand_x1_sg U11463 ( .A(n14014), .B(n14015), .X(n15215) );
  nand_x1_sg U11464 ( .A(\in[3][0][11] ), .B(n16736), .X(n14014) );
  nand_x1_sg U11465 ( .A(n14016), .B(n14017), .X(n15216) );
  nand_x1_sg U11466 ( .A(\in[3][0][12] ), .B(n16738), .X(n14016) );
  nand_x1_sg U11467 ( .A(n14032), .B(n14033), .X(n15224) );
  nand_x1_sg U11468 ( .A(\in[3][0][13] ), .B(n16739), .X(n14032) );
  nand_x1_sg U11469 ( .A(n14034), .B(n14035), .X(n15225) );
  nand_x1_sg U11470 ( .A(\in[3][0][14] ), .B(n16738), .X(n14034) );
  nand_x1_sg U11471 ( .A(n14026), .B(n14027), .X(n15221) );
  nand_x1_sg U11472 ( .A(\in[3][0][15] ), .B(n16736), .X(n14026) );
  nand_x1_sg U11473 ( .A(n14028), .B(n14029), .X(n15222) );
  nand_x1_sg U11474 ( .A(\in[3][0][16] ), .B(n16736), .X(n14028) );
  nand_x1_sg U11475 ( .A(n13996), .B(n13997), .X(n15206) );
  nand_x1_sg U11476 ( .A(\in[3][0][17] ), .B(n16737), .X(n13996) );
  nand_x1_sg U11477 ( .A(n13998), .B(n13999), .X(n15207) );
  nand_x1_sg U11478 ( .A(\in[3][0][18] ), .B(n16737), .X(n13998) );
  nand_x1_sg U11479 ( .A(n13990), .B(n13991), .X(n15203) );
  nand_x1_sg U11480 ( .A(\in[3][0][19] ), .B(n16737), .X(n13990) );
  nand_x1_sg U11481 ( .A(n13992), .B(n13993), .X(n15204) );
  nand_x1_sg U11482 ( .A(\in[3][1][0] ), .B(n16737), .X(n13992) );
  nand_x1_sg U11483 ( .A(n14008), .B(n14009), .X(n15212) );
  nand_x1_sg U11484 ( .A(\in[3][1][1] ), .B(n16736), .X(n14008) );
  nand_x1_sg U11485 ( .A(n14010), .B(n14011), .X(n15213) );
  nand_x1_sg U11486 ( .A(\in[3][1][2] ), .B(n16739), .X(n14010) );
  nand_x1_sg U11487 ( .A(n14002), .B(n14003), .X(n15209) );
  nand_x1_sg U11488 ( .A(\in[3][1][3] ), .B(n16737), .X(n14002) );
  nand_x1_sg U11489 ( .A(n14004), .B(n14005), .X(n15210) );
  nand_x1_sg U11490 ( .A(\in[3][1][4] ), .B(n16737), .X(n14004) );
  nand_x1_sg U11491 ( .A(n14068), .B(n14069), .X(n15242) );
  nand_x1_sg U11492 ( .A(\in[3][1][5] ), .B(n16738), .X(n14068) );
  nand_x1_sg U11493 ( .A(n14070), .B(n14071), .X(n15243) );
  nand_x1_sg U11494 ( .A(\in[3][1][6] ), .B(n16736), .X(n14070) );
  nand_x1_sg U11495 ( .A(n14062), .B(n14063), .X(n15239) );
  nand_x1_sg U11496 ( .A(\in[3][1][7] ), .B(n16739), .X(n14062) );
  nand_x1_sg U11497 ( .A(n14064), .B(n14065), .X(n15240) );
  nand_x1_sg U11498 ( .A(\in[3][1][8] ), .B(n16736), .X(n14064) );
  nand_x1_sg U11499 ( .A(n14080), .B(n14081), .X(n15248) );
  nand_x1_sg U11500 ( .A(\in[3][1][9] ), .B(n16736), .X(n14080) );
  nand_x1_sg U11501 ( .A(n14082), .B(n14083), .X(n15249) );
  nand_x1_sg U11502 ( .A(\in[3][1][10] ), .B(n16738), .X(n14082) );
  nand_x1_sg U11503 ( .A(n14074), .B(n14075), .X(n15245) );
  nand_x1_sg U11504 ( .A(\in[3][1][11] ), .B(n16737), .X(n14074) );
  nand_x1_sg U11505 ( .A(n14076), .B(n14077), .X(n15246) );
  nand_x1_sg U11506 ( .A(\in[3][1][12] ), .B(n16739), .X(n14076) );
  nand_x1_sg U11507 ( .A(n14044), .B(n14045), .X(n15230) );
  nand_x1_sg U11508 ( .A(\in[3][1][13] ), .B(n16737), .X(n14044) );
  nand_x1_sg U11509 ( .A(n14046), .B(n14047), .X(n15231) );
  nand_x1_sg U11510 ( .A(\in[3][1][14] ), .B(n16739), .X(n14046) );
  nand_x1_sg U11511 ( .A(n14038), .B(n14039), .X(n15227) );
  nand_x1_sg U11512 ( .A(\in[3][1][15] ), .B(n16736), .X(n14038) );
  nand_x1_sg U11513 ( .A(n14040), .B(n14041), .X(n15228) );
  nand_x1_sg U11514 ( .A(\in[3][1][16] ), .B(n16738), .X(n14040) );
  nand_x1_sg U11515 ( .A(n14056), .B(n14057), .X(n15236) );
  nand_x1_sg U11516 ( .A(\in[3][1][17] ), .B(n16738), .X(n14056) );
  nand_x1_sg U11517 ( .A(n14058), .B(n14059), .X(n15237) );
  nand_x1_sg U11518 ( .A(\in[3][1][18] ), .B(n16739), .X(n14058) );
  nand_x1_sg U11519 ( .A(n14050), .B(n14051), .X(n15233) );
  nand_x1_sg U11520 ( .A(\in[3][1][19] ), .B(n16736), .X(n14050) );
  nand_x1_sg U11521 ( .A(n14052), .B(n14053), .X(n15234) );
  nand_x1_sg U11522 ( .A(\in[3][2][0] ), .B(n16739), .X(n14052) );
  nand_x1_sg U11523 ( .A(n13924), .B(n13925), .X(n15170) );
  nand_x1_sg U11524 ( .A(\in[3][2][1] ), .B(n16736), .X(n13924) );
  nand_x1_sg U11525 ( .A(n13926), .B(n13927), .X(n15171) );
  nand_x1_sg U11526 ( .A(\in[3][2][2] ), .B(n16736), .X(n13926) );
  nand_x1_sg U11527 ( .A(n13918), .B(n13919), .X(n15167) );
  nand_x1_sg U11528 ( .A(\in[3][2][3] ), .B(n16737), .X(n13918) );
  nand_x1_sg U11529 ( .A(n13920), .B(n13921), .X(n15168) );
  nand_x1_sg U11530 ( .A(\in[3][2][4] ), .B(n16736), .X(n13920) );
  nand_x1_sg U11531 ( .A(n13936), .B(n13937), .X(n15176) );
  nand_x1_sg U11532 ( .A(\in[3][2][5] ), .B(n16736), .X(n13936) );
  nand_x1_sg U11533 ( .A(n13938), .B(n13939), .X(n15177) );
  nand_x1_sg U11534 ( .A(\in[3][2][6] ), .B(n16737), .X(n13938) );
  nand_x1_sg U11535 ( .A(n13930), .B(n13931), .X(n15173) );
  nand_x1_sg U11536 ( .A(\in[3][2][7] ), .B(n16736), .X(n13930) );
  nand_x1_sg U11537 ( .A(n13932), .B(n13933), .X(n15174) );
  nand_x1_sg U11538 ( .A(\in[3][2][8] ), .B(n16736), .X(n13932) );
  nand_x1_sg U11539 ( .A(n13900), .B(n13901), .X(n15158) );
  nand_x1_sg U11540 ( .A(\in[3][2][9] ), .B(n16738), .X(n13900) );
  nand_x1_sg U11541 ( .A(n13902), .B(n13903), .X(n15159) );
  nand_x1_sg U11542 ( .A(\in[3][2][10] ), .B(n16737), .X(n13902) );
  nand_x1_sg U11543 ( .A(n13894), .B(n13895), .X(n15155) );
  nand_x1_sg U11544 ( .A(\in[3][2][11] ), .B(n16738), .X(n13894) );
  nand_x1_sg U11545 ( .A(n13896), .B(n13897), .X(n15156) );
  nand_x1_sg U11546 ( .A(\in[3][2][12] ), .B(n16739), .X(n13896) );
  nand_x1_sg U11547 ( .A(n13912), .B(n13913), .X(n15164) );
  nand_x1_sg U11548 ( .A(\in[3][2][13] ), .B(n16737), .X(n13912) );
  nand_x1_sg U11549 ( .A(n13914), .B(n13915), .X(n15165) );
  nand_x1_sg U11550 ( .A(\in[3][2][14] ), .B(n16737), .X(n13914) );
  nand_x1_sg U11551 ( .A(n13906), .B(n13907), .X(n15161) );
  nand_x1_sg U11552 ( .A(\in[3][2][15] ), .B(n16737), .X(n13906) );
  nand_x1_sg U11553 ( .A(n13908), .B(n13909), .X(n15162) );
  nand_x1_sg U11554 ( .A(\in[3][2][16] ), .B(n16737), .X(n13908) );
  nand_x1_sg U11555 ( .A(n13972), .B(n13973), .X(n15194) );
  nand_x1_sg U11556 ( .A(\in[3][2][17] ), .B(n16739), .X(n13972) );
  nand_x1_sg U11557 ( .A(n13974), .B(n13975), .X(n15195) );
  nand_x1_sg U11558 ( .A(\in[3][2][18] ), .B(n16737), .X(n13974) );
  nand_x1_sg U11559 ( .A(n13966), .B(n13967), .X(n15191) );
  nand_x1_sg U11560 ( .A(\in[3][2][19] ), .B(n16736), .X(n13966) );
  nand_x1_sg U11561 ( .A(n13968), .B(n13969), .X(n15192) );
  nand_x1_sg U11562 ( .A(\in[3][3][0] ), .B(n16736), .X(n13968) );
  nand_x1_sg U11563 ( .A(n13984), .B(n13985), .X(n15200) );
  nand_x1_sg U11564 ( .A(\in[3][3][1] ), .B(n16739), .X(n13984) );
  nand_x1_sg U11565 ( .A(n13986), .B(n13987), .X(n15201) );
  nand_x1_sg U11566 ( .A(\in[3][3][2] ), .B(n16738), .X(n13986) );
  nand_x1_sg U11567 ( .A(n13978), .B(n13979), .X(n15197) );
  nand_x1_sg U11568 ( .A(\in[3][3][3] ), .B(n16738), .X(n13978) );
  nand_x1_sg U11569 ( .A(n13980), .B(n13981), .X(n15198) );
  nand_x1_sg U11570 ( .A(\in[3][3][4] ), .B(n16736), .X(n13980) );
  nand_x1_sg U11571 ( .A(n13948), .B(n13949), .X(n15182) );
  nand_x1_sg U11572 ( .A(\in[3][3][5] ), .B(n16739), .X(n13948) );
  nand_x1_sg U11573 ( .A(n13950), .B(n13951), .X(n15183) );
  nand_x1_sg U11574 ( .A(\in[3][3][6] ), .B(n16737), .X(n13950) );
  nand_x1_sg U11575 ( .A(n13942), .B(n13943), .X(n15179) );
  nand_x1_sg U11576 ( .A(\in[3][3][7] ), .B(n16737), .X(n13942) );
  nand_x1_sg U11577 ( .A(n13944), .B(n13945), .X(n15180) );
  nand_x1_sg U11578 ( .A(\in[3][3][8] ), .B(n16737), .X(n13944) );
  nand_x1_sg U11579 ( .A(n13960), .B(n13961), .X(n15188) );
  nand_x1_sg U11580 ( .A(\in[3][3][9] ), .B(n16739), .X(n13960) );
  nand_x1_sg U11581 ( .A(n13962), .B(n13963), .X(n15189) );
  nand_x1_sg U11582 ( .A(\in[3][3][10] ), .B(n16737), .X(n13962) );
  nand_x1_sg U11583 ( .A(n13954), .B(n13955), .X(n15185) );
  nand_x1_sg U11584 ( .A(\in[3][3][11] ), .B(n16737), .X(n13954) );
  nand_x1_sg U11585 ( .A(n13956), .B(n13957), .X(n15186) );
  nand_x1_sg U11586 ( .A(\in[3][3][12] ), .B(n16737), .X(n13956) );
  nand_x1_sg U11587 ( .A(n14212), .B(n14213), .X(n15314) );
  nand_x1_sg U11588 ( .A(\in[3][3][13] ), .B(n16737), .X(n14212) );
  nand_x1_sg U11589 ( .A(n14214), .B(n14215), .X(n15315) );
  nand_x1_sg U11590 ( .A(\in[3][3][14] ), .B(n16739), .X(n14214) );
  nand_x1_sg U11591 ( .A(n14206), .B(n14207), .X(n15311) );
  nand_x1_sg U11592 ( .A(\in[3][3][15] ), .B(n16739), .X(n14206) );
  nand_x1_sg U11593 ( .A(n14208), .B(n14209), .X(n15312) );
  nand_x1_sg U11594 ( .A(\in[3][3][16] ), .B(n16739), .X(n14208) );
  nand_x1_sg U11595 ( .A(n14224), .B(n14225), .X(n15320) );
  nand_x1_sg U11596 ( .A(\in[3][3][17] ), .B(n16739), .X(n14224) );
  nand_x1_sg U11597 ( .A(n14226), .B(n14227), .X(n15321) );
  nand_x1_sg U11598 ( .A(\in[3][3][18] ), .B(n16737), .X(n14226) );
  nand_x1_sg U11599 ( .A(n14218), .B(n14219), .X(n15317) );
  nand_x1_sg U11600 ( .A(\in[3][3][19] ), .B(n16736), .X(n14218) );
  nand_x1_sg U11601 ( .A(n16770), .B(n14473), .X(n15443) );
  nand_x1_sg U11602 ( .A(n14476), .B(n14477), .X(n15444) );
  inv_x4_sg U11603 ( .A(n15446), .X(n15449) );
  inv_x8_sg U11604 ( .A(n15449), .X(state[1]) );
  inv_x2_sg U11605 ( .A(\reg_in[3][3][19] ), .X(n16091) );
  inv_x2_sg U11606 ( .A(\reg_in[3][3][18] ), .X(n16093) );
  inv_x2_sg U11607 ( .A(\reg_in[3][3][17] ), .X(n16095) );
  inv_x2_sg U11608 ( .A(\reg_in[3][3][16] ), .X(n16097) );
  inv_x2_sg U11609 ( .A(\reg_in[3][3][15] ), .X(n16099) );
  inv_x2_sg U11610 ( .A(\reg_in[3][3][14] ), .X(n16101) );
  inv_x2_sg U11611 ( .A(\reg_in[3][3][13] ), .X(n16103) );
  inv_x2_sg U11612 ( .A(\reg_in[3][3][12] ), .X(n16105) );
  inv_x2_sg U11613 ( .A(\reg_in[3][3][11] ), .X(n16107) );
  inv_x2_sg U11614 ( .A(\reg_in[3][3][10] ), .X(n16109) );
  inv_x2_sg U11615 ( .A(\reg_in[3][3][9] ), .X(n16111) );
  inv_x2_sg U11616 ( .A(\reg_in[3][3][8] ), .X(n16113) );
  inv_x2_sg U11617 ( .A(\reg_in[3][3][7] ), .X(n16115) );
  inv_x2_sg U11618 ( .A(\reg_in[3][3][6] ), .X(n16117) );
  inv_x2_sg U11619 ( .A(\reg_in[3][3][5] ), .X(n16119) );
  inv_x2_sg U11620 ( .A(\reg_in[3][3][4] ), .X(n16121) );
  inv_x2_sg U11621 ( .A(\reg_in[3][3][3] ), .X(n16123) );
  inv_x2_sg U11622 ( .A(\reg_in[3][3][2] ), .X(n16125) );
  inv_x2_sg U11623 ( .A(\reg_in[3][3][1] ), .X(n16127) );
  inv_x2_sg U11624 ( .A(\reg_in[3][3][0] ), .X(n16129) );
  inv_x2_sg U11625 ( .A(\reg_in[3][2][19] ), .X(n16131) );
  inv_x2_sg U11626 ( .A(\reg_in[3][2][18] ), .X(n16133) );
  inv_x2_sg U11627 ( .A(\reg_in[3][2][17] ), .X(n16135) );
  inv_x2_sg U11628 ( .A(\reg_in[3][2][16] ), .X(n16137) );
  inv_x2_sg U11629 ( .A(\reg_in[3][2][15] ), .X(n16139) );
  inv_x2_sg U11630 ( .A(\reg_in[3][2][14] ), .X(n16141) );
  inv_x2_sg U11631 ( .A(\reg_in[3][2][13] ), .X(n16143) );
  inv_x2_sg U11632 ( .A(\reg_in[3][2][12] ), .X(n16145) );
  inv_x2_sg U11633 ( .A(\reg_in[3][2][11] ), .X(n16147) );
  inv_x2_sg U11634 ( .A(\reg_in[3][2][10] ), .X(n16149) );
  inv_x2_sg U11635 ( .A(\reg_in[3][2][9] ), .X(n16151) );
  inv_x2_sg U11636 ( .A(\reg_in[3][2][8] ), .X(n16153) );
  inv_x2_sg U11637 ( .A(\reg_in[3][2][7] ), .X(n16155) );
  inv_x2_sg U11638 ( .A(\reg_in[3][2][6] ), .X(n16157) );
  inv_x2_sg U11639 ( .A(\reg_in[3][2][5] ), .X(n16159) );
  inv_x2_sg U11640 ( .A(\reg_in[3][2][4] ), .X(n16161) );
  inv_x2_sg U11641 ( .A(\reg_in[3][2][3] ), .X(n16163) );
  inv_x2_sg U11642 ( .A(\reg_in[3][2][2] ), .X(n16165) );
  inv_x2_sg U11643 ( .A(\reg_in[3][2][1] ), .X(n16167) );
  inv_x2_sg U11644 ( .A(\reg_in[3][2][0] ), .X(n16169) );
  inv_x2_sg U11645 ( .A(\reg_in[3][1][19] ), .X(n16171) );
  inv_x2_sg U11646 ( .A(\reg_in[3][1][18] ), .X(n16173) );
  inv_x2_sg U11647 ( .A(\reg_in[3][1][17] ), .X(n16175) );
  inv_x2_sg U11648 ( .A(\reg_in[3][1][16] ), .X(n16177) );
  inv_x2_sg U11649 ( .A(\reg_in[3][1][15] ), .X(n16179) );
  inv_x2_sg U11650 ( .A(\reg_in[3][1][14] ), .X(n16181) );
  inv_x2_sg U11651 ( .A(\reg_in[3][1][13] ), .X(n16183) );
  inv_x2_sg U11652 ( .A(\reg_in[3][1][12] ), .X(n16185) );
  inv_x2_sg U11653 ( .A(\reg_in[3][1][11] ), .X(n16187) );
  inv_x2_sg U11654 ( .A(\reg_in[3][1][10] ), .X(n16189) );
  inv_x2_sg U11655 ( .A(\reg_in[3][1][9] ), .X(n16191) );
  inv_x2_sg U11656 ( .A(\reg_in[3][1][8] ), .X(n16193) );
  inv_x2_sg U11657 ( .A(\reg_in[3][1][7] ), .X(n16195) );
  inv_x2_sg U11658 ( .A(\reg_in[3][1][6] ), .X(n16197) );
  inv_x2_sg U11659 ( .A(\reg_in[3][1][5] ), .X(n16199) );
  inv_x2_sg U11660 ( .A(\reg_in[3][1][4] ), .X(n16201) );
  inv_x2_sg U11661 ( .A(\reg_in[3][1][3] ), .X(n16203) );
  inv_x2_sg U11662 ( .A(\reg_in[3][1][2] ), .X(n16205) );
  inv_x2_sg U11663 ( .A(\reg_in[3][1][1] ), .X(n16207) );
  inv_x2_sg U11664 ( .A(\reg_in[3][1][0] ), .X(n16209) );
  inv_x2_sg U11665 ( .A(\reg_in[3][0][19] ), .X(n16211) );
  inv_x2_sg U11666 ( .A(\reg_in[3][0][18] ), .X(n16213) );
  inv_x2_sg U11667 ( .A(\reg_in[3][0][17] ), .X(n16215) );
  inv_x2_sg U11668 ( .A(\reg_in[3][0][16] ), .X(n16217) );
  inv_x2_sg U11669 ( .A(\reg_in[3][0][15] ), .X(n16219) );
  inv_x2_sg U11670 ( .A(\reg_in[3][0][14] ), .X(n16221) );
  inv_x2_sg U11671 ( .A(\reg_in[3][0][13] ), .X(n16223) );
  inv_x2_sg U11672 ( .A(\reg_in[3][0][12] ), .X(n16225) );
  inv_x2_sg U11673 ( .A(\reg_in[3][0][11] ), .X(n16227) );
  inv_x2_sg U11674 ( .A(\reg_in[3][0][10] ), .X(n16229) );
  inv_x2_sg U11675 ( .A(\reg_in[3][0][9] ), .X(n16231) );
  inv_x2_sg U11676 ( .A(\reg_in[3][0][8] ), .X(n16233) );
  inv_x2_sg U11677 ( .A(\reg_in[3][0][7] ), .X(n16235) );
  inv_x2_sg U11678 ( .A(\reg_in[3][0][6] ), .X(n16237) );
  inv_x2_sg U11679 ( .A(\reg_in[3][0][5] ), .X(n16239) );
  inv_x2_sg U11680 ( .A(\reg_in[3][0][4] ), .X(n16241) );
  inv_x2_sg U11681 ( .A(\reg_in[3][0][3] ), .X(n16243) );
  inv_x2_sg U11682 ( .A(\reg_in[3][0][2] ), .X(n16245) );
  inv_x2_sg U11683 ( .A(\reg_in[3][0][1] ), .X(n16247) );
  inv_x2_sg U11684 ( .A(\reg_in[3][0][0] ), .X(n16249) );
  inv_x2_sg U11685 ( .A(\reg_in[2][3][19] ), .X(n16251) );
  inv_x2_sg U11686 ( .A(\reg_in[2][3][18] ), .X(n16253) );
  inv_x2_sg U11687 ( .A(\reg_in[2][3][17] ), .X(n16255) );
  inv_x2_sg U11688 ( .A(\reg_in[2][3][16] ), .X(n16257) );
  inv_x2_sg U11689 ( .A(\reg_in[2][3][15] ), .X(n16259) );
  inv_x2_sg U11690 ( .A(\reg_in[2][3][14] ), .X(n16261) );
  inv_x2_sg U11691 ( .A(\reg_in[2][3][13] ), .X(n16263) );
  inv_x2_sg U11692 ( .A(\reg_in[2][3][12] ), .X(n16265) );
  inv_x2_sg U11693 ( .A(\reg_in[2][3][11] ), .X(n16267) );
  inv_x2_sg U11694 ( .A(\reg_in[2][3][10] ), .X(n16269) );
  inv_x2_sg U11695 ( .A(\reg_in[2][3][9] ), .X(n16271) );
  inv_x2_sg U11696 ( .A(\reg_in[2][3][8] ), .X(n16273) );
  inv_x2_sg U11697 ( .A(\reg_in[2][3][7] ), .X(n16275) );
  inv_x2_sg U11698 ( .A(\reg_in[2][3][6] ), .X(n16277) );
  inv_x2_sg U11699 ( .A(\reg_in[2][3][5] ), .X(n16279) );
  inv_x2_sg U11700 ( .A(\reg_in[2][3][4] ), .X(n16281) );
  inv_x2_sg U11701 ( .A(\reg_in[2][3][3] ), .X(n16283) );
  inv_x2_sg U11702 ( .A(\reg_in[2][3][2] ), .X(n16285) );
  inv_x2_sg U11703 ( .A(\reg_in[2][3][1] ), .X(n16287) );
  inv_x2_sg U11704 ( .A(\reg_in[2][3][0] ), .X(n16289) );
  inv_x2_sg U11705 ( .A(\reg_in[2][2][19] ), .X(n16291) );
  inv_x2_sg U11706 ( .A(\reg_in[2][2][18] ), .X(n16293) );
  inv_x2_sg U11707 ( .A(\reg_in[2][2][17] ), .X(n16295) );
  inv_x2_sg U11708 ( .A(\reg_in[2][2][16] ), .X(n16297) );
  inv_x2_sg U11709 ( .A(\reg_in[2][2][15] ), .X(n16299) );
  inv_x2_sg U11710 ( .A(\reg_in[2][2][14] ), .X(n16301) );
  inv_x2_sg U11711 ( .A(\reg_in[2][2][13] ), .X(n16303) );
  inv_x2_sg U11712 ( .A(\reg_in[2][2][12] ), .X(n16305) );
  inv_x2_sg U11713 ( .A(\reg_in[2][2][11] ), .X(n16307) );
  inv_x2_sg U11714 ( .A(\reg_in[2][2][10] ), .X(n16309) );
  inv_x2_sg U11715 ( .A(\reg_in[2][2][9] ), .X(n16311) );
  inv_x2_sg U11716 ( .A(\reg_in[2][2][8] ), .X(n16313) );
  inv_x2_sg U11717 ( .A(\reg_in[2][2][7] ), .X(n16315) );
  inv_x2_sg U11718 ( .A(\reg_in[2][2][6] ), .X(n16317) );
  inv_x2_sg U11719 ( .A(\reg_in[2][2][5] ), .X(n16319) );
  inv_x2_sg U11720 ( .A(\reg_in[2][2][4] ), .X(n16321) );
  inv_x2_sg U11721 ( .A(\reg_in[2][2][3] ), .X(n16323) );
  inv_x2_sg U11722 ( .A(\reg_in[2][2][2] ), .X(n16325) );
  inv_x2_sg U11723 ( .A(\reg_in[2][2][1] ), .X(n16327) );
  inv_x2_sg U11724 ( .A(\reg_in[2][2][0] ), .X(n16329) );
  inv_x2_sg U11725 ( .A(\reg_in[2][1][19] ), .X(n16331) );
  inv_x2_sg U11726 ( .A(\reg_in[2][1][18] ), .X(n16333) );
  inv_x2_sg U11727 ( .A(\reg_in[2][1][17] ), .X(n16335) );
  inv_x2_sg U11728 ( .A(\reg_in[2][1][16] ), .X(n16337) );
  inv_x2_sg U11729 ( .A(\reg_in[2][1][15] ), .X(n16339) );
  inv_x2_sg U11730 ( .A(\reg_in[2][1][14] ), .X(n16341) );
  inv_x2_sg U11731 ( .A(\reg_in[2][1][13] ), .X(n16343) );
  inv_x2_sg U11732 ( .A(\reg_in[2][1][12] ), .X(n16345) );
  inv_x2_sg U11733 ( .A(\reg_in[2][1][11] ), .X(n16347) );
  inv_x2_sg U11734 ( .A(\reg_in[2][1][10] ), .X(n16349) );
  inv_x2_sg U11735 ( .A(\reg_in[2][1][9] ), .X(n16351) );
  inv_x2_sg U11736 ( .A(\reg_in[2][1][8] ), .X(n16353) );
  inv_x2_sg U11737 ( .A(\reg_in[2][1][7] ), .X(n16355) );
  inv_x2_sg U11738 ( .A(\reg_in[2][1][6] ), .X(n16357) );
  inv_x2_sg U11739 ( .A(\reg_in[2][1][5] ), .X(n16359) );
  inv_x2_sg U11740 ( .A(\reg_in[2][1][4] ), .X(n16361) );
  inv_x2_sg U11741 ( .A(\reg_in[2][1][3] ), .X(n16363) );
  inv_x2_sg U11742 ( .A(\reg_in[2][1][2] ), .X(n16365) );
  inv_x2_sg U11743 ( .A(\reg_in[2][1][1] ), .X(n16367) );
  inv_x2_sg U11744 ( .A(\reg_in[2][1][0] ), .X(n16369) );
  inv_x2_sg U11745 ( .A(\reg_in[2][0][19] ), .X(n16371) );
  inv_x2_sg U11746 ( .A(\reg_in[2][0][18] ), .X(n16373) );
  inv_x2_sg U11747 ( .A(\reg_in[2][0][17] ), .X(n16375) );
  inv_x2_sg U11748 ( .A(\reg_in[2][0][16] ), .X(n16377) );
  inv_x2_sg U11749 ( .A(\reg_in[2][0][15] ), .X(n16379) );
  inv_x2_sg U11750 ( .A(\reg_in[2][0][14] ), .X(n16381) );
  inv_x2_sg U11751 ( .A(\reg_in[2][0][13] ), .X(n16383) );
  inv_x2_sg U11752 ( .A(\reg_in[2][0][12] ), .X(n16385) );
  inv_x2_sg U11753 ( .A(\reg_in[2][0][11] ), .X(n16387) );
  inv_x2_sg U11754 ( .A(\reg_in[2][0][10] ), .X(n16389) );
  inv_x2_sg U11755 ( .A(\reg_in[2][0][9] ), .X(n16391) );
  inv_x2_sg U11756 ( .A(\reg_in[2][0][8] ), .X(n16393) );
  inv_x2_sg U11757 ( .A(\reg_in[2][0][7] ), .X(n16395) );
  inv_x2_sg U11758 ( .A(\reg_in[2][0][6] ), .X(n16397) );
  inv_x2_sg U11759 ( .A(\reg_in[2][0][5] ), .X(n16399) );
  inv_x2_sg U11760 ( .A(\reg_in[2][0][4] ), .X(n16401) );
  inv_x2_sg U11761 ( .A(\reg_in[2][0][3] ), .X(n16403) );
  inv_x2_sg U11762 ( .A(\reg_in[2][0][2] ), .X(n16405) );
  inv_x2_sg U11763 ( .A(\reg_in[2][0][1] ), .X(n16407) );
  inv_x2_sg U11764 ( .A(\reg_in[2][0][0] ), .X(n16409) );
  inv_x2_sg U11765 ( .A(\reg_in[1][3][19] ), .X(n16411) );
  inv_x2_sg U11766 ( .A(\reg_in[1][3][18] ), .X(n16413) );
  inv_x2_sg U11767 ( .A(\reg_in[1][3][17] ), .X(n16415) );
  inv_x2_sg U11768 ( .A(\reg_in[1][3][16] ), .X(n16417) );
  inv_x2_sg U11769 ( .A(\reg_in[1][3][15] ), .X(n16419) );
  inv_x2_sg U11770 ( .A(\reg_in[1][3][14] ), .X(n16421) );
  inv_x2_sg U11771 ( .A(\reg_in[1][3][13] ), .X(n16423) );
  inv_x2_sg U11772 ( .A(\reg_in[1][3][12] ), .X(n16425) );
  inv_x2_sg U11773 ( .A(\reg_in[1][3][11] ), .X(n16427) );
  inv_x2_sg U11774 ( .A(\reg_in[1][3][10] ), .X(n16429) );
  inv_x2_sg U11775 ( .A(\reg_in[1][3][9] ), .X(n16431) );
  inv_x2_sg U11776 ( .A(\reg_in[1][3][8] ), .X(n16433) );
  inv_x2_sg U11777 ( .A(\reg_in[1][3][7] ), .X(n16435) );
  inv_x2_sg U11778 ( .A(\reg_in[1][3][6] ), .X(n16437) );
  inv_x2_sg U11779 ( .A(\reg_in[1][3][5] ), .X(n16439) );
  inv_x2_sg U11780 ( .A(\reg_in[1][3][4] ), .X(n16441) );
  inv_x2_sg U11781 ( .A(\reg_in[1][3][3] ), .X(n16443) );
  inv_x2_sg U11782 ( .A(\reg_in[1][3][2] ), .X(n16445) );
  inv_x2_sg U11783 ( .A(\reg_in[1][3][1] ), .X(n16447) );
  inv_x2_sg U11784 ( .A(\reg_in[1][3][0] ), .X(n16449) );
  inv_x2_sg U11785 ( .A(\reg_in[1][2][19] ), .X(n16451) );
  inv_x2_sg U11786 ( .A(\reg_in[1][2][18] ), .X(n16453) );
  inv_x2_sg U11787 ( .A(\reg_in[1][2][17] ), .X(n16455) );
  inv_x2_sg U11788 ( .A(\reg_in[1][2][16] ), .X(n16457) );
  inv_x2_sg U11789 ( .A(\reg_in[1][2][15] ), .X(n16459) );
  inv_x2_sg U11790 ( .A(\reg_in[1][2][14] ), .X(n16461) );
  inv_x2_sg U11791 ( .A(\reg_in[1][2][13] ), .X(n16463) );
  inv_x2_sg U11792 ( .A(\reg_in[1][2][12] ), .X(n16465) );
  inv_x2_sg U11793 ( .A(\reg_in[1][2][11] ), .X(n16467) );
  inv_x2_sg U11794 ( .A(\reg_in[1][2][10] ), .X(n16469) );
  inv_x2_sg U11795 ( .A(\reg_in[1][2][9] ), .X(n16471) );
  inv_x2_sg U11796 ( .A(\reg_in[1][2][8] ), .X(n16473) );
  inv_x2_sg U11797 ( .A(\reg_in[1][2][7] ), .X(n16475) );
  inv_x2_sg U11798 ( .A(\reg_in[1][2][6] ), .X(n16477) );
  inv_x2_sg U11799 ( .A(\reg_in[1][2][5] ), .X(n16479) );
  inv_x2_sg U11800 ( .A(\reg_in[1][2][4] ), .X(n16481) );
  inv_x2_sg U11801 ( .A(\reg_in[1][2][3] ), .X(n16483) );
  inv_x2_sg U11802 ( .A(\reg_in[1][2][2] ), .X(n16485) );
  inv_x2_sg U11803 ( .A(\reg_in[1][2][1] ), .X(n16487) );
  inv_x2_sg U11804 ( .A(\reg_in[1][2][0] ), .X(n16489) );
  inv_x2_sg U11805 ( .A(\reg_in[1][1][19] ), .X(n16491) );
  inv_x2_sg U11806 ( .A(\reg_in[1][1][18] ), .X(n16493) );
  inv_x2_sg U11807 ( .A(\reg_in[1][1][17] ), .X(n16495) );
  inv_x2_sg U11808 ( .A(\reg_in[1][1][16] ), .X(n16497) );
  inv_x2_sg U11809 ( .A(\reg_in[1][1][15] ), .X(n16499) );
  inv_x2_sg U11810 ( .A(\reg_in[1][1][14] ), .X(n16501) );
  inv_x2_sg U11811 ( .A(\reg_in[1][1][13] ), .X(n16503) );
  inv_x2_sg U11812 ( .A(\reg_in[1][1][12] ), .X(n16505) );
  inv_x2_sg U11813 ( .A(\reg_in[1][1][11] ), .X(n16507) );
  inv_x2_sg U11814 ( .A(\reg_in[1][1][10] ), .X(n16509) );
  inv_x2_sg U11815 ( .A(\reg_in[1][1][9] ), .X(n16511) );
  inv_x2_sg U11816 ( .A(\reg_in[1][1][8] ), .X(n16513) );
  inv_x2_sg U11817 ( .A(\reg_in[1][1][7] ), .X(n16515) );
  inv_x2_sg U11818 ( .A(\reg_in[1][1][6] ), .X(n16517) );
  inv_x2_sg U11819 ( .A(\reg_in[1][1][5] ), .X(n16519) );
  inv_x2_sg U11820 ( .A(\reg_in[1][1][4] ), .X(n16521) );
  inv_x2_sg U11821 ( .A(\reg_in[1][1][3] ), .X(n16523) );
  inv_x2_sg U11822 ( .A(\reg_in[1][1][2] ), .X(n16525) );
  inv_x2_sg U11823 ( .A(\reg_in[1][1][1] ), .X(n16527) );
  inv_x2_sg U11824 ( .A(\reg_in[1][1][0] ), .X(n16529) );
  inv_x2_sg U11825 ( .A(\reg_in[1][0][19] ), .X(n16531) );
  inv_x2_sg U11826 ( .A(\reg_in[1][0][18] ), .X(n16533) );
  inv_x2_sg U11827 ( .A(\reg_in[1][0][17] ), .X(n16535) );
  inv_x2_sg U11828 ( .A(\reg_in[1][0][16] ), .X(n16537) );
  inv_x2_sg U11829 ( .A(\reg_in[1][0][15] ), .X(n16539) );
  inv_x2_sg U11830 ( .A(\reg_in[1][0][14] ), .X(n16541) );
  inv_x2_sg U11831 ( .A(\reg_in[1][0][13] ), .X(n16543) );
  inv_x2_sg U11832 ( .A(\reg_in[1][0][12] ), .X(n16545) );
  inv_x2_sg U11833 ( .A(\reg_in[1][0][11] ), .X(n16547) );
  inv_x2_sg U11834 ( .A(\reg_in[1][0][10] ), .X(n16549) );
  inv_x2_sg U11835 ( .A(\reg_in[1][0][9] ), .X(n16551) );
  inv_x2_sg U11836 ( .A(\reg_in[1][0][8] ), .X(n16553) );
  inv_x2_sg U11837 ( .A(\reg_in[1][0][7] ), .X(n16555) );
  inv_x2_sg U11838 ( .A(\reg_in[1][0][6] ), .X(n16557) );
  inv_x2_sg U11839 ( .A(\reg_in[1][0][5] ), .X(n16559) );
  inv_x2_sg U11840 ( .A(\reg_in[1][0][4] ), .X(n16561) );
  inv_x2_sg U11841 ( .A(\reg_in[1][0][3] ), .X(n16563) );
  inv_x2_sg U11842 ( .A(\reg_in[1][0][2] ), .X(n16565) );
  inv_x2_sg U11843 ( .A(\reg_in[1][0][1] ), .X(n16567) );
  inv_x2_sg U11844 ( .A(\reg_in[1][0][0] ), .X(n16569) );
  inv_x2_sg U11845 ( .A(\reg_in[0][3][19] ), .X(n16571) );
  inv_x2_sg U11846 ( .A(\reg_in[0][3][18] ), .X(n16573) );
  inv_x2_sg U11847 ( .A(\reg_in[0][3][17] ), .X(n16575) );
  inv_x2_sg U11848 ( .A(\reg_in[0][3][16] ), .X(n16577) );
  inv_x2_sg U11849 ( .A(\reg_in[0][3][15] ), .X(n16579) );
  inv_x2_sg U11850 ( .A(\reg_in[0][3][14] ), .X(n16581) );
  inv_x2_sg U11851 ( .A(\reg_in[0][3][13] ), .X(n16583) );
  inv_x2_sg U11852 ( .A(\reg_in[0][3][12] ), .X(n16585) );
  inv_x2_sg U11853 ( .A(\reg_in[0][3][11] ), .X(n16587) );
  inv_x2_sg U11854 ( .A(\reg_in[0][3][10] ), .X(n16589) );
  inv_x2_sg U11855 ( .A(\reg_in[0][3][9] ), .X(n16591) );
  inv_x2_sg U11856 ( .A(\reg_in[0][3][8] ), .X(n16593) );
  inv_x2_sg U11857 ( .A(\reg_in[0][3][7] ), .X(n16595) );
  inv_x2_sg U11858 ( .A(\reg_in[0][3][6] ), .X(n16597) );
  inv_x2_sg U11859 ( .A(\reg_in[0][3][5] ), .X(n16599) );
  inv_x2_sg U11860 ( .A(\reg_in[0][3][4] ), .X(n16601) );
  inv_x2_sg U11861 ( .A(\reg_in[0][3][3] ), .X(n16603) );
  inv_x2_sg U11862 ( .A(\reg_in[0][3][2] ), .X(n16605) );
  inv_x2_sg U11863 ( .A(\reg_in[0][3][1] ), .X(n16607) );
  inv_x2_sg U11864 ( .A(\reg_in[0][3][0] ), .X(n16609) );
  inv_x2_sg U11865 ( .A(\reg_in[0][2][19] ), .X(n16611) );
  inv_x2_sg U11866 ( .A(\reg_in[0][2][18] ), .X(n16613) );
  inv_x2_sg U11867 ( .A(\reg_in[0][2][17] ), .X(n16615) );
  inv_x2_sg U11868 ( .A(\reg_in[0][2][16] ), .X(n16617) );
  inv_x2_sg U11869 ( .A(\reg_in[0][2][15] ), .X(n16619) );
  inv_x2_sg U11870 ( .A(\reg_in[0][2][14] ), .X(n16621) );
  inv_x2_sg U11871 ( .A(\reg_in[0][2][13] ), .X(n16623) );
  inv_x2_sg U11872 ( .A(\reg_in[0][2][12] ), .X(n16625) );
  inv_x2_sg U11873 ( .A(\reg_in[0][2][11] ), .X(n16627) );
  inv_x2_sg U11874 ( .A(\reg_in[0][2][10] ), .X(n16629) );
  inv_x2_sg U11875 ( .A(\reg_in[0][2][9] ), .X(n16631) );
  inv_x2_sg U11876 ( .A(\reg_in[0][2][8] ), .X(n16633) );
  inv_x2_sg U11877 ( .A(\reg_in[0][2][7] ), .X(n16635) );
  inv_x2_sg U11878 ( .A(\reg_in[0][2][6] ), .X(n16637) );
  inv_x2_sg U11879 ( .A(\reg_in[0][2][5] ), .X(n16639) );
  inv_x2_sg U11880 ( .A(\reg_in[0][2][4] ), .X(n16641) );
  inv_x2_sg U11881 ( .A(\reg_in[0][2][3] ), .X(n16643) );
  inv_x2_sg U11882 ( .A(\reg_in[0][2][2] ), .X(n16645) );
  inv_x2_sg U11883 ( .A(\reg_in[0][2][1] ), .X(n16647) );
  inv_x2_sg U11884 ( .A(\reg_in[0][2][0] ), .X(n16649) );
  inv_x2_sg U11885 ( .A(\reg_in[0][1][19] ), .X(n16651) );
  inv_x2_sg U11886 ( .A(\reg_in[0][1][18] ), .X(n16653) );
  inv_x2_sg U11887 ( .A(\reg_in[0][1][17] ), .X(n16655) );
  inv_x2_sg U11888 ( .A(\reg_in[0][1][16] ), .X(n16657) );
  inv_x2_sg U11889 ( .A(\reg_in[0][1][15] ), .X(n16659) );
  inv_x2_sg U11890 ( .A(\reg_in[0][1][14] ), .X(n16661) );
  inv_x2_sg U11891 ( .A(\reg_in[0][1][13] ), .X(n16663) );
  inv_x2_sg U11892 ( .A(\reg_in[0][1][12] ), .X(n16665) );
  inv_x2_sg U11893 ( .A(\reg_in[0][1][11] ), .X(n16667) );
  inv_x2_sg U11894 ( .A(\reg_in[0][1][10] ), .X(n16669) );
  inv_x2_sg U11895 ( .A(\reg_in[0][1][9] ), .X(n16671) );
  inv_x2_sg U11896 ( .A(\reg_in[0][1][8] ), .X(n16673) );
  inv_x2_sg U11897 ( .A(\reg_in[0][1][7] ), .X(n16675) );
  inv_x2_sg U11898 ( .A(\reg_in[0][1][6] ), .X(n16677) );
  inv_x2_sg U11899 ( .A(\reg_in[0][1][5] ), .X(n16679) );
  inv_x2_sg U11900 ( .A(\reg_in[0][1][4] ), .X(n16681) );
  inv_x2_sg U11901 ( .A(\reg_in[0][1][3] ), .X(n16683) );
  inv_x2_sg U11902 ( .A(\reg_in[0][1][2] ), .X(n16685) );
  inv_x2_sg U11903 ( .A(\reg_in[0][1][1] ), .X(n16687) );
  inv_x2_sg U11904 ( .A(\reg_in[0][1][0] ), .X(n16689) );
  inv_x2_sg U11905 ( .A(\reg_in[0][0][19] ), .X(n16691) );
  inv_x2_sg U11906 ( .A(\reg_in[0][0][18] ), .X(n16693) );
  inv_x2_sg U11907 ( .A(\reg_in[0][0][17] ), .X(n16695) );
  inv_x2_sg U11908 ( .A(\reg_in[0][0][16] ), .X(n16697) );
  inv_x2_sg U11909 ( .A(\reg_in[0][0][15] ), .X(n16699) );
  inv_x2_sg U11910 ( .A(\reg_in[0][0][14] ), .X(n16701) );
  inv_x2_sg U11911 ( .A(\reg_in[0][0][13] ), .X(n16703) );
  inv_x2_sg U11912 ( .A(\reg_in[0][0][12] ), .X(n16705) );
  inv_x2_sg U11913 ( .A(\reg_in[0][0][11] ), .X(n16707) );
  inv_x2_sg U11914 ( .A(\reg_in[0][0][10] ), .X(n16709) );
  inv_x2_sg U11915 ( .A(\reg_in[0][0][9] ), .X(n16711) );
  inv_x2_sg U11916 ( .A(\reg_in[0][0][8] ), .X(n16713) );
  inv_x2_sg U11917 ( .A(\reg_in[0][0][7] ), .X(n16715) );
  inv_x2_sg U11918 ( .A(\reg_in[0][0][6] ), .X(n16717) );
  inv_x2_sg U11919 ( .A(\reg_in[0][0][5] ), .X(n16719) );
  inv_x2_sg U11920 ( .A(\reg_in[0][0][4] ), .X(n16721) );
  inv_x2_sg U11921 ( .A(\reg_in[0][0][3] ), .X(n16723) );
  inv_x2_sg U11922 ( .A(\reg_in[0][0][2] ), .X(n16725) );
  inv_x2_sg U11923 ( .A(\reg_in[0][0][1] ), .X(n16727) );
  inv_x2_sg U11924 ( .A(\reg_in[0][0][0] ), .X(n16729) );
  inv_x8_sg U11925 ( .A(state[1]), .X(n18399) );
  inv_x2_sg U11926 ( .A(n15451), .X(\out[3][3][19] ) );
  inv_x2_sg U11927 ( .A(n15453), .X(\out[3][3][18] ) );
  inv_x2_sg U11928 ( .A(n15455), .X(\out[3][3][17] ) );
  inv_x2_sg U11929 ( .A(n15457), .X(\out[3][3][16] ) );
  inv_x2_sg U11930 ( .A(n15459), .X(\out[3][3][15] ) );
  inv_x2_sg U11931 ( .A(n15461), .X(\out[3][3][14] ) );
  inv_x2_sg U11932 ( .A(n15463), .X(\out[3][3][13] ) );
  inv_x2_sg U11933 ( .A(n15465), .X(\out[3][3][12] ) );
  inv_x2_sg U11934 ( .A(n15467), .X(\out[3][3][11] ) );
  inv_x2_sg U11935 ( .A(n15469), .X(\out[3][3][10] ) );
  inv_x2_sg U11936 ( .A(n15471), .X(\out[3][3][9] ) );
  inv_x2_sg U11937 ( .A(n15473), .X(\out[3][3][8] ) );
  inv_x2_sg U11938 ( .A(n15475), .X(\out[3][3][7] ) );
  inv_x2_sg U11939 ( .A(n15477), .X(\out[3][3][6] ) );
  inv_x2_sg U11940 ( .A(n15479), .X(\out[3][3][5] ) );
  inv_x2_sg U11941 ( .A(n15481), .X(\out[3][3][4] ) );
  inv_x2_sg U11942 ( .A(n15483), .X(\out[3][3][3] ) );
  inv_x2_sg U11943 ( .A(n15485), .X(\out[3][3][2] ) );
  inv_x2_sg U11944 ( .A(n15487), .X(\out[3][3][1] ) );
  inv_x2_sg U11945 ( .A(n15489), .X(\out[3][3][0] ) );
  inv_x2_sg U11946 ( .A(n15491), .X(\out[3][2][19] ) );
  inv_x2_sg U11947 ( .A(n15493), .X(\out[3][2][18] ) );
  inv_x2_sg U11948 ( .A(n15495), .X(\out[3][2][17] ) );
  inv_x2_sg U11949 ( .A(n15497), .X(\out[3][2][16] ) );
  inv_x2_sg U11950 ( .A(n15499), .X(\out[3][2][15] ) );
  inv_x2_sg U11951 ( .A(n15501), .X(\out[3][2][14] ) );
  inv_x2_sg U11952 ( .A(n15503), .X(\out[3][2][13] ) );
  inv_x2_sg U11953 ( .A(n15505), .X(\out[3][2][12] ) );
  inv_x2_sg U11954 ( .A(n15507), .X(\out[3][2][11] ) );
  inv_x2_sg U11955 ( .A(n15509), .X(\out[3][2][10] ) );
  inv_x2_sg U11956 ( .A(n15511), .X(\out[3][2][9] ) );
  inv_x2_sg U11957 ( .A(n15513), .X(\out[3][2][8] ) );
  inv_x2_sg U11958 ( .A(n15515), .X(\out[3][2][7] ) );
  inv_x2_sg U11959 ( .A(n15517), .X(\out[3][2][6] ) );
  inv_x2_sg U11960 ( .A(n15519), .X(\out[3][2][5] ) );
  inv_x2_sg U11961 ( .A(n15521), .X(\out[3][2][4] ) );
  inv_x2_sg U11962 ( .A(n15523), .X(\out[3][2][3] ) );
  inv_x2_sg U11963 ( .A(n15525), .X(\out[3][2][2] ) );
  inv_x2_sg U11964 ( .A(n15527), .X(\out[3][2][1] ) );
  inv_x2_sg U11965 ( .A(n15529), .X(\out[3][2][0] ) );
  inv_x2_sg U11966 ( .A(n15531), .X(\out[3][1][19] ) );
  inv_x2_sg U11967 ( .A(n15533), .X(\out[3][1][18] ) );
  inv_x2_sg U11968 ( .A(n15535), .X(\out[3][1][17] ) );
  inv_x2_sg U11969 ( .A(n15537), .X(\out[3][1][16] ) );
  inv_x2_sg U11970 ( .A(n15539), .X(\out[3][1][15] ) );
  inv_x2_sg U11971 ( .A(n15541), .X(\out[3][1][14] ) );
  inv_x2_sg U11972 ( .A(n15543), .X(\out[3][1][13] ) );
  inv_x2_sg U11973 ( .A(n15545), .X(\out[3][1][12] ) );
  inv_x2_sg U11974 ( .A(n15547), .X(\out[3][1][11] ) );
  inv_x2_sg U11975 ( .A(n15549), .X(\out[3][1][10] ) );
  inv_x2_sg U11976 ( .A(n15551), .X(\out[3][1][9] ) );
  inv_x2_sg U11977 ( .A(n15553), .X(\out[3][1][8] ) );
  inv_x2_sg U11978 ( .A(n15555), .X(\out[3][1][7] ) );
  inv_x2_sg U11979 ( .A(n15557), .X(\out[3][1][6] ) );
  inv_x2_sg U11980 ( .A(n15559), .X(\out[3][1][5] ) );
  inv_x2_sg U11981 ( .A(n15561), .X(\out[3][1][4] ) );
  inv_x2_sg U11982 ( .A(n15563), .X(\out[3][1][3] ) );
  inv_x2_sg U11983 ( .A(n15565), .X(\out[3][1][2] ) );
  inv_x2_sg U11984 ( .A(n15567), .X(\out[3][1][1] ) );
  inv_x2_sg U11985 ( .A(n15569), .X(\out[3][1][0] ) );
  inv_x2_sg U11986 ( .A(n15571), .X(\out[3][0][19] ) );
  inv_x2_sg U11987 ( .A(n15573), .X(\out[3][0][18] ) );
  inv_x2_sg U11988 ( .A(n15575), .X(\out[3][0][17] ) );
  inv_x2_sg U11989 ( .A(n15577), .X(\out[3][0][16] ) );
  inv_x2_sg U11990 ( .A(n15579), .X(\out[3][0][15] ) );
  inv_x2_sg U11991 ( .A(n15581), .X(\out[3][0][14] ) );
  inv_x2_sg U11992 ( .A(n15583), .X(\out[3][0][13] ) );
  inv_x2_sg U11993 ( .A(n15585), .X(\out[3][0][12] ) );
  inv_x2_sg U11994 ( .A(n15587), .X(\out[3][0][11] ) );
  inv_x2_sg U11995 ( .A(n15589), .X(\out[3][0][10] ) );
  inv_x2_sg U11996 ( .A(n15591), .X(\out[3][0][9] ) );
  inv_x2_sg U11997 ( .A(n15593), .X(\out[3][0][8] ) );
  inv_x2_sg U11998 ( .A(n15595), .X(\out[3][0][7] ) );
  inv_x2_sg U11999 ( .A(n15597), .X(\out[3][0][6] ) );
  inv_x2_sg U12000 ( .A(n15599), .X(\out[3][0][5] ) );
  inv_x2_sg U12001 ( .A(n15601), .X(\out[3][0][4] ) );
  inv_x2_sg U12002 ( .A(n15603), .X(\out[3][0][3] ) );
  inv_x2_sg U12003 ( .A(n15605), .X(\out[3][0][2] ) );
  inv_x2_sg U12004 ( .A(n15607), .X(\out[3][0][1] ) );
  inv_x2_sg U12005 ( .A(n15609), .X(\out[3][0][0] ) );
  inv_x2_sg U12006 ( .A(n15611), .X(\out[2][3][19] ) );
  inv_x2_sg U12007 ( .A(n15613), .X(\out[2][3][18] ) );
  inv_x2_sg U12008 ( .A(n15615), .X(\out[2][3][17] ) );
  inv_x2_sg U12009 ( .A(n15617), .X(\out[2][3][16] ) );
  inv_x2_sg U12010 ( .A(n15619), .X(\out[2][3][15] ) );
  inv_x2_sg U12011 ( .A(n15621), .X(\out[2][3][14] ) );
  inv_x2_sg U12012 ( .A(n15623), .X(\out[2][3][13] ) );
  inv_x2_sg U12013 ( .A(n15625), .X(\out[2][3][12] ) );
  inv_x2_sg U12014 ( .A(n15627), .X(\out[2][3][11] ) );
  inv_x2_sg U12015 ( .A(n15629), .X(\out[2][3][10] ) );
  inv_x2_sg U12016 ( .A(n15631), .X(\out[2][3][9] ) );
  inv_x2_sg U12017 ( .A(n15633), .X(\out[2][3][8] ) );
  inv_x2_sg U12018 ( .A(n15635), .X(\out[2][3][7] ) );
  inv_x2_sg U12019 ( .A(n15637), .X(\out[2][3][6] ) );
  inv_x2_sg U12020 ( .A(n15639), .X(\out[2][3][5] ) );
  inv_x2_sg U12021 ( .A(n15641), .X(\out[2][3][4] ) );
  inv_x2_sg U12022 ( .A(n15643), .X(\out[2][3][3] ) );
  inv_x2_sg U12023 ( .A(n15645), .X(\out[2][3][2] ) );
  inv_x2_sg U12024 ( .A(n15647), .X(\out[2][3][1] ) );
  inv_x2_sg U12025 ( .A(n15649), .X(\out[2][3][0] ) );
  inv_x2_sg U12026 ( .A(n15651), .X(\out[2][2][19] ) );
  inv_x2_sg U12027 ( .A(n15653), .X(\out[2][2][18] ) );
  inv_x2_sg U12028 ( .A(n15655), .X(\out[2][2][17] ) );
  inv_x2_sg U12029 ( .A(n15657), .X(\out[2][2][16] ) );
  inv_x2_sg U12030 ( .A(n15659), .X(\out[2][2][15] ) );
  inv_x2_sg U12031 ( .A(n15661), .X(\out[2][2][14] ) );
  inv_x2_sg U12032 ( .A(n15663), .X(\out[2][2][13] ) );
  inv_x2_sg U12033 ( .A(n15665), .X(\out[2][2][12] ) );
  inv_x2_sg U12034 ( .A(n15667), .X(\out[2][2][11] ) );
  inv_x2_sg U12035 ( .A(n15669), .X(\out[2][2][10] ) );
  inv_x2_sg U12036 ( .A(n15671), .X(\out[2][2][9] ) );
  inv_x2_sg U12037 ( .A(n15673), .X(\out[2][2][8] ) );
  inv_x2_sg U12038 ( .A(n15675), .X(\out[2][2][7] ) );
  inv_x2_sg U12039 ( .A(n15677), .X(\out[2][2][6] ) );
  inv_x2_sg U12040 ( .A(n15679), .X(\out[2][2][5] ) );
  inv_x2_sg U12041 ( .A(n15681), .X(\out[2][2][4] ) );
  inv_x2_sg U12042 ( .A(n15683), .X(\out[2][2][3] ) );
  inv_x2_sg U12043 ( .A(n15685), .X(\out[2][2][2] ) );
  inv_x2_sg U12044 ( .A(n15687), .X(\out[2][2][1] ) );
  inv_x2_sg U12045 ( .A(n15689), .X(\out[2][2][0] ) );
  inv_x2_sg U12046 ( .A(n15691), .X(\out[2][1][19] ) );
  inv_x2_sg U12047 ( .A(n15693), .X(\out[2][1][18] ) );
  inv_x2_sg U12048 ( .A(n15695), .X(\out[2][1][17] ) );
  inv_x2_sg U12049 ( .A(n15697), .X(\out[2][1][16] ) );
  inv_x2_sg U12050 ( .A(n15699), .X(\out[2][1][15] ) );
  inv_x2_sg U12051 ( .A(n15701), .X(\out[2][1][14] ) );
  inv_x2_sg U12052 ( .A(n15703), .X(\out[2][1][13] ) );
  inv_x2_sg U12053 ( .A(n15705), .X(\out[2][1][12] ) );
  inv_x2_sg U12054 ( .A(n15707), .X(\out[2][1][11] ) );
  inv_x2_sg U12055 ( .A(n15709), .X(\out[2][1][10] ) );
  inv_x2_sg U12056 ( .A(n15711), .X(\out[2][1][9] ) );
  inv_x2_sg U12057 ( .A(n15713), .X(\out[2][1][8] ) );
  inv_x2_sg U12058 ( .A(n15715), .X(\out[2][1][7] ) );
  inv_x2_sg U12059 ( .A(n15717), .X(\out[2][1][6] ) );
  inv_x2_sg U12060 ( .A(n15719), .X(\out[2][1][5] ) );
  inv_x2_sg U12061 ( .A(n15721), .X(\out[2][1][4] ) );
  inv_x2_sg U12062 ( .A(n15723), .X(\out[2][1][3] ) );
  inv_x2_sg U12063 ( .A(n15725), .X(\out[2][1][2] ) );
  inv_x2_sg U12064 ( .A(n15727), .X(\out[2][1][1] ) );
  inv_x2_sg U12065 ( .A(n15729), .X(\out[2][1][0] ) );
  inv_x2_sg U12066 ( .A(n15731), .X(\out[2][0][19] ) );
  inv_x2_sg U12067 ( .A(n15733), .X(\out[2][0][18] ) );
  inv_x2_sg U12068 ( .A(n15735), .X(\out[2][0][17] ) );
  inv_x2_sg U12069 ( .A(n15737), .X(\out[2][0][16] ) );
  inv_x2_sg U12070 ( .A(n15739), .X(\out[2][0][15] ) );
  inv_x2_sg U12071 ( .A(n15741), .X(\out[2][0][14] ) );
  inv_x2_sg U12072 ( .A(n15743), .X(\out[2][0][13] ) );
  inv_x2_sg U12073 ( .A(n15745), .X(\out[2][0][12] ) );
  inv_x2_sg U12074 ( .A(n15747), .X(\out[2][0][11] ) );
  inv_x2_sg U12075 ( .A(n15749), .X(\out[2][0][10] ) );
  inv_x2_sg U12076 ( .A(n15751), .X(\out[2][0][9] ) );
  inv_x2_sg U12077 ( .A(n15753), .X(\out[2][0][8] ) );
  inv_x2_sg U12078 ( .A(n15755), .X(\out[2][0][7] ) );
  inv_x2_sg U12079 ( .A(n15757), .X(\out[2][0][6] ) );
  inv_x2_sg U12080 ( .A(n15759), .X(\out[2][0][5] ) );
  inv_x2_sg U12081 ( .A(n15761), .X(\out[2][0][4] ) );
  inv_x2_sg U12082 ( .A(n15763), .X(\out[2][0][3] ) );
  inv_x2_sg U12083 ( .A(n15765), .X(\out[2][0][2] ) );
  inv_x2_sg U12084 ( .A(n15767), .X(\out[2][0][1] ) );
  inv_x2_sg U12085 ( .A(n15769), .X(\out[2][0][0] ) );
  inv_x2_sg U12086 ( .A(n15771), .X(\out[1][3][19] ) );
  inv_x2_sg U12087 ( .A(n15773), .X(\out[1][3][18] ) );
  inv_x2_sg U12088 ( .A(n15775), .X(\out[1][3][17] ) );
  inv_x2_sg U12089 ( .A(n15777), .X(\out[1][3][16] ) );
  inv_x2_sg U12090 ( .A(n15779), .X(\out[1][3][15] ) );
  inv_x2_sg U12091 ( .A(n15781), .X(\out[1][3][14] ) );
  inv_x2_sg U12092 ( .A(n15783), .X(\out[1][3][13] ) );
  inv_x2_sg U12093 ( .A(n15785), .X(\out[1][3][12] ) );
  inv_x2_sg U12094 ( .A(n15787), .X(\out[1][3][11] ) );
  inv_x2_sg U12095 ( .A(n15789), .X(\out[1][3][10] ) );
  inv_x2_sg U12096 ( .A(n15791), .X(\out[1][3][9] ) );
  inv_x2_sg U12097 ( .A(n15793), .X(\out[1][3][8] ) );
  inv_x2_sg U12098 ( .A(n15795), .X(\out[1][3][7] ) );
  inv_x2_sg U12099 ( .A(n15797), .X(\out[1][3][6] ) );
  inv_x2_sg U12100 ( .A(n15799), .X(\out[1][3][5] ) );
  inv_x2_sg U12101 ( .A(n15801), .X(\out[1][3][4] ) );
  inv_x2_sg U12102 ( .A(n15803), .X(\out[1][3][3] ) );
  inv_x2_sg U12103 ( .A(n15805), .X(\out[1][3][2] ) );
  inv_x2_sg U12104 ( .A(n15807), .X(\out[1][3][1] ) );
  inv_x2_sg U12105 ( .A(n15809), .X(\out[1][3][0] ) );
  inv_x2_sg U12106 ( .A(n15811), .X(\out[1][2][19] ) );
  inv_x2_sg U12107 ( .A(n15813), .X(\out[1][2][18] ) );
  inv_x2_sg U12108 ( .A(n15815), .X(\out[1][2][17] ) );
  inv_x2_sg U12109 ( .A(n15817), .X(\out[1][2][16] ) );
  inv_x2_sg U12110 ( .A(n15819), .X(\out[1][2][15] ) );
  inv_x2_sg U12111 ( .A(n15821), .X(\out[1][2][14] ) );
  inv_x2_sg U12112 ( .A(n15823), .X(\out[1][2][13] ) );
  inv_x2_sg U12113 ( .A(n15825), .X(\out[1][2][12] ) );
  inv_x2_sg U12114 ( .A(n15827), .X(\out[1][2][11] ) );
  inv_x2_sg U12115 ( .A(n15829), .X(\out[1][2][10] ) );
  inv_x2_sg U12116 ( .A(n15831), .X(\out[1][2][9] ) );
  inv_x2_sg U12117 ( .A(n15833), .X(\out[1][2][8] ) );
  inv_x2_sg U12118 ( .A(n15835), .X(\out[1][2][7] ) );
  inv_x2_sg U12119 ( .A(n15837), .X(\out[1][2][6] ) );
  inv_x2_sg U12120 ( .A(n15839), .X(\out[1][2][5] ) );
  inv_x2_sg U12121 ( .A(n15841), .X(\out[1][2][4] ) );
  inv_x2_sg U12122 ( .A(n15843), .X(\out[1][2][3] ) );
  inv_x2_sg U12123 ( .A(n15845), .X(\out[1][2][2] ) );
  inv_x2_sg U12124 ( .A(n15847), .X(\out[1][2][1] ) );
  inv_x2_sg U12125 ( .A(n15849), .X(\out[1][2][0] ) );
  inv_x2_sg U12126 ( .A(n15851), .X(\out[1][1][19] ) );
  inv_x2_sg U12127 ( .A(n15853), .X(\out[1][1][18] ) );
  inv_x2_sg U12128 ( .A(n15855), .X(\out[1][1][17] ) );
  inv_x2_sg U12129 ( .A(n15857), .X(\out[1][1][16] ) );
  inv_x2_sg U12130 ( .A(n15859), .X(\out[1][1][15] ) );
  inv_x2_sg U12131 ( .A(n15861), .X(\out[1][1][14] ) );
  inv_x2_sg U12132 ( .A(n15863), .X(\out[1][1][13] ) );
  inv_x2_sg U12133 ( .A(n15865), .X(\out[1][1][12] ) );
  inv_x2_sg U12134 ( .A(n15867), .X(\out[1][1][11] ) );
  inv_x2_sg U12135 ( .A(n15869), .X(\out[1][1][10] ) );
  inv_x2_sg U12136 ( .A(n15871), .X(\out[1][1][9] ) );
  inv_x2_sg U12137 ( .A(n15873), .X(\out[1][1][8] ) );
  inv_x2_sg U12138 ( .A(n15875), .X(\out[1][1][7] ) );
  inv_x2_sg U12139 ( .A(n15877), .X(\out[1][1][6] ) );
  inv_x2_sg U12140 ( .A(n15879), .X(\out[1][1][5] ) );
  inv_x2_sg U12141 ( .A(n15881), .X(\out[1][1][4] ) );
  inv_x2_sg U12142 ( .A(n15883), .X(\out[1][1][3] ) );
  inv_x2_sg U12143 ( .A(n15885), .X(\out[1][1][2] ) );
  inv_x2_sg U12144 ( .A(n15887), .X(\out[1][1][1] ) );
  inv_x2_sg U12145 ( .A(n15889), .X(\out[1][1][0] ) );
  inv_x2_sg U12146 ( .A(n15891), .X(\out[1][0][19] ) );
  inv_x2_sg U12147 ( .A(n15893), .X(\out[1][0][18] ) );
  inv_x2_sg U12148 ( .A(n15895), .X(\out[1][0][17] ) );
  inv_x2_sg U12149 ( .A(n15897), .X(\out[1][0][16] ) );
  inv_x2_sg U12150 ( .A(n15899), .X(\out[1][0][15] ) );
  inv_x2_sg U12151 ( .A(n15901), .X(\out[1][0][14] ) );
  inv_x2_sg U12152 ( .A(n15903), .X(\out[1][0][13] ) );
  inv_x2_sg U12153 ( .A(n15905), .X(\out[1][0][12] ) );
  inv_x2_sg U12154 ( .A(n15907), .X(\out[1][0][11] ) );
  inv_x2_sg U12155 ( .A(n15909), .X(\out[1][0][10] ) );
  inv_x2_sg U12156 ( .A(n15911), .X(\out[1][0][9] ) );
  inv_x2_sg U12157 ( .A(n15913), .X(\out[1][0][8] ) );
  inv_x2_sg U12158 ( .A(n15915), .X(\out[1][0][7] ) );
  inv_x2_sg U12159 ( .A(n15917), .X(\out[1][0][6] ) );
  inv_x2_sg U12160 ( .A(n15919), .X(\out[1][0][5] ) );
  inv_x2_sg U12161 ( .A(n15921), .X(\out[1][0][4] ) );
  inv_x2_sg U12162 ( .A(n15923), .X(\out[1][0][3] ) );
  inv_x2_sg U12163 ( .A(n15925), .X(\out[1][0][2] ) );
  inv_x2_sg U12164 ( .A(n15927), .X(\out[1][0][1] ) );
  inv_x2_sg U12165 ( .A(n15929), .X(\out[1][0][0] ) );
  inv_x2_sg U12166 ( .A(n15931), .X(\out[0][3][19] ) );
  inv_x2_sg U12167 ( .A(n15933), .X(\out[0][3][18] ) );
  inv_x2_sg U12168 ( .A(n15935), .X(\out[0][3][17] ) );
  inv_x2_sg U12169 ( .A(n15937), .X(\out[0][3][16] ) );
  inv_x2_sg U12170 ( .A(n15939), .X(\out[0][3][15] ) );
  inv_x2_sg U12171 ( .A(n15941), .X(\out[0][3][14] ) );
  inv_x2_sg U12172 ( .A(n15943), .X(\out[0][3][13] ) );
  inv_x2_sg U12173 ( .A(n15945), .X(\out[0][3][12] ) );
  inv_x2_sg U12174 ( .A(n15947), .X(\out[0][3][11] ) );
  inv_x2_sg U12175 ( .A(n15949), .X(\out[0][3][10] ) );
  inv_x2_sg U12176 ( .A(n15951), .X(\out[0][3][9] ) );
  inv_x2_sg U12177 ( .A(n15953), .X(\out[0][3][8] ) );
  inv_x2_sg U12178 ( .A(n15955), .X(\out[0][3][7] ) );
  inv_x2_sg U12179 ( .A(n15957), .X(\out[0][3][6] ) );
  inv_x2_sg U12180 ( .A(n15959), .X(\out[0][3][5] ) );
  inv_x2_sg U12181 ( .A(n15961), .X(\out[0][3][4] ) );
  inv_x2_sg U12182 ( .A(n15963), .X(\out[0][3][3] ) );
  inv_x2_sg U12183 ( .A(n15965), .X(\out[0][3][2] ) );
  inv_x2_sg U12184 ( .A(n15967), .X(\out[0][3][1] ) );
  inv_x2_sg U12185 ( .A(n15969), .X(\out[0][3][0] ) );
  inv_x2_sg U12186 ( .A(n15971), .X(\out[0][2][19] ) );
  inv_x2_sg U12187 ( .A(n15973), .X(\out[0][2][18] ) );
  inv_x2_sg U12188 ( .A(n15975), .X(\out[0][2][17] ) );
  inv_x2_sg U12189 ( .A(n15977), .X(\out[0][2][16] ) );
  inv_x2_sg U12190 ( .A(n15979), .X(\out[0][2][15] ) );
  inv_x2_sg U12191 ( .A(n15981), .X(\out[0][2][14] ) );
  inv_x2_sg U12192 ( .A(n15983), .X(\out[0][2][13] ) );
  inv_x2_sg U12193 ( .A(n15985), .X(\out[0][2][12] ) );
  inv_x2_sg U12194 ( .A(n15987), .X(\out[0][2][11] ) );
  inv_x2_sg U12195 ( .A(n15989), .X(\out[0][2][10] ) );
  inv_x2_sg U12196 ( .A(n15991), .X(\out[0][2][9] ) );
  inv_x2_sg U12197 ( .A(n15993), .X(\out[0][2][8] ) );
  inv_x2_sg U12198 ( .A(n15995), .X(\out[0][2][7] ) );
  inv_x2_sg U12199 ( .A(n15997), .X(\out[0][2][6] ) );
  inv_x2_sg U12200 ( .A(n15999), .X(\out[0][2][5] ) );
  inv_x2_sg U12201 ( .A(n16001), .X(\out[0][2][4] ) );
  inv_x2_sg U12202 ( .A(n16003), .X(\out[0][2][3] ) );
  inv_x2_sg U12203 ( .A(n16005), .X(\out[0][2][2] ) );
  inv_x2_sg U12204 ( .A(n16007), .X(\out[0][2][1] ) );
  inv_x2_sg U12205 ( .A(n16009), .X(\out[0][2][0] ) );
  inv_x2_sg U12206 ( .A(n16011), .X(\out[0][1][19] ) );
  inv_x2_sg U12207 ( .A(n16013), .X(\out[0][1][18] ) );
  inv_x2_sg U12208 ( .A(n16015), .X(\out[0][1][17] ) );
  inv_x2_sg U12209 ( .A(n16017), .X(\out[0][1][16] ) );
  inv_x2_sg U12210 ( .A(n16019), .X(\out[0][1][15] ) );
  inv_x2_sg U12211 ( .A(n16021), .X(\out[0][1][14] ) );
  inv_x2_sg U12212 ( .A(n16023), .X(\out[0][1][13] ) );
  inv_x2_sg U12213 ( .A(n16025), .X(\out[0][1][12] ) );
  inv_x2_sg U12214 ( .A(n16027), .X(\out[0][1][11] ) );
  inv_x2_sg U12215 ( .A(n16029), .X(\out[0][1][10] ) );
  inv_x2_sg U12216 ( .A(n16031), .X(\out[0][1][9] ) );
  inv_x2_sg U12217 ( .A(n16033), .X(\out[0][1][8] ) );
  inv_x2_sg U12218 ( .A(n16035), .X(\out[0][1][7] ) );
  inv_x2_sg U12219 ( .A(n16037), .X(\out[0][1][6] ) );
  inv_x2_sg U12220 ( .A(n16039), .X(\out[0][1][5] ) );
  inv_x2_sg U12221 ( .A(n16041), .X(\out[0][1][4] ) );
  inv_x2_sg U12222 ( .A(n16043), .X(\out[0][1][3] ) );
  inv_x2_sg U12223 ( .A(n16045), .X(\out[0][1][2] ) );
  inv_x2_sg U12224 ( .A(n16047), .X(\out[0][1][1] ) );
  inv_x2_sg U12225 ( .A(n16049), .X(\out[0][1][0] ) );
  inv_x2_sg U12226 ( .A(n16051), .X(\out[0][0][19] ) );
  inv_x2_sg U12227 ( .A(n16053), .X(\out[0][0][18] ) );
  inv_x2_sg U12228 ( .A(n16055), .X(\out[0][0][17] ) );
  inv_x2_sg U12229 ( .A(n16057), .X(\out[0][0][16] ) );
  inv_x2_sg U12230 ( .A(n16059), .X(\out[0][0][15] ) );
  inv_x2_sg U12231 ( .A(n16061), .X(\out[0][0][14] ) );
  inv_x2_sg U12232 ( .A(n16063), .X(\out[0][0][13] ) );
  inv_x2_sg U12233 ( .A(n16065), .X(\out[0][0][12] ) );
  inv_x2_sg U12234 ( .A(n16067), .X(\out[0][0][11] ) );
  inv_x2_sg U12235 ( .A(n16069), .X(\out[0][0][10] ) );
  inv_x2_sg U12236 ( .A(n16071), .X(\out[0][0][9] ) );
  inv_x2_sg U12237 ( .A(n16073), .X(\out[0][0][8] ) );
  inv_x2_sg U12238 ( .A(n16075), .X(\out[0][0][7] ) );
  inv_x2_sg U12239 ( .A(n16077), .X(\out[0][0][6] ) );
  inv_x2_sg U12240 ( .A(n16079), .X(\out[0][0][5] ) );
  inv_x2_sg U12241 ( .A(n16081), .X(\out[0][0][4] ) );
  inv_x2_sg U12242 ( .A(n16083), .X(\out[0][0][3] ) );
  inv_x2_sg U12243 ( .A(n16085), .X(\out[0][0][2] ) );
  inv_x2_sg U12244 ( .A(n16087), .X(\out[0][0][1] ) );
  inv_x2_sg U12245 ( .A(n16089), .X(\out[0][0][0] ) );
  inv_x4_sg U12246 ( .A(n16091), .X(n16092) );
  inv_x4_sg U12247 ( .A(n16093), .X(n16094) );
  inv_x4_sg U12248 ( .A(n16095), .X(n16096) );
  inv_x4_sg U12249 ( .A(n16097), .X(n16098) );
  inv_x4_sg U12250 ( .A(n16099), .X(n16100) );
  inv_x4_sg U12251 ( .A(n16101), .X(n16102) );
  inv_x4_sg U12252 ( .A(n16103), .X(n16104) );
  inv_x4_sg U12253 ( .A(n16105), .X(n16106) );
  inv_x4_sg U12254 ( .A(n16107), .X(n16108) );
  inv_x4_sg U12255 ( .A(n16109), .X(n16110) );
  inv_x4_sg U12256 ( .A(n16111), .X(n16112) );
  inv_x4_sg U12257 ( .A(n16113), .X(n16114) );
  inv_x4_sg U12258 ( .A(n16115), .X(n16116) );
  inv_x4_sg U12259 ( .A(n16117), .X(n16118) );
  inv_x4_sg U12260 ( .A(n16119), .X(n16120) );
  inv_x4_sg U12261 ( .A(n16121), .X(n16122) );
  inv_x4_sg U12262 ( .A(n16123), .X(n16124) );
  inv_x4_sg U12263 ( .A(n16125), .X(n16126) );
  inv_x4_sg U12264 ( .A(n16127), .X(n16128) );
  inv_x4_sg U12265 ( .A(n16129), .X(n16130) );
  inv_x4_sg U12266 ( .A(n16131), .X(n16132) );
  inv_x4_sg U12267 ( .A(n16133), .X(n16134) );
  inv_x4_sg U12268 ( .A(n16135), .X(n16136) );
  inv_x4_sg U12269 ( .A(n16137), .X(n16138) );
  inv_x4_sg U12270 ( .A(n16139), .X(n16140) );
  inv_x4_sg U12271 ( .A(n16141), .X(n16142) );
  inv_x4_sg U12272 ( .A(n16143), .X(n16144) );
  inv_x4_sg U12273 ( .A(n16145), .X(n16146) );
  inv_x4_sg U12274 ( .A(n16147), .X(n16148) );
  inv_x4_sg U12275 ( .A(n16149), .X(n16150) );
  inv_x4_sg U12276 ( .A(n16151), .X(n16152) );
  inv_x4_sg U12277 ( .A(n16153), .X(n16154) );
  inv_x4_sg U12278 ( .A(n16155), .X(n16156) );
  inv_x4_sg U12279 ( .A(n16157), .X(n16158) );
  inv_x4_sg U12280 ( .A(n16159), .X(n16160) );
  inv_x4_sg U12281 ( .A(n16161), .X(n16162) );
  inv_x4_sg U12282 ( .A(n16163), .X(n16164) );
  inv_x4_sg U12283 ( .A(n16165), .X(n16166) );
  inv_x4_sg U12284 ( .A(n16167), .X(n16168) );
  inv_x4_sg U12285 ( .A(n16169), .X(n16170) );
  inv_x4_sg U12286 ( .A(n16171), .X(n16172) );
  inv_x4_sg U12287 ( .A(n16173), .X(n16174) );
  inv_x4_sg U12288 ( .A(n16175), .X(n16176) );
  inv_x4_sg U12289 ( .A(n16177), .X(n16178) );
  inv_x4_sg U12290 ( .A(n16179), .X(n16180) );
  inv_x4_sg U12291 ( .A(n16181), .X(n16182) );
  inv_x4_sg U12292 ( .A(n16183), .X(n16184) );
  inv_x4_sg U12293 ( .A(n16185), .X(n16186) );
  inv_x4_sg U12294 ( .A(n16187), .X(n16188) );
  inv_x4_sg U12295 ( .A(n16189), .X(n16190) );
  inv_x4_sg U12296 ( .A(n16191), .X(n16192) );
  inv_x4_sg U12297 ( .A(n16193), .X(n16194) );
  inv_x4_sg U12298 ( .A(n16195), .X(n16196) );
  inv_x4_sg U12299 ( .A(n16197), .X(n16198) );
  inv_x4_sg U12300 ( .A(n16199), .X(n16200) );
  inv_x4_sg U12301 ( .A(n16201), .X(n16202) );
  inv_x4_sg U12302 ( .A(n16203), .X(n16204) );
  inv_x4_sg U12303 ( .A(n16205), .X(n16206) );
  inv_x4_sg U12304 ( .A(n16207), .X(n16208) );
  inv_x4_sg U12305 ( .A(n16209), .X(n16210) );
  inv_x4_sg U12306 ( .A(n16211), .X(n16212) );
  inv_x4_sg U12307 ( .A(n16213), .X(n16214) );
  inv_x4_sg U12308 ( .A(n16215), .X(n16216) );
  inv_x4_sg U12309 ( .A(n16217), .X(n16218) );
  inv_x4_sg U12310 ( .A(n16219), .X(n16220) );
  inv_x4_sg U12311 ( .A(n16221), .X(n16222) );
  inv_x4_sg U12312 ( .A(n16223), .X(n16224) );
  inv_x4_sg U12313 ( .A(n16225), .X(n16226) );
  inv_x4_sg U12314 ( .A(n16227), .X(n16228) );
  inv_x4_sg U12315 ( .A(n16229), .X(n16230) );
  inv_x4_sg U12316 ( .A(n16231), .X(n16232) );
  inv_x4_sg U12317 ( .A(n16233), .X(n16234) );
  inv_x4_sg U12318 ( .A(n16235), .X(n16236) );
  inv_x4_sg U12319 ( .A(n16237), .X(n16238) );
  inv_x4_sg U12320 ( .A(n16239), .X(n16240) );
  inv_x4_sg U12321 ( .A(n16241), .X(n16242) );
  inv_x4_sg U12322 ( .A(n16243), .X(n16244) );
  inv_x4_sg U12323 ( .A(n16245), .X(n16246) );
  inv_x4_sg U12324 ( .A(n16247), .X(n16248) );
  inv_x4_sg U12325 ( .A(n16249), .X(n16250) );
  inv_x4_sg U12326 ( .A(n16251), .X(n16252) );
  inv_x4_sg U12327 ( .A(n16253), .X(n16254) );
  inv_x4_sg U12328 ( .A(n16255), .X(n16256) );
  inv_x4_sg U12329 ( .A(n16257), .X(n16258) );
  inv_x4_sg U12330 ( .A(n16259), .X(n16260) );
  inv_x4_sg U12331 ( .A(n16261), .X(n16262) );
  inv_x4_sg U12332 ( .A(n16263), .X(n16264) );
  inv_x4_sg U12333 ( .A(n16265), .X(n16266) );
  inv_x4_sg U12334 ( .A(n16267), .X(n16268) );
  inv_x4_sg U12335 ( .A(n16269), .X(n16270) );
  inv_x4_sg U12336 ( .A(n16271), .X(n16272) );
  inv_x4_sg U12337 ( .A(n16273), .X(n16274) );
  inv_x4_sg U12338 ( .A(n16275), .X(n16276) );
  inv_x4_sg U12339 ( .A(n16277), .X(n16278) );
  inv_x4_sg U12340 ( .A(n16279), .X(n16280) );
  inv_x4_sg U12341 ( .A(n16281), .X(n16282) );
  inv_x4_sg U12342 ( .A(n16283), .X(n16284) );
  inv_x4_sg U12343 ( .A(n16285), .X(n16286) );
  inv_x4_sg U12344 ( .A(n16287), .X(n16288) );
  inv_x4_sg U12345 ( .A(n16289), .X(n16290) );
  inv_x4_sg U12346 ( .A(n16291), .X(n16292) );
  inv_x4_sg U12347 ( .A(n16293), .X(n16294) );
  inv_x4_sg U12348 ( .A(n16295), .X(n16296) );
  inv_x4_sg U12349 ( .A(n16297), .X(n16298) );
  inv_x4_sg U12350 ( .A(n16299), .X(n16300) );
  inv_x4_sg U12351 ( .A(n16301), .X(n16302) );
  inv_x4_sg U12352 ( .A(n16303), .X(n16304) );
  inv_x4_sg U12353 ( .A(n16305), .X(n16306) );
  inv_x4_sg U12354 ( .A(n16307), .X(n16308) );
  inv_x4_sg U12355 ( .A(n16309), .X(n16310) );
  inv_x4_sg U12356 ( .A(n16311), .X(n16312) );
  inv_x4_sg U12357 ( .A(n16313), .X(n16314) );
  inv_x4_sg U12358 ( .A(n16315), .X(n16316) );
  inv_x4_sg U12359 ( .A(n16317), .X(n16318) );
  inv_x4_sg U12360 ( .A(n16319), .X(n16320) );
  inv_x4_sg U12361 ( .A(n16321), .X(n16322) );
  inv_x4_sg U12362 ( .A(n16323), .X(n16324) );
  inv_x4_sg U12363 ( .A(n16325), .X(n16326) );
  inv_x4_sg U12364 ( .A(n16327), .X(n16328) );
  inv_x4_sg U12365 ( .A(n16329), .X(n16330) );
  inv_x4_sg U12366 ( .A(n16331), .X(n16332) );
  inv_x4_sg U12367 ( .A(n16333), .X(n16334) );
  inv_x4_sg U12368 ( .A(n16335), .X(n16336) );
  inv_x4_sg U12369 ( .A(n16337), .X(n16338) );
  inv_x4_sg U12370 ( .A(n16339), .X(n16340) );
  inv_x4_sg U12371 ( .A(n16341), .X(n16342) );
  inv_x4_sg U12372 ( .A(n16343), .X(n16344) );
  inv_x4_sg U12373 ( .A(n16345), .X(n16346) );
  inv_x4_sg U12374 ( .A(n16347), .X(n16348) );
  inv_x4_sg U12375 ( .A(n16349), .X(n16350) );
  inv_x4_sg U12376 ( .A(n16351), .X(n16352) );
  inv_x4_sg U12377 ( .A(n16353), .X(n16354) );
  inv_x4_sg U12378 ( .A(n16355), .X(n16356) );
  inv_x4_sg U12379 ( .A(n16357), .X(n16358) );
  inv_x4_sg U12380 ( .A(n16359), .X(n16360) );
  inv_x4_sg U12381 ( .A(n16361), .X(n16362) );
  inv_x4_sg U12382 ( .A(n16363), .X(n16364) );
  inv_x4_sg U12383 ( .A(n16365), .X(n16366) );
  inv_x4_sg U12384 ( .A(n16367), .X(n16368) );
  inv_x4_sg U12385 ( .A(n16369), .X(n16370) );
  inv_x4_sg U12386 ( .A(n16371), .X(n16372) );
  inv_x4_sg U12387 ( .A(n16373), .X(n16374) );
  inv_x4_sg U12388 ( .A(n16375), .X(n16376) );
  inv_x4_sg U12389 ( .A(n16377), .X(n16378) );
  inv_x4_sg U12390 ( .A(n16379), .X(n16380) );
  inv_x4_sg U12391 ( .A(n16381), .X(n16382) );
  inv_x4_sg U12392 ( .A(n16383), .X(n16384) );
  inv_x4_sg U12393 ( .A(n16385), .X(n16386) );
  inv_x4_sg U12394 ( .A(n16387), .X(n16388) );
  inv_x4_sg U12395 ( .A(n16389), .X(n16390) );
  inv_x4_sg U12396 ( .A(n16391), .X(n16392) );
  inv_x4_sg U12397 ( .A(n16393), .X(n16394) );
  inv_x4_sg U12398 ( .A(n16395), .X(n16396) );
  inv_x4_sg U12399 ( .A(n16397), .X(n16398) );
  inv_x4_sg U12400 ( .A(n16399), .X(n16400) );
  inv_x4_sg U12401 ( .A(n16401), .X(n16402) );
  inv_x4_sg U12402 ( .A(n16403), .X(n16404) );
  inv_x4_sg U12403 ( .A(n16405), .X(n16406) );
  inv_x4_sg U12404 ( .A(n16407), .X(n16408) );
  inv_x4_sg U12405 ( .A(n16409), .X(n16410) );
  inv_x4_sg U12406 ( .A(n16411), .X(n16412) );
  inv_x4_sg U12407 ( .A(n16413), .X(n16414) );
  inv_x4_sg U12408 ( .A(n16415), .X(n16416) );
  inv_x4_sg U12409 ( .A(n16417), .X(n16418) );
  inv_x4_sg U12410 ( .A(n16419), .X(n16420) );
  inv_x4_sg U12411 ( .A(n16421), .X(n16422) );
  inv_x4_sg U12412 ( .A(n16423), .X(n16424) );
  inv_x4_sg U12413 ( .A(n16425), .X(n16426) );
  inv_x4_sg U12414 ( .A(n16427), .X(n16428) );
  inv_x4_sg U12415 ( .A(n16429), .X(n16430) );
  inv_x4_sg U12416 ( .A(n16431), .X(n16432) );
  inv_x4_sg U12417 ( .A(n16433), .X(n16434) );
  inv_x4_sg U12418 ( .A(n16435), .X(n16436) );
  inv_x4_sg U12419 ( .A(n16437), .X(n16438) );
  inv_x4_sg U12420 ( .A(n16439), .X(n16440) );
  inv_x4_sg U12421 ( .A(n16441), .X(n16442) );
  inv_x4_sg U12422 ( .A(n16443), .X(n16444) );
  inv_x4_sg U12423 ( .A(n16445), .X(n16446) );
  inv_x4_sg U12424 ( .A(n16447), .X(n16448) );
  inv_x4_sg U12425 ( .A(n16449), .X(n16450) );
  inv_x4_sg U12426 ( .A(n16451), .X(n16452) );
  inv_x4_sg U12427 ( .A(n16453), .X(n16454) );
  inv_x4_sg U12428 ( .A(n16455), .X(n16456) );
  inv_x4_sg U12429 ( .A(n16457), .X(n16458) );
  inv_x4_sg U12430 ( .A(n16459), .X(n16460) );
  inv_x4_sg U12431 ( .A(n16461), .X(n16462) );
  inv_x4_sg U12432 ( .A(n16463), .X(n16464) );
  inv_x4_sg U12433 ( .A(n16465), .X(n16466) );
  inv_x4_sg U12434 ( .A(n16467), .X(n16468) );
  inv_x4_sg U12435 ( .A(n16469), .X(n16470) );
  inv_x4_sg U12436 ( .A(n16471), .X(n16472) );
  inv_x4_sg U12437 ( .A(n16473), .X(n16474) );
  inv_x4_sg U12438 ( .A(n16475), .X(n16476) );
  inv_x4_sg U12439 ( .A(n16477), .X(n16478) );
  inv_x4_sg U12440 ( .A(n16479), .X(n16480) );
  inv_x4_sg U12441 ( .A(n16481), .X(n16482) );
  inv_x4_sg U12442 ( .A(n16483), .X(n16484) );
  inv_x4_sg U12443 ( .A(n16485), .X(n16486) );
  inv_x4_sg U12444 ( .A(n16487), .X(n16488) );
  inv_x4_sg U12445 ( .A(n16489), .X(n16490) );
  inv_x4_sg U12446 ( .A(n16491), .X(n16492) );
  inv_x4_sg U12447 ( .A(n16493), .X(n16494) );
  inv_x4_sg U12448 ( .A(n16495), .X(n16496) );
  inv_x4_sg U12449 ( .A(n16497), .X(n16498) );
  inv_x4_sg U12450 ( .A(n16499), .X(n16500) );
  inv_x4_sg U12451 ( .A(n16501), .X(n16502) );
  inv_x4_sg U12452 ( .A(n16503), .X(n16504) );
  inv_x4_sg U12453 ( .A(n16505), .X(n16506) );
  inv_x4_sg U12454 ( .A(n16507), .X(n16508) );
  inv_x4_sg U12455 ( .A(n16509), .X(n16510) );
  inv_x4_sg U12456 ( .A(n16511), .X(n16512) );
  inv_x4_sg U12457 ( .A(n16513), .X(n16514) );
  inv_x4_sg U12458 ( .A(n16515), .X(n16516) );
  inv_x4_sg U12459 ( .A(n16517), .X(n16518) );
  inv_x4_sg U12460 ( .A(n16519), .X(n16520) );
  inv_x4_sg U12461 ( .A(n16521), .X(n16522) );
  inv_x4_sg U12462 ( .A(n16523), .X(n16524) );
  inv_x4_sg U12463 ( .A(n16525), .X(n16526) );
  inv_x4_sg U12464 ( .A(n16527), .X(n16528) );
  inv_x4_sg U12465 ( .A(n16529), .X(n16530) );
  inv_x4_sg U12466 ( .A(n16531), .X(n16532) );
  inv_x4_sg U12467 ( .A(n16533), .X(n16534) );
  inv_x4_sg U12468 ( .A(n16535), .X(n16536) );
  inv_x4_sg U12469 ( .A(n16537), .X(n16538) );
  inv_x4_sg U12470 ( .A(n16539), .X(n16540) );
  inv_x4_sg U12471 ( .A(n16541), .X(n16542) );
  inv_x4_sg U12472 ( .A(n16543), .X(n16544) );
  inv_x4_sg U12473 ( .A(n16545), .X(n16546) );
  inv_x4_sg U12474 ( .A(n16547), .X(n16548) );
  inv_x4_sg U12475 ( .A(n16549), .X(n16550) );
  inv_x4_sg U12476 ( .A(n16551), .X(n16552) );
  inv_x4_sg U12477 ( .A(n16553), .X(n16554) );
  inv_x4_sg U12478 ( .A(n16555), .X(n16556) );
  inv_x4_sg U12479 ( .A(n16557), .X(n16558) );
  inv_x4_sg U12480 ( .A(n16559), .X(n16560) );
  inv_x4_sg U12481 ( .A(n16561), .X(n16562) );
  inv_x4_sg U12482 ( .A(n16563), .X(n16564) );
  inv_x4_sg U12483 ( .A(n16565), .X(n16566) );
  inv_x4_sg U12484 ( .A(n16567), .X(n16568) );
  inv_x4_sg U12485 ( .A(n16569), .X(n16570) );
  inv_x4_sg U12486 ( .A(n16571), .X(n16572) );
  inv_x4_sg U12487 ( .A(n16573), .X(n16574) );
  inv_x4_sg U12488 ( .A(n16575), .X(n16576) );
  inv_x4_sg U12489 ( .A(n16577), .X(n16578) );
  inv_x4_sg U12490 ( .A(n16579), .X(n16580) );
  inv_x4_sg U12491 ( .A(n16581), .X(n16582) );
  inv_x4_sg U12492 ( .A(n16583), .X(n16584) );
  inv_x4_sg U12493 ( .A(n16585), .X(n16586) );
  inv_x4_sg U12494 ( .A(n16587), .X(n16588) );
  inv_x4_sg U12495 ( .A(n16589), .X(n16590) );
  inv_x4_sg U12496 ( .A(n16591), .X(n16592) );
  inv_x4_sg U12497 ( .A(n16593), .X(n16594) );
  inv_x4_sg U12498 ( .A(n16595), .X(n16596) );
  inv_x4_sg U12499 ( .A(n16597), .X(n16598) );
  inv_x4_sg U12500 ( .A(n16599), .X(n16600) );
  inv_x4_sg U12501 ( .A(n16601), .X(n16602) );
  inv_x4_sg U12502 ( .A(n16603), .X(n16604) );
  inv_x4_sg U12503 ( .A(n16605), .X(n16606) );
  inv_x4_sg U12504 ( .A(n16607), .X(n16608) );
  inv_x4_sg U12505 ( .A(n16609), .X(n16610) );
  inv_x4_sg U12506 ( .A(n16611), .X(n16612) );
  inv_x4_sg U12507 ( .A(n16613), .X(n16614) );
  inv_x4_sg U12508 ( .A(n16615), .X(n16616) );
  inv_x4_sg U12509 ( .A(n16617), .X(n16618) );
  inv_x4_sg U12510 ( .A(n16619), .X(n16620) );
  inv_x4_sg U12511 ( .A(n16621), .X(n16622) );
  inv_x4_sg U12512 ( .A(n16623), .X(n16624) );
  inv_x4_sg U12513 ( .A(n16625), .X(n16626) );
  inv_x4_sg U12514 ( .A(n16627), .X(n16628) );
  inv_x4_sg U12515 ( .A(n16629), .X(n16630) );
  inv_x4_sg U12516 ( .A(n16631), .X(n16632) );
  inv_x4_sg U12517 ( .A(n16633), .X(n16634) );
  inv_x4_sg U12518 ( .A(n16635), .X(n16636) );
  inv_x4_sg U12519 ( .A(n16637), .X(n16638) );
  inv_x4_sg U12520 ( .A(n16639), .X(n16640) );
  inv_x4_sg U12521 ( .A(n16641), .X(n16642) );
  inv_x4_sg U12522 ( .A(n16643), .X(n16644) );
  inv_x4_sg U12523 ( .A(n16645), .X(n16646) );
  inv_x4_sg U12524 ( .A(n16647), .X(n16648) );
  inv_x4_sg U12525 ( .A(n16649), .X(n16650) );
  inv_x4_sg U12526 ( .A(n16651), .X(n16652) );
  inv_x4_sg U12527 ( .A(n16653), .X(n16654) );
  inv_x4_sg U12528 ( .A(n16655), .X(n16656) );
  inv_x4_sg U12529 ( .A(n16657), .X(n16658) );
  inv_x4_sg U12530 ( .A(n16659), .X(n16660) );
  inv_x4_sg U12531 ( .A(n16661), .X(n16662) );
  inv_x4_sg U12532 ( .A(n16663), .X(n16664) );
  inv_x4_sg U12533 ( .A(n16665), .X(n16666) );
  inv_x4_sg U12534 ( .A(n16667), .X(n16668) );
  inv_x4_sg U12535 ( .A(n16669), .X(n16670) );
  inv_x4_sg U12536 ( .A(n16671), .X(n16672) );
  inv_x4_sg U12537 ( .A(n16673), .X(n16674) );
  inv_x4_sg U12538 ( .A(n16675), .X(n16676) );
  inv_x4_sg U12539 ( .A(n16677), .X(n16678) );
  inv_x4_sg U12540 ( .A(n16679), .X(n16680) );
  inv_x4_sg U12541 ( .A(n16681), .X(n16682) );
  inv_x4_sg U12542 ( .A(n16683), .X(n16684) );
  inv_x4_sg U12543 ( .A(n16685), .X(n16686) );
  inv_x4_sg U12544 ( .A(n16687), .X(n16688) );
  inv_x4_sg U12545 ( .A(n16689), .X(n16690) );
  inv_x4_sg U12546 ( .A(n16691), .X(n16692) );
  inv_x4_sg U12547 ( .A(n16693), .X(n16694) );
  inv_x4_sg U12548 ( .A(n16695), .X(n16696) );
  inv_x4_sg U12549 ( .A(n16697), .X(n16698) );
  inv_x4_sg U12550 ( .A(n16699), .X(n16700) );
  inv_x4_sg U12551 ( .A(n16701), .X(n16702) );
  inv_x4_sg U12552 ( .A(n16703), .X(n16704) );
  inv_x4_sg U12553 ( .A(n16705), .X(n16706) );
  inv_x4_sg U12554 ( .A(n16707), .X(n16708) );
  inv_x4_sg U12555 ( .A(n16709), .X(n16710) );
  inv_x4_sg U12556 ( .A(n16711), .X(n16712) );
  inv_x4_sg U12557 ( .A(n16713), .X(n16714) );
  inv_x4_sg U12558 ( .A(n16715), .X(n16716) );
  inv_x4_sg U12559 ( .A(n16717), .X(n16718) );
  inv_x4_sg U12560 ( .A(n16719), .X(n16720) );
  inv_x4_sg U12561 ( .A(n16721), .X(n16722) );
  inv_x4_sg U12562 ( .A(n16723), .X(n16724) );
  inv_x4_sg U12563 ( .A(n16725), .X(n16726) );
  inv_x4_sg U12564 ( .A(n16727), .X(n16728) );
  inv_x4_sg U12565 ( .A(n16729), .X(n16730) );
  inv_x4_sg U12566 ( .A(n15448), .X(n16731) );
  inv_x8_sg U12567 ( .A(n16731), .X(state[0]) );
  nand_x2_sg U12568 ( .A(n16731), .B(n18399), .X(n14471) );
  nand_x1_sg U12569 ( .A(\out[0][3][4] ), .B(n16793), .X(n13379) );
  nand_x1_sg U12570 ( .A(\out[0][3][5] ), .B(n16785), .X(n13381) );
  nand_x1_sg U12571 ( .A(\out[0][3][6] ), .B(n16793), .X(n13373) );
  nand_x1_sg U12572 ( .A(\out[0][3][7] ), .B(n16793), .X(n13375) );
  nand_x1_sg U12573 ( .A(\out[0][3][8] ), .B(n16791), .X(n13391) );
  nand_x1_sg U12574 ( .A(\out[0][3][9] ), .B(n16789), .X(n13393) );
  nand_x1_sg U12575 ( .A(\out[0][3][10] ), .B(n16790), .X(n13385) );
  nand_x1_sg U12576 ( .A(\out[0][3][11] ), .B(n16788), .X(n13387) );
  nand_x1_sg U12577 ( .A(\out[0][3][12] ), .B(n16793), .X(n13355) );
  nand_x1_sg U12578 ( .A(\out[0][3][13] ), .B(n16793), .X(n13357) );
  nand_x1_sg U12579 ( .A(\out[0][3][14] ), .B(n16793), .X(n13349) );
  nand_x1_sg U12580 ( .A(\out[0][3][15] ), .B(n16793), .X(n13351) );
  nand_x1_sg U12581 ( .A(\out[0][3][16] ), .B(n16793), .X(n13367) );
  nand_x1_sg U12582 ( .A(\out[0][3][17] ), .B(n16793), .X(n13369) );
  nand_x1_sg U12583 ( .A(\out[0][3][18] ), .B(n16793), .X(n13361) );
  nand_x1_sg U12584 ( .A(\out[0][3][19] ), .B(n16793), .X(n13363) );
  nand_x1_sg U12585 ( .A(\out[1][0][0] ), .B(n16791), .X(n13427) );
  nand_x1_sg U12586 ( .A(\out[1][0][1] ), .B(n16785), .X(n13429) );
  nand_x1_sg U12587 ( .A(\out[1][0][2] ), .B(n16793), .X(n13421) );
  nand_x1_sg U12588 ( .A(\out[1][0][3] ), .B(n16789), .X(n13423) );
  nand_x1_sg U12589 ( .A(\out[1][0][4] ), .B(n16793), .X(n13439) );
  nand_x1_sg U12590 ( .A(\out[1][0][5] ), .B(n16786), .X(n13441) );
  nand_x1_sg U12591 ( .A(\out[1][0][6] ), .B(n16786), .X(n13433) );
  nand_x1_sg U12592 ( .A(\out[1][0][7] ), .B(n16793), .X(n13435) );
  nand_x1_sg U12593 ( .A(\out[1][0][8] ), .B(n16785), .X(n13403) );
  nand_x1_sg U12594 ( .A(\out[1][0][9] ), .B(n16784), .X(n13405) );
  nand_x1_sg U12595 ( .A(\out[1][0][10] ), .B(n16786), .X(n13397) );
  nand_x1_sg U12596 ( .A(\out[1][0][11] ), .B(n16784), .X(n13399) );
  nand_x1_sg U12597 ( .A(\out[1][0][12] ), .B(n16790), .X(n13415) );
  nand_x1_sg U12598 ( .A(\out[1][0][13] ), .B(n16788), .X(n13417) );
  nand_x1_sg U12599 ( .A(\out[1][0][14] ), .B(n16783), .X(n13409) );
  nand_x1_sg U12600 ( .A(\out[1][0][15] ), .B(n16783), .X(n13411) );
  nand_x1_sg U12601 ( .A(\out[1][1][12] ), .B(n16785), .X(n13331) );
  nand_x1_sg U12602 ( .A(\out[1][1][13] ), .B(n16793), .X(n13333) );
  nand_x1_sg U12603 ( .A(\out[1][1][14] ), .B(n16786), .X(n13325) );
  nand_x1_sg U12604 ( .A(\out[1][1][15] ), .B(n16784), .X(n13327) );
  nand_x1_sg U12605 ( .A(\out[1][1][16] ), .B(n16793), .X(n13343) );
  nand_x1_sg U12606 ( .A(\out[1][1][17] ), .B(n16793), .X(n13345) );
  nand_x1_sg U12607 ( .A(\out[1][1][18] ), .B(n16793), .X(n13337) );
  nand_x1_sg U12608 ( .A(\out[1][1][19] ), .B(n16793), .X(n13339) );
  nand_x1_sg U12609 ( .A(\out[1][2][4] ), .B(n16785), .X(n13319) );
  nand_x1_sg U12610 ( .A(\out[1][2][5] ), .B(n16786), .X(n13321) );
  nand_x1_sg U12611 ( .A(\out[1][2][8] ), .B(n16788), .X(n13571) );
  nand_x1_sg U12612 ( .A(\out[1][2][10] ), .B(n16784), .X(n13565) );
  nand_x1_sg U12613 ( .A(\out[1][2][11] ), .B(n16785), .X(n13567) );
  nand_x1_sg U12614 ( .A(\out[1][2][16] ), .B(n16786), .X(n13547) );
  nand_x1_sg U12615 ( .A(\out[1][2][17] ), .B(n16793), .X(n13549) );
  nand_x1_sg U12616 ( .A(\out[1][2][18] ), .B(n16786), .X(n13541) );
  nand_x1_sg U12617 ( .A(\out[1][2][19] ), .B(n16793), .X(n13543) );
  nand_x1_sg U12618 ( .A(\out[1][3][0] ), .B(n16786), .X(n13559) );
  nand_x1_sg U12619 ( .A(\out[1][3][1] ), .B(n16790), .X(n13561) );
  nand_x1_sg U12620 ( .A(\out[1][3][2] ), .B(n16790), .X(n13553) );
  nand_x1_sg U12621 ( .A(\out[1][3][3] ), .B(n16793), .X(n13555) );
  nand_x1_sg U12622 ( .A(\out[2][0][0] ), .B(n16793), .X(n13475) );
  nand_x1_sg U12623 ( .A(\out[2][0][1] ), .B(n16791), .X(n13477) );
  nand_x1_sg U12624 ( .A(\out[2][0][2] ), .B(n16791), .X(n13469) );
  nand_x1_sg U12625 ( .A(\out[2][0][3] ), .B(n16790), .X(n13471) );
  nand_x1_sg U12626 ( .A(\out[2][0][4] ), .B(n16789), .X(n13487) );
  nand_x1_sg U12627 ( .A(\out[2][0][5] ), .B(n16786), .X(n13489) );
  nand_x1_sg U12628 ( .A(\out[2][0][6] ), .B(n16789), .X(n13481) );
  nand_x1_sg U12629 ( .A(\out[2][0][7] ), .B(n16791), .X(n13483) );
  nand_x1_sg U12630 ( .A(\out[2][0][8] ), .B(n16788), .X(n13451) );
  nand_x1_sg U12631 ( .A(\out[2][0][9] ), .B(n16789), .X(n13453) );
  nand_x1_sg U12632 ( .A(\out[2][0][10] ), .B(n16791), .X(n13445) );
  nand_x1_sg U12633 ( .A(\out[2][0][11] ), .B(n16793), .X(n13447) );
  nand_x1_sg U12634 ( .A(\out[2][0][12] ), .B(n16788), .X(n13463) );
  nand_x1_sg U12635 ( .A(\out[2][0][13] ), .B(n16791), .X(n13465) );
  nand_x1_sg U12636 ( .A(\out[2][0][14] ), .B(n16785), .X(n13457) );
  nand_x1_sg U12637 ( .A(\out[2][0][15] ), .B(n16793), .X(n13459) );
  nand_x1_sg U12638 ( .A(\out[2][0][16] ), .B(n16788), .X(n13523) );
  nand_x1_sg U12639 ( .A(\out[2][0][17] ), .B(n16788), .X(n13525) );
  nand_x1_sg U12640 ( .A(\out[2][0][18] ), .B(n16789), .X(n13517) );
  nand_x1_sg U12641 ( .A(\out[2][0][19] ), .B(n16793), .X(n13519) );
  nand_x1_sg U12642 ( .A(\out[2][1][0] ), .B(n16783), .X(n13535) );
  nand_x1_sg U12643 ( .A(\out[2][1][1] ), .B(n16783), .X(n13537) );
  nand_x1_sg U12644 ( .A(\out[2][1][2] ), .B(n16784), .X(n13529) );
  nand_x1_sg U12645 ( .A(\out[2][1][3] ), .B(n16785), .X(n13531) );
  nand_x1_sg U12646 ( .A(\out[2][1][4] ), .B(n16785), .X(n13499) );
  nand_x1_sg U12647 ( .A(\out[2][1][5] ), .B(n16784), .X(n13501) );
  nand_x1_sg U12648 ( .A(\out[2][1][6] ), .B(n16790), .X(n13493) );
  nand_x1_sg U12649 ( .A(\out[2][1][7] ), .B(n16791), .X(n13495) );
  nand_x1_sg U12650 ( .A(\out[2][1][8] ), .B(n16793), .X(n13511) );
  nand_x1_sg U12651 ( .A(\out[2][1][9] ), .B(n16784), .X(n13513) );
  nand_x1_sg U12652 ( .A(\out[2][1][10] ), .B(n16789), .X(n13505) );
  nand_x1_sg U12653 ( .A(\out[2][1][11] ), .B(n16784), .X(n13507) );
  nand_x1_sg U12654 ( .A(\out[2][1][14] ), .B(n16793), .X(n13323) );
  nand_x1_sg U12655 ( .A(\out[2][1][18] ), .B(n16793), .X(n13347) );
  nand_x1_sg U12656 ( .A(\out[2][1][19] ), .B(n16793), .X(n13377) );
  nand_x1_sg U12657 ( .A(\out[2][2][0] ), .B(n16783), .X(n13479) );
  nand_x1_sg U12658 ( .A(\out[2][2][3] ), .B(n16784), .X(n13557) );
  nand_x1_sg U12659 ( .A(\out[2][2][8] ), .B(n16785), .X(n13401) );
  nand_x1_sg U12660 ( .A(\out[2][2][9] ), .B(n16793), .X(n13395) );
  nand_x1_sg U12661 ( .A(\out[2][2][11] ), .B(n16793), .X(n13365) );
  nand_x1_sg U12662 ( .A(\out[2][2][14] ), .B(n16783), .X(n13329) );
  nand_x1_sg U12663 ( .A(\out[2][3][4] ), .B(n16790), .X(n13515) );
  nand_x1_sg U12664 ( .A(\out[2][3][16] ), .B(n16789), .X(n13461) );
  nand_x1_sg U12665 ( .A(\out[2][3][17] ), .B(n16789), .X(n13497) );
  nand_x1_sg U12666 ( .A(\out[2][3][19] ), .B(n16793), .X(n13431) );
  nand_x1_sg U12667 ( .A(\out[3][0][16] ), .B(n16791), .X(n13503) );
  nand_x1_sg U12668 ( .A(\out[3][0][17] ), .B(n16793), .X(n13509) );
  nand_x1_sg U12669 ( .A(\out[3][1][0] ), .B(n16783), .X(n13521) );
  nand_x1_sg U12670 ( .A(\out[3][1][1] ), .B(n16786), .X(n13527) );
  nand_x1_sg U12671 ( .A(\out[3][1][2] ), .B(n16793), .X(n13533) );
  nand_x1_sg U12672 ( .A(\out[3][1][3] ), .B(n16783), .X(n13539) );
  nand_x1_sg U12673 ( .A(\out[3][1][4] ), .B(n16793), .X(n13467) );
  nand_x1_sg U12674 ( .A(\out[3][1][5] ), .B(n16788), .X(n13473) );
  nand_x1_sg U12675 ( .A(\out[3][1][6] ), .B(n16788), .X(n13485) );
  nand_x1_sg U12676 ( .A(\out[3][1][7] ), .B(n16790), .X(n13491) );
  nand_x1_sg U12677 ( .A(\out[3][1][8] ), .B(n16793), .X(n13437) );
  nand_x1_sg U12678 ( .A(\out[3][1][9] ), .B(n16793), .X(n13443) );
  nand_x1_sg U12679 ( .A(\out[3][1][10] ), .B(n16793), .X(n13449) );
  nand_x1_sg U12680 ( .A(\out[3][1][11] ), .B(n16789), .X(n13455) );
  nand_x1_sg U12681 ( .A(\out[3][2][0] ), .B(n16793), .X(n13545) );
  nand_x1_sg U12682 ( .A(\out[3][2][1] ), .B(n16793), .X(n13551) );
  nand_x1_sg U12683 ( .A(\out[3][2][2] ), .B(n16783), .X(n13563) );
  nand_x1_sg U12684 ( .A(\out[3][2][3] ), .B(n16790), .X(n13569) );
  nand_x1_sg U12685 ( .A(\out[3][3][4] ), .B(n16793), .X(n13383) );
  nand_x1_sg U12686 ( .A(\out[3][3][5] ), .B(n16793), .X(n13389) );
  nand_x1_sg U12687 ( .A(\out[3][3][6] ), .B(n16784), .X(n13407) );
  nand_x1_sg U12688 ( .A(\out[3][3][7] ), .B(n16793), .X(n13413) );
  nand_x1_sg U12689 ( .A(\out[3][3][8] ), .B(n16793), .X(n13353) );
  nand_x1_sg U12690 ( .A(\out[3][3][9] ), .B(n16793), .X(n13359) );
  nand_x1_sg U12691 ( .A(\out[3][3][10] ), .B(n16793), .X(n13419) );
  nand_x1_sg U12692 ( .A(\out[3][3][11] ), .B(n16782), .X(n13371) );
  nand_x1_sg U12693 ( .A(\out[3][3][15] ), .B(n16789), .X(n13317) );
  nand_x1_sg U12694 ( .A(\out[3][3][16] ), .B(n16793), .X(n13335) );
  nand_x1_sg U12695 ( .A(\out[3][3][17] ), .B(n16793), .X(n13341) );
  nand_x1_sg U12696 ( .A(\out[3][3][19] ), .B(n16783), .X(n13425) );
  nand_x1_sg U12697 ( .A(\out[0][0][0] ), .B(n16781), .X(n13765) );
  nand_x1_sg U12698 ( .A(\out[0][0][1] ), .B(n16790), .X(n13767) );
  nand_x1_sg U12699 ( .A(\out[0][0][2] ), .B(n16785), .X(n13759) );
  nand_x1_sg U12700 ( .A(\out[0][0][3] ), .B(n16784), .X(n13761) );
  nand_x1_sg U12701 ( .A(\out[0][0][4] ), .B(n16780), .X(n13777) );
  nand_x1_sg U12702 ( .A(\out[0][0][5] ), .B(n16788), .X(n13779) );
  nand_x1_sg U12703 ( .A(\out[0][0][6] ), .B(n16789), .X(n13771) );
  nand_x1_sg U12704 ( .A(\out[0][0][7] ), .B(n16783), .X(n13773) );
  nand_x1_sg U12705 ( .A(\out[0][0][8] ), .B(n16785), .X(n13741) );
  nand_x1_sg U12706 ( .A(\out[0][0][9] ), .B(n16784), .X(n13743) );
  nand_x1_sg U12707 ( .A(\out[0][0][10] ), .B(n16786), .X(n13735) );
  nand_x1_sg U12708 ( .A(\out[0][0][11] ), .B(n16785), .X(n13737) );
  nand_x1_sg U12709 ( .A(\out[0][0][12] ), .B(n16783), .X(n13753) );
  nand_x1_sg U12710 ( .A(\out[0][0][13] ), .B(n16780), .X(n13755) );
  nand_x1_sg U12711 ( .A(\out[0][0][14] ), .B(n16784), .X(n13747) );
  nand_x1_sg U12712 ( .A(\out[0][0][15] ), .B(n16781), .X(n13749) );
  nand_x1_sg U12713 ( .A(\out[0][0][16] ), .B(n16790), .X(n13813) );
  nand_x1_sg U12714 ( .A(\out[0][0][17] ), .B(n16790), .X(n13815) );
  nand_x1_sg U12715 ( .A(\out[0][0][18] ), .B(n16780), .X(n13807) );
  nand_x1_sg U12716 ( .A(\out[0][0][19] ), .B(n16780), .X(n13809) );
  nand_x1_sg U12717 ( .A(\out[0][1][0] ), .B(n16780), .X(n13825) );
  nand_x1_sg U12718 ( .A(\out[0][1][1] ), .B(n16780), .X(n13827) );
  nand_x1_sg U12719 ( .A(\out[0][1][2] ), .B(n16790), .X(n13819) );
  nand_x1_sg U12720 ( .A(\out[0][1][3] ), .B(n16780), .X(n13821) );
  nand_x1_sg U12721 ( .A(\out[0][1][4] ), .B(n16786), .X(n13789) );
  nand_x1_sg U12722 ( .A(\out[0][1][5] ), .B(n16790), .X(n13791) );
  nand_x1_sg U12723 ( .A(\out[0][1][6] ), .B(n16788), .X(n13783) );
  nand_x1_sg U12724 ( .A(\out[0][1][7] ), .B(n16780), .X(n13785) );
  nand_x1_sg U12725 ( .A(\out[0][1][8] ), .B(n16780), .X(n13801) );
  nand_x1_sg U12726 ( .A(\out[0][1][9] ), .B(n16790), .X(n13803) );
  nand_x1_sg U12727 ( .A(\out[0][1][10] ), .B(n16785), .X(n13795) );
  nand_x1_sg U12728 ( .A(\out[0][1][11] ), .B(n16780), .X(n13797) );
  nand_x1_sg U12729 ( .A(\out[0][1][12] ), .B(n16779), .X(n13669) );
  nand_x1_sg U12730 ( .A(\out[0][1][13] ), .B(n16779), .X(n13671) );
  nand_x1_sg U12731 ( .A(\out[0][1][14] ), .B(n16780), .X(n13663) );
  nand_x1_sg U12732 ( .A(\out[0][1][15] ), .B(n16780), .X(n13665) );
  nand_x1_sg U12733 ( .A(\out[0][1][16] ), .B(n16779), .X(n13681) );
  nand_x1_sg U12734 ( .A(\out[0][1][17] ), .B(n16779), .X(n13683) );
  nand_x1_sg U12735 ( .A(\out[0][1][18] ), .B(n16779), .X(n13675) );
  nand_x1_sg U12736 ( .A(\out[0][1][19] ), .B(n16779), .X(n13677) );
  nand_x1_sg U12737 ( .A(\out[0][2][0] ), .B(n16781), .X(n13645) );
  nand_x1_sg U12738 ( .A(\out[0][2][1] ), .B(n16781), .X(n13647) );
  nand_x1_sg U12739 ( .A(\out[0][2][2] ), .B(n16781), .X(n13639) );
  nand_x1_sg U12740 ( .A(\out[0][2][3] ), .B(n16781), .X(n13641) );
  nand_x1_sg U12741 ( .A(\out[0][2][4] ), .B(n16780), .X(n13657) );
  nand_x1_sg U12742 ( .A(\out[0][2][5] ), .B(n16780), .X(n13659) );
  nand_x1_sg U12743 ( .A(\out[0][2][6] ), .B(n16781), .X(n13651) );
  nand_x1_sg U12744 ( .A(\out[0][2][7] ), .B(n16780), .X(n13653) );
  nand_x1_sg U12745 ( .A(\out[0][2][8] ), .B(n16789), .X(n13717) );
  nand_x1_sg U12746 ( .A(\out[0][2][9] ), .B(n16789), .X(n13719) );
  nand_x1_sg U12747 ( .A(\out[0][2][10] ), .B(n16789), .X(n13711) );
  nand_x1_sg U12748 ( .A(\out[0][2][11] ), .B(n16782), .X(n13713) );
  nand_x1_sg U12749 ( .A(\out[0][2][12] ), .B(n16788), .X(n13729) );
  nand_x1_sg U12750 ( .A(\out[0][2][13] ), .B(n16785), .X(n13731) );
  nand_x1_sg U12751 ( .A(\out[0][2][14] ), .B(n16789), .X(n13723) );
  nand_x1_sg U12752 ( .A(\out[0][2][15] ), .B(n16786), .X(n13725) );
  nand_x1_sg U12753 ( .A(\out[0][2][16] ), .B(n16778), .X(n13693) );
  nand_x1_sg U12754 ( .A(\out[0][2][17] ), .B(n16778), .X(n13695) );
  nand_x1_sg U12755 ( .A(\out[0][2][18] ), .B(n16778), .X(n13687) );
  nand_x1_sg U12756 ( .A(\out[0][2][19] ), .B(n16778), .X(n13689) );
  nand_x1_sg U12757 ( .A(\out[0][3][0] ), .B(n16789), .X(n13705) );
  nand_x1_sg U12758 ( .A(\out[0][3][1] ), .B(n16779), .X(n13707) );
  nand_x1_sg U12759 ( .A(\out[0][3][2] ), .B(n16778), .X(n13699) );
  nand_x1_sg U12760 ( .A(\out[0][3][3] ), .B(n16778), .X(n13701) );
  nand_x1_sg U12761 ( .A(\out[1][2][9] ), .B(n16790), .X(n13573) );
  nand_x1_sg U12762 ( .A(\out[1][2][12] ), .B(n16788), .X(n13583) );
  nand_x1_sg U12763 ( .A(\out[1][2][13] ), .B(n16789), .X(n13585) );
  nand_x1_sg U12764 ( .A(\out[1][2][14] ), .B(n16780), .X(n13577) );
  nand_x1_sg U12765 ( .A(\out[1][2][15] ), .B(n16783), .X(n13579) );
  nand_x1_sg U12766 ( .A(\out[1][3][4] ), .B(n16779), .X(n13619) );
  nand_x1_sg U12767 ( .A(\out[1][3][5] ), .B(n16779), .X(n13621) );
  nand_x1_sg U12768 ( .A(\out[1][3][6] ), .B(n16778), .X(n13613) );
  nand_x1_sg U12769 ( .A(\out[1][3][7] ), .B(n16788), .X(n13615) );
  nand_x1_sg U12770 ( .A(\out[1][3][8] ), .B(n16788), .X(n13631) );
  nand_x1_sg U12771 ( .A(\out[1][3][9] ), .B(n16778), .X(n13633) );
  nand_x1_sg U12772 ( .A(\out[1][3][10] ), .B(n16791), .X(n13625) );
  nand_x1_sg U12773 ( .A(\out[1][3][11] ), .B(n16783), .X(n13627) );
  nand_x1_sg U12774 ( .A(\out[1][3][12] ), .B(n16782), .X(n13595) );
  nand_x1_sg U12775 ( .A(\out[1][3][13] ), .B(n16782), .X(n13597) );
  nand_x1_sg U12776 ( .A(\out[1][3][14] ), .B(n16782), .X(n13589) );
  nand_x1_sg U12777 ( .A(\out[1][3][15] ), .B(n16782), .X(n13591) );
  nand_x1_sg U12778 ( .A(\out[1][3][16] ), .B(n16788), .X(n13607) );
  nand_x1_sg U12779 ( .A(\out[1][3][17] ), .B(n16788), .X(n13609) );
  nand_x1_sg U12780 ( .A(\out[1][3][18] ), .B(n16782), .X(n13601) );
  nand_x1_sg U12781 ( .A(\out[1][3][19] ), .B(n16782), .X(n13603) );
  nand_x1_sg U12782 ( .A(\out[2][1][13] ), .B(n16788), .X(n13787) );
  nand_x1_sg U12783 ( .A(\out[2][1][15] ), .B(n16789), .X(n13635) );
  nand_x1_sg U12784 ( .A(\out[2][2][1] ), .B(n16778), .X(n13763) );
  nand_x1_sg U12785 ( .A(\out[2][2][2] ), .B(n16780), .X(n13781) );
  nand_x1_sg U12786 ( .A(\out[2][2][4] ), .B(n16778), .X(n13685) );
  nand_x1_sg U12787 ( .A(\out[2][2][12] ), .B(n16783), .X(n13745) );
  nand_x1_sg U12788 ( .A(\out[2][2][16] ), .B(n16781), .X(n13637) );
  nand_x1_sg U12789 ( .A(\out[2][2][17] ), .B(n16781), .X(n13643) );
  nand_x1_sg U12790 ( .A(\out[2][2][18] ), .B(n16786), .X(n13575) );
  nand_x1_sg U12791 ( .A(\out[2][2][19] ), .B(n16780), .X(n13811) );
  nand_x1_sg U12792 ( .A(\out[2][3][0] ), .B(n16778), .X(n13691) );
  nand_x1_sg U12793 ( .A(\out[2][3][1] ), .B(n16778), .X(n13697) );
  nand_x1_sg U12794 ( .A(\out[2][3][2] ), .B(n16785), .X(n13721) );
  nand_x1_sg U12795 ( .A(\out[2][3][3] ), .B(n16789), .X(n13775) );
  nand_x1_sg U12796 ( .A(\out[2][3][7] ), .B(n16780), .X(n13709) );
  nand_x1_sg U12797 ( .A(\out[2][3][8] ), .B(n16782), .X(n13605) );
  nand_x1_sg U12798 ( .A(\out[2][3][11] ), .B(n16790), .X(n13823) );
  nand_x1_sg U12799 ( .A(\out[3][0][0] ), .B(n16780), .X(n13655) );
  nand_x1_sg U12800 ( .A(\out[3][0][1] ), .B(n16780), .X(n13661) );
  nand_x1_sg U12801 ( .A(\out[3][0][2] ), .B(n16784), .X(n13727) );
  nand_x1_sg U12802 ( .A(\out[3][0][3] ), .B(n16779), .X(n13673) );
  nand_x1_sg U12803 ( .A(\out[3][0][4] ), .B(n16781), .X(n13703) );
  nand_x1_sg U12804 ( .A(\out[3][0][5] ), .B(n16780), .X(n13667) );
  nand_x1_sg U12805 ( .A(\out[3][0][6] ), .B(n16779), .X(n13679) );
  nand_x1_sg U12806 ( .A(\out[3][0][7] ), .B(n16784), .X(n13793) );
  nand_x1_sg U12807 ( .A(\out[3][0][8] ), .B(n16785), .X(n13581) );
  nand_x1_sg U12808 ( .A(\out[3][0][9] ), .B(n16780), .X(n13715) );
  nand_x1_sg U12809 ( .A(\out[3][0][11] ), .B(n16781), .X(n13649) );
  nand_x1_sg U12810 ( .A(\out[3][0][15] ), .B(n16788), .X(n13611) );
  nand_x1_sg U12811 ( .A(\out[3][1][12] ), .B(n16783), .X(n13617) );
  nand_x1_sg U12812 ( .A(\out[3][1][13] ), .B(n16782), .X(n13623) );
  nand_x1_sg U12813 ( .A(\out[3][1][15] ), .B(n16781), .X(n13629) );
  nand_x1_sg U12814 ( .A(\out[3][1][16] ), .B(n16784), .X(n13587) );
  nand_x1_sg U12815 ( .A(\out[3][1][17] ), .B(n16782), .X(n13593) );
  nand_x1_sg U12816 ( .A(\out[3][1][19] ), .B(n16782), .X(n13599) );
  nand_x1_sg U12817 ( .A(\out[3][2][10] ), .B(n16779), .X(n13757) );
  nand_x1_sg U12818 ( .A(\out[3][2][11] ), .B(n16786), .X(n13751) );
  nand_x1_sg U12819 ( .A(\out[3][2][16] ), .B(n16780), .X(n13799) );
  nand_x1_sg U12820 ( .A(\out[3][2][17] ), .B(n16790), .X(n13805) );
  nand_x1_sg U12821 ( .A(\out[3][2][19] ), .B(n16780), .X(n13817) );
  nand_x1_sg U12822 ( .A(\out[3][3][0] ), .B(n16784), .X(n13733) );
  nand_x1_sg U12823 ( .A(\out[3][3][1] ), .B(n16786), .X(n13739) );
  nand_x1_sg U12824 ( .A(\out[3][3][3] ), .B(n16786), .X(n13769) );
  nand_x1_sg U12825 ( .A(\out[1][0][16] ), .B(n16785), .X(n13283) );
  nand_x1_sg U12826 ( .A(\out[1][0][17] ), .B(n16784), .X(n13285) );
  nand_x1_sg U12827 ( .A(\out[1][0][18] ), .B(n16785), .X(n13277) );
  nand_x1_sg U12828 ( .A(\out[1][0][19] ), .B(n16785), .X(n13279) );
  nand_x1_sg U12829 ( .A(\out[1][1][0] ), .B(n16784), .X(n13295) );
  nand_x1_sg U12830 ( .A(\out[1][1][1] ), .B(n16784), .X(n13297) );
  nand_x1_sg U12831 ( .A(\out[1][1][2] ), .B(n16784), .X(n13289) );
  nand_x1_sg U12832 ( .A(\out[1][1][3] ), .B(n16784), .X(n13291) );
  nand_x1_sg U12833 ( .A(\out[1][1][4] ), .B(n16786), .X(n13259) );
  nand_x1_sg U12834 ( .A(\out[1][1][5] ), .B(n16786), .X(n13261) );
  nand_x1_sg U12835 ( .A(\out[1][1][6] ), .B(n16786), .X(n13253) );
  nand_x1_sg U12836 ( .A(\out[1][1][7] ), .B(n16786), .X(n13255) );
  nand_x1_sg U12837 ( .A(\out[1][1][8] ), .B(n16785), .X(n13271) );
  nand_x1_sg U12838 ( .A(\out[1][1][9] ), .B(n16785), .X(n13273) );
  nand_x1_sg U12839 ( .A(\out[1][1][10] ), .B(n16786), .X(n13265) );
  nand_x1_sg U12840 ( .A(\out[1][1][11] ), .B(n16786), .X(n13267) );
  nand_x1_sg U12841 ( .A(\out[1][2][0] ), .B(n16783), .X(n13307) );
  nand_x1_sg U12842 ( .A(\out[1][2][1] ), .B(n16783), .X(n13309) );
  nand_x1_sg U12843 ( .A(\out[1][2][2] ), .B(n16783), .X(n13301) );
  nand_x1_sg U12844 ( .A(\out[1][2][3] ), .B(n16783), .X(n13303) );
  nand_x1_sg U12845 ( .A(\out[1][2][6] ), .B(n16783), .X(n13313) );
  nand_x1_sg U12846 ( .A(\out[1][2][7] ), .B(n16783), .X(n13315) );
  nand_x1_sg U12847 ( .A(\out[2][1][12] ), .B(n16786), .X(n13257) );
  nand_x1_sg U12848 ( .A(\out[2][1][16] ), .B(n16788), .X(n13223) );
  nand_x1_sg U12849 ( .A(\out[2][1][17] ), .B(n16784), .X(n13299) );
  nand_x1_sg U12850 ( .A(\out[2][2][5] ), .B(n16790), .X(n13195) );
  nand_x1_sg U12851 ( .A(\out[2][2][6] ), .B(n16785), .X(n13281) );
  nand_x1_sg U12852 ( .A(\out[2][2][7] ), .B(n16791), .X(n13199) );
  nand_x1_sg U12853 ( .A(\out[2][2][10] ), .B(n16789), .X(n13197) );
  nand_x1_sg U12854 ( .A(\out[2][2][13] ), .B(n16783), .X(n13251) );
  nand_x1_sg U12855 ( .A(\out[2][2][15] ), .B(n16784), .X(n13293) );
  nand_x1_sg U12856 ( .A(\out[2][3][5] ), .B(n16791), .X(n13231) );
  nand_x1_sg U12857 ( .A(\out[2][3][6] ), .B(n16790), .X(n13209) );
  nand_x1_sg U12858 ( .A(\out[2][3][9] ), .B(n16789), .X(n13215) );
  nand_x1_sg U12859 ( .A(\out[2][3][10] ), .B(n16793), .X(n13211) );
  nand_x1_sg U12860 ( .A(\out[2][3][12] ), .B(n16790), .X(n13221) );
  nand_x1_sg U12861 ( .A(\out[2][3][13] ), .B(n16793), .X(n13213) );
  nand_x1_sg U12862 ( .A(\out[2][3][14] ), .B(n16790), .X(n13203) );
  nand_x1_sg U12863 ( .A(\out[2][3][15] ), .B(n16795), .X(n13205) );
  nand_x1_sg U12864 ( .A(\out[2][3][18] ), .B(n16791), .X(n13207) );
  nand_x1_sg U12865 ( .A(\out[3][0][10] ), .B(n16791), .X(n13229) );
  nand_x1_sg U12866 ( .A(\out[3][0][12] ), .B(n16791), .X(n13233) );
  nand_x1_sg U12867 ( .A(\out[3][0][13] ), .B(n16788), .X(n13239) );
  nand_x1_sg U12868 ( .A(\out[3][0][14] ), .B(n16789), .X(n13245) );
  nand_x1_sg U12869 ( .A(\out[3][0][18] ), .B(n16788), .X(n13217) );
  nand_x1_sg U12870 ( .A(\out[3][0][19] ), .B(n16790), .X(n13219) );
  nand_x1_sg U12871 ( .A(\out[3][1][14] ), .B(n16793), .X(n13247) );
  nand_x1_sg U12872 ( .A(\out[3][1][18] ), .B(n16793), .X(n13249) );
  nand_x1_sg U12873 ( .A(\out[3][2][4] ), .B(n16795), .X(n13241) );
  nand_x1_sg U12874 ( .A(\out[3][2][5] ), .B(n16793), .X(n13243) );
  nand_x1_sg U12875 ( .A(\out[3][2][6] ), .B(n16789), .X(n13235) );
  nand_x1_sg U12876 ( .A(\out[3][2][7] ), .B(n16793), .X(n13237) );
  nand_x1_sg U12877 ( .A(\out[3][2][8] ), .B(n16791), .X(n13187) );
  nand_x1_sg U12878 ( .A(\out[3][2][9] ), .B(n16788), .X(n13191) );
  nand_x1_sg U12879 ( .A(\out[3][2][12] ), .B(n16785), .X(n13269) );
  nand_x1_sg U12880 ( .A(\out[3][2][13] ), .B(n16785), .X(n13275) );
  nand_x1_sg U12881 ( .A(\out[3][2][14] ), .B(n16789), .X(n13193) );
  nand_x1_sg U12882 ( .A(\out[3][2][15] ), .B(n16784), .X(n13287) );
  nand_x1_sg U12883 ( .A(\out[3][2][18] ), .B(n16786), .X(n13263) );
  nand_x1_sg U12884 ( .A(\out[3][3][2] ), .B(n16790), .X(n13201) );
  nand_x1_sg U12885 ( .A(\out[3][3][12] ), .B(n16783), .X(n13305) );
  nand_x1_sg U12886 ( .A(\out[3][3][13] ), .B(n16783), .X(n13311) );
  nand_x1_sg U12887 ( .A(\out[3][3][14] ), .B(n16788), .X(n13227) );
  nand_x1_sg U12888 ( .A(\out[3][3][18] ), .B(n16788), .X(n13225) );
  nor_x1_sg U12889 ( .A(state[0]), .B(n18399), .X(n14481) );
  nand_x2_sg U12890 ( .A(n14472), .B(input_ready), .X(n14470) );
  nand_x1_sg U12891 ( .A(n16728), .B(n16748), .X(n14189) );
  nand_x1_sg U12892 ( .A(n16726), .B(n16748), .X(n14191) );
  nand_x1_sg U12893 ( .A(n16724), .B(n16748), .X(n14183) );
  nand_x1_sg U12894 ( .A(n16722), .B(n16748), .X(n14185) );
  nand_x1_sg U12895 ( .A(n16720), .B(n16747), .X(n14201) );
  nand_x1_sg U12896 ( .A(n16718), .B(n16747), .X(n14203) );
  nand_x1_sg U12897 ( .A(n16716), .B(n16748), .X(n14195) );
  nand_x1_sg U12898 ( .A(n16714), .B(n16748), .X(n14197) );
  nand_x1_sg U12899 ( .A(n16680), .B(n16745), .X(n14117) );
  nand_x1_sg U12900 ( .A(n16678), .B(n16752), .X(n14119) );
  nand_x1_sg U12901 ( .A(n16676), .B(n16746), .X(n14111) );
  nand_x1_sg U12902 ( .A(n16674), .B(n16751), .X(n14113) );
  nand_x1_sg U12903 ( .A(n16672), .B(n16752), .X(n14129) );
  nand_x1_sg U12904 ( .A(n16670), .B(n16752), .X(n14131) );
  nand_x1_sg U12905 ( .A(n16668), .B(n16752), .X(n14123) );
  nand_x1_sg U12906 ( .A(n16666), .B(n16752), .X(n14125) );
  nand_x1_sg U12907 ( .A(n16664), .B(n16748), .X(n14093) );
  nand_x1_sg U12908 ( .A(n16662), .B(n16748), .X(n14095) );
  nand_x1_sg U12909 ( .A(n16660), .B(n16747), .X(n14087) );
  nand_x1_sg U12910 ( .A(n16658), .B(n16753), .X(n14089) );
  nand_x1_sg U12911 ( .A(n16656), .B(n16745), .X(n14105) );
  nand_x1_sg U12912 ( .A(n16654), .B(n16745), .X(n14107) );
  nand_x1_sg U12913 ( .A(n16652), .B(n16754), .X(n14099) );
  nand_x1_sg U12914 ( .A(n16650), .B(n16755), .X(n14101) );
  nand_x1_sg U12915 ( .A(n16648), .B(n16750), .X(n14165) );
  nand_x1_sg U12916 ( .A(n16646), .B(n16749), .X(n14167) );
  nand_x1_sg U12917 ( .A(n16644), .B(n16750), .X(n14159) );
  nand_x1_sg U12918 ( .A(n16642), .B(n16750), .X(n14161) );
  nand_x1_sg U12919 ( .A(n16640), .B(n16749), .X(n14177) );
  nand_x1_sg U12920 ( .A(n16638), .B(n16749), .X(n14179) );
  nand_x1_sg U12921 ( .A(n16636), .B(n16749), .X(n14171) );
  nand_x1_sg U12922 ( .A(n16634), .B(n16749), .X(n14173) );
  nand_x1_sg U12923 ( .A(n16632), .B(n16751), .X(n14141) );
  nand_x1_sg U12924 ( .A(n16630), .B(n16751), .X(n14143) );
  nand_x1_sg U12925 ( .A(n16628), .B(n16751), .X(n14135) );
  nand_x1_sg U12926 ( .A(n16626), .B(n16751), .X(n14137) );
  nand_x1_sg U12927 ( .A(n16624), .B(n16750), .X(n14153) );
  nand_x1_sg U12928 ( .A(n16622), .B(n16750), .X(n14155) );
  nand_x1_sg U12929 ( .A(n16620), .B(n16751), .X(n14147) );
  nand_x1_sg U12930 ( .A(n16618), .B(n16751), .X(n14149) );
  nand_x1_sg U12931 ( .A(n16596), .B(n16755), .X(n13977) );
  nand_x1_sg U12932 ( .A(n16594), .B(n16752), .X(n14133) );
  nand_x1_sg U12933 ( .A(n16588), .B(n16757), .X(n14061) );
  nand_x1_sg U12934 ( .A(n16584), .B(n16748), .X(n14055) );
  nand_x1_sg U12935 ( .A(n16582), .B(n16750), .X(n14019) );
  nand_x1_sg U12936 ( .A(n16578), .B(n16751), .X(n14139) );
  nand_x1_sg U12937 ( .A(n16572), .B(n16745), .X(n13971) );
  nand_x1_sg U12938 ( .A(n16570), .B(n16748), .X(n13995) );
  nand_x1_sg U12939 ( .A(n16542), .B(n16755), .X(n13959) );
  nand_x1_sg U12940 ( .A(n16536), .B(n16747), .X(n14199) );
  nand_x1_sg U12941 ( .A(n16528), .B(n16750), .X(n14151) );
  nand_x1_sg U12942 ( .A(n16526), .B(n16749), .X(n14091) );
  nand_x1_sg U12943 ( .A(n16522), .B(n16749), .X(n14181) );
  nand_x1_sg U12944 ( .A(n16500), .B(n16757), .X(n14025) );
  nand_x1_sg U12945 ( .A(n16488), .B(n16748), .X(n14187) );
  nand_x1_sg U12946 ( .A(n16486), .B(n16748), .X(n14193) );
  nand_x1_sg U12947 ( .A(n16480), .B(n16747), .X(n14205) );
  nand_x1_sg U12948 ( .A(n16478), .B(n16747), .X(n14211) );
  nand_x1_sg U12949 ( .A(n16472), .B(n16752), .X(n14121) );
  nand_x1_sg U12950 ( .A(n16470), .B(n16752), .X(n14127) );
  nand_x1_sg U12951 ( .A(n16466), .B(n16751), .X(n14145) );
  nand_x1_sg U12952 ( .A(n16464), .B(n16750), .X(n14097) );
  nand_x1_sg U12953 ( .A(n16462), .B(n16746), .X(n14103) );
  nand_x1_sg U12954 ( .A(n16460), .B(n16752), .X(n14109) );
  nand_x1_sg U12955 ( .A(n16458), .B(n16745), .X(n14115) );
  nand_x1_sg U12956 ( .A(n16456), .B(n16748), .X(n14013) );
  nand_x1_sg U12957 ( .A(n16454), .B(n16746), .X(n13989) );
  nand_x1_sg U12958 ( .A(n16440), .B(n16750), .X(n14157) );
  nand_x1_sg U12959 ( .A(n16438), .B(n16750), .X(n14163) );
  nand_x1_sg U12960 ( .A(n16436), .B(n16749), .X(n14169) );
  nand_x1_sg U12961 ( .A(n16434), .B(n16749), .X(n14175) );
  nand_x1_sg U12962 ( .A(n16392), .B(n16757), .X(n14043) );
  nand_x1_sg U12963 ( .A(n16390), .B(n16753), .X(n14049) );
  nand_x1_sg U12964 ( .A(n16388), .B(n16750), .X(n14073) );
  nand_x1_sg U12965 ( .A(n16386), .B(n16752), .X(n14079) );
  nand_x1_sg U12966 ( .A(n16384), .B(n16757), .X(n14001) );
  nand_x1_sg U12967 ( .A(n16382), .B(n16747), .X(n14007) );
  nand_x1_sg U12968 ( .A(n16380), .B(n16757), .X(n14031) );
  nand_x1_sg U12969 ( .A(n16378), .B(n16749), .X(n14037) );
  nand_x1_sg U12970 ( .A(n16370), .B(n16757), .X(n13965) );
  nand_x1_sg U12971 ( .A(n16368), .B(n16749), .X(n14067) );
  nand_x1_sg U12972 ( .A(n16366), .B(n16752), .X(n13983) );
  nand_x1_sg U12973 ( .A(n16362), .B(n16757), .X(n14085) );
  nand_x1_sg U12974 ( .A(n16232), .B(n16749), .X(n14021) );
  nand_x1_sg U12975 ( .A(n16230), .B(n16753), .X(n14023) );
  nand_x1_sg U12976 ( .A(n16228), .B(n16752), .X(n14015) );
  nand_x1_sg U12977 ( .A(n16226), .B(n16751), .X(n14017) );
  nand_x1_sg U12978 ( .A(n16224), .B(n16754), .X(n14033) );
  nand_x1_sg U12979 ( .A(n16222), .B(n16755), .X(n14035) );
  nand_x1_sg U12980 ( .A(n16220), .B(n16757), .X(n14027) );
  nand_x1_sg U12981 ( .A(n16218), .B(n16757), .X(n14029) );
  nand_x1_sg U12982 ( .A(n16216), .B(n16746), .X(n13997) );
  nand_x1_sg U12983 ( .A(n16214), .B(n16749), .X(n13999) );
  nand_x1_sg U12984 ( .A(n16212), .B(n16757), .X(n13991) );
  nand_x1_sg U12985 ( .A(n16210), .B(n16747), .X(n13993) );
  nand_x1_sg U12986 ( .A(n16208), .B(n16757), .X(n14009) );
  nand_x1_sg U12987 ( .A(n16206), .B(n16753), .X(n14011) );
  nand_x1_sg U12988 ( .A(n16204), .B(n16757), .X(n14003) );
  nand_x1_sg U12989 ( .A(n16202), .B(n16757), .X(n14005) );
  nand_x1_sg U12990 ( .A(n16200), .B(n16753), .X(n14069) );
  nand_x1_sg U12991 ( .A(n16198), .B(n16751), .X(n14071) );
  nand_x1_sg U12992 ( .A(n16196), .B(n16754), .X(n14063) );
  nand_x1_sg U12993 ( .A(n16194), .B(n16755), .X(n14065) );
  nand_x1_sg U12994 ( .A(n16192), .B(n16757), .X(n14081) );
  nand_x1_sg U12995 ( .A(n16190), .B(n16751), .X(n14083) );
  nand_x1_sg U12996 ( .A(n16188), .B(n16754), .X(n14075) );
  nand_x1_sg U12997 ( .A(n16186), .B(n16749), .X(n14077) );
  nand_x1_sg U12998 ( .A(n16184), .B(n16754), .X(n14045) );
  nand_x1_sg U12999 ( .A(n16182), .B(n16757), .X(n14047) );
  nand_x1_sg U13000 ( .A(n16180), .B(n16750), .X(n14039) );
  nand_x1_sg U13001 ( .A(n16178), .B(n16757), .X(n14041) );
  nand_x1_sg U13002 ( .A(n16176), .B(n16752), .X(n14057) );
  nand_x1_sg U13003 ( .A(n16174), .B(n16757), .X(n14059) );
  nand_x1_sg U13004 ( .A(n16172), .B(n16746), .X(n14051) );
  nand_x1_sg U13005 ( .A(n16170), .B(n16750), .X(n14053) );
  nand_x1_sg U13006 ( .A(n16136), .B(n16757), .X(n13973) );
  nand_x1_sg U13007 ( .A(n16134), .B(n16751), .X(n13975) );
  nand_x1_sg U13008 ( .A(n16132), .B(n16755), .X(n13967) );
  nand_x1_sg U13009 ( .A(n16130), .B(n16757), .X(n13969) );
  nand_x1_sg U13010 ( .A(n16128), .B(n16752), .X(n13985) );
  nand_x1_sg U13011 ( .A(n16126), .B(n16747), .X(n13987) );
  nand_x1_sg U13012 ( .A(n16124), .B(n16755), .X(n13979) );
  nand_x1_sg U13013 ( .A(n16122), .B(n16750), .X(n13981) );
  nand_x1_sg U13014 ( .A(n16112), .B(n16755), .X(n13961) );
  nand_x1_sg U13015 ( .A(n16110), .B(n16748), .X(n13963) );
  nand_x1_sg U13016 ( .A(n16104), .B(n16747), .X(n14213) );
  nand_x1_sg U13017 ( .A(n16100), .B(n16747), .X(n14207) );
  nand_x1_sg U13018 ( .A(n16098), .B(n16747), .X(n14209) );
  nand_x1_sg U13019 ( .A(n16730), .B(n16751), .X(n14221) );
  nand_x1_sg U13020 ( .A(n16712), .B(n16746), .X(n14261) );
  nand_x1_sg U13021 ( .A(n16710), .B(n16745), .X(n14263) );
  nand_x1_sg U13022 ( .A(n16708), .B(n16745), .X(n14255) );
  nand_x1_sg U13023 ( .A(n16706), .B(n16747), .X(n14257) );
  nand_x1_sg U13024 ( .A(n16704), .B(n16745), .X(n14273) );
  nand_x1_sg U13025 ( .A(n16702), .B(n16745), .X(n14275) );
  nand_x1_sg U13026 ( .A(n16700), .B(n16745), .X(n14267) );
  nand_x1_sg U13027 ( .A(n16698), .B(n16745), .X(n14269) );
  nand_x1_sg U13028 ( .A(n16696), .B(n16746), .X(n14237) );
  nand_x1_sg U13029 ( .A(n16694), .B(n16746), .X(n14239) );
  nand_x1_sg U13030 ( .A(n16692), .B(n16746), .X(n14231) );
  nand_x1_sg U13031 ( .A(n16690), .B(n16746), .X(n14233) );
  nand_x1_sg U13032 ( .A(n16688), .B(n16748), .X(n14249) );
  nand_x1_sg U13033 ( .A(n16686), .B(n16749), .X(n14251) );
  nand_x1_sg U13034 ( .A(n16684), .B(n16746), .X(n14243) );
  nand_x1_sg U13035 ( .A(n16682), .B(n16746), .X(n14245) );
  nand_x1_sg U13036 ( .A(n16614), .B(n16755), .X(n14279) );
  nand_x1_sg U13037 ( .A(n16612), .B(n16754), .X(n14393) );
  nand_x1_sg U13038 ( .A(n16610), .B(n16745), .X(n14277) );
  nand_x1_sg U13039 ( .A(n16604), .B(n16753), .X(n14447) );
  nand_x1_sg U13040 ( .A(n16600), .B(n16752), .X(n14217) );
  nand_x1_sg U13041 ( .A(n16598), .B(n16748), .X(n14291) );
  nand_x1_sg U13042 ( .A(n16592), .B(n16757), .X(n14327) );
  nand_x1_sg U13043 ( .A(n16568), .B(n16752), .X(n14303) );
  nand_x1_sg U13044 ( .A(n16566), .B(n16755), .X(n14321) );
  nand_x1_sg U13045 ( .A(n16564), .B(n16746), .X(n14235) );
  nand_x1_sg U13046 ( .A(n16562), .B(n16757), .X(n14453) );
  nand_x1_sg U13047 ( .A(n16560), .B(n16754), .X(n14333) );
  nand_x1_sg U13048 ( .A(n16558), .B(n16753), .X(n14339) );
  nand_x1_sg U13049 ( .A(n16556), .B(n16753), .X(n14345) );
  nand_x1_sg U13050 ( .A(n16554), .B(n16748), .X(n14363) );
  nand_x1_sg U13051 ( .A(n16544), .B(n16750), .X(n14253) );
  nand_x1_sg U13052 ( .A(n16538), .B(n16745), .X(n14465) );
  nand_x1_sg U13053 ( .A(n16520), .B(n16751), .X(n14375) );
  nand_x1_sg U13054 ( .A(n16518), .B(n16755), .X(n14381) );
  nand_x1_sg U13055 ( .A(n16516), .B(n16753), .X(n14423) );
  nand_x1_sg U13056 ( .A(n16514), .B(n16757), .X(n14387) );
  nand_x1_sg U13057 ( .A(n16512), .B(n16751), .X(n14417) );
  nand_x1_sg U13058 ( .A(n16510), .B(n16750), .X(n14309) );
  nand_x1_sg U13059 ( .A(n16508), .B(n16751), .X(n14351) );
  nand_x1_sg U13060 ( .A(n16506), .B(n16752), .X(n14357) );
  nand_x1_sg U13061 ( .A(n16504), .B(n16750), .X(n14411) );
  nand_x1_sg U13062 ( .A(n16502), .B(n16749), .X(n14369) );
  nand_x1_sg U13063 ( .A(n16498), .B(n16754), .X(n14429) );
  nand_x1_sg U13064 ( .A(n16492), .B(n16745), .X(n14271) );
  nand_x1_sg U13065 ( .A(n16484), .B(n16746), .X(n14223) );
  nand_x1_sg U13066 ( .A(n16482), .B(n16753), .X(n14229) );
  nand_x1_sg U13067 ( .A(n16448), .B(n16746), .X(n14241) );
  nand_x1_sg U13068 ( .A(n16446), .B(n16746), .X(n14247) );
  nand_x1_sg U13069 ( .A(n16444), .B(n16754), .X(n14259) );
  nand_x1_sg U13070 ( .A(n16442), .B(n16745), .X(n14265) );
  nand_x1_sg U13071 ( .A(n16420), .B(n16746), .X(n14399) );
  nand_x1_sg U13072 ( .A(n16418), .B(n16752), .X(n14405) );
  nand_x1_sg U13073 ( .A(n16408), .B(n16757), .X(n14285) );
  nand_x1_sg U13074 ( .A(n16406), .B(n16749), .X(n14297) );
  nand_x1_sg U13075 ( .A(n16402), .B(n16754), .X(n14315) );
  nand_x1_sg U13076 ( .A(n16400), .B(n16757), .X(n14435) );
  nand_x1_sg U13077 ( .A(n16398), .B(n16754), .X(n14441) );
  nand_x1_sg U13078 ( .A(n16394), .B(n16757), .X(n14459) );
  nand_x1_sg U13079 ( .A(n16360), .B(n16752), .X(n14407) );
  nand_x1_sg U13080 ( .A(n16358), .B(n16750), .X(n14409) );
  nand_x1_sg U13081 ( .A(n16356), .B(n16745), .X(n14401) );
  nand_x1_sg U13082 ( .A(n16354), .B(n16745), .X(n14403) );
  nand_x1_sg U13083 ( .A(n16352), .B(n16755), .X(n14419) );
  nand_x1_sg U13084 ( .A(n16350), .B(n16757), .X(n14421) );
  nand_x1_sg U13085 ( .A(n16348), .B(n16745), .X(n14413) );
  nand_x1_sg U13086 ( .A(n16346), .B(n16747), .X(n14415) );
  nand_x1_sg U13087 ( .A(n16344), .B(n16752), .X(n14383) );
  nand_x1_sg U13088 ( .A(n16342), .B(n16746), .X(n14385) );
  nand_x1_sg U13089 ( .A(n16340), .B(n16757), .X(n14377) );
  nand_x1_sg U13090 ( .A(n16338), .B(n16748), .X(n14379) );
  nand_x1_sg U13091 ( .A(n16336), .B(n16746), .X(n14395) );
  nand_x1_sg U13092 ( .A(n16334), .B(n16751), .X(n14397) );
  nand_x1_sg U13093 ( .A(n16332), .B(n16747), .X(n14389) );
  nand_x1_sg U13094 ( .A(n16330), .B(n16745), .X(n14391) );
  nand_x1_sg U13095 ( .A(n16328), .B(n16751), .X(n14455) );
  nand_x1_sg U13096 ( .A(n16326), .B(n16752), .X(n14457) );
  nand_x1_sg U13097 ( .A(n16324), .B(n16753), .X(n14449) );
  nand_x1_sg U13098 ( .A(n16322), .B(n16752), .X(n14451) );
  nand_x1_sg U13099 ( .A(n16320), .B(n16748), .X(n14467) );
  nand_x1_sg U13100 ( .A(n16318), .B(n16757), .X(n14469) );
  nand_x1_sg U13101 ( .A(n16316), .B(n16745), .X(n14461) );
  nand_x1_sg U13102 ( .A(n16314), .B(n16755), .X(n14463) );
  nand_x1_sg U13103 ( .A(n16312), .B(n16757), .X(n14431) );
  nand_x1_sg U13104 ( .A(n16310), .B(n16746), .X(n14433) );
  nand_x1_sg U13105 ( .A(n16308), .B(n16750), .X(n14425) );
  nand_x1_sg U13106 ( .A(n16306), .B(n16748), .X(n14427) );
  nand_x1_sg U13107 ( .A(n16304), .B(n16751), .X(n14443) );
  nand_x1_sg U13108 ( .A(n16302), .B(n16757), .X(n14445) );
  nand_x1_sg U13109 ( .A(n16300), .B(n16749), .X(n14437) );
  nand_x1_sg U13110 ( .A(n16298), .B(n16747), .X(n14439) );
  nand_x1_sg U13111 ( .A(n16296), .B(n16753), .X(n14311) );
  nand_x1_sg U13112 ( .A(n16294), .B(n16757), .X(n14313) );
  nand_x1_sg U13113 ( .A(n16292), .B(n16757), .X(n14305) );
  nand_x1_sg U13114 ( .A(n16290), .B(n16748), .X(n14307) );
  nand_x1_sg U13115 ( .A(n16288), .B(n16745), .X(n14323) );
  nand_x1_sg U13116 ( .A(n16286), .B(n16751), .X(n14325) );
  nand_x1_sg U13117 ( .A(n16284), .B(n16755), .X(n14317) );
  nand_x1_sg U13118 ( .A(n16282), .B(n16749), .X(n14319) );
  nand_x1_sg U13119 ( .A(n16280), .B(n16753), .X(n14287) );
  nand_x1_sg U13120 ( .A(n16278), .B(n16749), .X(n14289) );
  nand_x1_sg U13121 ( .A(n16276), .B(n16754), .X(n14281) );
  nand_x1_sg U13122 ( .A(n16274), .B(n16757), .X(n14283) );
  nand_x1_sg U13123 ( .A(n16272), .B(n16747), .X(n14299) );
  nand_x1_sg U13124 ( .A(n16270), .B(n16753), .X(n14301) );
  nand_x1_sg U13125 ( .A(n16268), .B(n16750), .X(n14293) );
  nand_x1_sg U13126 ( .A(n16266), .B(n16754), .X(n14295) );
  nand_x1_sg U13127 ( .A(n16264), .B(n16748), .X(n14359) );
  nand_x1_sg U13128 ( .A(n16262), .B(n16749), .X(n14361) );
  nand_x1_sg U13129 ( .A(n16260), .B(n16750), .X(n14353) );
  nand_x1_sg U13130 ( .A(n16258), .B(n16754), .X(n14355) );
  nand_x1_sg U13131 ( .A(n16256), .B(n16747), .X(n14371) );
  nand_x1_sg U13132 ( .A(n16254), .B(n16757), .X(n14373) );
  nand_x1_sg U13133 ( .A(n16252), .B(n16755), .X(n14365) );
  nand_x1_sg U13134 ( .A(n16250), .B(n16746), .X(n14367) );
  nand_x1_sg U13135 ( .A(n16248), .B(n16757), .X(n14335) );
  nand_x1_sg U13136 ( .A(n16246), .B(n16747), .X(n14337) );
  nand_x1_sg U13137 ( .A(n16244), .B(n16747), .X(n14329) );
  nand_x1_sg U13138 ( .A(n16242), .B(n16748), .X(n14331) );
  nand_x1_sg U13139 ( .A(n16240), .B(n16750), .X(n14347) );
  nand_x1_sg U13140 ( .A(n16238), .B(n16746), .X(n14349) );
  nand_x1_sg U13141 ( .A(n16236), .B(n16750), .X(n14341) );
  nand_x1_sg U13142 ( .A(n16234), .B(n16753), .X(n14343) );
  nand_x1_sg U13143 ( .A(n16102), .B(n16755), .X(n14215) );
  nand_x1_sg U13144 ( .A(n16096), .B(n16751), .X(n14225) );
  nand_x1_sg U13145 ( .A(n16094), .B(n16752), .X(n14227) );
  nand_x1_sg U13146 ( .A(n16092), .B(n16746), .X(n14219) );
  nand_x1_sg U13147 ( .A(n16616), .B(n16749), .X(n13899) );
  nand_x1_sg U13148 ( .A(n16608), .B(n16753), .X(n13865) );
  nand_x1_sg U13149 ( .A(n16606), .B(n16755), .X(n13845) );
  nand_x1_sg U13150 ( .A(n16602), .B(n16753), .X(n13893) );
  nand_x1_sg U13151 ( .A(n16590), .B(n16755), .X(n13837) );
  nand_x1_sg U13152 ( .A(n16586), .B(n16755), .X(n13841) );
  nand_x1_sg U13153 ( .A(n16580), .B(n16755), .X(n13839) );
  nand_x1_sg U13154 ( .A(n16576), .B(n16757), .X(n13941) );
  nand_x1_sg U13155 ( .A(n16574), .B(n16747), .X(n13923) );
  nand_x1_sg U13156 ( .A(n16552), .B(n16753), .X(n13873) );
  nand_x1_sg U13157 ( .A(n16550), .B(n16753), .X(n13871) );
  nand_x1_sg U13158 ( .A(n16548), .B(n16754), .X(n13851) );
  nand_x1_sg U13159 ( .A(n16546), .B(n16754), .X(n13857) );
  nand_x1_sg U13160 ( .A(n16540), .B(n16754), .X(n13853) );
  nand_x1_sg U13161 ( .A(n16534), .B(n16754), .X(n13855) );
  nand_x1_sg U13162 ( .A(n16532), .B(n16754), .X(n13847) );
  nand_x1_sg U13163 ( .A(n16530), .B(n16753), .X(n13875) );
  nand_x1_sg U13164 ( .A(n16524), .B(n16754), .X(n13849) );
  nand_x1_sg U13165 ( .A(n16496), .B(n16754), .X(n13881) );
  nand_x1_sg U13166 ( .A(n16494), .B(n16754), .X(n13859) );
  nand_x1_sg U13167 ( .A(n16490), .B(n16755), .X(n13891) );
  nand_x1_sg U13168 ( .A(n16476), .B(n16755), .X(n13829) );
  nand_x1_sg U13169 ( .A(n16474), .B(n16755), .X(n13833) );
  nand_x1_sg U13170 ( .A(n16468), .B(n16755), .X(n13835) );
  nand_x1_sg U13171 ( .A(n16452), .B(n16754), .X(n13861) );
  nand_x1_sg U13172 ( .A(n16450), .B(n16753), .X(n13863) );
  nand_x1_sg U13173 ( .A(n16432), .B(n16745), .X(n13883) );
  nand_x1_sg U13174 ( .A(n16430), .B(n16747), .X(n13885) );
  nand_x1_sg U13175 ( .A(n16428), .B(n16753), .X(n13877) );
  nand_x1_sg U13176 ( .A(n16426), .B(n16747), .X(n13879) );
  nand_x1_sg U13177 ( .A(n16424), .B(n16748), .X(n13887) );
  nand_x1_sg U13178 ( .A(n16422), .B(n16755), .X(n13843) );
  nand_x1_sg U13179 ( .A(n16416), .B(n16749), .X(n13889) );
  nand_x1_sg U13180 ( .A(n16414), .B(n16753), .X(n13917) );
  nand_x1_sg U13181 ( .A(n16412), .B(n16757), .X(n13929) );
  nand_x1_sg U13182 ( .A(n16410), .B(n16757), .X(n13935) );
  nand_x1_sg U13183 ( .A(n16404), .B(n16751), .X(n13905) );
  nand_x1_sg U13184 ( .A(n16396), .B(n16757), .X(n13911) );
  nand_x1_sg U13185 ( .A(n16376), .B(n16754), .X(n13947) );
  nand_x1_sg U13186 ( .A(n16374), .B(n16757), .X(n13953) );
  nand_x1_sg U13187 ( .A(n16372), .B(n16753), .X(n13869) );
  nand_x1_sg U13188 ( .A(n16364), .B(n16753), .X(n13867) );
  nand_x1_sg U13189 ( .A(n16168), .B(n16757), .X(n13925) );
  nand_x1_sg U13190 ( .A(n16166), .B(n16757), .X(n13927) );
  nand_x1_sg U13191 ( .A(n16164), .B(n16745), .X(n13919) );
  nand_x1_sg U13192 ( .A(n16162), .B(n16748), .X(n13921) );
  nand_x1_sg U13193 ( .A(n16160), .B(n16759), .X(n13937) );
  nand_x1_sg U13194 ( .A(n16158), .B(n16745), .X(n13939) );
  nand_x1_sg U13195 ( .A(n16156), .B(n16746), .X(n13931) );
  nand_x1_sg U13196 ( .A(n16154), .B(n16757), .X(n13933) );
  nand_x1_sg U13197 ( .A(n16152), .B(n16750), .X(n13901) );
  nand_x1_sg U13198 ( .A(n16150), .B(n16757), .X(n13903) );
  nand_x1_sg U13199 ( .A(n16148), .B(n16757), .X(n13895) );
  nand_x1_sg U13200 ( .A(n16146), .B(n16759), .X(n13897) );
  nand_x1_sg U13201 ( .A(n16144), .B(n16757), .X(n13913) );
  nand_x1_sg U13202 ( .A(n16142), .B(n16757), .X(n13915) );
  nand_x1_sg U13203 ( .A(n16140), .B(n16757), .X(n13907) );
  nand_x1_sg U13204 ( .A(n16138), .B(n16757), .X(n13909) );
  nand_x1_sg U13205 ( .A(n16120), .B(n16751), .X(n13949) );
  nand_x1_sg U13206 ( .A(n16118), .B(n16752), .X(n13951) );
  nand_x1_sg U13207 ( .A(n16116), .B(n16749), .X(n13943) );
  nand_x1_sg U13208 ( .A(n16114), .B(n16757), .X(n13945) );
  nand_x1_sg U13209 ( .A(n16108), .B(n16747), .X(n13955) );
  nand_x1_sg U13210 ( .A(n16106), .B(n16747), .X(n13957) );
  nand_x1_sg U13211 ( .A(n14474), .B(state[1]), .X(n14473) );
  nand_x1_sg U13212 ( .A(n18399), .B(input_ready), .X(n14482) );
  nand_x1_sg U13213 ( .A(n14474), .B(state[0]), .X(n14476) );
  nand_x1_sg U13214 ( .A(n14478), .B(n14472), .X(n14477) );
  nor_x1_sg U13215 ( .A(n16734), .B(n14474), .X(n14478) );
  nor_x1_sg U13216 ( .A(n16730), .B(n16733), .X(n3869) );
  nor_x1_sg U13217 ( .A(n16728), .B(n16733), .X(n5145) );
  nor_x1_sg U13218 ( .A(n16726), .B(n16733), .X(n5141) );
  nor_x1_sg U13219 ( .A(n16724), .B(n16733), .X(n5137) );
  nor_x1_sg U13220 ( .A(n16722), .B(n16733), .X(n5133) );
  nor_x1_sg U13221 ( .A(n16720), .B(n16733), .X(n5129) );
  nor_x1_sg U13222 ( .A(n16718), .B(n16733), .X(n5125) );
  nor_x1_sg U13223 ( .A(n16716), .B(n16733), .X(n5121) );
  nor_x1_sg U13224 ( .A(n16714), .B(n16733), .X(n5117) );
  nor_x1_sg U13225 ( .A(n16712), .B(n16733), .X(n5113) );
  nor_x1_sg U13226 ( .A(n16710), .B(n16733), .X(n5109) );
  nor_x1_sg U13227 ( .A(n16708), .B(n16733), .X(n5105) );
  nor_x1_sg U13228 ( .A(n16706), .B(n16733), .X(n5101) );
  nor_x1_sg U13229 ( .A(n16704), .B(n16733), .X(n5097) );
  nor_x1_sg U13230 ( .A(n16702), .B(n16733), .X(n5093) );
  nor_x1_sg U13231 ( .A(n16700), .B(n16733), .X(n5089) );
  nor_x1_sg U13232 ( .A(n16698), .B(n16733), .X(n5085) );
  nor_x1_sg U13233 ( .A(n16696), .B(n16733), .X(n5081) );
  nor_x1_sg U13234 ( .A(n16694), .B(n16733), .X(n5077) );
  nor_x1_sg U13235 ( .A(n16692), .B(n16733), .X(n5073) );
  nor_x1_sg U13236 ( .A(n16570), .B(n16733), .X(n5069) );
  nor_x1_sg U13237 ( .A(n16568), .B(n16733), .X(n5065) );
  nor_x1_sg U13238 ( .A(n16566), .B(n16733), .X(n5061) );
  nor_x1_sg U13239 ( .A(n16564), .B(n16733), .X(n5057) );
  nor_x1_sg U13240 ( .A(n16562), .B(n16733), .X(n5053) );
  nor_x1_sg U13241 ( .A(n16560), .B(n16733), .X(n5049) );
  nor_x1_sg U13242 ( .A(n16558), .B(n16733), .X(n5045) );
  nor_x1_sg U13243 ( .A(n16556), .B(n16733), .X(n5041) );
  nor_x1_sg U13244 ( .A(n16554), .B(n16733), .X(n5037) );
  nor_x1_sg U13245 ( .A(n16552), .B(n16733), .X(n5033) );
  nor_x1_sg U13246 ( .A(n16550), .B(n16733), .X(n5029) );
  nor_x1_sg U13247 ( .A(n16548), .B(n16733), .X(n5025) );
  nor_x1_sg U13248 ( .A(n16546), .B(n16733), .X(n5021) );
  nor_x1_sg U13249 ( .A(n16544), .B(n16733), .X(n5017) );
  nor_x1_sg U13250 ( .A(n16542), .B(n16733), .X(n5013) );
  nor_x1_sg U13251 ( .A(n16540), .B(n16733), .X(n5009) );
  nor_x1_sg U13252 ( .A(n16538), .B(n16733), .X(n5005) );
  nor_x1_sg U13253 ( .A(n16536), .B(n16733), .X(n5001) );
  nor_x1_sg U13254 ( .A(n16534), .B(n16733), .X(n4997) );
  nor_x1_sg U13255 ( .A(n16532), .B(n16733), .X(n4993) );
  nor_x1_sg U13256 ( .A(n16410), .B(n16733), .X(n4989) );
  nor_x1_sg U13257 ( .A(n16408), .B(n16733), .X(n4985) );
  nor_x1_sg U13258 ( .A(n16406), .B(n16733), .X(n4981) );
  nor_x1_sg U13259 ( .A(n16404), .B(n16733), .X(n4977) );
  nor_x1_sg U13260 ( .A(n16402), .B(n16733), .X(n4973) );
  nor_x1_sg U13261 ( .A(n16400), .B(n16733), .X(n4969) );
  nor_x1_sg U13262 ( .A(n16398), .B(n16733), .X(n4965) );
  nor_x1_sg U13263 ( .A(n16396), .B(n16733), .X(n4961) );
  nor_x1_sg U13264 ( .A(n16394), .B(n16733), .X(n4957) );
  nor_x1_sg U13265 ( .A(n16392), .B(n16733), .X(n4953) );
  nor_x1_sg U13266 ( .A(n16390), .B(n16733), .X(n4949) );
  nor_x1_sg U13267 ( .A(n16388), .B(n16733), .X(n4945) );
  nor_x1_sg U13268 ( .A(n16386), .B(n16733), .X(n4941) );
  nor_x1_sg U13269 ( .A(n16384), .B(n16733), .X(n4937) );
  nor_x1_sg U13270 ( .A(n16382), .B(n16733), .X(n4933) );
  nor_x1_sg U13271 ( .A(n16380), .B(n16733), .X(n4929) );
  nor_x1_sg U13272 ( .A(n16378), .B(n16733), .X(n4925) );
  nor_x1_sg U13273 ( .A(n16376), .B(n16733), .X(n4921) );
  nor_x1_sg U13274 ( .A(n16374), .B(n16733), .X(n4917) );
  nor_x1_sg U13275 ( .A(n16372), .B(n16733), .X(n4913) );
  nor_x1_sg U13276 ( .A(n16250), .B(n16733), .X(n4909) );
  nor_x1_sg U13277 ( .A(n16248), .B(n16733), .X(n4905) );
  nor_x1_sg U13278 ( .A(n16246), .B(n16733), .X(n4901) );
  nor_x1_sg U13279 ( .A(n16244), .B(n16733), .X(n4897) );
  nor_x1_sg U13280 ( .A(n16242), .B(n16733), .X(n4893) );
  nor_x1_sg U13281 ( .A(n16240), .B(n16733), .X(n4889) );
  nor_x1_sg U13282 ( .A(n16238), .B(n16733), .X(n4885) );
  nor_x1_sg U13283 ( .A(n16236), .B(n16733), .X(n4881) );
  nor_x1_sg U13284 ( .A(n16234), .B(n16733), .X(n4877) );
  nor_x1_sg U13285 ( .A(n16232), .B(n16733), .X(n4873) );
  nor_x1_sg U13286 ( .A(n16230), .B(n16733), .X(n4869) );
  nor_x1_sg U13287 ( .A(n16228), .B(n16733), .X(n4865) );
  nor_x1_sg U13288 ( .A(n16226), .B(n16733), .X(n4861) );
  nor_x1_sg U13289 ( .A(n16224), .B(n16733), .X(n4857) );
  nor_x1_sg U13290 ( .A(n16222), .B(n16733), .X(n4853) );
  nor_x1_sg U13291 ( .A(n16220), .B(n16733), .X(n4849) );
  nor_x1_sg U13292 ( .A(n16218), .B(n16733), .X(n4845) );
  nor_x1_sg U13293 ( .A(n16216), .B(n16733), .X(n4841) );
  nor_x1_sg U13294 ( .A(n16214), .B(n16733), .X(n4837) );
  nor_x1_sg U13295 ( .A(n16212), .B(n16733), .X(n4833) );
  nor_x1_sg U13296 ( .A(n16690), .B(n16733), .X(n4829) );
  nor_x1_sg U13297 ( .A(n16688), .B(n16733), .X(n4825) );
  nor_x1_sg U13298 ( .A(n16686), .B(n16733), .X(n4821) );
  nor_x1_sg U13299 ( .A(n16684), .B(n16733), .X(n4817) );
  nor_x1_sg U13300 ( .A(n16682), .B(n16733), .X(n4813) );
  nor_x1_sg U13301 ( .A(n16680), .B(n16733), .X(n4809) );
  nor_x1_sg U13302 ( .A(n16678), .B(n16733), .X(n4805) );
  nor_x1_sg U13303 ( .A(n16676), .B(n16733), .X(n4801) );
  nor_x1_sg U13304 ( .A(n16674), .B(n16733), .X(n4797) );
  nor_x1_sg U13305 ( .A(n16672), .B(n16733), .X(n4793) );
  nor_x1_sg U13306 ( .A(n16670), .B(n16733), .X(n4789) );
  nor_x1_sg U13307 ( .A(n16668), .B(n16733), .X(n4785) );
  nor_x1_sg U13308 ( .A(n16666), .B(n16733), .X(n4781) );
  nor_x1_sg U13309 ( .A(n16664), .B(n16733), .X(n4777) );
  nor_x1_sg U13310 ( .A(n16662), .B(n16733), .X(n4773) );
  nor_x1_sg U13311 ( .A(n16660), .B(n16733), .X(n4769) );
  nor_x1_sg U13312 ( .A(n16658), .B(n16733), .X(n4765) );
  nor_x1_sg U13313 ( .A(n16656), .B(n16733), .X(n4761) );
  nor_x1_sg U13314 ( .A(n16654), .B(n16733), .X(n4757) );
  nor_x1_sg U13315 ( .A(n16652), .B(n16733), .X(n4753) );
  nor_x1_sg U13316 ( .A(n16530), .B(n16733), .X(n4749) );
  nor_x1_sg U13317 ( .A(n16528), .B(n16733), .X(n4745) );
  nor_x1_sg U13318 ( .A(n16526), .B(n16733), .X(n4741) );
  nor_x1_sg U13319 ( .A(n16524), .B(n16733), .X(n4737) );
  nor_x1_sg U13320 ( .A(n16522), .B(n16733), .X(n4733) );
  nor_x1_sg U13321 ( .A(n16520), .B(n16733), .X(n4729) );
  nor_x1_sg U13322 ( .A(n16518), .B(n16733), .X(n4725) );
  nor_x1_sg U13323 ( .A(n16516), .B(n16733), .X(n4721) );
  nor_x1_sg U13324 ( .A(n16514), .B(n16733), .X(n4717) );
  nor_x1_sg U13325 ( .A(n16512), .B(n16733), .X(n4713) );
  nor_x1_sg U13326 ( .A(n16510), .B(n16733), .X(n4709) );
  nor_x1_sg U13327 ( .A(n16508), .B(n16733), .X(n4705) );
  nor_x1_sg U13328 ( .A(n16506), .B(n16733), .X(n4701) );
  nor_x1_sg U13329 ( .A(n16504), .B(n16733), .X(n4697) );
  nor_x1_sg U13330 ( .A(n16502), .B(n16733), .X(n4693) );
  nor_x1_sg U13331 ( .A(n16500), .B(n16733), .X(n4689) );
  nor_x1_sg U13332 ( .A(n16498), .B(n16733), .X(n4685) );
  nor_x1_sg U13333 ( .A(n16496), .B(n16733), .X(n4681) );
  nor_x1_sg U13334 ( .A(n16494), .B(n16733), .X(n4677) );
  nor_x1_sg U13335 ( .A(n16492), .B(n16733), .X(n4673) );
  nor_x1_sg U13336 ( .A(n16370), .B(n16733), .X(n4669) );
  nor_x1_sg U13337 ( .A(n16368), .B(n16733), .X(n4665) );
  nor_x1_sg U13338 ( .A(n16366), .B(n16733), .X(n4661) );
  nor_x1_sg U13339 ( .A(n16364), .B(n16733), .X(n4657) );
  nor_x1_sg U13340 ( .A(n16362), .B(n16733), .X(n4653) );
  nor_x1_sg U13341 ( .A(n16360), .B(n16733), .X(n4649) );
  nor_x1_sg U13342 ( .A(n16358), .B(n16733), .X(n4645) );
  nor_x1_sg U13343 ( .A(n16356), .B(n16733), .X(n4641) );
  nor_x1_sg U13344 ( .A(n16354), .B(n16733), .X(n4637) );
  nor_x1_sg U13345 ( .A(n16352), .B(n16733), .X(n4633) );
  nor_x1_sg U13346 ( .A(n16350), .B(n16733), .X(n4629) );
  nor_x1_sg U13347 ( .A(n16348), .B(n16733), .X(n4625) );
  nor_x1_sg U13348 ( .A(n16346), .B(n16733), .X(n4621) );
  nor_x1_sg U13349 ( .A(n16344), .B(n16733), .X(n4617) );
  nor_x1_sg U13350 ( .A(n16342), .B(n16733), .X(n4613) );
  nor_x1_sg U13351 ( .A(n16340), .B(n16733), .X(n4609) );
  nor_x1_sg U13352 ( .A(n16338), .B(n16733), .X(n4605) );
  nor_x1_sg U13353 ( .A(n16336), .B(n16733), .X(n4601) );
  nor_x1_sg U13354 ( .A(n16334), .B(n16733), .X(n4597) );
  nor_x1_sg U13355 ( .A(n16332), .B(n16733), .X(n4593) );
  nor_x1_sg U13356 ( .A(n16210), .B(n16733), .X(n4589) );
  nor_x1_sg U13357 ( .A(n16208), .B(n16733), .X(n4585) );
  nor_x1_sg U13358 ( .A(n16206), .B(n16733), .X(n4581) );
  nor_x1_sg U13359 ( .A(n16204), .B(n16733), .X(n4577) );
  nor_x1_sg U13360 ( .A(n16202), .B(n16733), .X(n4573) );
  nor_x1_sg U13361 ( .A(n16200), .B(n16733), .X(n4569) );
  nor_x1_sg U13362 ( .A(n16198), .B(n16733), .X(n4565) );
  nor_x1_sg U13363 ( .A(n16196), .B(n16733), .X(n4561) );
  nor_x1_sg U13364 ( .A(n16194), .B(n16733), .X(n4557) );
  nor_x1_sg U13365 ( .A(n16192), .B(n16733), .X(n4553) );
  nor_x1_sg U13366 ( .A(n16190), .B(n16733), .X(n4549) );
  nor_x1_sg U13367 ( .A(n16188), .B(n16733), .X(n4545) );
  nor_x1_sg U13368 ( .A(n16186), .B(n16733), .X(n4541) );
  nor_x1_sg U13369 ( .A(n16184), .B(n16733), .X(n4537) );
  nor_x1_sg U13370 ( .A(n16182), .B(n16733), .X(n4533) );
  nor_x1_sg U13371 ( .A(n16180), .B(n16733), .X(n4529) );
  nor_x1_sg U13372 ( .A(n16178), .B(n16733), .X(n4525) );
  nor_x1_sg U13373 ( .A(n16176), .B(n16733), .X(n4521) );
  nor_x1_sg U13374 ( .A(n16174), .B(n16733), .X(n4517) );
  nor_x1_sg U13375 ( .A(n16172), .B(n16733), .X(n4513) );
  nor_x1_sg U13376 ( .A(n16650), .B(n16733), .X(n4509) );
  nor_x1_sg U13377 ( .A(n16648), .B(n16733), .X(n4505) );
  nor_x1_sg U13378 ( .A(n16646), .B(n16733), .X(n4501) );
  nor_x1_sg U13379 ( .A(n16644), .B(n16733), .X(n4497) );
  nor_x1_sg U13380 ( .A(n16642), .B(n16733), .X(n4493) );
  nor_x1_sg U13381 ( .A(n16640), .B(n16733), .X(n4489) );
  nor_x1_sg U13382 ( .A(n16638), .B(n16733), .X(n4485) );
  nor_x1_sg U13383 ( .A(n16636), .B(n16733), .X(n4481) );
  nor_x1_sg U13384 ( .A(n16634), .B(n16733), .X(n4477) );
  nor_x1_sg U13385 ( .A(n16632), .B(n16733), .X(n4473) );
  nor_x1_sg U13386 ( .A(n16630), .B(n16733), .X(n4469) );
  nor_x1_sg U13387 ( .A(n16628), .B(n16733), .X(n4465) );
  nor_x1_sg U13388 ( .A(n16626), .B(n16733), .X(n4461) );
  nor_x1_sg U13389 ( .A(n16624), .B(n16733), .X(n4457) );
  nor_x1_sg U13390 ( .A(n16622), .B(n16733), .X(n4453) );
  nor_x1_sg U13391 ( .A(n16620), .B(n16733), .X(n4449) );
  nor_x1_sg U13392 ( .A(n16618), .B(n16733), .X(n4445) );
  nor_x1_sg U13393 ( .A(n16616), .B(n16733), .X(n4441) );
  nor_x1_sg U13394 ( .A(n16614), .B(n16733), .X(n4437) );
  nor_x1_sg U13395 ( .A(n16612), .B(n16733), .X(n4433) );
  nor_x1_sg U13396 ( .A(n16490), .B(n16733), .X(n4429) );
  nor_x1_sg U13397 ( .A(n16488), .B(n16733), .X(n4425) );
  nor_x1_sg U13398 ( .A(n16486), .B(n16733), .X(n4421) );
  nor_x1_sg U13399 ( .A(n16484), .B(n16733), .X(n4417) );
  nor_x1_sg U13400 ( .A(n16482), .B(n16733), .X(n4413) );
  nor_x1_sg U13401 ( .A(n16480), .B(n16733), .X(n4409) );
  nor_x1_sg U13402 ( .A(n16478), .B(n16733), .X(n4405) );
  nor_x1_sg U13403 ( .A(n16476), .B(n16733), .X(n4401) );
  nor_x1_sg U13404 ( .A(n16474), .B(n16733), .X(n4397) );
  nor_x1_sg U13405 ( .A(n16472), .B(n16733), .X(n4393) );
  nor_x1_sg U13406 ( .A(n16470), .B(n16733), .X(n4389) );
  nor_x1_sg U13407 ( .A(n16468), .B(n16733), .X(n4385) );
  nor_x1_sg U13408 ( .A(n16466), .B(n16733), .X(n4381) );
  nor_x1_sg U13409 ( .A(n16464), .B(n16733), .X(n4377) );
  nor_x1_sg U13410 ( .A(n16462), .B(n16733), .X(n4373) );
  nor_x1_sg U13411 ( .A(n16460), .B(n16733), .X(n4369) );
  nor_x1_sg U13412 ( .A(n16458), .B(n16733), .X(n4365) );
  nor_x1_sg U13413 ( .A(n16456), .B(n16733), .X(n4361) );
  nor_x1_sg U13414 ( .A(n16454), .B(n16733), .X(n4357) );
  nor_x1_sg U13415 ( .A(n16452), .B(n16733), .X(n4353) );
  nor_x1_sg U13416 ( .A(n16330), .B(n16733), .X(n4349) );
  nor_x1_sg U13417 ( .A(n16328), .B(n16733), .X(n4345) );
  nor_x1_sg U13418 ( .A(n16326), .B(n16733), .X(n4341) );
  nor_x1_sg U13419 ( .A(n16324), .B(n16733), .X(n4337) );
  nor_x1_sg U13420 ( .A(n16322), .B(n16733), .X(n4333) );
  nor_x1_sg U13421 ( .A(n16320), .B(n16733), .X(n4329) );
  nor_x1_sg U13422 ( .A(n16318), .B(n16733), .X(n4325) );
  nor_x1_sg U13423 ( .A(n16316), .B(n16733), .X(n4321) );
  nor_x1_sg U13424 ( .A(n16314), .B(n16733), .X(n4317) );
  nor_x1_sg U13425 ( .A(n16312), .B(n16733), .X(n4313) );
  nor_x1_sg U13426 ( .A(n16310), .B(n16733), .X(n4309) );
  nor_x1_sg U13427 ( .A(n16308), .B(n16733), .X(n4305) );
  nor_x1_sg U13428 ( .A(n16306), .B(n16733), .X(n4301) );
  nor_x1_sg U13429 ( .A(n16304), .B(n16733), .X(n4297) );
  nor_x1_sg U13430 ( .A(n16302), .B(n16733), .X(n4293) );
  nor_x1_sg U13431 ( .A(n16300), .B(n16733), .X(n4289) );
  nor_x1_sg U13432 ( .A(n16298), .B(n16733), .X(n4285) );
  nor_x1_sg U13433 ( .A(n16296), .B(n16733), .X(n4281) );
  nor_x1_sg U13434 ( .A(n16294), .B(n16733), .X(n4277) );
  nor_x1_sg U13435 ( .A(n16292), .B(n16733), .X(n4273) );
  nor_x1_sg U13436 ( .A(n16170), .B(n16733), .X(n4269) );
  nor_x1_sg U13437 ( .A(n16168), .B(n16733), .X(n4265) );
  nor_x1_sg U13438 ( .A(n16166), .B(n16733), .X(n4261) );
  nor_x1_sg U13439 ( .A(n16164), .B(n16733), .X(n4257) );
  nor_x1_sg U13440 ( .A(n16162), .B(n16733), .X(n4253) );
  nor_x1_sg U13441 ( .A(n16160), .B(n16733), .X(n4249) );
  nor_x1_sg U13442 ( .A(n16158), .B(n16733), .X(n4245) );
  nor_x1_sg U13443 ( .A(n16156), .B(n16733), .X(n4241) );
  nor_x1_sg U13444 ( .A(n16154), .B(n16733), .X(n4237) );
  nor_x1_sg U13445 ( .A(n16152), .B(n16733), .X(n4233) );
  nor_x1_sg U13446 ( .A(n16150), .B(n16733), .X(n4229) );
  nor_x1_sg U13447 ( .A(n16148), .B(n16733), .X(n4225) );
  nor_x1_sg U13448 ( .A(n16146), .B(n16733), .X(n4221) );
  nor_x1_sg U13449 ( .A(n16144), .B(n16733), .X(n4217) );
  nor_x1_sg U13450 ( .A(n16142), .B(n16733), .X(n4213) );
  nor_x1_sg U13451 ( .A(n16140), .B(n16733), .X(n4209) );
  nor_x1_sg U13452 ( .A(n16138), .B(n16733), .X(n4205) );
  nor_x1_sg U13453 ( .A(n16136), .B(n16733), .X(n4201) );
  nor_x1_sg U13454 ( .A(n16134), .B(n16733), .X(n4197) );
  nor_x1_sg U13455 ( .A(n16132), .B(n16733), .X(n4193) );
  nor_x1_sg U13456 ( .A(n16610), .B(n16733), .X(n4189) );
  nor_x1_sg U13457 ( .A(n16608), .B(n16733), .X(n4185) );
  nor_x1_sg U13458 ( .A(n16606), .B(n16733), .X(n4181) );
  nor_x1_sg U13459 ( .A(n16604), .B(n16733), .X(n4177) );
  nor_x1_sg U13460 ( .A(n16602), .B(n16733), .X(n4173) );
  nor_x1_sg U13461 ( .A(n16600), .B(n16733), .X(n4169) );
  nor_x1_sg U13462 ( .A(n16598), .B(n16733), .X(n4165) );
  nor_x1_sg U13463 ( .A(n16596), .B(n16733), .X(n4161) );
  nor_x1_sg U13464 ( .A(n16594), .B(n16733), .X(n4157) );
  nor_x1_sg U13465 ( .A(n16592), .B(n16733), .X(n4153) );
  nor_x1_sg U13466 ( .A(n16590), .B(n16733), .X(n4149) );
  nor_x1_sg U13467 ( .A(n16588), .B(n16733), .X(n4145) );
  nor_x1_sg U13468 ( .A(n16586), .B(n16733), .X(n4141) );
  nor_x1_sg U13469 ( .A(n16584), .B(n16733), .X(n4137) );
  nor_x1_sg U13470 ( .A(n16582), .B(n16733), .X(n4133) );
  nor_x1_sg U13471 ( .A(n16580), .B(n16733), .X(n4129) );
  nor_x1_sg U13472 ( .A(n16578), .B(n16733), .X(n4125) );
  nor_x1_sg U13473 ( .A(n16576), .B(n16733), .X(n4121) );
  nor_x1_sg U13474 ( .A(n16574), .B(n16733), .X(n4117) );
  nor_x1_sg U13475 ( .A(n16572), .B(n16733), .X(n4113) );
  nor_x1_sg U13476 ( .A(n16450), .B(n16733), .X(n4109) );
  nor_x1_sg U13477 ( .A(n16448), .B(n16733), .X(n4105) );
  nor_x1_sg U13478 ( .A(n16446), .B(n16733), .X(n4101) );
  nor_x1_sg U13479 ( .A(n16444), .B(n16733), .X(n4097) );
  nor_x1_sg U13480 ( .A(n16442), .B(n16733), .X(n4093) );
  nor_x1_sg U13481 ( .A(n16440), .B(n16733), .X(n4089) );
  nor_x1_sg U13482 ( .A(n16438), .B(n16733), .X(n4085) );
  nor_x1_sg U13483 ( .A(n16436), .B(n16733), .X(n4081) );
  nor_x1_sg U13484 ( .A(n16434), .B(n16733), .X(n4077) );
  nor_x1_sg U13485 ( .A(n16432), .B(n16733), .X(n4073) );
  nor_x1_sg U13486 ( .A(n16430), .B(n16733), .X(n4069) );
  nor_x1_sg U13487 ( .A(n16428), .B(n16733), .X(n4065) );
  nor_x1_sg U13488 ( .A(n16426), .B(n16733), .X(n4061) );
  nor_x1_sg U13489 ( .A(n16424), .B(n16733), .X(n4057) );
  nor_x1_sg U13490 ( .A(n16422), .B(n16733), .X(n4053) );
  nor_x1_sg U13491 ( .A(n16420), .B(n16733), .X(n4049) );
  nor_x1_sg U13492 ( .A(n16418), .B(n16733), .X(n4045) );
  nor_x1_sg U13493 ( .A(n16416), .B(n16733), .X(n4041) );
  nor_x1_sg U13494 ( .A(n16414), .B(n16733), .X(n4037) );
  nor_x1_sg U13495 ( .A(n16412), .B(n16733), .X(n4033) );
  nor_x1_sg U13496 ( .A(n16290), .B(n16733), .X(n4029) );
  nor_x1_sg U13497 ( .A(n16288), .B(n16733), .X(n4025) );
  nor_x1_sg U13498 ( .A(n16286), .B(n16733), .X(n4021) );
  nor_x1_sg U13499 ( .A(n16284), .B(n16733), .X(n4017) );
  nor_x1_sg U13500 ( .A(n16282), .B(n16733), .X(n4013) );
  nor_x1_sg U13501 ( .A(n16280), .B(n16733), .X(n4009) );
  nor_x1_sg U13502 ( .A(n16278), .B(n16733), .X(n4005) );
  nor_x1_sg U13503 ( .A(n16276), .B(n16733), .X(n4001) );
  nor_x1_sg U13504 ( .A(n16274), .B(n16733), .X(n3997) );
  nor_x1_sg U13505 ( .A(n16272), .B(n16733), .X(n3993) );
  nor_x1_sg U13506 ( .A(n16270), .B(n16733), .X(n3989) );
  nor_x1_sg U13507 ( .A(n16268), .B(n16733), .X(n3985) );
  nor_x1_sg U13508 ( .A(n16266), .B(n16733), .X(n3981) );
  nor_x1_sg U13509 ( .A(n16264), .B(n16733), .X(n3977) );
  nor_x1_sg U13510 ( .A(n16262), .B(n16733), .X(n3973) );
  nor_x1_sg U13511 ( .A(n16260), .B(n16733), .X(n3969) );
  nor_x1_sg U13512 ( .A(n16258), .B(n16733), .X(n3965) );
  nor_x1_sg U13513 ( .A(n16256), .B(n16733), .X(n3961) );
  nor_x1_sg U13514 ( .A(n16254), .B(n16733), .X(n3957) );
  nor_x1_sg U13515 ( .A(n16252), .B(n16733), .X(n3953) );
  nor_x1_sg U13516 ( .A(n16130), .B(n16733), .X(n3949) );
  nor_x1_sg U13517 ( .A(n16128), .B(n16733), .X(n3945) );
  nor_x1_sg U13518 ( .A(n16126), .B(n16733), .X(n3941) );
  nor_x1_sg U13519 ( .A(n16124), .B(n16733), .X(n3937) );
  nor_x1_sg U13520 ( .A(n16122), .B(n16733), .X(n3933) );
  nor_x1_sg U13521 ( .A(n16120), .B(n16733), .X(n3929) );
  nor_x1_sg U13522 ( .A(n16118), .B(n16733), .X(n3925) );
  nor_x1_sg U13523 ( .A(n16116), .B(n16733), .X(n3921) );
  nor_x1_sg U13524 ( .A(n16114), .B(n16733), .X(n3917) );
  nor_x1_sg U13525 ( .A(n16112), .B(n16733), .X(n3913) );
  nor_x1_sg U13526 ( .A(n16110), .B(n16733), .X(n3909) );
  nor_x1_sg U13527 ( .A(n16108), .B(n16733), .X(n3905) );
  nor_x1_sg U13528 ( .A(n16106), .B(n16733), .X(n3901) );
  nor_x1_sg U13529 ( .A(n16104), .B(n16733), .X(n3897) );
  nor_x1_sg U13530 ( .A(n16102), .B(n16733), .X(n3893) );
  nor_x1_sg U13531 ( .A(n16100), .B(n16733), .X(n3889) );
  nor_x1_sg U13532 ( .A(n16098), .B(n16733), .X(n3885) );
  nor_x1_sg U13533 ( .A(n16096), .B(n16733), .X(n3881) );
  nor_x1_sg U13534 ( .A(n16094), .B(n16733), .X(n3877) );
  nor_x1_sg U13535 ( .A(n16092), .B(n16733), .X(n3873) );
  nand_x1_sg U13536 ( .A(n16735), .B(n16730), .X(n12859) );
  nand_x1_sg U13537 ( .A(n16735), .B(n16728), .X(n12540) );
  nand_x1_sg U13538 ( .A(n16735), .B(n16726), .X(n12541) );
  nand_x1_sg U13539 ( .A(n16735), .B(n16724), .X(n12542) );
  nand_x1_sg U13540 ( .A(n16735), .B(n16722), .X(n12543) );
  nand_x1_sg U13541 ( .A(n16735), .B(n16720), .X(n12544) );
  nand_x1_sg U13542 ( .A(n16735), .B(n16718), .X(n12545) );
  nand_x1_sg U13543 ( .A(n16735), .B(n16716), .X(n12546) );
  nand_x1_sg U13544 ( .A(n16735), .B(n16714), .X(n12547) );
  nand_x1_sg U13545 ( .A(n16735), .B(n16712), .X(n12548) );
  nand_x1_sg U13546 ( .A(n16735), .B(n16710), .X(n12549) );
  nand_x1_sg U13547 ( .A(n16735), .B(n16708), .X(n12550) );
  nand_x1_sg U13548 ( .A(n16735), .B(n16706), .X(n12551) );
  nand_x1_sg U13549 ( .A(n16735), .B(n16704), .X(n12552) );
  nand_x1_sg U13550 ( .A(n16735), .B(n16702), .X(n12553) );
  nand_x1_sg U13551 ( .A(n16735), .B(n16700), .X(n12554) );
  nand_x1_sg U13552 ( .A(n16735), .B(n16698), .X(n12555) );
  nand_x1_sg U13553 ( .A(n16735), .B(n16696), .X(n12556) );
  nand_x1_sg U13554 ( .A(n16735), .B(n16694), .X(n12557) );
  nand_x1_sg U13555 ( .A(n16735), .B(n16692), .X(n12558) );
  nand_x1_sg U13556 ( .A(n16735), .B(n16570), .X(n12559) );
  nand_x1_sg U13557 ( .A(n16735), .B(n16568), .X(n12560) );
  nand_x1_sg U13558 ( .A(n16735), .B(n16566), .X(n12561) );
  nand_x1_sg U13559 ( .A(n16735), .B(n16564), .X(n12562) );
  nand_x1_sg U13560 ( .A(n16735), .B(n16562), .X(n12563) );
  nand_x1_sg U13561 ( .A(n16735), .B(n16560), .X(n12564) );
  nand_x1_sg U13562 ( .A(n16735), .B(n16558), .X(n12565) );
  nand_x1_sg U13563 ( .A(n16735), .B(n16556), .X(n12566) );
  nand_x1_sg U13564 ( .A(n16735), .B(n16554), .X(n12567) );
  nand_x1_sg U13565 ( .A(n16735), .B(n16552), .X(n12568) );
  nand_x1_sg U13566 ( .A(n16735), .B(n16550), .X(n12569) );
  nand_x1_sg U13567 ( .A(n16735), .B(n16548), .X(n12570) );
  nand_x1_sg U13568 ( .A(n16735), .B(n16546), .X(n12571) );
  nand_x1_sg U13569 ( .A(n16735), .B(n16544), .X(n12572) );
  nand_x1_sg U13570 ( .A(n16735), .B(n16542), .X(n12573) );
  nand_x1_sg U13571 ( .A(n16735), .B(n16540), .X(n12574) );
  nand_x1_sg U13572 ( .A(n16735), .B(n16538), .X(n12575) );
  nand_x1_sg U13573 ( .A(n16735), .B(n16536), .X(n12576) );
  nand_x1_sg U13574 ( .A(n16735), .B(n16534), .X(n12577) );
  nand_x1_sg U13575 ( .A(n16735), .B(n16532), .X(n12578) );
  nand_x1_sg U13576 ( .A(n16735), .B(n16410), .X(n12579) );
  nand_x1_sg U13577 ( .A(n16735), .B(n16408), .X(n12580) );
  nand_x1_sg U13578 ( .A(n16735), .B(n16406), .X(n12581) );
  nand_x1_sg U13579 ( .A(n16735), .B(n16404), .X(n12582) );
  nand_x1_sg U13580 ( .A(n16735), .B(n16402), .X(n12583) );
  nand_x1_sg U13581 ( .A(n16735), .B(n16400), .X(n12584) );
  nand_x1_sg U13582 ( .A(n16735), .B(n16398), .X(n12585) );
  nand_x1_sg U13583 ( .A(n16735), .B(n16396), .X(n12586) );
  nand_x1_sg U13584 ( .A(n16735), .B(n16394), .X(n12587) );
  nand_x1_sg U13585 ( .A(n16735), .B(n16392), .X(n12588) );
  nand_x1_sg U13586 ( .A(n16735), .B(n16390), .X(n12589) );
  nand_x1_sg U13587 ( .A(n16735), .B(n16388), .X(n12590) );
  nand_x1_sg U13588 ( .A(n16735), .B(n16386), .X(n12591) );
  nand_x1_sg U13589 ( .A(n16735), .B(n16384), .X(n12592) );
  nand_x1_sg U13590 ( .A(n16735), .B(n16382), .X(n12593) );
  nand_x1_sg U13591 ( .A(n16735), .B(n16380), .X(n12594) );
  nand_x1_sg U13592 ( .A(n16735), .B(n16378), .X(n12595) );
  nand_x1_sg U13593 ( .A(n16735), .B(n16376), .X(n12596) );
  nand_x1_sg U13594 ( .A(n16735), .B(n16374), .X(n12597) );
  nand_x1_sg U13595 ( .A(n16735), .B(n16372), .X(n12598) );
  nand_x1_sg U13596 ( .A(n16735), .B(n16250), .X(n12599) );
  nand_x1_sg U13597 ( .A(n16735), .B(n16248), .X(n12600) );
  nand_x1_sg U13598 ( .A(n16735), .B(n16246), .X(n12601) );
  nand_x1_sg U13599 ( .A(n16735), .B(n16244), .X(n12602) );
  nand_x1_sg U13600 ( .A(n16735), .B(n16242), .X(n12603) );
  nand_x1_sg U13601 ( .A(n16735), .B(n16240), .X(n12604) );
  nand_x1_sg U13602 ( .A(n16735), .B(n16238), .X(n12605) );
  nand_x1_sg U13603 ( .A(n16735), .B(n16236), .X(n12606) );
  nand_x1_sg U13604 ( .A(n16735), .B(n16234), .X(n12607) );
  nand_x1_sg U13605 ( .A(n16735), .B(n16232), .X(n12608) );
  nand_x1_sg U13606 ( .A(n16735), .B(n16230), .X(n12609) );
  nand_x1_sg U13607 ( .A(n16735), .B(n16228), .X(n12610) );
  nand_x1_sg U13608 ( .A(n16735), .B(n16226), .X(n12611) );
  nand_x1_sg U13609 ( .A(n16735), .B(n16224), .X(n12612) );
  nand_x1_sg U13610 ( .A(n16735), .B(n16222), .X(n12613) );
  nand_x1_sg U13611 ( .A(n16735), .B(n16220), .X(n12614) );
  nand_x1_sg U13612 ( .A(n16735), .B(n16218), .X(n12615) );
  nand_x1_sg U13613 ( .A(n16735), .B(n16216), .X(n12616) );
  nand_x1_sg U13614 ( .A(n16735), .B(n16214), .X(n12617) );
  nand_x1_sg U13615 ( .A(n16735), .B(n16212), .X(n12618) );
  nand_x1_sg U13616 ( .A(n16735), .B(n16690), .X(n12619) );
  nand_x1_sg U13617 ( .A(n16735), .B(n16688), .X(n12620) );
  nand_x1_sg U13618 ( .A(n16735), .B(n16686), .X(n12621) );
  nand_x1_sg U13619 ( .A(n16735), .B(n16684), .X(n12622) );
  nand_x1_sg U13620 ( .A(n16735), .B(n16682), .X(n12623) );
  nand_x1_sg U13621 ( .A(n16735), .B(n16680), .X(n12624) );
  nand_x1_sg U13622 ( .A(n16735), .B(n16678), .X(n12625) );
  nand_x1_sg U13623 ( .A(n16735), .B(n16676), .X(n12626) );
  nand_x1_sg U13624 ( .A(n16735), .B(n16674), .X(n12627) );
  nand_x1_sg U13625 ( .A(n16735), .B(n16672), .X(n12628) );
  nand_x1_sg U13626 ( .A(n16735), .B(n16670), .X(n12629) );
  nand_x1_sg U13627 ( .A(n16735), .B(n16668), .X(n12630) );
  nand_x1_sg U13628 ( .A(n16735), .B(n16666), .X(n12631) );
  nand_x1_sg U13629 ( .A(n16735), .B(n16664), .X(n12632) );
  nand_x1_sg U13630 ( .A(n16735), .B(n16662), .X(n12633) );
  nand_x1_sg U13631 ( .A(n16735), .B(n16660), .X(n12634) );
  nand_x1_sg U13632 ( .A(n16735), .B(n16658), .X(n12635) );
  nand_x1_sg U13633 ( .A(n16735), .B(n16656), .X(n12636) );
  nand_x1_sg U13634 ( .A(n16735), .B(n16654), .X(n12637) );
  nand_x1_sg U13635 ( .A(n16735), .B(n16652), .X(n12638) );
  nand_x1_sg U13636 ( .A(n16735), .B(n16530), .X(n12639) );
  nand_x1_sg U13637 ( .A(n16735), .B(n16528), .X(n12640) );
  nand_x1_sg U13638 ( .A(n16735), .B(n16526), .X(n12641) );
  nand_x1_sg U13639 ( .A(n16735), .B(n16524), .X(n12642) );
  nand_x1_sg U13640 ( .A(n16735), .B(n16522), .X(n12643) );
  nand_x1_sg U13641 ( .A(n16735), .B(n16520), .X(n12644) );
  nand_x1_sg U13642 ( .A(n16735), .B(n16518), .X(n12645) );
  nand_x1_sg U13643 ( .A(n16735), .B(n16516), .X(n12646) );
  nand_x1_sg U13644 ( .A(n16735), .B(n16514), .X(n12647) );
  nand_x1_sg U13645 ( .A(n16734), .B(n16512), .X(n12648) );
  nand_x1_sg U13646 ( .A(n16735), .B(n16510), .X(n12649) );
  nand_x1_sg U13647 ( .A(n16735), .B(n16508), .X(n12650) );
  nand_x1_sg U13648 ( .A(n16735), .B(n16506), .X(n12651) );
  nand_x1_sg U13649 ( .A(n16735), .B(n16504), .X(n12652) );
  nand_x1_sg U13650 ( .A(n16735), .B(n16502), .X(n12653) );
  nand_x1_sg U13651 ( .A(n16735), .B(n16500), .X(n12654) );
  nand_x1_sg U13652 ( .A(n16735), .B(n16498), .X(n12655) );
  nand_x1_sg U13653 ( .A(n16735), .B(n16496), .X(n12656) );
  nand_x1_sg U13654 ( .A(n16735), .B(n16494), .X(n12657) );
  nand_x1_sg U13655 ( .A(n16735), .B(n16492), .X(n12658) );
  nand_x1_sg U13656 ( .A(n16735), .B(n16370), .X(n12659) );
  nand_x1_sg U13657 ( .A(n16735), .B(n16368), .X(n12660) );
  nand_x1_sg U13658 ( .A(n16735), .B(n16366), .X(n12661) );
  nand_x1_sg U13659 ( .A(n16735), .B(n16364), .X(n12662) );
  nand_x1_sg U13660 ( .A(n16735), .B(n16362), .X(n12663) );
  nand_x1_sg U13661 ( .A(n16735), .B(n16360), .X(n12664) );
  nand_x1_sg U13662 ( .A(n16735), .B(n16358), .X(n12665) );
  nand_x1_sg U13663 ( .A(n16735), .B(n16356), .X(n12666) );
  nand_x1_sg U13664 ( .A(n16735), .B(n16354), .X(n12667) );
  nand_x1_sg U13665 ( .A(n16734), .B(n16352), .X(n12668) );
  nand_x1_sg U13666 ( .A(n16735), .B(n16350), .X(n12669) );
  nand_x1_sg U13667 ( .A(n16735), .B(n16348), .X(n12670) );
  nand_x1_sg U13668 ( .A(n16735), .B(n16346), .X(n12671) );
  nand_x1_sg U13669 ( .A(n16735), .B(n16344), .X(n12672) );
  nand_x1_sg U13670 ( .A(n16735), .B(n16342), .X(n12673) );
  nand_x1_sg U13671 ( .A(n16735), .B(n16340), .X(n12674) );
  nand_x1_sg U13672 ( .A(n16735), .B(n16338), .X(n12675) );
  nand_x1_sg U13673 ( .A(n16735), .B(n16336), .X(n12676) );
  nand_x1_sg U13674 ( .A(n16735), .B(n16334), .X(n12677) );
  nand_x1_sg U13675 ( .A(n16735), .B(n16332), .X(n12678) );
  nand_x1_sg U13676 ( .A(n16735), .B(n16210), .X(n12679) );
  nand_x1_sg U13677 ( .A(n16735), .B(n16208), .X(n12680) );
  nand_x1_sg U13678 ( .A(n16735), .B(n16206), .X(n12681) );
  nand_x1_sg U13679 ( .A(n16735), .B(n16204), .X(n12682) );
  nand_x1_sg U13680 ( .A(n16735), .B(n16202), .X(n12683) );
  nand_x1_sg U13681 ( .A(n16735), .B(n16200), .X(n12684) );
  nand_x1_sg U13682 ( .A(n16735), .B(n16198), .X(n12685) );
  nand_x1_sg U13683 ( .A(n16735), .B(n16196), .X(n12686) );
  nand_x1_sg U13684 ( .A(n16735), .B(n16194), .X(n12687) );
  nand_x1_sg U13685 ( .A(n16735), .B(n16192), .X(n12688) );
  nand_x1_sg U13686 ( .A(n16735), .B(n16190), .X(n12689) );
  nand_x1_sg U13687 ( .A(n16735), .B(n16188), .X(n12690) );
  nand_x1_sg U13688 ( .A(n16735), .B(n16186), .X(n12691) );
  nand_x1_sg U13689 ( .A(n16735), .B(n16184), .X(n12692) );
  nand_x1_sg U13690 ( .A(n16735), .B(n16182), .X(n12693) );
  nand_x1_sg U13691 ( .A(n16735), .B(n16180), .X(n12694) );
  nand_x1_sg U13692 ( .A(n16735), .B(n16178), .X(n12695) );
  nand_x1_sg U13693 ( .A(n16735), .B(n16176), .X(n12696) );
  nand_x1_sg U13694 ( .A(n16735), .B(n16174), .X(n12697) );
  nand_x1_sg U13695 ( .A(n16735), .B(n16172), .X(n12698) );
  nand_x1_sg U13696 ( .A(n16735), .B(n16650), .X(n12699) );
  nand_x1_sg U13697 ( .A(n16735), .B(n16648), .X(n12700) );
  nand_x1_sg U13698 ( .A(n16735), .B(n16646), .X(n12701) );
  nand_x1_sg U13699 ( .A(n16735), .B(n16644), .X(n12702) );
  nand_x1_sg U13700 ( .A(n16735), .B(n16642), .X(n12703) );
  nand_x1_sg U13701 ( .A(n16735), .B(n16640), .X(n12704) );
  nand_x1_sg U13702 ( .A(n16735), .B(n16638), .X(n12705) );
  nand_x1_sg U13703 ( .A(n16735), .B(n16636), .X(n12706) );
  nand_x1_sg U13704 ( .A(n16735), .B(n16634), .X(n12707) );
  nand_x1_sg U13705 ( .A(n16735), .B(n16632), .X(n12708) );
  nand_x1_sg U13706 ( .A(n16735), .B(n16630), .X(n12709) );
  nand_x1_sg U13707 ( .A(n16735), .B(n16628), .X(n12710) );
  nand_x1_sg U13708 ( .A(n16735), .B(n16626), .X(n12711) );
  nand_x1_sg U13709 ( .A(n16735), .B(n16624), .X(n12712) );
  nand_x1_sg U13710 ( .A(n16735), .B(n16622), .X(n12713) );
  nand_x1_sg U13711 ( .A(n16735), .B(n16620), .X(n12714) );
  nand_x1_sg U13712 ( .A(n16735), .B(n16618), .X(n12715) );
  nand_x1_sg U13713 ( .A(n16735), .B(n16616), .X(n12716) );
  nand_x1_sg U13714 ( .A(n16735), .B(n16614), .X(n12717) );
  nand_x1_sg U13715 ( .A(n16735), .B(n16612), .X(n12718) );
  nand_x1_sg U13716 ( .A(n16735), .B(n16490), .X(n12719) );
  nand_x1_sg U13717 ( .A(n16735), .B(n16488), .X(n12720) );
  nand_x1_sg U13718 ( .A(n16734), .B(n16486), .X(n12721) );
  nand_x1_sg U13719 ( .A(n16735), .B(n16484), .X(n12722) );
  nand_x1_sg U13720 ( .A(n16735), .B(n16482), .X(n12723) );
  nand_x1_sg U13721 ( .A(n16735), .B(n16480), .X(n12724) );
  nand_x1_sg U13722 ( .A(n16735), .B(n16478), .X(n12725) );
  nand_x1_sg U13723 ( .A(n16735), .B(n16476), .X(n12726) );
  nand_x1_sg U13724 ( .A(n16735), .B(n16474), .X(n12727) );
  nand_x1_sg U13725 ( .A(n16735), .B(n16472), .X(n12728) );
  nand_x1_sg U13726 ( .A(n16735), .B(n16470), .X(n12729) );
  nand_x1_sg U13727 ( .A(n16735), .B(n16468), .X(n12730) );
  nand_x1_sg U13728 ( .A(n16735), .B(n16466), .X(n12731) );
  nand_x1_sg U13729 ( .A(n16735), .B(n16464), .X(n12732) );
  nand_x1_sg U13730 ( .A(n16735), .B(n16462), .X(n12733) );
  nand_x1_sg U13731 ( .A(n16735), .B(n16460), .X(n12734) );
  nand_x1_sg U13732 ( .A(n16735), .B(n16458), .X(n12735) );
  nand_x1_sg U13733 ( .A(n16735), .B(n16456), .X(n12736) );
  nand_x1_sg U13734 ( .A(n16735), .B(n16454), .X(n12737) );
  nand_x1_sg U13735 ( .A(n16735), .B(n16452), .X(n12738) );
  nand_x1_sg U13736 ( .A(n16735), .B(n16330), .X(n12739) );
  nand_x1_sg U13737 ( .A(n16735), .B(n16328), .X(n12740) );
  nand_x1_sg U13738 ( .A(n16734), .B(n16326), .X(n12741) );
  nand_x1_sg U13739 ( .A(n16735), .B(n16324), .X(n12742) );
  nand_x1_sg U13740 ( .A(n16735), .B(n16322), .X(n12743) );
  nand_x1_sg U13741 ( .A(n16735), .B(n16320), .X(n12744) );
  nand_x1_sg U13742 ( .A(n16735), .B(n16318), .X(n12745) );
  nand_x1_sg U13743 ( .A(n16735), .B(n16316), .X(n12746) );
  nand_x1_sg U13744 ( .A(n16735), .B(n16314), .X(n12747) );
  nand_x1_sg U13745 ( .A(n16735), .B(n16312), .X(n12748) );
  nand_x1_sg U13746 ( .A(n16735), .B(n16310), .X(n12749) );
  nand_x1_sg U13747 ( .A(n16735), .B(n16308), .X(n12750) );
  nand_x1_sg U13748 ( .A(n16735), .B(n16306), .X(n12751) );
  nand_x1_sg U13749 ( .A(n16735), .B(n16304), .X(n12752) );
  nand_x1_sg U13750 ( .A(n16735), .B(n16302), .X(n12753) );
  nand_x1_sg U13751 ( .A(n16735), .B(n16300), .X(n12754) );
  nand_x1_sg U13752 ( .A(n16735), .B(n16298), .X(n12755) );
  nand_x1_sg U13753 ( .A(n16735), .B(n16296), .X(n12756) );
  nand_x1_sg U13754 ( .A(n16735), .B(n16294), .X(n12757) );
  nand_x1_sg U13755 ( .A(n16735), .B(n16292), .X(n12758) );
  nand_x1_sg U13756 ( .A(n16735), .B(n16170), .X(n12759) );
  nand_x1_sg U13757 ( .A(n16735), .B(n16168), .X(n12760) );
  nand_x1_sg U13758 ( .A(n16735), .B(n16166), .X(n12761) );
  nand_x1_sg U13759 ( .A(n16735), .B(n16164), .X(n12762) );
  nand_x1_sg U13760 ( .A(n16735), .B(n16162), .X(n12763) );
  nand_x1_sg U13761 ( .A(n16735), .B(n16160), .X(n12764) );
  nand_x1_sg U13762 ( .A(n16735), .B(n16158), .X(n12765) );
  nand_x1_sg U13763 ( .A(n16735), .B(n16156), .X(n12766) );
  nand_x1_sg U13764 ( .A(n16735), .B(n16154), .X(n12767) );
  nand_x1_sg U13765 ( .A(n16735), .B(n16152), .X(n12768) );
  nand_x1_sg U13766 ( .A(n16735), .B(n16150), .X(n12769) );
  nand_x1_sg U13767 ( .A(n16735), .B(n16148), .X(n12770) );
  nand_x1_sg U13768 ( .A(n16735), .B(n16146), .X(n12771) );
  nand_x1_sg U13769 ( .A(n16735), .B(n16144), .X(n12772) );
  nand_x1_sg U13770 ( .A(n16735), .B(n16142), .X(n12773) );
  nand_x1_sg U13771 ( .A(n16735), .B(n16140), .X(n12774) );
  nand_x1_sg U13772 ( .A(n16735), .B(n16138), .X(n12775) );
  nand_x1_sg U13773 ( .A(n16735), .B(n16136), .X(n12776) );
  nand_x1_sg U13774 ( .A(n16735), .B(n16134), .X(n12777) );
  nand_x1_sg U13775 ( .A(n16735), .B(n16132), .X(n12778) );
  nand_x1_sg U13776 ( .A(n16735), .B(n16610), .X(n12779) );
  nand_x1_sg U13777 ( .A(n16735), .B(n16608), .X(n12780) );
  nand_x1_sg U13778 ( .A(n16735), .B(n16606), .X(n12781) );
  nand_x1_sg U13779 ( .A(n16735), .B(n16604), .X(n12782) );
  nand_x1_sg U13780 ( .A(n16735), .B(n16602), .X(n12783) );
  nand_x1_sg U13781 ( .A(n16735), .B(n16600), .X(n12784) );
  nand_x1_sg U13782 ( .A(n16735), .B(n16598), .X(n12785) );
  nand_x1_sg U13783 ( .A(n16735), .B(n16596), .X(n12786) );
  nand_x1_sg U13784 ( .A(n16735), .B(n16594), .X(n12787) );
  nand_x1_sg U13785 ( .A(n16735), .B(n16592), .X(n12788) );
  nand_x1_sg U13786 ( .A(n16735), .B(n16590), .X(n12789) );
  nand_x1_sg U13787 ( .A(n16735), .B(n16588), .X(n12790) );
  nand_x1_sg U13788 ( .A(n16735), .B(n16586), .X(n12791) );
  nand_x1_sg U13789 ( .A(n16735), .B(n16584), .X(n12792) );
  nand_x1_sg U13790 ( .A(n16735), .B(n16582), .X(n12793) );
  nand_x1_sg U13791 ( .A(n16735), .B(n16580), .X(n12794) );
  nand_x1_sg U13792 ( .A(n16735), .B(n16578), .X(n12795) );
  nand_x1_sg U13793 ( .A(n16735), .B(n16576), .X(n12796) );
  nand_x1_sg U13794 ( .A(n16735), .B(n16574), .X(n12797) );
  nand_x1_sg U13795 ( .A(n16735), .B(n16572), .X(n12798) );
  nand_x1_sg U13796 ( .A(n16735), .B(n16450), .X(n12799) );
  nand_x1_sg U13797 ( .A(n16735), .B(n16448), .X(n12800) );
  nand_x1_sg U13798 ( .A(n16735), .B(n16446), .X(n12801) );
  nand_x1_sg U13799 ( .A(n16735), .B(n16444), .X(n12802) );
  nand_x1_sg U13800 ( .A(n16735), .B(n16442), .X(n12803) );
  nand_x1_sg U13801 ( .A(n16735), .B(n16440), .X(n12804) );
  nand_x1_sg U13802 ( .A(n16735), .B(n16438), .X(n12805) );
  nand_x1_sg U13803 ( .A(n16735), .B(n16436), .X(n12806) );
  nand_x1_sg U13804 ( .A(n16735), .B(n16434), .X(n12807) );
  nand_x1_sg U13805 ( .A(n16735), .B(n16432), .X(n12808) );
  nand_x1_sg U13806 ( .A(n16735), .B(n16430), .X(n12809) );
  nand_x1_sg U13807 ( .A(n16735), .B(n16428), .X(n12810) );
  nand_x1_sg U13808 ( .A(n16735), .B(n16426), .X(n12811) );
  nand_x1_sg U13809 ( .A(n16735), .B(n16424), .X(n12812) );
  nand_x1_sg U13810 ( .A(n16735), .B(n16422), .X(n12813) );
  nand_x1_sg U13811 ( .A(n16735), .B(n16420), .X(n12814) );
  nand_x1_sg U13812 ( .A(n16735), .B(n16418), .X(n12815) );
  nand_x1_sg U13813 ( .A(n16735), .B(n16416), .X(n12816) );
  nand_x1_sg U13814 ( .A(n16735), .B(n16414), .X(n12817) );
  nand_x1_sg U13815 ( .A(n16735), .B(n16412), .X(n12818) );
  nand_x1_sg U13816 ( .A(n16735), .B(n16290), .X(n12819) );
  nand_x1_sg U13817 ( .A(n16735), .B(n16288), .X(n12820) );
  nand_x1_sg U13818 ( .A(n16735), .B(n16286), .X(n12821) );
  nand_x1_sg U13819 ( .A(n16735), .B(n16284), .X(n12822) );
  nand_x1_sg U13820 ( .A(n16735), .B(n16282), .X(n12823) );
  nand_x1_sg U13821 ( .A(n16735), .B(n16280), .X(n12824) );
  nand_x1_sg U13822 ( .A(n16735), .B(n16278), .X(n12825) );
  nand_x1_sg U13823 ( .A(n16735), .B(n16276), .X(n12826) );
  nand_x1_sg U13824 ( .A(n16735), .B(n16274), .X(n12827) );
  nand_x1_sg U13825 ( .A(n16735), .B(n16272), .X(n12828) );
  nand_x1_sg U13826 ( .A(n16735), .B(n16270), .X(n12829) );
  nand_x1_sg U13827 ( .A(n16735), .B(n16268), .X(n12830) );
  nand_x1_sg U13828 ( .A(n16735), .B(n16266), .X(n12831) );
  nand_x1_sg U13829 ( .A(n16735), .B(n16264), .X(n12832) );
  nand_x1_sg U13830 ( .A(n16735), .B(n16262), .X(n12833) );
  nand_x1_sg U13831 ( .A(n16735), .B(n16260), .X(n12834) );
  nand_x1_sg U13832 ( .A(n16735), .B(n16258), .X(n12835) );
  nand_x1_sg U13833 ( .A(n16735), .B(n16256), .X(n12836) );
  nand_x1_sg U13834 ( .A(n16735), .B(n16254), .X(n12837) );
  nand_x1_sg U13835 ( .A(n16735), .B(n16252), .X(n12838) );
  nand_x1_sg U13836 ( .A(n16735), .B(n16130), .X(n12839) );
  nand_x1_sg U13837 ( .A(n16735), .B(n16128), .X(n12840) );
  nand_x1_sg U13838 ( .A(n16735), .B(n16126), .X(n12841) );
  nand_x1_sg U13839 ( .A(n16735), .B(n16124), .X(n12842) );
  nand_x1_sg U13840 ( .A(n16735), .B(n16122), .X(n12843) );
  nand_x1_sg U13841 ( .A(n16735), .B(n16120), .X(n12844) );
  nand_x1_sg U13842 ( .A(n16735), .B(n16118), .X(n12845) );
  nand_x1_sg U13843 ( .A(n16735), .B(n16116), .X(n12846) );
  nand_x1_sg U13844 ( .A(n16735), .B(n16114), .X(n12847) );
  nand_x1_sg U13845 ( .A(n16735), .B(n16112), .X(n12848) );
  nand_x1_sg U13846 ( .A(n16735), .B(n16110), .X(n12849) );
  nand_x1_sg U13847 ( .A(n16735), .B(n16108), .X(n12850) );
  nand_x1_sg U13848 ( .A(n16735), .B(n16106), .X(n12851) );
  nand_x1_sg U13849 ( .A(n16735), .B(n16104), .X(n12852) );
  nand_x1_sg U13850 ( .A(n16735), .B(n16102), .X(n12853) );
  nand_x1_sg U13851 ( .A(n16735), .B(n16100), .X(n12854) );
  nand_x1_sg U13852 ( .A(n16735), .B(n16098), .X(n12855) );
  nand_x1_sg U13853 ( .A(n16735), .B(n16096), .X(n12856) );
  nand_x1_sg U13854 ( .A(n16735), .B(n16094), .X(n12857) );
  nand_x1_sg U13855 ( .A(n16735), .B(n16092), .X(n12858) );
  inv_x8_sg U13856 ( .A(n16734), .X(n16733) );
  inv_x8_sg U13857 ( .A(n14475), .X(n16734) );
  inv_x8_sg U13858 ( .A(n16733), .X(n16735) );
  inv_x8_sg U13859 ( .A(n16740), .X(n16736) );
  inv_x8_sg U13860 ( .A(n16740), .X(n16737) );
  inv_x8_sg U13861 ( .A(n16740), .X(n16738) );
  inv_x8_sg U13862 ( .A(n16740), .X(n16739) );
  inv_x8_sg U13863 ( .A(n16741), .X(n16740) );
  inv_x8_sg U13864 ( .A(n16742), .X(n16741) );
  inv_x8_sg U13865 ( .A(n16756), .X(n16745) );
  inv_x8_sg U13866 ( .A(n16756), .X(n16746) );
  inv_x8_sg U13867 ( .A(n16756), .X(n16747) );
  inv_x8_sg U13868 ( .A(n16756), .X(n16748) );
  inv_x8_sg U13869 ( .A(n16756), .X(n16749) );
  inv_x8_sg U13870 ( .A(n16756), .X(n16750) );
  inv_x8_sg U13871 ( .A(n16756), .X(n16751) );
  inv_x8_sg U13872 ( .A(n16756), .X(n16752) );
  inv_x8_sg U13873 ( .A(n16756), .X(n16753) );
  inv_x8_sg U13874 ( .A(n16756), .X(n16754) );
  inv_x8_sg U13875 ( .A(n16756), .X(n16755) );
  inv_x8_sg U13876 ( .A(n16757), .X(n16756) );
  inv_x8_sg U13877 ( .A(n16758), .X(n16757) );
  inv_x8_sg U13878 ( .A(n16773), .X(n16761) );
  inv_x8_sg U13879 ( .A(n16770), .X(n16762) );
  inv_x8_sg U13880 ( .A(n16770), .X(n16763) );
  inv_x8_sg U13881 ( .A(n16770), .X(n16764) );
  inv_x8_sg U13882 ( .A(n16770), .X(n16765) );
  inv_x8_sg U13883 ( .A(n16770), .X(n16766) );
  inv_x8_sg U13884 ( .A(n16770), .X(n16767) );
  inv_x8_sg U13885 ( .A(n16770), .X(n16768) );
  inv_x8_sg U13886 ( .A(n16770), .X(n16769) );
  inv_x8_sg U13887 ( .A(n16772), .X(n16770) );
  inv_x8_sg U13888 ( .A(n16773), .X(n16771) );
  inv_x8_sg U13889 ( .A(n16773), .X(n16772) );
  inv_x8_sg U13890 ( .A(n16774), .X(n16773) );
  inv_x8_sg U13891 ( .A(n16775), .X(n16774) );
  inv_x8_sg U13892 ( .A(n16787), .X(n16778) );
  inv_x8_sg U13893 ( .A(n16787), .X(n16779) );
  inv_x8_sg U13894 ( .A(n16792), .X(n16780) );
  inv_x8_sg U13895 ( .A(n16787), .X(n16781) );
  inv_x8_sg U13896 ( .A(n16787), .X(n16782) );
  inv_x8_sg U13897 ( .A(n16792), .X(n16783) );
  inv_x8_sg U13898 ( .A(n16792), .X(n16784) );
  inv_x8_sg U13899 ( .A(n16792), .X(n16785) );
  inv_x8_sg U13900 ( .A(n16792), .X(n16786) );
  inv_x8_sg U13901 ( .A(n16791), .X(n16787) );
  inv_x8_sg U13902 ( .A(n16792), .X(n16788) );
  inv_x8_sg U13903 ( .A(n16792), .X(n16789) );
  inv_x8_sg U13904 ( .A(n16792), .X(n16790) );
  inv_x8_sg U13905 ( .A(n16792), .X(n16791) );
  inv_x8_sg U13906 ( .A(n16793), .X(n16792) );
  inv_x8_sg U13907 ( .A(n16794), .X(n16793) );
endmodule

