
module sparsity ( clk, reset, i_0, i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, 
        i_10, i_11, i_12, i_13, i_14, i_15, w_0, w_1, w_2, w_3, w_4, w_5, w_6, 
        w_7, w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15, i_mask, w_mask, 
        input_ready, output_taken, oi_0, oi_1, oi_2, oi_3, oi_4, oi_5, oi_6, 
        oi_7, oi_8, oi_9, oi_10, oi_11, oi_12, oi_13, oi_14, oi_15, ow_0, ow_1, 
        ow_2, ow_3, ow_4, ow_5, ow_6, ow_7, ow_8, ow_9, ow_10, ow_11, ow_12, 
        ow_13, ow_14, ow_15, o_mask, state, input_taken );
  input [19:0] i_0;
  input [19:0] i_1;
  input [19:0] i_2;
  input [19:0] i_3;
  input [19:0] i_4;
  input [19:0] i_5;
  input [19:0] i_6;
  input [19:0] i_7;
  input [19:0] i_8;
  input [19:0] i_9;
  input [19:0] i_10;
  input [19:0] i_11;
  input [19:0] i_12;
  input [19:0] i_13;
  input [19:0] i_14;
  input [19:0] i_15;
  input [19:0] w_0;
  input [19:0] w_1;
  input [19:0] w_2;
  input [19:0] w_3;
  input [19:0] w_4;
  input [19:0] w_5;
  input [19:0] w_6;
  input [19:0] w_7;
  input [19:0] w_8;
  input [19:0] w_9;
  input [19:0] w_10;
  input [19:0] w_11;
  input [19:0] w_12;
  input [19:0] w_13;
  input [19:0] w_14;
  input [19:0] w_15;
  input [31:0] i_mask;
  input [31:0] w_mask;
  output [19:0] oi_0;
  output [19:0] oi_1;
  output [19:0] oi_2;
  output [19:0] oi_3;
  output [19:0] oi_4;
  output [19:0] oi_5;
  output [19:0] oi_6;
  output [19:0] oi_7;
  output [19:0] oi_8;
  output [19:0] oi_9;
  output [19:0] oi_10;
  output [19:0] oi_11;
  output [19:0] oi_12;
  output [19:0] oi_13;
  output [19:0] oi_14;
  output [19:0] oi_15;
  output [19:0] ow_0;
  output [19:0] ow_1;
  output [19:0] ow_2;
  output [19:0] ow_3;
  output [19:0] ow_4;
  output [19:0] ow_5;
  output [19:0] ow_6;
  output [19:0] ow_7;
  output [19:0] ow_8;
  output [19:0] ow_9;
  output [19:0] ow_10;
  output [19:0] ow_11;
  output [19:0] ow_12;
  output [19:0] ow_13;
  output [19:0] ow_14;
  output [19:0] ow_15;
  output [31:0] o_mask;
  output [1:0] state;
  input clk, reset, input_ready, output_taken;
  output input_taken;
  wire   mask_input_ready, mask_output_filter_input_taken, delayed_input_ready,
         filter_input_ready, filter_output_shifter_input_taken, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, \mask_0/n774 , \mask_0/n773 ,
         \mask_0/n772 , \mask_0/n771 , \mask_0/n770 , \mask_0/n769 ,
         \mask_0/n768 , \mask_0/n767 , \mask_0/n766 , \mask_0/n765 ,
         \mask_0/n764 , \mask_0/n763 , \mask_0/n762 , \mask_0/n761 ,
         \mask_0/n760 , \mask_0/n759 , \mask_0/n758 , \mask_0/n757 ,
         \mask_0/n756 , \mask_0/n755 , \mask_0/n754 , \mask_0/n753 ,
         \mask_0/n752 , \mask_0/n751 , \mask_0/n750 , \mask_0/n749 ,
         \mask_0/n748 , \mask_0/n747 , \mask_0/n746 , \mask_0/n745 ,
         \mask_0/n744 , \mask_0/n743 , \mask_0/n742 , \mask_0/n741 ,
         \mask_0/n740 , \mask_0/n739 , \mask_0/n738 , \mask_0/n737 ,
         \mask_0/n736 , \mask_0/n735 , \mask_0/n734 , \mask_0/n733 ,
         \mask_0/n732 , \mask_0/n731 , \mask_0/n730 , \mask_0/n729 ,
         \mask_0/n728 , \mask_0/n727 , \mask_0/n726 , \mask_0/n725 ,
         \mask_0/n724 , \mask_0/n723 , \mask_0/n722 , \mask_0/n721 ,
         \mask_0/n720 , \mask_0/n719 , \mask_0/n718 , \mask_0/n717 ,
         \mask_0/n716 , \mask_0/n715 , \mask_0/n714 , \mask_0/n713 ,
         \mask_0/n712 , \mask_0/n711 , \mask_0/n710 , \mask_0/n709 ,
         \mask_0/n708 , \mask_0/n707 , \mask_0/n706 , \mask_0/n705 ,
         \mask_0/n704 , \mask_0/n703 , \mask_0/n702 , \mask_0/n701 ,
         \mask_0/n700 , \mask_0/n699 , \mask_0/n698 , \mask_0/n697 ,
         \mask_0/n696 , \mask_0/n695 , \mask_0/n694 , \mask_0/n693 ,
         \mask_0/n692 , \mask_0/n691 , \mask_0/n690 , \mask_0/n689 ,
         \mask_0/n688 , \mask_0/n687 , \mask_0/n686 , \mask_0/n685 ,
         \mask_0/n684 , \mask_0/n683 , \mask_0/n682 , \mask_0/n681 ,
         \mask_0/n680 , \mask_0/n679 , \mask_0/n678 , \mask_0/n677 ,
         \mask_0/n676 , \mask_0/n675 , \mask_0/n674 , \mask_0/n673 ,
         \mask_0/n672 , \mask_0/n671 , \mask_0/n670 , \mask_0/n669 ,
         \mask_0/n668 , \mask_0/n667 , \mask_0/n666 , \mask_0/n665 ,
         \mask_0/n664 , \mask_0/n663 , \mask_0/n662 , \mask_0/n661 ,
         \mask_0/n660 , \mask_0/n659 , \mask_0/n658 , \mask_0/n657 ,
         \mask_0/n656 , \mask_0/n655 , \mask_0/n654 , \mask_0/n653 ,
         \mask_0/n652 , \mask_0/n651 , \mask_0/n650 , \mask_0/n649 ,
         \mask_0/n648 , \mask_0/n647 , \mask_0/n646 , \mask_0/n645 ,
         \mask_0/n644 , \mask_0/n643 , \mask_0/n642 , \mask_0/n641 ,
         \mask_0/n640 , \mask_0/n639 , \mask_0/n638 , \mask_0/n637 ,
         \mask_0/n636 , \mask_0/n635 , \mask_0/n634 , \mask_0/n633 ,
         \mask_0/n632 , \mask_0/n631 , \mask_0/n630 , \mask_0/n629 ,
         \mask_0/n628 , \mask_0/n627 , \mask_0/n626 , \mask_0/n625 ,
         \mask_0/n624 , \mask_0/n623 , \mask_0/n622 , \mask_0/n621 ,
         \mask_0/n620 , \mask_0/n619 , \mask_0/n618 , \mask_0/n617 ,
         \mask_0/n616 , \mask_0/n615 , \mask_0/n614 , \mask_0/n613 ,
         \mask_0/n612 , \mask_0/n611 , \mask_0/reg_ww_mask[0] ,
         \mask_0/reg_ww_mask[1] , \mask_0/reg_ww_mask[2] ,
         \mask_0/reg_ww_mask[3] , \mask_0/reg_ww_mask[4] ,
         \mask_0/reg_ww_mask[5] , \mask_0/reg_ww_mask[6] ,
         \mask_0/reg_ww_mask[7] , \mask_0/reg_ww_mask[8] ,
         \mask_0/reg_ww_mask[9] , \mask_0/reg_ww_mask[10] ,
         \mask_0/reg_ww_mask[11] , \mask_0/reg_ww_mask[12] ,
         \mask_0/reg_ww_mask[13] , \mask_0/reg_ww_mask[14] ,
         \mask_0/reg_ww_mask[15] , \mask_0/reg_ww_mask[16] ,
         \mask_0/reg_ww_mask[17] , \mask_0/reg_ww_mask[18] ,
         \mask_0/reg_ww_mask[19] , \mask_0/reg_ww_mask[20] ,
         \mask_0/reg_ww_mask[21] , \mask_0/reg_ww_mask[22] ,
         \mask_0/reg_ww_mask[23] , \mask_0/reg_ww_mask[24] ,
         \mask_0/reg_ww_mask[25] , \mask_0/reg_ww_mask[26] ,
         \mask_0/reg_ww_mask[27] , \mask_0/reg_ww_mask[28] ,
         \mask_0/reg_ww_mask[29] , \mask_0/reg_ww_mask[30] ,
         \mask_0/reg_ww_mask[31] , \mask_0/reg_ii_mask[0] ,
         \mask_0/reg_ii_mask[1] , \mask_0/reg_ii_mask[2] ,
         \mask_0/reg_ii_mask[3] , \mask_0/reg_ii_mask[4] ,
         \mask_0/reg_ii_mask[5] , \mask_0/reg_ii_mask[6] ,
         \mask_0/reg_ii_mask[7] , \mask_0/reg_ii_mask[8] ,
         \mask_0/reg_ii_mask[9] , \mask_0/reg_ii_mask[10] ,
         \mask_0/reg_ii_mask[11] , \mask_0/reg_ii_mask[12] ,
         \mask_0/reg_ii_mask[13] , \mask_0/reg_ii_mask[14] ,
         \mask_0/reg_ii_mask[15] , \mask_0/reg_ii_mask[16] ,
         \mask_0/reg_ii_mask[17] , \mask_0/reg_ii_mask[18] ,
         \mask_0/reg_ii_mask[19] , \mask_0/reg_ii_mask[20] ,
         \mask_0/reg_ii_mask[21] , \mask_0/reg_ii_mask[22] ,
         \mask_0/reg_ii_mask[23] , \mask_0/reg_ii_mask[24] ,
         \mask_0/reg_ii_mask[25] , \mask_0/reg_ii_mask[26] ,
         \mask_0/reg_ii_mask[27] , \mask_0/reg_ii_mask[28] ,
         \mask_0/reg_ii_mask[29] , \mask_0/reg_ii_mask[30] ,
         \mask_0/reg_ii_mask[31] , \mask_0/counter[0] , \mask_0/counter[1] ,
         \mask_0/reg_w_mask[0] , \mask_0/reg_w_mask[1] ,
         \mask_0/reg_w_mask[2] , \mask_0/reg_w_mask[3] ,
         \mask_0/reg_w_mask[4] , \mask_0/reg_w_mask[5] ,
         \mask_0/reg_w_mask[6] , \mask_0/reg_w_mask[7] ,
         \mask_0/reg_w_mask[8] , \mask_0/reg_w_mask[9] ,
         \mask_0/reg_w_mask[10] , \mask_0/reg_w_mask[11] ,
         \mask_0/reg_w_mask[12] , \mask_0/reg_w_mask[13] ,
         \mask_0/reg_w_mask[14] , \mask_0/reg_w_mask[15] ,
         \mask_0/reg_w_mask[16] , \mask_0/reg_w_mask[17] ,
         \mask_0/reg_w_mask[18] , \mask_0/reg_w_mask[19] ,
         \mask_0/reg_w_mask[20] , \mask_0/reg_w_mask[21] ,
         \mask_0/reg_w_mask[22] , \mask_0/reg_w_mask[23] ,
         \mask_0/reg_w_mask[24] , \mask_0/reg_w_mask[25] ,
         \mask_0/reg_w_mask[26] , \mask_0/reg_w_mask[27] ,
         \mask_0/reg_w_mask[28] , \mask_0/reg_w_mask[29] ,
         \mask_0/reg_w_mask[30] , \mask_0/reg_w_mask[31] ,
         \mask_0/reg_i_mask[0] , \mask_0/reg_i_mask[1] ,
         \mask_0/reg_i_mask[2] , \mask_0/reg_i_mask[3] ,
         \mask_0/reg_i_mask[4] , \mask_0/reg_i_mask[5] ,
         \mask_0/reg_i_mask[6] , \mask_0/reg_i_mask[7] ,
         \mask_0/reg_i_mask[8] , \mask_0/reg_i_mask[9] ,
         \mask_0/reg_i_mask[10] , \mask_0/reg_i_mask[11] ,
         \mask_0/reg_i_mask[12] , \mask_0/reg_i_mask[13] ,
         \mask_0/reg_i_mask[14] , \mask_0/reg_i_mask[15] ,
         \mask_0/reg_i_mask[16] , \mask_0/reg_i_mask[17] ,
         \mask_0/reg_i_mask[18] , \mask_0/reg_i_mask[19] ,
         \mask_0/reg_i_mask[20] , \mask_0/reg_i_mask[21] ,
         \mask_0/reg_i_mask[22] , \mask_0/reg_i_mask[23] ,
         \mask_0/reg_i_mask[24] , \mask_0/reg_i_mask[25] ,
         \mask_0/reg_i_mask[26] , \mask_0/reg_i_mask[27] ,
         \mask_0/reg_i_mask[28] , \mask_0/reg_i_mask[29] ,
         \mask_0/reg_i_mask[30] , \mask_0/reg_i_mask[31] , \mask_0/state[0] ,
         \mask_0/state[1] , \filter_0/n9635 , \filter_0/n9634 ,
         \filter_0/n9633 , \filter_0/n9632 , \filter_0/n9631 ,
         \filter_0/n9630 , \filter_0/n9629 , \filter_0/n9628 ,
         \filter_0/n9627 , \filter_0/n9626 , \filter_0/n9625 ,
         \filter_0/n9624 , \filter_0/n9623 , \filter_0/n9622 ,
         \filter_0/n9621 , \filter_0/n9620 , \filter_0/n9619 ,
         \filter_0/n9618 , \filter_0/n9617 , \filter_0/n9616 ,
         \filter_0/n9615 , \filter_0/n9614 , \filter_0/n9613 ,
         \filter_0/n9612 , \filter_0/n9611 , \filter_0/n9610 ,
         \filter_0/n9609 , \filter_0/n9608 , \filter_0/n9607 ,
         \filter_0/n9606 , \filter_0/n9605 , \filter_0/n9604 ,
         \filter_0/n9603 , \filter_0/n9602 , \filter_0/n9601 ,
         \filter_0/n9600 , \filter_0/n9599 , \filter_0/n9598 ,
         \filter_0/n9597 , \filter_0/n9596 , \filter_0/n9595 ,
         \filter_0/n9594 , \filter_0/n9593 , \filter_0/n9592 ,
         \filter_0/n9591 , \filter_0/n9590 , \filter_0/n9589 ,
         \filter_0/n9588 , \filter_0/n9587 , \filter_0/n9586 ,
         \filter_0/n9585 , \filter_0/n9584 , \filter_0/n9583 ,
         \filter_0/n9582 , \filter_0/n9581 , \filter_0/n9580 ,
         \filter_0/n9579 , \filter_0/n9578 , \filter_0/n9577 ,
         \filter_0/n9576 , \filter_0/n9575 , \filter_0/n9574 ,
         \filter_0/n9573 , \filter_0/n9572 , \filter_0/n9571 ,
         \filter_0/n9570 , \filter_0/n9569 , \filter_0/n9568 ,
         \filter_0/n9567 , \filter_0/n9566 , \filter_0/n9565 ,
         \filter_0/n9564 , \filter_0/n9563 , \filter_0/n9562 ,
         \filter_0/n9561 , \filter_0/n9560 , \filter_0/n9559 ,
         \filter_0/n9558 , \filter_0/n9557 , \filter_0/n9556 ,
         \filter_0/n9555 , \filter_0/n9554 , \filter_0/n9553 ,
         \filter_0/n9552 , \filter_0/n9551 , \filter_0/n9550 ,
         \filter_0/n9549 , \filter_0/n9548 , \filter_0/n9547 ,
         \filter_0/n9546 , \filter_0/n9545 , \filter_0/n9544 ,
         \filter_0/n9543 , \filter_0/n9542 , \filter_0/n9541 ,
         \filter_0/n9540 , \filter_0/n9539 , \filter_0/n9538 ,
         \filter_0/n9537 , \filter_0/n9536 , \filter_0/n9535 ,
         \filter_0/n9534 , \filter_0/n9533 , \filter_0/n9532 ,
         \filter_0/n9531 , \filter_0/n9530 , \filter_0/n9529 ,
         \filter_0/n9528 , \filter_0/n9527 , \filter_0/n9526 ,
         \filter_0/n9525 , \filter_0/n9524 , \filter_0/n9523 ,
         \filter_0/n9522 , \filter_0/n9521 , \filter_0/n9520 ,
         \filter_0/n9519 , \filter_0/n9518 , \filter_0/n9517 ,
         \filter_0/n9516 , \filter_0/n9515 , \filter_0/n9514 ,
         \filter_0/n9513 , \filter_0/n9512 , \filter_0/n9511 ,
         \filter_0/n9510 , \filter_0/n9509 , \filter_0/n9508 ,
         \filter_0/n9507 , \filter_0/n9506 , \filter_0/n9505 ,
         \filter_0/n9504 , \filter_0/n9503 , \filter_0/n9502 ,
         \filter_0/n9501 , \filter_0/n9500 , \filter_0/n9499 ,
         \filter_0/n9498 , \filter_0/n9497 , \filter_0/n9496 ,
         \filter_0/n9495 , \filter_0/n9494 , \filter_0/n9493 ,
         \filter_0/n9492 , \filter_0/n9491 , \filter_0/n9490 ,
         \filter_0/n9489 , \filter_0/n9488 , \filter_0/n9487 ,
         \filter_0/n9486 , \filter_0/n9485 , \filter_0/n9484 ,
         \filter_0/n9483 , \filter_0/n9482 , \filter_0/n9481 ,
         \filter_0/n9480 , \filter_0/n9479 , \filter_0/n9478 ,
         \filter_0/n9477 , \filter_0/n9476 , \filter_0/n9475 ,
         \filter_0/n9474 , \filter_0/n9473 , \filter_0/n9472 ,
         \filter_0/n9471 , \filter_0/n9470 , \filter_0/n9469 ,
         \filter_0/n9468 , \filter_0/n9467 , \filter_0/n9466 ,
         \filter_0/n9465 , \filter_0/n9464 , \filter_0/n9463 ,
         \filter_0/n9462 , \filter_0/n9461 , \filter_0/n9460 ,
         \filter_0/n9459 , \filter_0/n9458 , \filter_0/n9457 ,
         \filter_0/n9456 , \filter_0/n9455 , \filter_0/n9454 ,
         \filter_0/n9453 , \filter_0/n9452 , \filter_0/n9451 ,
         \filter_0/n9450 , \filter_0/n9449 , \filter_0/n9448 ,
         \filter_0/n9447 , \filter_0/n9446 , \filter_0/n9445 ,
         \filter_0/n9444 , \filter_0/n9443 , \filter_0/n9442 ,
         \filter_0/n9441 , \filter_0/n9440 , \filter_0/n9439 ,
         \filter_0/n9438 , \filter_0/n9437 , \filter_0/n9436 ,
         \filter_0/n9435 , \filter_0/n9434 , \filter_0/n9433 ,
         \filter_0/n9432 , \filter_0/n9431 , \filter_0/n9430 ,
         \filter_0/n9429 , \filter_0/n9428 , \filter_0/n9427 ,
         \filter_0/n9426 , \filter_0/n9425 , \filter_0/n9424 ,
         \filter_0/n9423 , \filter_0/n9422 , \filter_0/n9421 ,
         \filter_0/n9420 , \filter_0/n9419 , \filter_0/n9418 ,
         \filter_0/n9417 , \filter_0/n9416 , \filter_0/n9415 ,
         \filter_0/n9414 , \filter_0/n9413 , \filter_0/n9412 ,
         \filter_0/n9411 , \filter_0/n9410 , \filter_0/n9409 ,
         \filter_0/n9408 , \filter_0/n9407 , \filter_0/n9406 ,
         \filter_0/n9405 , \filter_0/n9404 , \filter_0/n9403 ,
         \filter_0/n9402 , \filter_0/n9401 , \filter_0/n9400 ,
         \filter_0/n9399 , \filter_0/n9398 , \filter_0/n9397 ,
         \filter_0/n9396 , \filter_0/n9395 , \filter_0/n9394 ,
         \filter_0/n9393 , \filter_0/n9392 , \filter_0/n9391 ,
         \filter_0/n9390 , \filter_0/n9389 , \filter_0/n9388 ,
         \filter_0/n9387 , \filter_0/n9386 , \filter_0/n9385 ,
         \filter_0/n9384 , \filter_0/n9383 , \filter_0/n9382 ,
         \filter_0/n9381 , \filter_0/n9380 , \filter_0/n9379 ,
         \filter_0/n9378 , \filter_0/n9377 , \filter_0/n9376 ,
         \filter_0/n9375 , \filter_0/n9374 , \filter_0/n9373 ,
         \filter_0/n9372 , \filter_0/n9371 , \filter_0/n9370 ,
         \filter_0/n9369 , \filter_0/n9368 , \filter_0/n9367 ,
         \filter_0/n9366 , \filter_0/n9365 , \filter_0/n9364 ,
         \filter_0/n9363 , \filter_0/n9362 , \filter_0/n9361 ,
         \filter_0/n9360 , \filter_0/n9359 , \filter_0/n9358 ,
         \filter_0/n9357 , \filter_0/n9356 , \filter_0/n9355 ,
         \filter_0/n9354 , \filter_0/n9353 , \filter_0/n9352 ,
         \filter_0/n9351 , \filter_0/n9350 , \filter_0/n9349 ,
         \filter_0/n9348 , \filter_0/n9347 , \filter_0/n9346 ,
         \filter_0/n9345 , \filter_0/n9344 , \filter_0/n9343 ,
         \filter_0/n9342 , \filter_0/n9341 , \filter_0/n9340 ,
         \filter_0/n9339 , \filter_0/n9338 , \filter_0/n9337 ,
         \filter_0/n9336 , \filter_0/n9335 , \filter_0/n9334 ,
         \filter_0/n9333 , \filter_0/n9332 , \filter_0/n9331 ,
         \filter_0/n9330 , \filter_0/n9329 , \filter_0/n9328 ,
         \filter_0/n9327 , \filter_0/n9326 , \filter_0/n9325 ,
         \filter_0/n9324 , \filter_0/n9323 , \filter_0/n9322 ,
         \filter_0/n9321 , \filter_0/n9320 , \filter_0/n9319 ,
         \filter_0/n9318 , \filter_0/n9317 , \filter_0/n9316 ,
         \filter_0/n9315 , \filter_0/n9314 , \filter_0/n9313 ,
         \filter_0/n9312 , \filter_0/n9311 , \filter_0/n9310 ,
         \filter_0/n9309 , \filter_0/n9308 , \filter_0/n9307 ,
         \filter_0/n9306 , \filter_0/n9305 , \filter_0/n9304 ,
         \filter_0/n9303 , \filter_0/n9302 , \filter_0/n9301 ,
         \filter_0/n9300 , \filter_0/n9299 , \filter_0/n9298 ,
         \filter_0/n9297 , \filter_0/n9296 , \filter_0/n9295 ,
         \filter_0/n9294 , \filter_0/n9293 , \filter_0/n9292 ,
         \filter_0/n9291 , \filter_0/n9290 , \filter_0/n9289 ,
         \filter_0/n9288 , \filter_0/n9287 , \filter_0/n9286 ,
         \filter_0/n9285 , \filter_0/n9284 , \filter_0/n9283 ,
         \filter_0/n9282 , \filter_0/n9281 , \filter_0/n9280 ,
         \filter_0/n9279 , \filter_0/n9278 , \filter_0/n9277 ,
         \filter_0/n9276 , \filter_0/n9275 , \filter_0/n9274 ,
         \filter_0/n9273 , \filter_0/n9272 , \filter_0/n9271 ,
         \filter_0/n9270 , \filter_0/n9269 , \filter_0/n9268 ,
         \filter_0/n9267 , \filter_0/n9266 , \filter_0/n9265 ,
         \filter_0/n9264 , \filter_0/n9263 , \filter_0/n9262 ,
         \filter_0/n9261 , \filter_0/n9260 , \filter_0/n9259 ,
         \filter_0/n9258 , \filter_0/n9257 , \filter_0/n9256 ,
         \filter_0/n9255 , \filter_0/n9254 , \filter_0/n9253 ,
         \filter_0/n9252 , \filter_0/n9251 , \filter_0/n9250 ,
         \filter_0/n9249 , \filter_0/n9248 , \filter_0/n9247 ,
         \filter_0/n9246 , \filter_0/n9245 , \filter_0/n9244 ,
         \filter_0/n9243 , \filter_0/n9242 , \filter_0/n9241 ,
         \filter_0/n9240 , \filter_0/n9239 , \filter_0/n9238 ,
         \filter_0/n9237 , \filter_0/n9236 , \filter_0/n9235 ,
         \filter_0/n9234 , \filter_0/n9233 , \filter_0/n9232 ,
         \filter_0/n9231 , \filter_0/n9230 , \filter_0/n9229 ,
         \filter_0/n9228 , \filter_0/n9227 , \filter_0/n9226 ,
         \filter_0/n9225 , \filter_0/n9224 , \filter_0/n9223 ,
         \filter_0/n9222 , \filter_0/n9221 , \filter_0/n9220 ,
         \filter_0/n9219 , \filter_0/n9218 , \filter_0/n9217 ,
         \filter_0/n9216 , \filter_0/n9215 , \filter_0/n9214 ,
         \filter_0/n9213 , \filter_0/n9212 , \filter_0/n9211 ,
         \filter_0/n9210 , \filter_0/n9209 , \filter_0/n9208 ,
         \filter_0/n9207 , \filter_0/n9206 , \filter_0/n9205 ,
         \filter_0/n9204 , \filter_0/n9203 , \filter_0/n9202 ,
         \filter_0/n9201 , \filter_0/n9200 , \filter_0/n9199 ,
         \filter_0/n9198 , \filter_0/n9197 , \filter_0/n9196 ,
         \filter_0/n9195 , \filter_0/n9194 , \filter_0/n9193 ,
         \filter_0/n9192 , \filter_0/n9191 , \filter_0/n9190 ,
         \filter_0/n9189 , \filter_0/n9188 , \filter_0/n9187 ,
         \filter_0/n9186 , \filter_0/n9185 , \filter_0/n9184 ,
         \filter_0/n9183 , \filter_0/n9182 , \filter_0/n9181 ,
         \filter_0/n9180 , \filter_0/n9179 , \filter_0/n9178 ,
         \filter_0/n9177 , \filter_0/n9176 , \filter_0/n9175 ,
         \filter_0/n9174 , \filter_0/n9173 , \filter_0/n9172 ,
         \filter_0/n9171 , \filter_0/n9170 , \filter_0/n9169 ,
         \filter_0/n9168 , \filter_0/n9167 , \filter_0/n9166 ,
         \filter_0/n9165 , \filter_0/n9164 , \filter_0/n9163 ,
         \filter_0/n9162 , \filter_0/n9161 , \filter_0/n9160 ,
         \filter_0/n9159 , \filter_0/n9158 , \filter_0/n9157 ,
         \filter_0/n9156 , \filter_0/n9155 , \filter_0/n9154 ,
         \filter_0/n9153 , \filter_0/n9152 , \filter_0/n9151 ,
         \filter_0/n9150 , \filter_0/n9149 , \filter_0/n9148 ,
         \filter_0/n9147 , \filter_0/n9146 , \filter_0/n9145 ,
         \filter_0/n9144 , \filter_0/n9143 , \filter_0/n9142 ,
         \filter_0/n9141 , \filter_0/n9140 , \filter_0/n9139 ,
         \filter_0/n9138 , \filter_0/n9137 , \filter_0/n9136 ,
         \filter_0/n9135 , \filter_0/n9134 , \filter_0/n9133 ,
         \filter_0/n9132 , \filter_0/n9131 , \filter_0/n9130 ,
         \filter_0/n9129 , \filter_0/n9128 , \filter_0/n9127 ,
         \filter_0/n9126 , \filter_0/n9125 , \filter_0/n9124 ,
         \filter_0/n9123 , \filter_0/n9122 , \filter_0/n9121 ,
         \filter_0/n9120 , \filter_0/n9119 , \filter_0/n9118 ,
         \filter_0/n9117 , \filter_0/n9116 , \filter_0/n9115 ,
         \filter_0/n9114 , \filter_0/n9113 , \filter_0/n9112 ,
         \filter_0/n9111 , \filter_0/n9110 , \filter_0/n9109 ,
         \filter_0/n9108 , \filter_0/n9107 , \filter_0/n9106 ,
         \filter_0/n9105 , \filter_0/n9104 , \filter_0/n9103 ,
         \filter_0/n9102 , \filter_0/n9101 , \filter_0/n9100 ,
         \filter_0/n9099 , \filter_0/n9098 , \filter_0/n9097 ,
         \filter_0/n9096 , \filter_0/n9095 , \filter_0/n9094 ,
         \filter_0/n9093 , \filter_0/n9092 , \filter_0/n9091 ,
         \filter_0/n9090 , \filter_0/n9089 , \filter_0/n9088 ,
         \filter_0/n9087 , \filter_0/n9086 , \filter_0/n9085 ,
         \filter_0/n9084 , \filter_0/n9083 , \filter_0/n9082 ,
         \filter_0/n9081 , \filter_0/n9080 , \filter_0/n9079 ,
         \filter_0/n9078 , \filter_0/n9077 , \filter_0/n9076 ,
         \filter_0/n9075 , \filter_0/n9074 , \filter_0/n9073 ,
         \filter_0/n9072 , \filter_0/n9071 , \filter_0/n9070 ,
         \filter_0/n9069 , \filter_0/n9068 , \filter_0/n9067 ,
         \filter_0/n9066 , \filter_0/n9065 , \filter_0/n9064 ,
         \filter_0/n9063 , \filter_0/n9062 , \filter_0/n9061 ,
         \filter_0/n9060 , \filter_0/n9059 , \filter_0/n9058 ,
         \filter_0/n9057 , \filter_0/n9056 , \filter_0/n9055 ,
         \filter_0/n9054 , \filter_0/n9053 , \filter_0/n9052 ,
         \filter_0/n9051 , \filter_0/n9050 , \filter_0/n9049 ,
         \filter_0/n9048 , \filter_0/n9047 , \filter_0/n9046 ,
         \filter_0/n9045 , \filter_0/n9044 , \filter_0/n9043 ,
         \filter_0/n9042 , \filter_0/n9041 , \filter_0/n9040 ,
         \filter_0/n9039 , \filter_0/n9038 , \filter_0/n9037 ,
         \filter_0/n9036 , \filter_0/n9035 , \filter_0/n9034 ,
         \filter_0/n9033 , \filter_0/n9032 , \filter_0/n9031 ,
         \filter_0/n9030 , \filter_0/n9029 , \filter_0/n9028 ,
         \filter_0/n9027 , \filter_0/n9026 , \filter_0/n9025 ,
         \filter_0/n9024 , \filter_0/n9023 , \filter_0/n9022 ,
         \filter_0/n9021 , \filter_0/n9020 , \filter_0/n9019 ,
         \filter_0/n9018 , \filter_0/n9017 , \filter_0/n9016 ,
         \filter_0/n9015 , \filter_0/n9014 , \filter_0/n9013 ,
         \filter_0/n9012 , \filter_0/n9011 , \filter_0/n9010 ,
         \filter_0/n9009 , \filter_0/n9008 , \filter_0/n9007 ,
         \filter_0/n9006 , \filter_0/n9005 , \filter_0/n9004 ,
         \filter_0/n9003 , \filter_0/n9002 , \filter_0/n9001 ,
         \filter_0/n9000 , \filter_0/n8999 , \filter_0/n8998 ,
         \filter_0/n8997 , \filter_0/n8996 , \filter_0/n8995 ,
         \filter_0/n8994 , \filter_0/n8993 , \filter_0/n8992 ,
         \filter_0/n8991 , \filter_0/n8990 , \filter_0/n8989 ,
         \filter_0/n8988 , \filter_0/n8987 , \filter_0/n8986 ,
         \filter_0/n8985 , \filter_0/n8984 , \filter_0/n8983 ,
         \filter_0/n8982 , \filter_0/n8981 , \filter_0/n8980 ,
         \filter_0/n8979 , \filter_0/n8978 , \filter_0/n8977 ,
         \filter_0/n8976 , \filter_0/n8975 , \filter_0/n8974 ,
         \filter_0/n8973 , \filter_0/n8972 , \filter_0/n8971 ,
         \filter_0/n8970 , \filter_0/n8969 , \filter_0/n8968 ,
         \filter_0/n8967 , \filter_0/n8966 , \filter_0/n8965 ,
         \filter_0/n8964 , \filter_0/n8963 , \filter_0/n8962 ,
         \filter_0/n8961 , \filter_0/n8960 , \filter_0/n8959 ,
         \filter_0/n8958 , \filter_0/n8957 , \filter_0/n8956 ,
         \filter_0/n8955 , \filter_0/n8954 , \filter_0/n8953 ,
         \filter_0/n8952 , \filter_0/n8951 , \filter_0/n8950 ,
         \filter_0/n8949 , \filter_0/n8948 , \filter_0/n8947 ,
         \filter_0/n8946 , \filter_0/n8945 , \filter_0/n8944 ,
         \filter_0/n8943 , \filter_0/n8942 , \filter_0/n8941 ,
         \filter_0/n8940 , \filter_0/n8939 , \filter_0/n8938 ,
         \filter_0/n8937 , \filter_0/n8936 , \filter_0/n8935 ,
         \filter_0/n8934 , \filter_0/n8933 , \filter_0/n8932 ,
         \filter_0/n8931 , \filter_0/n8930 , \filter_0/n8929 ,
         \filter_0/n8928 , \filter_0/n8927 , \filter_0/n8926 ,
         \filter_0/n8925 , \filter_0/n8924 , \filter_0/n8923 ,
         \filter_0/n8922 , \filter_0/n8921 , \filter_0/n8920 ,
         \filter_0/n8919 , \filter_0/n8918 , \filter_0/n8917 ,
         \filter_0/n8916 , \filter_0/n8915 , \filter_0/n8914 ,
         \filter_0/n8913 , \filter_0/n8912 , \filter_0/n8911 ,
         \filter_0/n8910 , \filter_0/n8909 , \filter_0/n8908 ,
         \filter_0/n8907 , \filter_0/n8906 , \filter_0/n8905 ,
         \filter_0/n8904 , \filter_0/n8903 , \filter_0/n8902 ,
         \filter_0/n8901 , \filter_0/n8900 , \filter_0/n8899 ,
         \filter_0/n8898 , \filter_0/n8897 , \filter_0/n8896 ,
         \filter_0/n8895 , \filter_0/n8894 , \filter_0/n8893 ,
         \filter_0/n8892 , \filter_0/n8891 , \filter_0/n8890 ,
         \filter_0/n8889 , \filter_0/n8888 , \filter_0/n8887 ,
         \filter_0/n8886 , \filter_0/n8885 , \filter_0/n8884 ,
         \filter_0/n8883 , \filter_0/n8882 , \filter_0/n8881 ,
         \filter_0/n8880 , \filter_0/n8879 , \filter_0/n8878 ,
         \filter_0/n8877 , \filter_0/n8876 , \filter_0/n8875 ,
         \filter_0/n8874 , \filter_0/n8873 , \filter_0/n8872 ,
         \filter_0/n8871 , \filter_0/n8870 , \filter_0/n8869 ,
         \filter_0/n8868 , \filter_0/n8867 , \filter_0/n8866 ,
         \filter_0/n8865 , \filter_0/n8864 , \filter_0/n8863 ,
         \filter_0/n8862 , \filter_0/n8861 , \filter_0/n8860 ,
         \filter_0/n8859 , \filter_0/n8858 , \filter_0/n8857 ,
         \filter_0/n8856 , \filter_0/n8855 , \filter_0/n8854 ,
         \filter_0/n8853 , \filter_0/n8852 , \filter_0/n8851 ,
         \filter_0/n8850 , \filter_0/n8849 , \filter_0/n8848 ,
         \filter_0/n8847 , \filter_0/n8846 , \filter_0/n8845 ,
         \filter_0/n8844 , \filter_0/n8843 , \filter_0/n8842 ,
         \filter_0/n8841 , \filter_0/n8840 , \filter_0/n8839 ,
         \filter_0/n8838 , \filter_0/n8837 , \filter_0/n8836 ,
         \filter_0/n8835 , \filter_0/n8834 , \filter_0/n8833 ,
         \filter_0/n8832 , \filter_0/n8831 , \filter_0/n8830 ,
         \filter_0/n8829 , \filter_0/n8828 , \filter_0/n8827 ,
         \filter_0/n8826 , \filter_0/n8825 , \filter_0/n8824 ,
         \filter_0/n8823 , \filter_0/n8822 , \filter_0/n8821 ,
         \filter_0/n8820 , \filter_0/n8819 , \filter_0/n8818 ,
         \filter_0/n8817 , \filter_0/n8816 , \filter_0/n8815 ,
         \filter_0/n8814 , \filter_0/n8813 , \filter_0/n8812 ,
         \filter_0/n8811 , \filter_0/n8810 , \filter_0/n8809 ,
         \filter_0/n8808 , \filter_0/n8807 , \filter_0/n8806 ,
         \filter_0/n8805 , \filter_0/n8804 , \filter_0/n8803 ,
         \filter_0/n8802 , \filter_0/n8801 , \filter_0/n8800 ,
         \filter_0/n8799 , \filter_0/n8798 , \filter_0/n8797 ,
         \filter_0/n8796 , \filter_0/n8795 , \filter_0/n8794 ,
         \filter_0/n8793 , \filter_0/n8792 , \filter_0/n8791 ,
         \filter_0/n8790 , \filter_0/n8789 , \filter_0/n8788 ,
         \filter_0/n8787 , \filter_0/n8786 , \filter_0/n8785 ,
         \filter_0/n8784 , \filter_0/n8783 , \filter_0/n8782 ,
         \filter_0/n8781 , \filter_0/n8780 , \filter_0/n8779 ,
         \filter_0/n8778 , \filter_0/n8777 , \filter_0/n8776 ,
         \filter_0/n8775 , \filter_0/n8774 , \filter_0/n8773 ,
         \filter_0/n8772 , \filter_0/n8771 , \filter_0/n8770 ,
         \filter_0/n8769 , \filter_0/n8768 , \filter_0/n8767 ,
         \filter_0/n8766 , \filter_0/n8765 , \filter_0/n8764 ,
         \filter_0/n8763 , \filter_0/n8762 , \filter_0/n8761 ,
         \filter_0/n8760 , \filter_0/n8759 , \filter_0/n8758 ,
         \filter_0/n8757 , \filter_0/n8756 , \filter_0/n8755 ,
         \filter_0/n8754 , \filter_0/n8753 , \filter_0/n8752 ,
         \filter_0/n8751 , \filter_0/n8750 , \filter_0/n8749 ,
         \filter_0/n8748 , \filter_0/n8747 , \filter_0/n8746 ,
         \filter_0/n8745 , \filter_0/n8744 , \filter_0/n8743 ,
         \filter_0/n8742 , \filter_0/n8741 , \filter_0/n8740 ,
         \filter_0/n8739 , \filter_0/n8738 , \filter_0/n8737 ,
         \filter_0/n8736 , \filter_0/n8735 , \filter_0/n8734 ,
         \filter_0/n8733 , \filter_0/n8732 , \filter_0/n8731 ,
         \filter_0/n8730 , \filter_0/n8729 , \filter_0/n8728 ,
         \filter_0/n8727 , \filter_0/n8726 , \filter_0/n8725 ,
         \filter_0/n8724 , \filter_0/n8723 , \filter_0/n8722 ,
         \filter_0/n8721 , \filter_0/n8720 , \filter_0/n8719 ,
         \filter_0/n8718 , \filter_0/n8717 , \filter_0/n8716 ,
         \filter_0/n8715 , \filter_0/n8714 , \filter_0/n8713 ,
         \filter_0/n8712 , \filter_0/n8711 , \filter_0/n8710 ,
         \filter_0/n8709 , \filter_0/n8708 , \filter_0/n8707 ,
         \filter_0/n8706 , \filter_0/n8705 , \filter_0/n8704 ,
         \filter_0/n8703 , \filter_0/n8702 , \filter_0/n8701 ,
         \filter_0/n8700 , \filter_0/n8699 , \filter_0/n8698 ,
         \filter_0/n8697 , \filter_0/n8696 , \filter_0/n8695 ,
         \filter_0/n8694 , \filter_0/n8693 , \filter_0/n8692 ,
         \filter_0/n8691 , \filter_0/n8690 , \filter_0/n8689 ,
         \filter_0/n8688 , \filter_0/n8687 , \filter_0/n8686 ,
         \filter_0/n8685 , \filter_0/n8684 , \filter_0/n8683 ,
         \filter_0/n8682 , \filter_0/n8681 , \filter_0/n8680 ,
         \filter_0/n8679 , \filter_0/n8678 , \filter_0/n8677 ,
         \filter_0/n8676 , \filter_0/n8675 , \filter_0/n8674 ,
         \filter_0/n8673 , \filter_0/n8672 , \filter_0/n8671 ,
         \filter_0/n8670 , \filter_0/n8669 , \filter_0/n8668 ,
         \filter_0/n8667 , \filter_0/n8666 , \filter_0/n8665 ,
         \filter_0/n8664 , \filter_0/n8663 , \filter_0/n8662 ,
         \filter_0/n8661 , \filter_0/n8660 , \filter_0/n8659 ,
         \filter_0/n8658 , \filter_0/n8657 , \filter_0/n8656 ,
         \filter_0/n8655 , \filter_0/n8654 , \filter_0/n8653 ,
         \filter_0/n8652 , \filter_0/n8651 , \filter_0/n8650 ,
         \filter_0/n8649 , \filter_0/n8648 , \filter_0/n8647 ,
         \filter_0/n8646 , \filter_0/n8645 , \filter_0/n8644 ,
         \filter_0/n8643 , \filter_0/n8642 , \filter_0/n8641 ,
         \filter_0/n8640 , \filter_0/n8639 , \filter_0/n8638 ,
         \filter_0/n8637 , \filter_0/n8636 , \filter_0/n8635 ,
         \filter_0/n8634 , \filter_0/n8633 , \filter_0/n8632 ,
         \filter_0/n8631 , \filter_0/n8630 , \filter_0/n8629 ,
         \filter_0/n8628 , \filter_0/n8627 , \filter_0/n8626 ,
         \filter_0/n8625 , \filter_0/n8624 , \filter_0/n8623 ,
         \filter_0/n8622 , \filter_0/n8621 , \filter_0/n8620 ,
         \filter_0/n8619 , \filter_0/n8618 , \filter_0/n8617 ,
         \filter_0/n8616 , \filter_0/n8615 , \filter_0/n8614 ,
         \filter_0/n8613 , \filter_0/n8612 , \filter_0/n8611 ,
         \filter_0/n8610 , \filter_0/n8609 , \filter_0/n8608 ,
         \filter_0/n8607 , \filter_0/n8606 , \filter_0/n8605 ,
         \filter_0/n8604 , \filter_0/n8603 , \filter_0/n8602 ,
         \filter_0/n8601 , \filter_0/n8600 , \filter_0/n8599 ,
         \filter_0/n8598 , \filter_0/n8597 , \filter_0/n8596 ,
         \filter_0/n8595 , \filter_0/n8594 , \filter_0/n8593 ,
         \filter_0/n8592 , \filter_0/n8591 , \filter_0/n8590 ,
         \filter_0/n8589 , \filter_0/n8588 , \filter_0/n8587 ,
         \filter_0/n8586 , \filter_0/n8585 , \filter_0/n8584 ,
         \filter_0/n8583 , \filter_0/n8582 , \filter_0/n8581 ,
         \filter_0/n8580 , \filter_0/n8579 , \filter_0/n8578 ,
         \filter_0/n8577 , \filter_0/n8576 , \filter_0/n8575 ,
         \filter_0/n8574 , \filter_0/n8573 , \filter_0/n8572 ,
         \filter_0/n8571 , \filter_0/n8570 , \filter_0/n8569 ,
         \filter_0/n8568 , \filter_0/n8567 , \filter_0/n8566 ,
         \filter_0/n8565 , \filter_0/n8564 , \filter_0/n8563 ,
         \filter_0/n8562 , \filter_0/n8561 , \filter_0/n8560 ,
         \filter_0/n8559 , \filter_0/n8558 , \filter_0/n8557 ,
         \filter_0/n8556 , \filter_0/n8555 , \filter_0/n8554 ,
         \filter_0/n8553 , \filter_0/n8552 , \filter_0/n8551 ,
         \filter_0/n8550 , \filter_0/n8549 , \filter_0/n8548 ,
         \filter_0/n8547 , \filter_0/n8546 , \filter_0/n8545 ,
         \filter_0/n8544 , \filter_0/n8543 , \filter_0/n8542 ,
         \filter_0/n8541 , \filter_0/n8540 , \filter_0/n8539 ,
         \filter_0/n8538 , \filter_0/n8537 , \filter_0/n8536 ,
         \filter_0/n8535 , \filter_0/n8534 , \filter_0/n8533 ,
         \filter_0/n8532 , \filter_0/n8531 , \filter_0/n8530 ,
         \filter_0/n8529 , \filter_0/n8528 , \filter_0/n8527 ,
         \filter_0/n8526 , \filter_0/n8525 , \filter_0/n8524 ,
         \filter_0/n8523 , \filter_0/n8522 , \filter_0/n8521 ,
         \filter_0/n8520 , \filter_0/n8519 , \filter_0/n8518 ,
         \filter_0/n8517 , \filter_0/n8516 , \filter_0/n8515 ,
         \filter_0/n8514 , \filter_0/n8513 , \filter_0/n8512 ,
         \filter_0/n8511 , \filter_0/n8510 , \filter_0/n8509 ,
         \filter_0/n8508 , \filter_0/n8507 , \filter_0/n8506 ,
         \filter_0/n8505 , \filter_0/n8504 , \filter_0/n8503 ,
         \filter_0/n8502 , \filter_0/n8501 , \filter_0/n8500 ,
         \filter_0/n8499 , \filter_0/n8498 , \filter_0/n8497 ,
         \filter_0/n8496 , \filter_0/n8495 , \filter_0/n8494 ,
         \filter_0/n8493 , \filter_0/n8492 , \filter_0/n8491 ,
         \filter_0/n8490 , \filter_0/n8489 , \filter_0/n8488 ,
         \filter_0/n8487 , \filter_0/n8486 , \filter_0/n8485 ,
         \filter_0/n8484 , \filter_0/n8483 , \filter_0/n8482 ,
         \filter_0/n8481 , \filter_0/n8480 , \filter_0/n8479 ,
         \filter_0/n8478 , \filter_0/n8477 , \filter_0/n8476 ,
         \filter_0/n8475 , \filter_0/n8474 , \filter_0/n8473 ,
         \filter_0/n8472 , \filter_0/n8471 , \filter_0/n8470 ,
         \filter_0/n8469 , \filter_0/n8468 , \filter_0/n8467 ,
         \filter_0/n8466 , \filter_0/n8465 , \filter_0/n8464 ,
         \filter_0/n8463 , \filter_0/n8462 , \filter_0/n8461 ,
         \filter_0/n8460 , \filter_0/n8459 , \filter_0/n8458 ,
         \filter_0/n8457 , \filter_0/n8456 , \filter_0/n8455 ,
         \filter_0/n8454 , \filter_0/n8453 , \filter_0/n8452 ,
         \filter_0/n8451 , \filter_0/n8450 , \filter_0/n8449 ,
         \filter_0/n8448 , \filter_0/n8447 , \filter_0/n8446 ,
         \filter_0/n8445 , \filter_0/n8444 , \filter_0/n8443 ,
         \filter_0/n8442 , \filter_0/n8441 , \filter_0/n8440 ,
         \filter_0/n8439 , \filter_0/n8438 , \filter_0/n8437 ,
         \filter_0/n8436 , \filter_0/n8435 , \filter_0/n8434 ,
         \filter_0/n8433 , \filter_0/n8432 , \filter_0/n8431 ,
         \filter_0/n8430 , \filter_0/n8429 , \filter_0/n8428 ,
         \filter_0/n8427 , \filter_0/n8426 , \filter_0/n8425 ,
         \filter_0/n8424 , \filter_0/n8423 , \filter_0/n8422 ,
         \filter_0/n8421 , \filter_0/n8420 , \filter_0/n8419 ,
         \filter_0/n8418 , \filter_0/n8417 , \filter_0/n8416 ,
         \filter_0/n8415 , \filter_0/n8414 , \filter_0/n8413 ,
         \filter_0/n8412 , \filter_0/n8411 , \filter_0/n8410 ,
         \filter_0/n8409 , \filter_0/n8408 , \filter_0/n8407 ,
         \filter_0/n8406 , \filter_0/n8405 , \filter_0/n8404 ,
         \filter_0/n8403 , \filter_0/n8402 , \filter_0/n8401 ,
         \filter_0/n8400 , \filter_0/n8399 , \filter_0/n8398 ,
         \filter_0/n8397 , \filter_0/n8396 , \filter_0/n8395 ,
         \filter_0/n8394 , \filter_0/n8393 , \filter_0/n8392 ,
         \filter_0/n8391 , \filter_0/n8390 , \filter_0/n8389 ,
         \filter_0/n8388 , \filter_0/n8387 , \filter_0/n8386 ,
         \filter_0/n8385 , \filter_0/n8384 , \filter_0/n8383 ,
         \filter_0/n8382 , \filter_0/n8381 , \filter_0/n8380 ,
         \filter_0/n8379 , \filter_0/n8378 , \filter_0/n8377 ,
         \filter_0/n8376 , \filter_0/n8375 , \filter_0/n8374 ,
         \filter_0/n8373 , \filter_0/n8372 , \filter_0/n8371 ,
         \filter_0/n8370 , \filter_0/n8369 , \filter_0/n8368 ,
         \filter_0/n8367 , \filter_0/n8366 , \filter_0/n8365 ,
         \filter_0/n8364 , \filter_0/n8363 , \filter_0/n8362 ,
         \filter_0/n8361 , \filter_0/n8360 , \filter_0/n8359 ,
         \filter_0/n8358 , \filter_0/n8357 , \filter_0/n8356 ,
         \filter_0/n8355 , \filter_0/n8354 , \filter_0/n8353 ,
         \filter_0/n8352 , \filter_0/n8351 , \filter_0/n8350 ,
         \filter_0/n8349 , \filter_0/n8348 , \filter_0/n8347 ,
         \filter_0/n8346 , \filter_0/n8345 , \filter_0/n8344 ,
         \filter_0/n8343 , \filter_0/n8342 , \filter_0/n8341 ,
         \filter_0/n8340 , \filter_0/n8339 , \filter_0/n8338 ,
         \filter_0/n8337 , \filter_0/n8336 , \filter_0/n8335 ,
         \filter_0/n8334 , \filter_0/n8333 , \filter_0/n8332 ,
         \filter_0/n8331 , \filter_0/n8330 , \filter_0/n8329 ,
         \filter_0/n8328 , \filter_0/n8327 , \filter_0/n8326 ,
         \filter_0/n8325 , \filter_0/n8324 , \filter_0/n8323 ,
         \filter_0/n8322 , \filter_0/n8321 , \filter_0/n8320 ,
         \filter_0/n8319 , \filter_0/n8318 , \filter_0/n8317 ,
         \filter_0/n8316 , \filter_0/n8315 , \filter_0/n8314 ,
         \filter_0/n8313 , \filter_0/n8312 , \filter_0/n8311 ,
         \filter_0/n8310 , \filter_0/n8309 , \filter_0/n8308 ,
         \filter_0/n8307 , \filter_0/n8306 , \filter_0/n8305 ,
         \filter_0/n8304 , \filter_0/n8303 , \filter_0/n8302 ,
         \filter_0/n8301 , \filter_0/n8300 , \filter_0/n8299 ,
         \filter_0/n8298 , \filter_0/n8297 , \filter_0/n8296 ,
         \filter_0/n8295 , \filter_0/n8294 , \filter_0/n8293 ,
         \filter_0/n8292 , \filter_0/n8291 , \filter_0/n8290 ,
         \filter_0/n8289 , \filter_0/n8288 , \filter_0/n8287 ,
         \filter_0/n8286 , \filter_0/n8285 , \filter_0/n8284 ,
         \filter_0/n8283 , \filter_0/n8282 , \filter_0/n8281 ,
         \filter_0/n8280 , \filter_0/n8279 , \filter_0/n8278 ,
         \filter_0/n8277 , \filter_0/n8276 , \filter_0/n8275 ,
         \filter_0/n8274 , \filter_0/n8273 , \filter_0/n8272 ,
         \filter_0/n8271 , \filter_0/n8270 , \filter_0/n8269 ,
         \filter_0/n8268 , \filter_0/n8267 , \filter_0/n8266 ,
         \filter_0/n8265 , \filter_0/n8264 , \filter_0/n8263 ,
         \filter_0/n8262 , \filter_0/n8261 , \filter_0/n8260 ,
         \filter_0/n8259 , \filter_0/n8258 , \filter_0/n8257 ,
         \filter_0/n8256 , \filter_0/n8255 , \filter_0/n8254 ,
         \filter_0/n8253 , \filter_0/n8252 , \filter_0/n8251 ,
         \filter_0/n8250 , \filter_0/n8249 , \filter_0/n8248 ,
         \filter_0/n8247 , \filter_0/n8246 , \filter_0/n8245 ,
         \filter_0/n8244 , \filter_0/n8243 , \filter_0/n8242 ,
         \filter_0/n8241 , \filter_0/n8240 , \filter_0/n8239 ,
         \filter_0/n8238 , \filter_0/n8237 , \filter_0/n8236 ,
         \filter_0/n8235 , \filter_0/n8234 , \filter_0/n8233 ,
         \filter_0/n8232 , \filter_0/n8231 , \filter_0/n8230 ,
         \filter_0/n8229 , \filter_0/n8228 , \filter_0/n8227 ,
         \filter_0/n8226 , \filter_0/n8225 , \filter_0/n8224 ,
         \filter_0/n8223 , \filter_0/n8222 , \filter_0/n8221 ,
         \filter_0/n8220 , \filter_0/n8219 , \filter_0/n8218 ,
         \filter_0/n8217 , \filter_0/n8216 , \filter_0/n8215 ,
         \filter_0/n8214 , \filter_0/n8213 , \filter_0/n8212 ,
         \filter_0/n8211 , \filter_0/n8210 , \filter_0/n8209 ,
         \filter_0/n8208 , \filter_0/n8207 , \filter_0/n8206 ,
         \filter_0/n8205 , \filter_0/n8204 , \filter_0/n8203 ,
         \filter_0/n8202 , \filter_0/n8201 , \filter_0/n8200 ,
         \filter_0/n8199 , \filter_0/n8198 , \filter_0/n8197 ,
         \filter_0/n8196 , \filter_0/n8195 , \filter_0/n8194 ,
         \filter_0/n8193 , \filter_0/n8192 , \filter_0/n8191 ,
         \filter_0/n8190 , \filter_0/n8189 , \filter_0/n8188 ,
         \filter_0/n8187 , \filter_0/n8186 , \filter_0/n8185 ,
         \filter_0/n8184 , \filter_0/n8183 , \filter_0/n8182 ,
         \filter_0/n8181 , \filter_0/n8180 , \filter_0/n8179 ,
         \filter_0/n8178 , \filter_0/n8177 , \filter_0/n8176 ,
         \filter_0/n8175 , \filter_0/n8174 , \filter_0/n8173 ,
         \filter_0/n8172 , \filter_0/n8171 , \filter_0/n8170 ,
         \filter_0/n8169 , \filter_0/n8168 , \filter_0/n8167 ,
         \filter_0/n8166 , \filter_0/n8165 , \filter_0/n8164 ,
         \filter_0/n8163 , \filter_0/n8162 , \filter_0/n8161 ,
         \filter_0/n8160 , \filter_0/n8159 , \filter_0/n8158 ,
         \filter_0/n8157 , \filter_0/n8156 , \filter_0/n8155 ,
         \filter_0/n8154 , \filter_0/n8153 , \filter_0/n8152 ,
         \filter_0/n8151 , \filter_0/n8150 , \filter_0/n8149 ,
         \filter_0/n8148 , \filter_0/n8147 , \filter_0/n8146 ,
         \filter_0/n8145 , \filter_0/n8144 , \filter_0/n8143 ,
         \filter_0/n8142 , \filter_0/n8141 , \filter_0/n8140 ,
         \filter_0/n8139 , \filter_0/n8138 , \filter_0/n8137 ,
         \filter_0/n8136 , \filter_0/n8135 , \filter_0/n8134 ,
         \filter_0/n8133 , \filter_0/n8132 , \filter_0/n8131 ,
         \filter_0/n8130 , \filter_0/n8129 , \filter_0/n8128 ,
         \filter_0/n8127 , \filter_0/n8126 , \filter_0/n8125 ,
         \filter_0/n8124 , \filter_0/n8123 , \filter_0/n8122 ,
         \filter_0/n8121 , \filter_0/n8120 , \filter_0/n8119 ,
         \filter_0/n8118 , \filter_0/n8117 , \filter_0/n8116 ,
         \filter_0/n8115 , \filter_0/n8114 , \filter_0/n8113 ,
         \filter_0/n8112 , \filter_0/n8111 , \filter_0/n8110 ,
         \filter_0/n8109 , \filter_0/n8108 , \filter_0/n8107 ,
         \filter_0/n8106 , \filter_0/n8105 , \filter_0/n8104 ,
         \filter_0/n8103 , \filter_0/n8102 , \filter_0/n8101 ,
         \filter_0/n8100 , \filter_0/n8099 , \filter_0/n8098 ,
         \filter_0/n8097 , \filter_0/n8096 , \filter_0/n8095 ,
         \filter_0/n8094 , \filter_0/n8093 , \filter_0/n8092 ,
         \filter_0/n8091 , \filter_0/n8090 , \filter_0/n8089 ,
         \filter_0/n8088 , \filter_0/n8087 , \filter_0/n8086 ,
         \filter_0/n8085 , \filter_0/n8084 , \filter_0/n8083 ,
         \filter_0/n8082 , \filter_0/n8081 , \filter_0/n8080 ,
         \filter_0/n8079 , \filter_0/n8078 , \filter_0/n8077 ,
         \filter_0/n8076 , \filter_0/n8075 , \filter_0/n8074 ,
         \filter_0/n8073 , \filter_0/n8072 , \filter_0/n8071 ,
         \filter_0/n8070 , \filter_0/n8069 , \filter_0/n8068 ,
         \filter_0/n8067 , \filter_0/n8066 , \filter_0/n8065 ,
         \filter_0/n8064 , \filter_0/n8063 , \filter_0/n8062 ,
         \filter_0/n8061 , \filter_0/n8060 , \filter_0/n8059 ,
         \filter_0/n8058 , \filter_0/n8057 , \filter_0/n8056 ,
         \filter_0/n8055 , \filter_0/n8054 , \filter_0/n8053 ,
         \filter_0/n8052 , \filter_0/n8051 , \filter_0/n8050 ,
         \filter_0/n8049 , \filter_0/n8048 , \filter_0/n8047 ,
         \filter_0/n8046 , \filter_0/n8045 , \filter_0/n8044 ,
         \filter_0/n8043 , \filter_0/n8042 , \filter_0/n8041 ,
         \filter_0/n8040 , \filter_0/n8039 , \filter_0/n8038 ,
         \filter_0/n8037 , \filter_0/n8036 , \filter_0/n8035 ,
         \filter_0/n8034 , \filter_0/n8033 , \filter_0/n8032 ,
         \filter_0/n8031 , \filter_0/n8030 , \filter_0/n8029 ,
         \filter_0/n8028 , \filter_0/n8027 , \filter_0/n8026 ,
         \filter_0/n8025 , \filter_0/n8024 , \filter_0/n8023 ,
         \filter_0/n8022 , \filter_0/n8021 , \filter_0/n8020 ,
         \filter_0/n8019 , \filter_0/n8018 , \filter_0/n8017 ,
         \filter_0/n8016 , \filter_0/n8015 , \filter_0/n8014 ,
         \filter_0/n8013 , \filter_0/n8012 , \filter_0/n8011 ,
         \filter_0/n8010 , \filter_0/n8009 , \filter_0/n8008 ,
         \filter_0/n8007 , \filter_0/n8006 , \filter_0/n8005 ,
         \filter_0/n8004 , \filter_0/n8003 , \filter_0/n8002 ,
         \filter_0/n8001 , \filter_0/n8000 , \filter_0/n7999 ,
         \filter_0/n7998 , \filter_0/n7997 , \filter_0/n7996 ,
         \filter_0/n7995 , \filter_0/n7994 , \filter_0/n7993 ,
         \filter_0/n7992 , \filter_0/n7991 , \filter_0/n7990 ,
         \filter_0/n7989 , \filter_0/n7988 , \filter_0/n7987 ,
         \filter_0/n7986 , \filter_0/n7985 , \filter_0/n7984 ,
         \filter_0/n7983 , \filter_0/n7982 , \filter_0/n7981 ,
         \filter_0/n7980 , \filter_0/n7979 , \filter_0/n7978 ,
         \filter_0/n7977 , \filter_0/n7976 , \filter_0/n7975 ,
         \filter_0/n7974 , \filter_0/n7973 , \filter_0/n7972 ,
         \filter_0/n7971 , \filter_0/n7970 , \filter_0/n7969 ,
         \filter_0/n7968 , \filter_0/n7967 , \filter_0/n7966 ,
         \filter_0/n7965 , \filter_0/n7964 , \filter_0/n7963 ,
         \filter_0/n7962 , \filter_0/n7961 , \filter_0/n7960 ,
         \filter_0/n7959 , \filter_0/n7958 , \filter_0/n7957 ,
         \filter_0/n7956 , \filter_0/n7955 , \filter_0/n7954 ,
         \filter_0/n7953 , \filter_0/n7952 , \filter_0/n7951 ,
         \filter_0/n7950 , \filter_0/n7949 , \filter_0/n7948 ,
         \filter_0/n7947 , \filter_0/n7946 , \filter_0/n7945 ,
         \filter_0/n7944 , \filter_0/n7943 , \filter_0/n7942 ,
         \filter_0/n7941 , \filter_0/n7940 , \filter_0/n7939 ,
         \filter_0/n7938 , \filter_0/n7937 , \filter_0/n7936 ,
         \filter_0/n7935 , \filter_0/n7934 , \filter_0/n7933 ,
         \filter_0/n7932 , \filter_0/n7931 , \filter_0/n7930 ,
         \filter_0/n7929 , \filter_0/n7928 , \filter_0/n7927 ,
         \filter_0/n7926 , \filter_0/n7925 , \filter_0/n7924 ,
         \filter_0/n7923 , \filter_0/n7922 , \filter_0/n7921 ,
         \filter_0/n7920 , \filter_0/n7919 , \filter_0/n7918 ,
         \filter_0/n7917 , \filter_0/n7916 , \filter_0/n7915 ,
         \filter_0/n7914 , \filter_0/n7913 , \filter_0/n7912 ,
         \filter_0/n7911 , \filter_0/n7910 , \filter_0/n7909 ,
         \filter_0/n7908 , \filter_0/n7907 , \filter_0/n7906 ,
         \filter_0/n7905 , \filter_0/n7904 , \filter_0/n7903 ,
         \filter_0/n7902 , \filter_0/n7901 , \filter_0/n7900 ,
         \filter_0/n7899 , \filter_0/n7898 , \filter_0/n7897 ,
         \filter_0/n7896 , \filter_0/n7895 , \filter_0/n7894 ,
         \filter_0/n7893 , \filter_0/n7892 , \filter_0/n7891 ,
         \filter_0/n7890 , \filter_0/n7889 , \filter_0/n7888 ,
         \filter_0/n7887 , \filter_0/n7886 , \filter_0/n7885 ,
         \filter_0/n7884 , \filter_0/n7883 , \filter_0/n7882 ,
         \filter_0/n7881 , \filter_0/n7880 , \filter_0/n7879 ,
         \filter_0/n7878 , \filter_0/n7877 , \filter_0/n7876 ,
         \filter_0/n7875 , \filter_0/n7874 , \filter_0/n7873 ,
         \filter_0/n7872 , \filter_0/n7871 , \filter_0/n7870 ,
         \filter_0/n7869 , \filter_0/n7868 , \filter_0/n7867 ,
         \filter_0/n7866 , \filter_0/n7865 , \filter_0/n7864 ,
         \filter_0/n7863 , \filter_0/n7862 , \filter_0/n7861 ,
         \filter_0/n7860 , \filter_0/n7859 , \filter_0/n7858 ,
         \filter_0/n7857 , \filter_0/n7856 , \filter_0/n7855 ,
         \filter_0/n7854 , \filter_0/n7853 , \filter_0/n7852 ,
         \filter_0/n7851 , \filter_0/n7850 , \filter_0/n7849 ,
         \filter_0/n7848 , \filter_0/n7847 , \filter_0/n7846 ,
         \filter_0/n7845 , \filter_0/n7844 , \filter_0/n7843 ,
         \filter_0/n7842 , \filter_0/n7841 , \filter_0/n7840 ,
         \filter_0/n7839 , \filter_0/n7838 , \filter_0/n7837 ,
         \filter_0/n7836 , \filter_0/n7835 , \filter_0/n7834 ,
         \filter_0/n7833 , \filter_0/n7832 , \filter_0/n7831 ,
         \filter_0/n7830 , \filter_0/n7829 , \filter_0/n7828 ,
         \filter_0/n7827 , \filter_0/n7826 , \filter_0/n7825 ,
         \filter_0/n7824 , \filter_0/n7823 , \filter_0/n7822 ,
         \filter_0/n7821 , \filter_0/n7820 , \filter_0/n7819 ,
         \filter_0/n7818 , \filter_0/n7817 , \filter_0/n7816 ,
         \filter_0/n7815 , \filter_0/n7814 , \filter_0/n7813 ,
         \filter_0/n7812 , \filter_0/n7811 , \filter_0/n7810 ,
         \filter_0/n7809 , \filter_0/n7808 , \filter_0/n7807 ,
         \filter_0/n7806 , \filter_0/n7805 , \filter_0/n7804 ,
         \filter_0/n7803 , \filter_0/n7802 , \filter_0/n7801 ,
         \filter_0/n7800 , \filter_0/n7799 , \filter_0/n7798 ,
         \filter_0/n7797 , \filter_0/n7796 , \filter_0/n7795 ,
         \filter_0/n7794 , \filter_0/n7793 , \filter_0/n7792 ,
         \filter_0/n7791 , \filter_0/n7790 , \filter_0/n7789 ,
         \filter_0/n7788 , \filter_0/n7787 , \filter_0/n7786 ,
         \filter_0/n7785 , \filter_0/n7784 , \filter_0/n7783 ,
         \filter_0/n7782 , \filter_0/n7781 , \filter_0/n7780 ,
         \filter_0/n7779 , \filter_0/n7778 , \filter_0/n7777 ,
         \filter_0/n7776 , \filter_0/n7775 , \filter_0/n7774 ,
         \filter_0/n7773 , \filter_0/n7772 , \filter_0/n7771 ,
         \filter_0/n7770 , \filter_0/n7769 , \filter_0/n7768 ,
         \filter_0/n7767 , \filter_0/n7766 , \filter_0/n7765 ,
         \filter_0/n7764 , \filter_0/n7763 , \filter_0/n7762 ,
         \filter_0/n7761 , \filter_0/n7760 , \filter_0/n7759 ,
         \filter_0/n7758 , \filter_0/n7757 , \filter_0/n7756 ,
         \filter_0/n7755 , \filter_0/n7754 , \filter_0/n7753 ,
         \filter_0/n7752 , \filter_0/n7751 , \filter_0/n7750 ,
         \filter_0/n7749 , \filter_0/n7748 , \filter_0/n7747 ,
         \filter_0/n7746 , \filter_0/n7745 , \filter_0/n7744 ,
         \filter_0/n7743 , \filter_0/n7742 , \filter_0/n7741 ,
         \filter_0/n7740 , \filter_0/n7739 , \filter_0/n7738 ,
         \filter_0/n7737 , \filter_0/n7736 , \filter_0/n7735 ,
         \filter_0/n7734 , \filter_0/n7733 , \filter_0/n7732 ,
         \filter_0/n7731 , \filter_0/n7730 , \filter_0/n7729 ,
         \filter_0/n7728 , \filter_0/n7727 , \filter_0/n7726 ,
         \filter_0/n7725 , \filter_0/n7724 , \filter_0/n7723 ,
         \filter_0/n7722 , \filter_0/n7721 , \filter_0/n7720 ,
         \filter_0/n7719 , \filter_0/n7718 , \filter_0/n7717 ,
         \filter_0/n7716 , \filter_0/n7715 , \filter_0/n7714 ,
         \filter_0/n7713 , \filter_0/n7712 , \filter_0/n7711 ,
         \filter_0/n7710 , \filter_0/n7709 , \filter_0/n7708 ,
         \filter_0/n7707 , \filter_0/n7706 , \filter_0/n7705 ,
         \filter_0/n7704 , \filter_0/n7703 , \filter_0/n7702 ,
         \filter_0/n7701 , \filter_0/n7700 , \filter_0/n7699 ,
         \filter_0/n7698 , \filter_0/n7697 , \filter_0/n7696 ,
         \filter_0/n7695 , \filter_0/n7694 , \filter_0/n7693 ,
         \filter_0/n7692 , \filter_0/n7691 , \filter_0/n7690 ,
         \filter_0/n7689 , \filter_0/n7688 , \filter_0/n7687 ,
         \filter_0/n7686 , \filter_0/n7685 , \filter_0/n7684 ,
         \filter_0/n7683 , \filter_0/n7682 , \filter_0/n7681 ,
         \filter_0/n7680 , \filter_0/n7679 , \filter_0/n7678 ,
         \filter_0/n7677 , \filter_0/n7676 , \filter_0/n7675 ,
         \filter_0/n7674 , \filter_0/n7673 , \filter_0/n7672 ,
         \filter_0/n7671 , \filter_0/n7670 , \filter_0/n7669 ,
         \filter_0/n7668 , \filter_0/n7667 , \filter_0/n7666 ,
         \filter_0/n7665 , \filter_0/n7664 , \filter_0/n7663 ,
         \filter_0/n7662 , \filter_0/n7661 , \filter_0/n7660 ,
         \filter_0/n7659 , \filter_0/n7658 , \filter_0/n7657 ,
         \filter_0/n7656 , \filter_0/n7655 , \filter_0/n7654 ,
         \filter_0/n7653 , \filter_0/n7652 , \filter_0/n7651 ,
         \filter_0/n7650 , \filter_0/n7649 , \filter_0/n7648 ,
         \filter_0/n7647 , \filter_0/n7646 , \filter_0/n7645 ,
         \filter_0/n7644 , \filter_0/n7643 , \filter_0/n7642 ,
         \filter_0/n7641 , \filter_0/n7640 , \filter_0/n7639 ,
         \filter_0/n7638 , \filter_0/n7637 , \filter_0/n7636 ,
         \filter_0/n7635 , \filter_0/n7634 , \filter_0/n7633 ,
         \filter_0/n7632 , \filter_0/n7631 , \filter_0/n7630 ,
         \filter_0/n7629 , \filter_0/n7628 , \filter_0/n7627 ,
         \filter_0/n7626 , \filter_0/n7625 , \filter_0/n7624 ,
         \filter_0/n7623 , \filter_0/n7622 , \filter_0/n7621 ,
         \filter_0/n7620 , \filter_0/n7619 , \filter_0/n7618 ,
         \filter_0/n7617 , \filter_0/n7616 , \filter_0/n7615 ,
         \filter_0/n7614 , \filter_0/n7613 , \filter_0/n7612 ,
         \filter_0/n7611 , \filter_0/n7610 , \filter_0/n7609 ,
         \filter_0/n7608 , \filter_0/n7607 , \filter_0/n7606 ,
         \filter_0/n7605 , \filter_0/n7604 , \filter_0/n7603 ,
         \filter_0/n7602 , \filter_0/n7601 , \filter_0/n7600 ,
         \filter_0/n7599 , \filter_0/n7598 , \filter_0/n7597 ,
         \filter_0/n7596 , \filter_0/n7595 , \filter_0/n7594 ,
         \filter_0/n7593 , \filter_0/n7592 , \filter_0/n7591 ,
         \filter_0/N1845 , \filter_0/w_pointer[0] , \filter_0/w_pointer[1] ,
         \filter_0/w_pointer[2] , \filter_0/w_pointer[3] ,
         \filter_0/i_pointer[0] , \filter_0/i_pointer[1] ,
         \filter_0/i_pointer[2] , \filter_0/i_pointer[3] ,
         \filter_0/reg_xor_w_mask[0] , \filter_0/reg_xor_w_mask[1] ,
         \filter_0/reg_xor_w_mask[2] , \filter_0/reg_xor_w_mask[3] ,
         \filter_0/reg_xor_w_mask[4] , \filter_0/reg_xor_w_mask[5] ,
         \filter_0/reg_xor_w_mask[6] , \filter_0/reg_xor_w_mask[7] ,
         \filter_0/reg_xor_w_mask[8] , \filter_0/reg_xor_w_mask[9] ,
         \filter_0/reg_xor_w_mask[10] , \filter_0/reg_xor_w_mask[11] ,
         \filter_0/reg_xor_w_mask[12] , \filter_0/reg_xor_w_mask[13] ,
         \filter_0/reg_xor_w_mask[14] , \filter_0/reg_xor_w_mask[15] ,
         \filter_0/reg_xor_w_mask[16] , \filter_0/reg_xor_w_mask[17] ,
         \filter_0/reg_xor_w_mask[18] , \filter_0/reg_xor_w_mask[19] ,
         \filter_0/reg_xor_w_mask[20] , \filter_0/reg_xor_w_mask[21] ,
         \filter_0/reg_xor_w_mask[22] , \filter_0/reg_xor_w_mask[23] ,
         \filter_0/reg_xor_w_mask[24] , \filter_0/reg_xor_w_mask[25] ,
         \filter_0/reg_xor_w_mask[26] , \filter_0/reg_xor_w_mask[27] ,
         \filter_0/reg_xor_w_mask[28] , \filter_0/reg_xor_w_mask[29] ,
         \filter_0/reg_xor_w_mask[30] , \filter_0/reg_xor_w_mask[31] ,
         \filter_0/reg_xor_i_mask[0] , \filter_0/reg_xor_i_mask[1] ,
         \filter_0/reg_xor_i_mask[2] , \filter_0/reg_xor_i_mask[3] ,
         \filter_0/reg_xor_i_mask[4] , \filter_0/reg_xor_i_mask[5] ,
         \filter_0/reg_xor_i_mask[6] , \filter_0/reg_xor_i_mask[7] ,
         \filter_0/reg_xor_i_mask[8] , \filter_0/reg_xor_i_mask[9] ,
         \filter_0/reg_xor_i_mask[10] , \filter_0/reg_xor_i_mask[11] ,
         \filter_0/reg_xor_i_mask[12] , \filter_0/reg_xor_i_mask[13] ,
         \filter_0/reg_xor_i_mask[14] , \filter_0/reg_xor_i_mask[15] ,
         \filter_0/reg_xor_i_mask[16] , \filter_0/reg_xor_i_mask[17] ,
         \filter_0/reg_xor_i_mask[18] , \filter_0/reg_xor_i_mask[19] ,
         \filter_0/reg_xor_i_mask[20] , \filter_0/reg_xor_i_mask[21] ,
         \filter_0/reg_xor_i_mask[22] , \filter_0/reg_xor_i_mask[23] ,
         \filter_0/reg_xor_i_mask[24] , \filter_0/reg_xor_i_mask[25] ,
         \filter_0/reg_xor_i_mask[26] , \filter_0/reg_xor_i_mask[27] ,
         \filter_0/reg_xor_i_mask[28] , \filter_0/reg_xor_i_mask[29] ,
         \filter_0/reg_xor_i_mask[30] , \filter_0/reg_xor_i_mask[31] ,
         \filter_0/reg_o_mask[0] , \filter_0/reg_o_mask[1] ,
         \filter_0/reg_o_mask[2] , \filter_0/reg_o_mask[3] ,
         \filter_0/reg_o_mask[4] , \filter_0/reg_o_mask[5] ,
         \filter_0/reg_o_mask[6] , \filter_0/reg_o_mask[7] ,
         \filter_0/reg_o_mask[8] , \filter_0/reg_o_mask[9] ,
         \filter_0/reg_o_mask[10] , \filter_0/reg_o_mask[11] ,
         \filter_0/reg_o_mask[12] , \filter_0/reg_o_mask[13] ,
         \filter_0/reg_o_mask[14] , \filter_0/reg_o_mask[15] ,
         \filter_0/reg_o_mask[16] , \filter_0/reg_o_mask[17] ,
         \filter_0/reg_o_mask[18] , \filter_0/reg_o_mask[19] ,
         \filter_0/reg_o_mask[20] , \filter_0/reg_o_mask[21] ,
         \filter_0/reg_o_mask[22] , \filter_0/reg_o_mask[23] ,
         \filter_0/reg_o_mask[24] , \filter_0/reg_o_mask[25] ,
         \filter_0/reg_o_mask[26] , \filter_0/reg_o_mask[27] ,
         \filter_0/reg_o_mask[28] , \filter_0/reg_o_mask[29] ,
         \filter_0/reg_o_mask[30] , \filter_0/reg_o_mask[31] ,
         \filter_0/reg_w_15[0] , \filter_0/reg_w_15[1] ,
         \filter_0/reg_w_15[2] , \filter_0/reg_w_15[3] ,
         \filter_0/reg_w_15[4] , \filter_0/reg_w_15[5] ,
         \filter_0/reg_w_15[6] , \filter_0/reg_w_15[7] ,
         \filter_0/reg_w_15[8] , \filter_0/reg_w_15[9] ,
         \filter_0/reg_w_15[10] , \filter_0/reg_w_15[11] ,
         \filter_0/reg_w_15[12] , \filter_0/reg_w_15[13] ,
         \filter_0/reg_w_15[14] , \filter_0/reg_w_15[15] ,
         \filter_0/reg_w_15[16] , \filter_0/reg_w_15[17] ,
         \filter_0/reg_w_15[18] , \filter_0/reg_w_15[19] ,
         \filter_0/reg_w_14[0] , \filter_0/reg_w_14[1] ,
         \filter_0/reg_w_14[2] , \filter_0/reg_w_14[3] ,
         \filter_0/reg_w_14[4] , \filter_0/reg_w_14[5] ,
         \filter_0/reg_w_14[6] , \filter_0/reg_w_14[7] ,
         \filter_0/reg_w_14[8] , \filter_0/reg_w_14[9] ,
         \filter_0/reg_w_14[10] , \filter_0/reg_w_14[11] ,
         \filter_0/reg_w_14[12] , \filter_0/reg_w_14[13] ,
         \filter_0/reg_w_14[14] , \filter_0/reg_w_14[15] ,
         \filter_0/reg_w_14[16] , \filter_0/reg_w_14[17] ,
         \filter_0/reg_w_14[18] , \filter_0/reg_w_14[19] ,
         \filter_0/reg_w_13[0] , \filter_0/reg_w_13[1] ,
         \filter_0/reg_w_13[2] , \filter_0/reg_w_13[3] ,
         \filter_0/reg_w_13[4] , \filter_0/reg_w_13[5] ,
         \filter_0/reg_w_13[6] , \filter_0/reg_w_13[7] ,
         \filter_0/reg_w_13[8] , \filter_0/reg_w_13[9] ,
         \filter_0/reg_w_13[10] , \filter_0/reg_w_13[11] ,
         \filter_0/reg_w_13[12] , \filter_0/reg_w_13[13] ,
         \filter_0/reg_w_13[14] , \filter_0/reg_w_13[15] ,
         \filter_0/reg_w_13[16] , \filter_0/reg_w_13[17] ,
         \filter_0/reg_w_13[18] , \filter_0/reg_w_13[19] ,
         \filter_0/reg_w_12[0] , \filter_0/reg_w_12[1] ,
         \filter_0/reg_w_12[2] , \filter_0/reg_w_12[3] ,
         \filter_0/reg_w_12[4] , \filter_0/reg_w_12[5] ,
         \filter_0/reg_w_12[6] , \filter_0/reg_w_12[7] ,
         \filter_0/reg_w_12[8] , \filter_0/reg_w_12[9] ,
         \filter_0/reg_w_12[10] , \filter_0/reg_w_12[11] ,
         \filter_0/reg_w_12[12] , \filter_0/reg_w_12[13] ,
         \filter_0/reg_w_12[14] , \filter_0/reg_w_12[15] ,
         \filter_0/reg_w_12[16] , \filter_0/reg_w_12[17] ,
         \filter_0/reg_w_12[18] , \filter_0/reg_w_12[19] ,
         \filter_0/reg_w_11[0] , \filter_0/reg_w_11[1] ,
         \filter_0/reg_w_11[2] , \filter_0/reg_w_11[3] ,
         \filter_0/reg_w_11[4] , \filter_0/reg_w_11[5] ,
         \filter_0/reg_w_11[6] , \filter_0/reg_w_11[7] ,
         \filter_0/reg_w_11[8] , \filter_0/reg_w_11[9] ,
         \filter_0/reg_w_11[10] , \filter_0/reg_w_11[11] ,
         \filter_0/reg_w_11[12] , \filter_0/reg_w_11[13] ,
         \filter_0/reg_w_11[14] , \filter_0/reg_w_11[15] ,
         \filter_0/reg_w_11[16] , \filter_0/reg_w_11[17] ,
         \filter_0/reg_w_11[18] , \filter_0/reg_w_11[19] ,
         \filter_0/reg_w_10[0] , \filter_0/reg_w_10[1] ,
         \filter_0/reg_w_10[2] , \filter_0/reg_w_10[3] ,
         \filter_0/reg_w_10[4] , \filter_0/reg_w_10[5] ,
         \filter_0/reg_w_10[6] , \filter_0/reg_w_10[7] ,
         \filter_0/reg_w_10[8] , \filter_0/reg_w_10[9] ,
         \filter_0/reg_w_10[10] , \filter_0/reg_w_10[11] ,
         \filter_0/reg_w_10[12] , \filter_0/reg_w_10[13] ,
         \filter_0/reg_w_10[14] , \filter_0/reg_w_10[15] ,
         \filter_0/reg_w_10[16] , \filter_0/reg_w_10[17] ,
         \filter_0/reg_w_10[18] , \filter_0/reg_w_10[19] ,
         \filter_0/reg_w_9[0] , \filter_0/reg_w_9[1] , \filter_0/reg_w_9[2] ,
         \filter_0/reg_w_9[3] , \filter_0/reg_w_9[4] , \filter_0/reg_w_9[5] ,
         \filter_0/reg_w_9[6] , \filter_0/reg_w_9[7] , \filter_0/reg_w_9[8] ,
         \filter_0/reg_w_9[9] , \filter_0/reg_w_9[10] , \filter_0/reg_w_9[11] ,
         \filter_0/reg_w_9[12] , \filter_0/reg_w_9[13] ,
         \filter_0/reg_w_9[14] , \filter_0/reg_w_9[15] ,
         \filter_0/reg_w_9[16] , \filter_0/reg_w_9[17] ,
         \filter_0/reg_w_9[18] , \filter_0/reg_w_9[19] , \filter_0/reg_w_8[0] ,
         \filter_0/reg_w_8[1] , \filter_0/reg_w_8[2] , \filter_0/reg_w_8[3] ,
         \filter_0/reg_w_8[4] , \filter_0/reg_w_8[5] , \filter_0/reg_w_8[6] ,
         \filter_0/reg_w_8[7] , \filter_0/reg_w_8[8] , \filter_0/reg_w_8[9] ,
         \filter_0/reg_w_8[10] , \filter_0/reg_w_8[11] ,
         \filter_0/reg_w_8[12] , \filter_0/reg_w_8[13] ,
         \filter_0/reg_w_8[14] , \filter_0/reg_w_8[15] ,
         \filter_0/reg_w_8[16] , \filter_0/reg_w_8[17] ,
         \filter_0/reg_w_8[18] , \filter_0/reg_w_8[19] , \filter_0/reg_w_7[0] ,
         \filter_0/reg_w_7[1] , \filter_0/reg_w_7[2] , \filter_0/reg_w_7[3] ,
         \filter_0/reg_w_7[4] , \filter_0/reg_w_7[5] , \filter_0/reg_w_7[6] ,
         \filter_0/reg_w_7[7] , \filter_0/reg_w_7[8] , \filter_0/reg_w_7[9] ,
         \filter_0/reg_w_7[10] , \filter_0/reg_w_7[11] ,
         \filter_0/reg_w_7[12] , \filter_0/reg_w_7[13] ,
         \filter_0/reg_w_7[14] , \filter_0/reg_w_7[15] ,
         \filter_0/reg_w_7[16] , \filter_0/reg_w_7[17] ,
         \filter_0/reg_w_7[18] , \filter_0/reg_w_7[19] , \filter_0/reg_w_6[0] ,
         \filter_0/reg_w_6[1] , \filter_0/reg_w_6[2] , \filter_0/reg_w_6[3] ,
         \filter_0/reg_w_6[4] , \filter_0/reg_w_6[5] , \filter_0/reg_w_6[6] ,
         \filter_0/reg_w_6[7] , \filter_0/reg_w_6[8] , \filter_0/reg_w_6[9] ,
         \filter_0/reg_w_6[10] , \filter_0/reg_w_6[11] ,
         \filter_0/reg_w_6[12] , \filter_0/reg_w_6[13] ,
         \filter_0/reg_w_6[14] , \filter_0/reg_w_6[15] ,
         \filter_0/reg_w_6[16] , \filter_0/reg_w_6[17] ,
         \filter_0/reg_w_6[18] , \filter_0/reg_w_6[19] , \filter_0/reg_w_5[0] ,
         \filter_0/reg_w_5[1] , \filter_0/reg_w_5[2] , \filter_0/reg_w_5[3] ,
         \filter_0/reg_w_5[4] , \filter_0/reg_w_5[5] , \filter_0/reg_w_5[6] ,
         \filter_0/reg_w_5[7] , \filter_0/reg_w_5[8] , \filter_0/reg_w_5[9] ,
         \filter_0/reg_w_5[10] , \filter_0/reg_w_5[11] ,
         \filter_0/reg_w_5[12] , \filter_0/reg_w_5[13] ,
         \filter_0/reg_w_5[14] , \filter_0/reg_w_5[15] ,
         \filter_0/reg_w_5[16] , \filter_0/reg_w_5[17] ,
         \filter_0/reg_w_5[18] , \filter_0/reg_w_5[19] , \filter_0/reg_w_4[0] ,
         \filter_0/reg_w_4[1] , \filter_0/reg_w_4[2] , \filter_0/reg_w_4[3] ,
         \filter_0/reg_w_4[4] , \filter_0/reg_w_4[5] , \filter_0/reg_w_4[6] ,
         \filter_0/reg_w_4[7] , \filter_0/reg_w_4[8] , \filter_0/reg_w_4[9] ,
         \filter_0/reg_w_4[10] , \filter_0/reg_w_4[11] ,
         \filter_0/reg_w_4[12] , \filter_0/reg_w_4[13] ,
         \filter_0/reg_w_4[14] , \filter_0/reg_w_4[15] ,
         \filter_0/reg_w_4[16] , \filter_0/reg_w_4[17] ,
         \filter_0/reg_w_4[18] , \filter_0/reg_w_4[19] , \filter_0/reg_w_3[0] ,
         \filter_0/reg_w_3[1] , \filter_0/reg_w_3[2] , \filter_0/reg_w_3[3] ,
         \filter_0/reg_w_3[4] , \filter_0/reg_w_3[5] , \filter_0/reg_w_3[6] ,
         \filter_0/reg_w_3[7] , \filter_0/reg_w_3[8] , \filter_0/reg_w_3[9] ,
         \filter_0/reg_w_3[10] , \filter_0/reg_w_3[11] ,
         \filter_0/reg_w_3[12] , \filter_0/reg_w_3[13] ,
         \filter_0/reg_w_3[14] , \filter_0/reg_w_3[15] ,
         \filter_0/reg_w_3[16] , \filter_0/reg_w_3[17] ,
         \filter_0/reg_w_3[18] , \filter_0/reg_w_3[19] , \filter_0/reg_w_2[0] ,
         \filter_0/reg_w_2[1] , \filter_0/reg_w_2[2] , \filter_0/reg_w_2[3] ,
         \filter_0/reg_w_2[4] , \filter_0/reg_w_2[5] , \filter_0/reg_w_2[6] ,
         \filter_0/reg_w_2[7] , \filter_0/reg_w_2[8] , \filter_0/reg_w_2[9] ,
         \filter_0/reg_w_2[10] , \filter_0/reg_w_2[11] ,
         \filter_0/reg_w_2[12] , \filter_0/reg_w_2[13] ,
         \filter_0/reg_w_2[14] , \filter_0/reg_w_2[15] ,
         \filter_0/reg_w_2[16] , \filter_0/reg_w_2[17] ,
         \filter_0/reg_w_2[18] , \filter_0/reg_w_2[19] , \filter_0/reg_w_1[0] ,
         \filter_0/reg_w_1[1] , \filter_0/reg_w_1[2] , \filter_0/reg_w_1[3] ,
         \filter_0/reg_w_1[4] , \filter_0/reg_w_1[5] , \filter_0/reg_w_1[6] ,
         \filter_0/reg_w_1[7] , \filter_0/reg_w_1[8] , \filter_0/reg_w_1[9] ,
         \filter_0/reg_w_1[10] , \filter_0/reg_w_1[11] ,
         \filter_0/reg_w_1[12] , \filter_0/reg_w_1[13] ,
         \filter_0/reg_w_1[14] , \filter_0/reg_w_1[15] ,
         \filter_0/reg_w_1[16] , \filter_0/reg_w_1[17] ,
         \filter_0/reg_w_1[18] , \filter_0/reg_w_1[19] , \filter_0/reg_w_0[0] ,
         \filter_0/reg_w_0[1] , \filter_0/reg_w_0[2] , \filter_0/reg_w_0[3] ,
         \filter_0/reg_w_0[4] , \filter_0/reg_w_0[5] , \filter_0/reg_w_0[6] ,
         \filter_0/reg_w_0[7] , \filter_0/reg_w_0[8] , \filter_0/reg_w_0[9] ,
         \filter_0/reg_w_0[10] , \filter_0/reg_w_0[11] ,
         \filter_0/reg_w_0[12] , \filter_0/reg_w_0[13] ,
         \filter_0/reg_w_0[14] , \filter_0/reg_w_0[15] ,
         \filter_0/reg_w_0[16] , \filter_0/reg_w_0[17] ,
         \filter_0/reg_w_0[18] , \filter_0/reg_w_0[19] ,
         \filter_0/reg_i_15[0] , \filter_0/reg_i_15[1] ,
         \filter_0/reg_i_15[2] , \filter_0/reg_i_15[3] ,
         \filter_0/reg_i_15[4] , \filter_0/reg_i_15[5] ,
         \filter_0/reg_i_15[6] , \filter_0/reg_i_15[7] ,
         \filter_0/reg_i_15[8] , \filter_0/reg_i_15[9] ,
         \filter_0/reg_i_15[10] , \filter_0/reg_i_15[11] ,
         \filter_0/reg_i_15[12] , \filter_0/reg_i_15[13] ,
         \filter_0/reg_i_15[14] , \filter_0/reg_i_15[15] ,
         \filter_0/reg_i_15[16] , \filter_0/reg_i_15[17] ,
         \filter_0/reg_i_15[18] , \filter_0/reg_i_15[19] ,
         \filter_0/reg_i_14[0] , \filter_0/reg_i_14[1] ,
         \filter_0/reg_i_14[2] , \filter_0/reg_i_14[3] ,
         \filter_0/reg_i_14[4] , \filter_0/reg_i_14[5] ,
         \filter_0/reg_i_14[6] , \filter_0/reg_i_14[7] ,
         \filter_0/reg_i_14[8] , \filter_0/reg_i_14[9] ,
         \filter_0/reg_i_14[10] , \filter_0/reg_i_14[11] ,
         \filter_0/reg_i_14[12] , \filter_0/reg_i_14[13] ,
         \filter_0/reg_i_14[14] , \filter_0/reg_i_14[15] ,
         \filter_0/reg_i_14[16] , \filter_0/reg_i_14[17] ,
         \filter_0/reg_i_14[18] , \filter_0/reg_i_14[19] ,
         \filter_0/reg_i_13[0] , \filter_0/reg_i_13[1] ,
         \filter_0/reg_i_13[2] , \filter_0/reg_i_13[3] ,
         \filter_0/reg_i_13[4] , \filter_0/reg_i_13[5] ,
         \filter_0/reg_i_13[6] , \filter_0/reg_i_13[7] ,
         \filter_0/reg_i_13[8] , \filter_0/reg_i_13[9] ,
         \filter_0/reg_i_13[10] , \filter_0/reg_i_13[11] ,
         \filter_0/reg_i_13[12] , \filter_0/reg_i_13[13] ,
         \filter_0/reg_i_13[14] , \filter_0/reg_i_13[15] ,
         \filter_0/reg_i_13[16] , \filter_0/reg_i_13[17] ,
         \filter_0/reg_i_13[18] , \filter_0/reg_i_13[19] ,
         \filter_0/reg_i_12[0] , \filter_0/reg_i_12[1] ,
         \filter_0/reg_i_12[2] , \filter_0/reg_i_12[3] ,
         \filter_0/reg_i_12[4] , \filter_0/reg_i_12[5] ,
         \filter_0/reg_i_12[6] , \filter_0/reg_i_12[7] ,
         \filter_0/reg_i_12[8] , \filter_0/reg_i_12[9] ,
         \filter_0/reg_i_12[10] , \filter_0/reg_i_12[11] ,
         \filter_0/reg_i_12[12] , \filter_0/reg_i_12[13] ,
         \filter_0/reg_i_12[14] , \filter_0/reg_i_12[15] ,
         \filter_0/reg_i_12[16] , \filter_0/reg_i_12[17] ,
         \filter_0/reg_i_12[18] , \filter_0/reg_i_12[19] ,
         \filter_0/reg_i_11[0] , \filter_0/reg_i_11[1] ,
         \filter_0/reg_i_11[2] , \filter_0/reg_i_11[3] ,
         \filter_0/reg_i_11[4] , \filter_0/reg_i_11[5] ,
         \filter_0/reg_i_11[6] , \filter_0/reg_i_11[7] ,
         \filter_0/reg_i_11[8] , \filter_0/reg_i_11[9] ,
         \filter_0/reg_i_11[10] , \filter_0/reg_i_11[11] ,
         \filter_0/reg_i_11[12] , \filter_0/reg_i_11[13] ,
         \filter_0/reg_i_11[14] , \filter_0/reg_i_11[15] ,
         \filter_0/reg_i_11[16] , \filter_0/reg_i_11[17] ,
         \filter_0/reg_i_11[18] , \filter_0/reg_i_11[19] ,
         \filter_0/reg_i_10[0] , \filter_0/reg_i_10[1] ,
         \filter_0/reg_i_10[2] , \filter_0/reg_i_10[3] ,
         \filter_0/reg_i_10[4] , \filter_0/reg_i_10[5] ,
         \filter_0/reg_i_10[6] , \filter_0/reg_i_10[7] ,
         \filter_0/reg_i_10[8] , \filter_0/reg_i_10[9] ,
         \filter_0/reg_i_10[10] , \filter_0/reg_i_10[11] ,
         \filter_0/reg_i_10[12] , \filter_0/reg_i_10[13] ,
         \filter_0/reg_i_10[14] , \filter_0/reg_i_10[15] ,
         \filter_0/reg_i_10[16] , \filter_0/reg_i_10[17] ,
         \filter_0/reg_i_10[18] , \filter_0/reg_i_10[19] ,
         \filter_0/reg_i_9[0] , \filter_0/reg_i_9[1] , \filter_0/reg_i_9[2] ,
         \filter_0/reg_i_9[3] , \filter_0/reg_i_9[4] , \filter_0/reg_i_9[5] ,
         \filter_0/reg_i_9[6] , \filter_0/reg_i_9[7] , \filter_0/reg_i_9[8] ,
         \filter_0/reg_i_9[9] , \filter_0/reg_i_9[10] , \filter_0/reg_i_9[11] ,
         \filter_0/reg_i_9[12] , \filter_0/reg_i_9[13] ,
         \filter_0/reg_i_9[14] , \filter_0/reg_i_9[15] ,
         \filter_0/reg_i_9[16] , \filter_0/reg_i_9[17] ,
         \filter_0/reg_i_9[18] , \filter_0/reg_i_9[19] , \filter_0/reg_i_8[0] ,
         \filter_0/reg_i_8[1] , \filter_0/reg_i_8[2] , \filter_0/reg_i_8[3] ,
         \filter_0/reg_i_8[4] , \filter_0/reg_i_8[5] , \filter_0/reg_i_8[6] ,
         \filter_0/reg_i_8[7] , \filter_0/reg_i_8[8] , \filter_0/reg_i_8[9] ,
         \filter_0/reg_i_8[10] , \filter_0/reg_i_8[11] ,
         \filter_0/reg_i_8[12] , \filter_0/reg_i_8[13] ,
         \filter_0/reg_i_8[14] , \filter_0/reg_i_8[15] ,
         \filter_0/reg_i_8[16] , \filter_0/reg_i_8[17] ,
         \filter_0/reg_i_8[18] , \filter_0/reg_i_8[19] , \filter_0/reg_i_7[0] ,
         \filter_0/reg_i_7[1] , \filter_0/reg_i_7[2] , \filter_0/reg_i_7[3] ,
         \filter_0/reg_i_7[4] , \filter_0/reg_i_7[5] , \filter_0/reg_i_7[6] ,
         \filter_0/reg_i_7[7] , \filter_0/reg_i_7[8] , \filter_0/reg_i_7[9] ,
         \filter_0/reg_i_7[10] , \filter_0/reg_i_7[11] ,
         \filter_0/reg_i_7[12] , \filter_0/reg_i_7[13] ,
         \filter_0/reg_i_7[14] , \filter_0/reg_i_7[15] ,
         \filter_0/reg_i_7[16] , \filter_0/reg_i_7[17] ,
         \filter_0/reg_i_7[18] , \filter_0/reg_i_7[19] , \filter_0/reg_i_6[0] ,
         \filter_0/reg_i_6[1] , \filter_0/reg_i_6[2] , \filter_0/reg_i_6[3] ,
         \filter_0/reg_i_6[4] , \filter_0/reg_i_6[5] , \filter_0/reg_i_6[6] ,
         \filter_0/reg_i_6[7] , \filter_0/reg_i_6[8] , \filter_0/reg_i_6[9] ,
         \filter_0/reg_i_6[10] , \filter_0/reg_i_6[11] ,
         \filter_0/reg_i_6[12] , \filter_0/reg_i_6[13] ,
         \filter_0/reg_i_6[14] , \filter_0/reg_i_6[15] ,
         \filter_0/reg_i_6[16] , \filter_0/reg_i_6[17] ,
         \filter_0/reg_i_6[18] , \filter_0/reg_i_6[19] , \filter_0/reg_i_5[0] ,
         \filter_0/reg_i_5[1] , \filter_0/reg_i_5[2] , \filter_0/reg_i_5[3] ,
         \filter_0/reg_i_5[4] , \filter_0/reg_i_5[5] , \filter_0/reg_i_5[6] ,
         \filter_0/reg_i_5[7] , \filter_0/reg_i_5[8] , \filter_0/reg_i_5[9] ,
         \filter_0/reg_i_5[10] , \filter_0/reg_i_5[11] ,
         \filter_0/reg_i_5[12] , \filter_0/reg_i_5[13] ,
         \filter_0/reg_i_5[14] , \filter_0/reg_i_5[15] ,
         \filter_0/reg_i_5[16] , \filter_0/reg_i_5[17] ,
         \filter_0/reg_i_5[18] , \filter_0/reg_i_5[19] , \filter_0/reg_i_4[0] ,
         \filter_0/reg_i_4[1] , \filter_0/reg_i_4[2] , \filter_0/reg_i_4[3] ,
         \filter_0/reg_i_4[4] , \filter_0/reg_i_4[5] , \filter_0/reg_i_4[6] ,
         \filter_0/reg_i_4[7] , \filter_0/reg_i_4[8] , \filter_0/reg_i_4[9] ,
         \filter_0/reg_i_4[10] , \filter_0/reg_i_4[11] ,
         \filter_0/reg_i_4[12] , \filter_0/reg_i_4[13] ,
         \filter_0/reg_i_4[14] , \filter_0/reg_i_4[15] ,
         \filter_0/reg_i_4[16] , \filter_0/reg_i_4[17] ,
         \filter_0/reg_i_4[18] , \filter_0/reg_i_4[19] , \filter_0/reg_i_3[0] ,
         \filter_0/reg_i_3[1] , \filter_0/reg_i_3[2] , \filter_0/reg_i_3[3] ,
         \filter_0/reg_i_3[4] , \filter_0/reg_i_3[5] , \filter_0/reg_i_3[6] ,
         \filter_0/reg_i_3[7] , \filter_0/reg_i_3[8] , \filter_0/reg_i_3[9] ,
         \filter_0/reg_i_3[10] , \filter_0/reg_i_3[11] ,
         \filter_0/reg_i_3[12] , \filter_0/reg_i_3[13] ,
         \filter_0/reg_i_3[14] , \filter_0/reg_i_3[15] ,
         \filter_0/reg_i_3[16] , \filter_0/reg_i_3[17] ,
         \filter_0/reg_i_3[18] , \filter_0/reg_i_3[19] , \filter_0/reg_i_2[0] ,
         \filter_0/reg_i_2[1] , \filter_0/reg_i_2[2] , \filter_0/reg_i_2[3] ,
         \filter_0/reg_i_2[4] , \filter_0/reg_i_2[5] , \filter_0/reg_i_2[6] ,
         \filter_0/reg_i_2[7] , \filter_0/reg_i_2[8] , \filter_0/reg_i_2[9] ,
         \filter_0/reg_i_2[10] , \filter_0/reg_i_2[11] ,
         \filter_0/reg_i_2[12] , \filter_0/reg_i_2[13] ,
         \filter_0/reg_i_2[14] , \filter_0/reg_i_2[15] ,
         \filter_0/reg_i_2[16] , \filter_0/reg_i_2[17] ,
         \filter_0/reg_i_2[18] , \filter_0/reg_i_2[19] , \filter_0/reg_i_1[0] ,
         \filter_0/reg_i_1[1] , \filter_0/reg_i_1[2] , \filter_0/reg_i_1[3] ,
         \filter_0/reg_i_1[4] , \filter_0/reg_i_1[5] , \filter_0/reg_i_1[6] ,
         \filter_0/reg_i_1[7] , \filter_0/reg_i_1[8] , \filter_0/reg_i_1[9] ,
         \filter_0/reg_i_1[10] , \filter_0/reg_i_1[11] ,
         \filter_0/reg_i_1[12] , \filter_0/reg_i_1[13] ,
         \filter_0/reg_i_1[14] , \filter_0/reg_i_1[15] ,
         \filter_0/reg_i_1[16] , \filter_0/reg_i_1[17] ,
         \filter_0/reg_i_1[18] , \filter_0/reg_i_1[19] , \filter_0/reg_i_0[0] ,
         \filter_0/reg_i_0[1] , \filter_0/reg_i_0[2] , \filter_0/reg_i_0[3] ,
         \filter_0/reg_i_0[4] , \filter_0/reg_i_0[5] , \filter_0/reg_i_0[6] ,
         \filter_0/reg_i_0[7] , \filter_0/reg_i_0[8] , \filter_0/reg_i_0[9] ,
         \filter_0/reg_i_0[10] , \filter_0/reg_i_0[11] ,
         \filter_0/reg_i_0[12] , \filter_0/reg_i_0[13] ,
         \filter_0/reg_i_0[14] , \filter_0/reg_i_0[15] ,
         \filter_0/reg_i_0[16] , \filter_0/reg_i_0[17] ,
         \filter_0/reg_i_0[18] , \filter_0/reg_i_0[19] , \filter_0/done ,
         \filter_0/N16 , \filter_0/N15 , \filter_0/N14 , \filter_0/N13 ,
         \filter_0/N12 , \shifter_0/n10886 , \shifter_0/n10885 ,
         \shifter_0/n10884 , \shifter_0/n10883 , \shifter_0/n10882 ,
         \shifter_0/n10881 , \shifter_0/n10880 , \shifter_0/n10879 ,
         \shifter_0/n10878 , \shifter_0/n10877 , \shifter_0/n10876 ,
         \shifter_0/n10875 , \shifter_0/n10874 , \shifter_0/n10873 ,
         \shifter_0/n10872 , \shifter_0/n10871 , \shifter_0/n10870 ,
         \shifter_0/n10869 , \shifter_0/n10868 , \shifter_0/n10867 ,
         \shifter_0/n10866 , \shifter_0/n10865 , \shifter_0/n10864 ,
         \shifter_0/n10863 , \shifter_0/n10862 , \shifter_0/n10861 ,
         \shifter_0/n10860 , \shifter_0/n10859 , \shifter_0/n10858 ,
         \shifter_0/n10857 , \shifter_0/n10856 , \shifter_0/n10855 ,
         \shifter_0/n10854 , \shifter_0/n10853 , \shifter_0/n10852 ,
         \shifter_0/n10851 , \shifter_0/n10850 , \shifter_0/n10849 ,
         \shifter_0/n10848 , \shifter_0/n10847 , \shifter_0/n10846 ,
         \shifter_0/n10845 , \shifter_0/n10844 , \shifter_0/n10843 ,
         \shifter_0/n10842 , \shifter_0/n10841 , \shifter_0/n10840 ,
         \shifter_0/n10839 , \shifter_0/n10838 , \shifter_0/n10837 ,
         \shifter_0/n10836 , \shifter_0/n10835 , \shifter_0/n10834 ,
         \shifter_0/n10833 , \shifter_0/n10832 , \shifter_0/n10831 ,
         \shifter_0/n10830 , \shifter_0/n10829 , \shifter_0/n10828 ,
         \shifter_0/n10827 , \shifter_0/n10826 , \shifter_0/n10825 ,
         \shifter_0/n10824 , \shifter_0/n10823 , \shifter_0/n10822 ,
         \shifter_0/n10821 , \shifter_0/n10820 , \shifter_0/n10819 ,
         \shifter_0/n10818 , \shifter_0/n10817 , \shifter_0/n10816 ,
         \shifter_0/n10815 , \shifter_0/n10814 , \shifter_0/n10813 ,
         \shifter_0/n10812 , \shifter_0/n10811 , \shifter_0/n10810 ,
         \shifter_0/n10809 , \shifter_0/n10808 , \shifter_0/n10807 ,
         \shifter_0/n10806 , \shifter_0/n10805 , \shifter_0/n10804 ,
         \shifter_0/n10803 , \shifter_0/n10802 , \shifter_0/n10801 ,
         \shifter_0/n10800 , \shifter_0/n10799 , \shifter_0/n10798 ,
         \shifter_0/n10797 , \shifter_0/n10796 , \shifter_0/n10795 ,
         \shifter_0/n10794 , \shifter_0/n10793 , \shifter_0/n10792 ,
         \shifter_0/n10791 , \shifter_0/n10790 , \shifter_0/n10789 ,
         \shifter_0/n10788 , \shifter_0/n10787 , \shifter_0/n10786 ,
         \shifter_0/n10785 , \shifter_0/n10784 , \shifter_0/n10783 ,
         \shifter_0/n10782 , \shifter_0/n10781 , \shifter_0/n10780 ,
         \shifter_0/n10779 , \shifter_0/n10778 , \shifter_0/n10777 ,
         \shifter_0/n10776 , \shifter_0/n10775 , \shifter_0/n10774 ,
         \shifter_0/n10773 , \shifter_0/n10772 , \shifter_0/n10771 ,
         \shifter_0/n10770 , \shifter_0/n10769 , \shifter_0/n10768 ,
         \shifter_0/n10767 , \shifter_0/n10766 , \shifter_0/n10765 ,
         \shifter_0/n10764 , \shifter_0/n10763 , \shifter_0/n10762 ,
         \shifter_0/n10761 , \shifter_0/n10760 , \shifter_0/n10759 ,
         \shifter_0/n10758 , \shifter_0/n10757 , \shifter_0/n10756 ,
         \shifter_0/n10755 , \shifter_0/n10754 , \shifter_0/n10753 ,
         \shifter_0/n10752 , \shifter_0/n10751 , \shifter_0/n10750 ,
         \shifter_0/n10749 , \shifter_0/n10748 , \shifter_0/n10747 ,
         \shifter_0/n10746 , \shifter_0/n10745 , \shifter_0/n10744 ,
         \shifter_0/n10743 , \shifter_0/n10742 , \shifter_0/n10741 ,
         \shifter_0/n10740 , \shifter_0/n10739 , \shifter_0/n10738 ,
         \shifter_0/n10737 , \shifter_0/n10736 , \shifter_0/n10735 ,
         \shifter_0/n10734 , \shifter_0/n10733 , \shifter_0/n10732 ,
         \shifter_0/n10731 , \shifter_0/n10730 , \shifter_0/n10729 ,
         \shifter_0/n10728 , \shifter_0/n10727 , \shifter_0/n10726 ,
         \shifter_0/n10725 , \shifter_0/n10724 , \shifter_0/n10723 ,
         \shifter_0/n10722 , \shifter_0/n10721 , \shifter_0/n10720 ,
         \shifter_0/n10719 , \shifter_0/n10718 , \shifter_0/n10717 ,
         \shifter_0/n10716 , \shifter_0/n10715 , \shifter_0/n10714 ,
         \shifter_0/n10713 , \shifter_0/n10712 , \shifter_0/n10711 ,
         \shifter_0/n10710 , \shifter_0/n10709 , \shifter_0/n10708 ,
         \shifter_0/n10707 , \shifter_0/n10706 , \shifter_0/n10705 ,
         \shifter_0/n10704 , \shifter_0/n10703 , \shifter_0/n10702 ,
         \shifter_0/n10701 , \shifter_0/n10700 , \shifter_0/n10699 ,
         \shifter_0/n10698 , \shifter_0/n10697 , \shifter_0/n10696 ,
         \shifter_0/n10695 , \shifter_0/n10694 , \shifter_0/n10693 ,
         \shifter_0/n10692 , \shifter_0/n10691 , \shifter_0/n10690 ,
         \shifter_0/n10689 , \shifter_0/n10688 , \shifter_0/n10687 ,
         \shifter_0/n10686 , \shifter_0/n10685 , \shifter_0/n10684 ,
         \shifter_0/n10683 , \shifter_0/n10682 , \shifter_0/n10681 ,
         \shifter_0/n10680 , \shifter_0/n10679 , \shifter_0/n10678 ,
         \shifter_0/n10677 , \shifter_0/n10676 , \shifter_0/n10675 ,
         \shifter_0/n10674 , \shifter_0/n10673 , \shifter_0/n10672 ,
         \shifter_0/n10671 , \shifter_0/n10670 , \shifter_0/n10669 ,
         \shifter_0/n10668 , \shifter_0/n10667 , \shifter_0/n10666 ,
         \shifter_0/n10665 , \shifter_0/n10664 , \shifter_0/n10663 ,
         \shifter_0/n10662 , \shifter_0/n10661 , \shifter_0/n10660 ,
         \shifter_0/n10659 , \shifter_0/n10658 , \shifter_0/n10657 ,
         \shifter_0/n10656 , \shifter_0/n10655 , \shifter_0/n10654 ,
         \shifter_0/n10653 , \shifter_0/n10652 , \shifter_0/n10651 ,
         \shifter_0/n10650 , \shifter_0/n10649 , \shifter_0/n10648 ,
         \shifter_0/n10647 , \shifter_0/n10646 , \shifter_0/n10645 ,
         \shifter_0/n10644 , \shifter_0/n10643 , \shifter_0/n10642 ,
         \shifter_0/n10641 , \shifter_0/n10640 , \shifter_0/n10639 ,
         \shifter_0/n10638 , \shifter_0/n10637 , \shifter_0/n10636 ,
         \shifter_0/n10635 , \shifter_0/n10634 , \shifter_0/n10633 ,
         \shifter_0/n10632 , \shifter_0/n10631 , \shifter_0/n10630 ,
         \shifter_0/n10629 , \shifter_0/n10628 , \shifter_0/n10627 ,
         \shifter_0/n10626 , \shifter_0/n10625 , \shifter_0/n10624 ,
         \shifter_0/n10623 , \shifter_0/n10622 , \shifter_0/n10621 ,
         \shifter_0/n10620 , \shifter_0/n10619 , \shifter_0/n10618 ,
         \shifter_0/n10617 , \shifter_0/n10616 , \shifter_0/n10615 ,
         \shifter_0/n10614 , \shifter_0/n10613 , \shifter_0/n10612 ,
         \shifter_0/n10611 , \shifter_0/n10610 , \shifter_0/n10609 ,
         \shifter_0/n10608 , \shifter_0/n10607 , \shifter_0/n10606 ,
         \shifter_0/n10605 , \shifter_0/n10604 , \shifter_0/n10603 ,
         \shifter_0/n10602 , \shifter_0/n10601 , \shifter_0/n10600 ,
         \shifter_0/n10599 , \shifter_0/n10598 , \shifter_0/n10597 ,
         \shifter_0/n10596 , \shifter_0/n10595 , \shifter_0/n10594 ,
         \shifter_0/n10593 , \shifter_0/n10592 , \shifter_0/n10591 ,
         \shifter_0/n10590 , \shifter_0/n10589 , \shifter_0/n10588 ,
         \shifter_0/n10587 , \shifter_0/n10586 , \shifter_0/n10585 ,
         \shifter_0/n10584 , \shifter_0/n10583 , \shifter_0/n10582 ,
         \shifter_0/n10581 , \shifter_0/n10580 , \shifter_0/n10579 ,
         \shifter_0/n10578 , \shifter_0/n10577 , \shifter_0/n10576 ,
         \shifter_0/n10575 , \shifter_0/n10574 , \shifter_0/n10573 ,
         \shifter_0/n10572 , \shifter_0/n10571 , \shifter_0/n10570 ,
         \shifter_0/n10569 , \shifter_0/n10568 , \shifter_0/n10567 ,
         \shifter_0/n10566 , \shifter_0/n10565 , \shifter_0/n10564 ,
         \shifter_0/n10563 , \shifter_0/n10562 , \shifter_0/n10561 ,
         \shifter_0/n10560 , \shifter_0/n10559 , \shifter_0/n10558 ,
         \shifter_0/n10557 , \shifter_0/n10556 , \shifter_0/n10555 ,
         \shifter_0/n10554 , \shifter_0/n10553 , \shifter_0/n10552 ,
         \shifter_0/n10551 , \shifter_0/n10550 , \shifter_0/n10549 ,
         \shifter_0/n10548 , \shifter_0/n10547 , \shifter_0/n10546 ,
         \shifter_0/n10545 , \shifter_0/n10544 , \shifter_0/n10543 ,
         \shifter_0/n10542 , \shifter_0/n10541 , \shifter_0/n10540 ,
         \shifter_0/n10539 , \shifter_0/n10538 , \shifter_0/n10537 ,
         \shifter_0/n10536 , \shifter_0/n10535 , \shifter_0/n10534 ,
         \shifter_0/n10533 , \shifter_0/n10532 , \shifter_0/n10531 ,
         \shifter_0/n10530 , \shifter_0/n10529 , \shifter_0/n10528 ,
         \shifter_0/n10527 , \shifter_0/n10526 , \shifter_0/n10525 ,
         \shifter_0/n10524 , \shifter_0/n10523 , \shifter_0/n10522 ,
         \shifter_0/n10521 , \shifter_0/n10520 , \shifter_0/n10519 ,
         \shifter_0/n10518 , \shifter_0/n10517 , \shifter_0/n10516 ,
         \shifter_0/n10515 , \shifter_0/n10514 , \shifter_0/n10513 ,
         \shifter_0/n10512 , \shifter_0/n10511 , \shifter_0/n10510 ,
         \shifter_0/n10509 , \shifter_0/n10508 , \shifter_0/n10507 ,
         \shifter_0/n10506 , \shifter_0/n10505 , \shifter_0/n10504 ,
         \shifter_0/n10503 , \shifter_0/n10502 , \shifter_0/n10501 ,
         \shifter_0/n10500 , \shifter_0/n10499 , \shifter_0/n10498 ,
         \shifter_0/n10497 , \shifter_0/n10496 , \shifter_0/n10495 ,
         \shifter_0/n10494 , \shifter_0/n10493 , \shifter_0/n10492 ,
         \shifter_0/n10491 , \shifter_0/n10490 , \shifter_0/n10489 ,
         \shifter_0/n10488 , \shifter_0/n10487 , \shifter_0/n10486 ,
         \shifter_0/n10485 , \shifter_0/n10484 , \shifter_0/n10483 ,
         \shifter_0/n10482 , \shifter_0/n10481 , \shifter_0/n10480 ,
         \shifter_0/n10479 , \shifter_0/n10478 , \shifter_0/n10477 ,
         \shifter_0/n10476 , \shifter_0/n10475 , \shifter_0/n10474 ,
         \shifter_0/n10473 , \shifter_0/n10472 , \shifter_0/n10471 ,
         \shifter_0/n10470 , \shifter_0/n10469 , \shifter_0/n10468 ,
         \shifter_0/n10467 , \shifter_0/n10466 , \shifter_0/n10465 ,
         \shifter_0/n10464 , \shifter_0/n10463 , \shifter_0/n10462 ,
         \shifter_0/n10461 , \shifter_0/n10460 , \shifter_0/n10459 ,
         \shifter_0/n10458 , \shifter_0/n10457 , \shifter_0/n10456 ,
         \shifter_0/n10455 , \shifter_0/n10454 , \shifter_0/n10453 ,
         \shifter_0/n10452 , \shifter_0/n10451 , \shifter_0/n10450 ,
         \shifter_0/n10449 , \shifter_0/n10448 , \shifter_0/n10447 ,
         \shifter_0/n10446 , \shifter_0/n10445 , \shifter_0/n10444 ,
         \shifter_0/n10443 , \shifter_0/n10442 , \shifter_0/n10441 ,
         \shifter_0/n10440 , \shifter_0/n10439 , \shifter_0/n10438 ,
         \shifter_0/n10437 , \shifter_0/n10436 , \shifter_0/n10435 ,
         \shifter_0/n10434 , \shifter_0/n10433 , \shifter_0/n10432 ,
         \shifter_0/n10431 , \shifter_0/n10430 , \shifter_0/n10429 ,
         \shifter_0/n10428 , \shifter_0/n10427 , \shifter_0/n10426 ,
         \shifter_0/n10425 , \shifter_0/n10424 , \shifter_0/n10423 ,
         \shifter_0/n10422 , \shifter_0/n10421 , \shifter_0/n10420 ,
         \shifter_0/n10419 , \shifter_0/n10418 , \shifter_0/n10417 ,
         \shifter_0/n10416 , \shifter_0/n10415 , \shifter_0/n10414 ,
         \shifter_0/n10413 , \shifter_0/n10412 , \shifter_0/n10411 ,
         \shifter_0/n10410 , \shifter_0/n10409 , \shifter_0/n10408 ,
         \shifter_0/n10407 , \shifter_0/n10406 , \shifter_0/n10405 ,
         \shifter_0/n10404 , \shifter_0/n10403 , \shifter_0/n10402 ,
         \shifter_0/n10401 , \shifter_0/n10400 , \shifter_0/n10399 ,
         \shifter_0/n10398 , \shifter_0/n10397 , \shifter_0/n10396 ,
         \shifter_0/n10395 , \shifter_0/n10394 , \shifter_0/n10393 ,
         \shifter_0/n10392 , \shifter_0/n10391 , \shifter_0/n10390 ,
         \shifter_0/n10389 , \shifter_0/n10388 , \shifter_0/n10387 ,
         \shifter_0/n10386 , \shifter_0/n10385 , \shifter_0/n10384 ,
         \shifter_0/n10383 , \shifter_0/n10382 , \shifter_0/n10381 ,
         \shifter_0/n10380 , \shifter_0/n10379 , \shifter_0/n10378 ,
         \shifter_0/n10377 , \shifter_0/n10376 , \shifter_0/n10375 ,
         \shifter_0/n10374 , \shifter_0/n10373 , \shifter_0/n10372 ,
         \shifter_0/n10371 , \shifter_0/n10370 , \shifter_0/n10369 ,
         \shifter_0/n10368 , \shifter_0/n10367 , \shifter_0/n10366 ,
         \shifter_0/n10365 , \shifter_0/n10364 , \shifter_0/n10363 ,
         \shifter_0/n10362 , \shifter_0/n10361 , \shifter_0/n10360 ,
         \shifter_0/n10359 , \shifter_0/n10358 , \shifter_0/n10357 ,
         \shifter_0/n10356 , \shifter_0/n10355 , \shifter_0/n10354 ,
         \shifter_0/n10353 , \shifter_0/n10352 , \shifter_0/n10351 ,
         \shifter_0/n10350 , \shifter_0/n10349 , \shifter_0/n10348 ,
         \shifter_0/n10347 , \shifter_0/n10346 , \shifter_0/n10345 ,
         \shifter_0/n10344 , \shifter_0/n10343 , \shifter_0/n10342 ,
         \shifter_0/n10341 , \shifter_0/n10340 , \shifter_0/n10339 ,
         \shifter_0/n10338 , \shifter_0/n10337 , \shifter_0/n10336 ,
         \shifter_0/n10335 , \shifter_0/n10334 , \shifter_0/n10333 ,
         \shifter_0/n10332 , \shifter_0/n10331 , \shifter_0/n10330 ,
         \shifter_0/n10329 , \shifter_0/n10328 , \shifter_0/n10327 ,
         \shifter_0/n10326 , \shifter_0/n10325 , \shifter_0/n10324 ,
         \shifter_0/n10323 , \shifter_0/n10322 , \shifter_0/n10321 ,
         \shifter_0/n10320 , \shifter_0/n10319 , \shifter_0/n10318 ,
         \shifter_0/n10317 , \shifter_0/n10316 , \shifter_0/n10315 ,
         \shifter_0/n10314 , \shifter_0/n10313 , \shifter_0/n10312 ,
         \shifter_0/n10311 , \shifter_0/n10310 , \shifter_0/n10309 ,
         \shifter_0/n10308 , \shifter_0/n10307 , \shifter_0/n10306 ,
         \shifter_0/n10305 , \shifter_0/n10304 , \shifter_0/n10303 ,
         \shifter_0/n10302 , \shifter_0/n10301 , \shifter_0/n10300 ,
         \shifter_0/n10299 , \shifter_0/n10298 , \shifter_0/n10297 ,
         \shifter_0/n10296 , \shifter_0/n10295 , \shifter_0/n10294 ,
         \shifter_0/n10293 , \shifter_0/n10292 , \shifter_0/n10291 ,
         \shifter_0/n10290 , \shifter_0/n10289 , \shifter_0/n10288 ,
         \shifter_0/n10287 , \shifter_0/n10286 , \shifter_0/n10285 ,
         \shifter_0/n10284 , \shifter_0/n10283 , \shifter_0/n10282 ,
         \shifter_0/n10281 , \shifter_0/n10280 , \shifter_0/n10279 ,
         \shifter_0/n10278 , \shifter_0/n10277 , \shifter_0/n10276 ,
         \shifter_0/n10275 , \shifter_0/n10274 , \shifter_0/n10273 ,
         \shifter_0/n10272 , \shifter_0/n10271 , \shifter_0/n10270 ,
         \shifter_0/n10269 , \shifter_0/n10268 , \shifter_0/n10267 ,
         \shifter_0/n10266 , \shifter_0/n10265 , \shifter_0/n10264 ,
         \shifter_0/n10263 , \shifter_0/n10262 , \shifter_0/n10261 ,
         \shifter_0/n10260 , \shifter_0/n10259 , \shifter_0/n10258 ,
         \shifter_0/n10257 , \shifter_0/n10256 , \shifter_0/n10255 ,
         \shifter_0/n10254 , \shifter_0/n10253 , \shifter_0/n10252 ,
         \shifter_0/n10251 , \shifter_0/n10250 , \shifter_0/n10249 ,
         \shifter_0/n10248 , \shifter_0/n10247 , \shifter_0/n10246 ,
         \shifter_0/n10245 , \shifter_0/n10244 , \shifter_0/n10243 ,
         \shifter_0/n10242 , \shifter_0/n10241 , \shifter_0/n10240 ,
         \shifter_0/n10239 , \shifter_0/n10238 , \shifter_0/n10237 ,
         \shifter_0/n10236 , \shifter_0/n10235 , \shifter_0/n10234 ,
         \shifter_0/n10233 , \shifter_0/n10232 , \shifter_0/n10231 ,
         \shifter_0/n10230 , \shifter_0/n10229 , \shifter_0/n10228 ,
         \shifter_0/n10227 , \shifter_0/n10226 , \shifter_0/n10225 ,
         \shifter_0/n10224 , \shifter_0/n10223 , \shifter_0/n10222 ,
         \shifter_0/n10221 , \shifter_0/n10220 , \shifter_0/n10219 ,
         \shifter_0/n10218 , \shifter_0/n10217 , \shifter_0/n10216 ,
         \shifter_0/n10215 , \shifter_0/n10214 , \shifter_0/n10213 ,
         \shifter_0/n10212 , \shifter_0/n10211 , \shifter_0/n10210 ,
         \shifter_0/n10209 , \shifter_0/n10208 , \shifter_0/n10207 ,
         \shifter_0/n10206 , \shifter_0/n10205 , \shifter_0/n10204 ,
         \shifter_0/n10203 , \shifter_0/n10202 , \shifter_0/n10201 ,
         \shifter_0/n10200 , \shifter_0/n10199 , \shifter_0/n10198 ,
         \shifter_0/n10197 , \shifter_0/n10196 , \shifter_0/n10195 ,
         \shifter_0/n10194 , \shifter_0/n10193 , \shifter_0/n10192 ,
         \shifter_0/n10191 , \shifter_0/n10190 , \shifter_0/n10189 ,
         \shifter_0/n10188 , \shifter_0/n10187 , \shifter_0/n10186 ,
         \shifter_0/n10185 , \shifter_0/n10184 , \shifter_0/n10183 ,
         \shifter_0/n10182 , \shifter_0/n10181 , \shifter_0/n10180 ,
         \shifter_0/n10179 , \shifter_0/n10178 , \shifter_0/n10177 ,
         \shifter_0/n10176 , \shifter_0/n10175 , \shifter_0/n10174 ,
         \shifter_0/n10173 , \shifter_0/n10172 , \shifter_0/n10171 ,
         \shifter_0/n10170 , \shifter_0/n10169 , \shifter_0/n10168 ,
         \shifter_0/n10167 , \shifter_0/n10166 , \shifter_0/n10165 ,
         \shifter_0/n10164 , \shifter_0/n10163 , \shifter_0/n10162 ,
         \shifter_0/n10161 , \shifter_0/n10160 , \shifter_0/n10159 ,
         \shifter_0/n10158 , \shifter_0/n10157 , \shifter_0/n10156 ,
         \shifter_0/n10155 , \shifter_0/n10154 , \shifter_0/n10153 ,
         \shifter_0/n10152 , \shifter_0/n10151 , \shifter_0/n10150 ,
         \shifter_0/n10149 , \shifter_0/n10148 , \shifter_0/n10147 ,
         \shifter_0/n10146 , \shifter_0/n10145 , \shifter_0/n10144 ,
         \shifter_0/n10143 , \shifter_0/n10142 , \shifter_0/n10141 ,
         \shifter_0/n10140 , \shifter_0/n10139 , \shifter_0/n10138 ,
         \shifter_0/n10137 , \shifter_0/n10136 , \shifter_0/n10135 ,
         \shifter_0/n10134 , \shifter_0/n10133 , \shifter_0/n10132 ,
         \shifter_0/n10131 , \shifter_0/n10130 , \shifter_0/n10129 ,
         \shifter_0/n10128 , \shifter_0/n10127 , \shifter_0/n10126 ,
         \shifter_0/n10125 , \shifter_0/n10124 , \shifter_0/n10123 ,
         \shifter_0/n10122 , \shifter_0/n10121 , \shifter_0/n10120 ,
         \shifter_0/n10119 , \shifter_0/n10118 , \shifter_0/n10117 ,
         \shifter_0/n10116 , \shifter_0/n10115 , \shifter_0/n10114 ,
         \shifter_0/n10113 , \shifter_0/n10112 , \shifter_0/n10111 ,
         \shifter_0/n10110 , \shifter_0/n10109 , \shifter_0/n10108 ,
         \shifter_0/n10107 , \shifter_0/n10106 , \shifter_0/n10105 ,
         \shifter_0/n10104 , \shifter_0/n10103 , \shifter_0/n10102 ,
         \shifter_0/n10101 , \shifter_0/n10100 , \shifter_0/n10099 ,
         \shifter_0/n10098 , \shifter_0/n10097 , \shifter_0/n10096 ,
         \shifter_0/n10095 , \shifter_0/n10094 , \shifter_0/n10093 ,
         \shifter_0/n10092 , \shifter_0/n10091 , \shifter_0/n10090 ,
         \shifter_0/n10089 , \shifter_0/n10088 , \shifter_0/n10087 ,
         \shifter_0/n10086 , \shifter_0/n10085 , \shifter_0/n10084 ,
         \shifter_0/n10083 , \shifter_0/n10082 , \shifter_0/n10081 ,
         \shifter_0/n10080 , \shifter_0/n10079 , \shifter_0/n10078 ,
         \shifter_0/n10077 , \shifter_0/n10076 , \shifter_0/n10075 ,
         \shifter_0/n10074 , \shifter_0/n10073 , \shifter_0/n10072 ,
         \shifter_0/n10071 , \shifter_0/n10070 , \shifter_0/n10069 ,
         \shifter_0/n10068 , \shifter_0/n10067 , \shifter_0/n10066 ,
         \shifter_0/n10065 , \shifter_0/n10064 , \shifter_0/n10063 ,
         \shifter_0/n10062 , \shifter_0/n10061 , \shifter_0/n10060 ,
         \shifter_0/n10059 , \shifter_0/n10058 , \shifter_0/n10057 ,
         \shifter_0/n10056 , \shifter_0/n10055 , \shifter_0/n10054 ,
         \shifter_0/n10053 , \shifter_0/n10052 , \shifter_0/n10051 ,
         \shifter_0/n10050 , \shifter_0/n10049 , \shifter_0/n10048 ,
         \shifter_0/n10047 , \shifter_0/n10046 , \shifter_0/n10045 ,
         \shifter_0/n10044 , \shifter_0/n10043 , \shifter_0/n10042 ,
         \shifter_0/n10041 , \shifter_0/n10040 , \shifter_0/n10039 ,
         \shifter_0/n10038 , \shifter_0/n10037 , \shifter_0/n10036 ,
         \shifter_0/n10035 , \shifter_0/n10034 , \shifter_0/n10033 ,
         \shifter_0/n10032 , \shifter_0/n10031 , \shifter_0/n10030 ,
         \shifter_0/n10029 , \shifter_0/n10028 , \shifter_0/n10027 ,
         \shifter_0/n10026 , \shifter_0/n10025 , \shifter_0/n10024 ,
         \shifter_0/n10023 , \shifter_0/n10022 , \shifter_0/n10021 ,
         \shifter_0/n10020 , \shifter_0/n10019 , \shifter_0/n10018 ,
         \shifter_0/n10017 , \shifter_0/n10016 , \shifter_0/n10015 ,
         \shifter_0/n10014 , \shifter_0/n10013 , \shifter_0/n10012 ,
         \shifter_0/n10011 , \shifter_0/n10010 , \shifter_0/n10009 ,
         \shifter_0/n10008 , \shifter_0/n10007 , \shifter_0/n10006 ,
         \shifter_0/n10005 , \shifter_0/n10004 , \shifter_0/n10003 ,
         \shifter_0/n10002 , \shifter_0/n10001 , \shifter_0/n10000 ,
         \shifter_0/n9999 , \shifter_0/n9998 , \shifter_0/n9997 ,
         \shifter_0/n9996 , \shifter_0/n9995 , \shifter_0/n9994 ,
         \shifter_0/n9993 , \shifter_0/n9992 , \shifter_0/n9991 ,
         \shifter_0/n9990 , \shifter_0/n9989 , \shifter_0/n9988 ,
         \shifter_0/n9987 , \shifter_0/n9986 , \shifter_0/n9985 ,
         \shifter_0/n9984 , \shifter_0/n9983 , \shifter_0/n9982 ,
         \shifter_0/n9981 , \shifter_0/n9980 , \shifter_0/n9979 ,
         \shifter_0/n9978 , \shifter_0/n9977 , \shifter_0/n9976 ,
         \shifter_0/n9975 , \shifter_0/n9974 , \shifter_0/n9973 ,
         \shifter_0/n9972 , \shifter_0/n9971 , \shifter_0/n9970 ,
         \shifter_0/n9969 , \shifter_0/n9968 , \shifter_0/n9967 ,
         \shifter_0/n9966 , \shifter_0/n9965 , \shifter_0/n9964 ,
         \shifter_0/n9963 , \shifter_0/n9962 , \shifter_0/n9961 ,
         \shifter_0/n9960 , \shifter_0/n9959 , \shifter_0/n9958 ,
         \shifter_0/n9957 , \shifter_0/n9956 , \shifter_0/n9955 ,
         \shifter_0/n9954 , \shifter_0/n9953 , \shifter_0/n9952 ,
         \shifter_0/n9951 , \shifter_0/n9950 , \shifter_0/n9949 ,
         \shifter_0/n9948 , \shifter_0/n9947 , \shifter_0/n9946 ,
         \shifter_0/n9945 , \shifter_0/n9944 , \shifter_0/n9943 ,
         \shifter_0/n9942 , \shifter_0/n9941 , \shifter_0/n9940 ,
         \shifter_0/n9939 , \shifter_0/n9938 , \shifter_0/n9937 ,
         \shifter_0/n9936 , \shifter_0/n9935 , \shifter_0/n9934 ,
         \shifter_0/n9933 , \shifter_0/n9932 , \shifter_0/n9931 ,
         \shifter_0/n9930 , \shifter_0/n9929 , \shifter_0/n9928 ,
         \shifter_0/n9927 , \shifter_0/n9926 , \shifter_0/n9925 ,
         \shifter_0/n9924 , \shifter_0/n9923 , \shifter_0/n9922 ,
         \shifter_0/n9921 , \shifter_0/n9920 , \shifter_0/n9919 ,
         \shifter_0/n9918 , \shifter_0/n9917 , \shifter_0/n9916 ,
         \shifter_0/n9915 , \shifter_0/n9914 , \shifter_0/n9913 ,
         \shifter_0/n9912 , \shifter_0/n9911 , \shifter_0/n9910 ,
         \shifter_0/n9909 , \shifter_0/n9908 , \shifter_0/n9907 ,
         \shifter_0/n9906 , \shifter_0/n9905 , \shifter_0/n9904 ,
         \shifter_0/n9903 , \shifter_0/n9902 , \shifter_0/n9901 ,
         \shifter_0/n9900 , \shifter_0/n9899 , \shifter_0/n9898 ,
         \shifter_0/n9897 , \shifter_0/n9896 , \shifter_0/n9895 ,
         \shifter_0/n9894 , \shifter_0/n9893 , \shifter_0/n9892 ,
         \shifter_0/n9891 , \shifter_0/n9890 , \shifter_0/n9889 ,
         \shifter_0/n9888 , \shifter_0/n9887 , \shifter_0/n9886 ,
         \shifter_0/n9885 , \shifter_0/n9884 , \shifter_0/n9883 ,
         \shifter_0/n9882 , \shifter_0/n9881 , \shifter_0/n9880 ,
         \shifter_0/n9879 , \shifter_0/n9878 , \shifter_0/n9877 ,
         \shifter_0/n9876 , \shifter_0/n9875 , \shifter_0/n9874 ,
         \shifter_0/n9873 , \shifter_0/n9872 , \shifter_0/n9871 ,
         \shifter_0/n9870 , \shifter_0/n9869 , \shifter_0/n9868 ,
         \shifter_0/n9867 , \shifter_0/n9866 , \shifter_0/n9865 ,
         \shifter_0/n9864 , \shifter_0/n9863 , \shifter_0/n9862 ,
         \shifter_0/n9861 , \shifter_0/n9860 , \shifter_0/n9859 ,
         \shifter_0/n9858 , \shifter_0/n9857 , \shifter_0/n9856 ,
         \shifter_0/n9855 , \shifter_0/n9854 , \shifter_0/n9853 ,
         \shifter_0/n9852 , \shifter_0/n9851 , \shifter_0/n9850 ,
         \shifter_0/n9849 , \shifter_0/n9848 , \shifter_0/n9847 ,
         \shifter_0/n9846 , \shifter_0/n9845 , \shifter_0/n9844 ,
         \shifter_0/n9843 , \shifter_0/n9842 , \shifter_0/n9841 ,
         \shifter_0/n9840 , \shifter_0/n9839 , \shifter_0/n9838 ,
         \shifter_0/n9837 , \shifter_0/n9836 , \shifter_0/n9835 ,
         \shifter_0/n9834 , \shifter_0/n9833 , \shifter_0/n9832 ,
         \shifter_0/n9831 , \shifter_0/n9830 , \shifter_0/n9829 ,
         \shifter_0/n9828 , \shifter_0/n9827 , \shifter_0/n9826 ,
         \shifter_0/n9825 , \shifter_0/n9824 , \shifter_0/n9823 ,
         \shifter_0/n9822 , \shifter_0/n9821 , \shifter_0/n9820 ,
         \shifter_0/n9819 , \shifter_0/n9818 , \shifter_0/n9817 ,
         \shifter_0/n9816 , \shifter_0/n9815 , \shifter_0/n9814 ,
         \shifter_0/n9813 , \shifter_0/n9812 , \shifter_0/n9811 ,
         \shifter_0/n9810 , \shifter_0/n9809 , \shifter_0/n9808 ,
         \shifter_0/n9807 , \shifter_0/n9806 , \shifter_0/n9805 ,
         \shifter_0/n9804 , \shifter_0/n9803 , \shifter_0/n9802 ,
         \shifter_0/n9801 , \shifter_0/n9800 , \shifter_0/n9799 ,
         \shifter_0/n9798 , \shifter_0/n9797 , \shifter_0/n9796 ,
         \shifter_0/n9795 , \shifter_0/n9794 , \shifter_0/n9793 ,
         \shifter_0/n9792 , \shifter_0/n9791 , \shifter_0/n9790 ,
         \shifter_0/n9789 , \shifter_0/n9788 , \shifter_0/n9787 ,
         \shifter_0/n9786 , \shifter_0/n9785 , \shifter_0/n9784 ,
         \shifter_0/n9783 , \shifter_0/n9782 , \shifter_0/n9781 ,
         \shifter_0/n9780 , \shifter_0/n9779 , \shifter_0/n9778 ,
         \shifter_0/n9777 , \shifter_0/n9776 , \shifter_0/n9775 ,
         \shifter_0/n9774 , \shifter_0/n9773 , \shifter_0/n9772 ,
         \shifter_0/n9771 , \shifter_0/n9770 , \shifter_0/n9769 ,
         \shifter_0/n9768 , \shifter_0/n9767 , \shifter_0/n9766 ,
         \shifter_0/n9765 , \shifter_0/n9764 , \shifter_0/n9763 ,
         \shifter_0/n9762 , \shifter_0/n9761 , \shifter_0/n9760 ,
         \shifter_0/n9759 , \shifter_0/n9758 , \shifter_0/n9757 ,
         \shifter_0/n9756 , \shifter_0/n9755 , \shifter_0/n9754 ,
         \shifter_0/n9753 , \shifter_0/n9752 , \shifter_0/n9751 ,
         \shifter_0/n9750 , \shifter_0/n9749 , \shifter_0/n9748 ,
         \shifter_0/n9747 , \shifter_0/n9746 , \shifter_0/n9745 ,
         \shifter_0/n9744 , \shifter_0/n9743 , \shifter_0/n9742 ,
         \shifter_0/n9741 , \shifter_0/n9740 , \shifter_0/n9739 ,
         \shifter_0/n9738 , \shifter_0/n9737 , \shifter_0/n9736 ,
         \shifter_0/n9735 , \shifter_0/n9734 , \shifter_0/n9733 ,
         \shifter_0/n9732 , \shifter_0/n9731 , \shifter_0/n9730 ,
         \shifter_0/n9729 , \shifter_0/n9728 , \shifter_0/n9727 ,
         \shifter_0/n9726 , \shifter_0/n9725 , \shifter_0/n9724 ,
         \shifter_0/n9723 , \shifter_0/n9722 , \shifter_0/n9721 ,
         \shifter_0/n9720 , \shifter_0/n9719 , \shifter_0/n9718 ,
         \shifter_0/n9717 , \shifter_0/n9716 , \shifter_0/n9715 ,
         \shifter_0/n9714 , \shifter_0/n9713 , \shifter_0/n9712 ,
         \shifter_0/n9711 , \shifter_0/n9710 , \shifter_0/n9709 ,
         \shifter_0/n9708 , \shifter_0/n9707 , \shifter_0/n9706 ,
         \shifter_0/n9705 , \shifter_0/n9704 , \shifter_0/n9703 ,
         \shifter_0/n9702 , \shifter_0/n9701 , \shifter_0/n9700 ,
         \shifter_0/n9699 , \shifter_0/n9698 , \shifter_0/n9697 ,
         \shifter_0/n9696 , \shifter_0/n9695 , \shifter_0/n9694 ,
         \shifter_0/n9693 , \shifter_0/n9692 , \shifter_0/n9691 ,
         \shifter_0/n9690 , \shifter_0/n9689 , \shifter_0/n9688 ,
         \shifter_0/n9687 , \shifter_0/n9686 , \shifter_0/n9685 ,
         \shifter_0/n9684 , \shifter_0/n9683 , \shifter_0/n9682 ,
         \shifter_0/n9681 , \shifter_0/n9680 , \shifter_0/n9679 ,
         \shifter_0/n9678 , \shifter_0/n9677 , \shifter_0/n9676 ,
         \shifter_0/n9675 , \shifter_0/n9674 , \shifter_0/n9673 ,
         \shifter_0/n9672 , \shifter_0/n9671 , \shifter_0/n9670 ,
         \shifter_0/n9669 , \shifter_0/n9668 , \shifter_0/n9667 ,
         \shifter_0/n9666 , \shifter_0/n9665 , \shifter_0/n9664 ,
         \shifter_0/n9663 , \shifter_0/n9662 , \shifter_0/n9661 ,
         \shifter_0/n9660 , \shifter_0/n9659 , \shifter_0/n9658 ,
         \shifter_0/n9657 , \shifter_0/n9656 , \shifter_0/n9655 ,
         \shifter_0/n9654 , \shifter_0/n9653 , \shifter_0/n9652 ,
         \shifter_0/n9651 , \shifter_0/n9650 , \shifter_0/n9649 ,
         \shifter_0/n9648 , \shifter_0/n9647 , \shifter_0/n9646 ,
         \shifter_0/n9645 , \shifter_0/n9644 , \shifter_0/n9643 ,
         \shifter_0/n9642 , \shifter_0/n9641 , \shifter_0/n9640 ,
         \shifter_0/n9639 , \shifter_0/n9638 , \shifter_0/n9637 ,
         \shifter_0/n9636 , \shifter_0/n9635 , \shifter_0/n9634 ,
         \shifter_0/n9633 , \shifter_0/n9632 , \shifter_0/n9631 ,
         \shifter_0/n9630 , \shifter_0/n9629 , \shifter_0/n9628 ,
         \shifter_0/n9627 , \shifter_0/n9626 , \shifter_0/n9625 ,
         \shifter_0/n9624 , \shifter_0/n9623 , \shifter_0/n9622 ,
         \shifter_0/n9621 , \shifter_0/n9620 , \shifter_0/n9619 ,
         \shifter_0/n9618 , \shifter_0/n9617 , \shifter_0/n9616 ,
         \shifter_0/n9615 , \shifter_0/n9614 , \shifter_0/n9613 ,
         \shifter_0/n9612 , \shifter_0/n9611 , \shifter_0/n9610 ,
         \shifter_0/n9609 , \shifter_0/n9608 , \shifter_0/n9607 ,
         \shifter_0/n9606 , \shifter_0/n9605 , \shifter_0/n9604 ,
         \shifter_0/n9603 , \shifter_0/n9602 , \shifter_0/n9601 ,
         \shifter_0/n9600 , \shifter_0/n9599 , \shifter_0/n9598 ,
         \shifter_0/n9597 , \shifter_0/n9596 , \shifter_0/n9595 ,
         \shifter_0/n9594 , \shifter_0/n9593 , \shifter_0/n9592 ,
         \shifter_0/n9591 , \shifter_0/n9590 , \shifter_0/n9589 ,
         \shifter_0/n9588 , \shifter_0/n9587 , \shifter_0/n9586 ,
         \shifter_0/n9585 , \shifter_0/n9584 , \shifter_0/n9583 ,
         \shifter_0/n9582 , \shifter_0/n9581 , \shifter_0/n9580 ,
         \shifter_0/n9579 , \shifter_0/n9578 , \shifter_0/n9577 ,
         \shifter_0/n9576 , \shifter_0/n9575 , \shifter_0/n9574 ,
         \shifter_0/n9573 , \shifter_0/n9572 , \shifter_0/n9571 ,
         \shifter_0/n9570 , \shifter_0/n9569 , \shifter_0/n9568 ,
         \shifter_0/n9567 , \shifter_0/n9566 , \shifter_0/n9565 ,
         \shifter_0/n9564 , \shifter_0/n9563 , \shifter_0/n9562 ,
         \shifter_0/n9561 , \shifter_0/n9560 , \shifter_0/n9559 ,
         \shifter_0/n9558 , \shifter_0/n9557 , \shifter_0/n9556 ,
         \shifter_0/n9555 , \shifter_0/n9554 , \shifter_0/n9553 ,
         \shifter_0/n9552 , \shifter_0/n9551 , \shifter_0/n9550 ,
         \shifter_0/n9549 , \shifter_0/n9548 , \shifter_0/n9547 ,
         \shifter_0/n9546 , \shifter_0/n9545 , \shifter_0/n9544 ,
         \shifter_0/n9543 , \shifter_0/n9542 , \shifter_0/n9541 ,
         \shifter_0/n9540 , \shifter_0/n9539 , \shifter_0/n9538 ,
         \shifter_0/n9537 , \shifter_0/n9536 , \shifter_0/n9535 ,
         \shifter_0/n9534 , \shifter_0/n9533 , \shifter_0/n9532 ,
         \shifter_0/n9531 , \shifter_0/n9530 , \shifter_0/n9529 ,
         \shifter_0/n9528 , \shifter_0/n9527 , \shifter_0/n9526 ,
         \shifter_0/n9525 , \shifter_0/n9524 , \shifter_0/n9523 ,
         \shifter_0/n9522 , \shifter_0/n9521 , \shifter_0/n9520 ,
         \shifter_0/n9519 , \shifter_0/n9518 , \shifter_0/n9517 ,
         \shifter_0/n9516 , \shifter_0/n9515 , \shifter_0/n9514 ,
         \shifter_0/n9513 , \shifter_0/n9512 , \shifter_0/n9511 ,
         \shifter_0/n9510 , \shifter_0/n9509 , \shifter_0/n9508 ,
         \shifter_0/n9507 , \shifter_0/n9506 , \shifter_0/n9505 ,
         \shifter_0/n9504 , \shifter_0/n9503 , \shifter_0/n9502 ,
         \shifter_0/n9501 , \shifter_0/n9500 , \shifter_0/n9499 ,
         \shifter_0/n9498 , \shifter_0/n9497 , \shifter_0/n9496 ,
         \shifter_0/n9495 , \shifter_0/n9494 , \shifter_0/n9493 ,
         \shifter_0/n9492 , \shifter_0/n9491 , \shifter_0/n9490 ,
         \shifter_0/n9489 , \shifter_0/n9488 , \shifter_0/n9487 ,
         \shifter_0/n9486 , \shifter_0/n9485 , \shifter_0/n9484 ,
         \shifter_0/n9483 , \shifter_0/n9482 , \shifter_0/n9481 ,
         \shifter_0/n9480 , \shifter_0/n9479 , \shifter_0/n9478 ,
         \shifter_0/n9477 , \shifter_0/n9476 , \shifter_0/n9475 ,
         \shifter_0/n9474 , \shifter_0/n9473 , \shifter_0/n9472 ,
         \shifter_0/n9471 , \shifter_0/n9470 , \shifter_0/n9469 ,
         \shifter_0/n9468 , \shifter_0/n9467 , \shifter_0/n9466 ,
         \shifter_0/n9465 , \shifter_0/n9464 , \shifter_0/n9463 ,
         \shifter_0/n9462 , \shifter_0/n9461 , \shifter_0/n9460 ,
         \shifter_0/n9459 , \shifter_0/n9458 , \shifter_0/n9457 ,
         \shifter_0/n9456 , \shifter_0/n9455 , \shifter_0/n9454 ,
         \shifter_0/n9453 , \shifter_0/n9452 , \shifter_0/n9451 ,
         \shifter_0/n9450 , \shifter_0/n9449 , \shifter_0/n9448 ,
         \shifter_0/n9447 , \shifter_0/n9446 , \shifter_0/n9445 ,
         \shifter_0/n9444 , \shifter_0/n9443 , \shifter_0/n9442 ,
         \shifter_0/n9441 , \shifter_0/n9440 , \shifter_0/n9439 ,
         \shifter_0/n9438 , \shifter_0/n9437 , \shifter_0/n9436 ,
         \shifter_0/n9435 , \shifter_0/n9434 , \shifter_0/n9433 ,
         \shifter_0/n9432 , \shifter_0/n9431 , \shifter_0/n9430 ,
         \shifter_0/n9429 , \shifter_0/n9428 , \shifter_0/n9427 ,
         \shifter_0/n9426 , \shifter_0/n9425 , \shifter_0/n9424 ,
         \shifter_0/n9423 , \shifter_0/n9422 , \shifter_0/n9421 ,
         \shifter_0/n9420 , \shifter_0/n9419 , \shifter_0/n9418 ,
         \shifter_0/n9417 , \shifter_0/n9416 , \shifter_0/n9415 ,
         \shifter_0/n9414 , \shifter_0/n9413 , \shifter_0/n9412 ,
         \shifter_0/n9411 , \shifter_0/n9410 , \shifter_0/n9409 ,
         \shifter_0/n9408 , \shifter_0/n9407 , \shifter_0/n9406 ,
         \shifter_0/n9405 , \shifter_0/n9404 , \shifter_0/n9403 ,
         \shifter_0/n9402 , \shifter_0/n9401 , \shifter_0/n9400 ,
         \shifter_0/n9399 , \shifter_0/n9398 , \shifter_0/n9397 ,
         \shifter_0/n9396 , \shifter_0/n9395 , \shifter_0/n9394 ,
         \shifter_0/n9393 , \shifter_0/n9392 , \shifter_0/n9391 ,
         \shifter_0/n9390 , \shifter_0/n9389 , \shifter_0/n9388 ,
         \shifter_0/n9387 , \shifter_0/n9386 , \shifter_0/n9385 ,
         \shifter_0/n9384 , \shifter_0/n9383 , \shifter_0/n9382 ,
         \shifter_0/n9381 , \shifter_0/n9380 , \shifter_0/n9379 ,
         \shifter_0/n9378 , \shifter_0/n9377 , \shifter_0/n9376 ,
         \shifter_0/n9375 , \shifter_0/n9374 , \shifter_0/n9373 ,
         \shifter_0/n9372 , \shifter_0/n9371 , \shifter_0/n9370 ,
         \shifter_0/n9369 , \shifter_0/n9368 , \shifter_0/n9367 ,
         \shifter_0/n9366 , \shifter_0/n9365 , \shifter_0/n9364 ,
         \shifter_0/n9363 , \shifter_0/n9362 , \shifter_0/n9361 ,
         \shifter_0/n9360 , \shifter_0/n9359 , \shifter_0/n9358 ,
         \shifter_0/n9357 , \shifter_0/n9356 , \shifter_0/n9355 ,
         \shifter_0/n9354 , \shifter_0/n9353 , \shifter_0/n9352 ,
         \shifter_0/n9351 , \shifter_0/n9350 , \shifter_0/n9349 ,
         \shifter_0/n9348 , \shifter_0/n9347 , \shifter_0/n9346 ,
         \shifter_0/n9345 , \shifter_0/n9344 , \shifter_0/n9343 ,
         \shifter_0/n9342 , \shifter_0/n9341 , \shifter_0/n9340 ,
         \shifter_0/n9339 , \shifter_0/n9338 , \shifter_0/n9337 ,
         \shifter_0/n9336 , \shifter_0/n9335 , \shifter_0/n9334 ,
         \shifter_0/n9333 , \shifter_0/n9332 , \shifter_0/n9331 ,
         \shifter_0/n9330 , \shifter_0/n9329 , \shifter_0/n9328 ,
         \shifter_0/n9327 , \shifter_0/n9326 , \shifter_0/n9325 ,
         \shifter_0/n9324 , \shifter_0/n9323 , \shifter_0/n9322 ,
         \shifter_0/n9321 , \shifter_0/n9320 , \shifter_0/n9319 ,
         \shifter_0/n9318 , \shifter_0/n9317 , \shifter_0/n9316 ,
         \shifter_0/n9315 , \shifter_0/n9314 , \shifter_0/n9313 ,
         \shifter_0/n9312 , \shifter_0/n9311 , \shifter_0/n9310 ,
         \shifter_0/n9309 , \shifter_0/n9308 , \shifter_0/n9307 ,
         \shifter_0/n9306 , \shifter_0/n9305 , \shifter_0/n9304 ,
         \shifter_0/n9303 , \shifter_0/n9302 , \shifter_0/n9301 ,
         \shifter_0/n9300 , \shifter_0/n9299 , \shifter_0/n9298 ,
         \shifter_0/n9297 , \shifter_0/n9296 , \shifter_0/n9295 ,
         \shifter_0/n9294 , \shifter_0/n9293 , \shifter_0/n9292 ,
         \shifter_0/n9291 , \shifter_0/n9290 , \shifter_0/n9289 ,
         \shifter_0/n9288 , \shifter_0/n9287 , \shifter_0/n9286 ,
         \shifter_0/n9285 , \shifter_0/n9284 , \shifter_0/n9283 ,
         \shifter_0/n9282 , \shifter_0/n9281 , \shifter_0/n9280 ,
         \shifter_0/n9279 , \shifter_0/n9278 , \shifter_0/n9277 ,
         \shifter_0/n9276 , \shifter_0/n9275 , \shifter_0/n9274 ,
         \shifter_0/n9273 , \shifter_0/n9272 , \shifter_0/n9271 ,
         \shifter_0/n9270 , \shifter_0/n9269 , \shifter_0/n9268 ,
         \shifter_0/n9267 , \shifter_0/n9266 , \shifter_0/n9265 ,
         \shifter_0/n9264 , \shifter_0/n9263 , \shifter_0/n9262 ,
         \shifter_0/n9261 , \shifter_0/n9260 , \shifter_0/n9259 ,
         \shifter_0/n9258 , \shifter_0/n9257 , \shifter_0/n9256 ,
         \shifter_0/n9255 , \shifter_0/n9254 , \shifter_0/n9253 ,
         \shifter_0/n9252 , \shifter_0/n9251 , \shifter_0/n9250 ,
         \shifter_0/n9249 , \shifter_0/n9248 , \shifter_0/n9247 ,
         \shifter_0/n9246 , \shifter_0/n9245 , \shifter_0/n9244 ,
         \shifter_0/n9243 , \shifter_0/n9242 , \shifter_0/n9241 ,
         \shifter_0/n9240 , \shifter_0/n9239 , \shifter_0/n9238 ,
         \shifter_0/n9237 , \shifter_0/n9236 , \shifter_0/n9235 ,
         \shifter_0/n9234 , \shifter_0/n9233 , \shifter_0/n9232 ,
         \shifter_0/n9231 , \shifter_0/n9230 , \shifter_0/n9229 ,
         \shifter_0/n9228 , \shifter_0/n9227 , \shifter_0/n9226 ,
         \shifter_0/n9225 , \shifter_0/n9224 , \shifter_0/n9223 ,
         \shifter_0/n9222 , \shifter_0/n9221 , \shifter_0/n9220 ,
         \shifter_0/n9219 , \shifter_0/n9218 , \shifter_0/n9217 ,
         \shifter_0/n9216 , \shifter_0/n9215 , \shifter_0/n9214 ,
         \shifter_0/n9213 , \shifter_0/n9212 , \shifter_0/n9211 ,
         \shifter_0/n9210 , \shifter_0/n9209 , \shifter_0/n9208 ,
         \shifter_0/n9207 , \shifter_0/n9206 , \shifter_0/n9205 ,
         \shifter_0/n9204 , \shifter_0/n9203 , \shifter_0/n9202 ,
         \shifter_0/n9201 , \shifter_0/n9200 , \shifter_0/n9199 ,
         \shifter_0/n9198 , \shifter_0/n9197 , \shifter_0/n9196 ,
         \shifter_0/n9195 , \shifter_0/n9194 , \shifter_0/n9193 ,
         \shifter_0/n9192 , \shifter_0/n9191 , \shifter_0/n9190 ,
         \shifter_0/n9189 , \shifter_0/n9188 , \shifter_0/n9187 ,
         \shifter_0/n9186 , \shifter_0/n9185 , \shifter_0/n9184 ,
         \shifter_0/n9183 , \shifter_0/n9182 , \shifter_0/n9181 ,
         \shifter_0/n9180 , \shifter_0/n9179 , \shifter_0/n9178 ,
         \shifter_0/n9177 , \shifter_0/n9176 , \shifter_0/n9175 ,
         \shifter_0/n9174 , \shifter_0/n9173 , \shifter_0/n9172 ,
         \shifter_0/n9171 , \shifter_0/n9170 , \shifter_0/n9169 ,
         \shifter_0/n9168 , \shifter_0/n9167 , \shifter_0/n9166 ,
         \shifter_0/n9165 , \shifter_0/n9164 , \shifter_0/n9163 ,
         \shifter_0/n9162 , \shifter_0/n9161 , \shifter_0/n9160 ,
         \shifter_0/n9159 , \shifter_0/n9158 , \shifter_0/n9157 ,
         \shifter_0/n9156 , \shifter_0/n9155 , \shifter_0/n9154 ,
         \shifter_0/n9153 , \shifter_0/n9152 , \shifter_0/n9151 ,
         \shifter_0/n9150 , \shifter_0/n9149 , \shifter_0/n9148 ,
         \shifter_0/n9147 , \shifter_0/n9146 , \shifter_0/n9145 ,
         \shifter_0/n9144 , \shifter_0/n9143 , \shifter_0/n9142 ,
         \shifter_0/n9141 , \shifter_0/n9140 , \shifter_0/n9139 ,
         \shifter_0/n9138 , \shifter_0/n9137 , \shifter_0/n9136 ,
         \shifter_0/n9135 , \shifter_0/n9134 , \shifter_0/n9133 ,
         \shifter_0/n9132 , \shifter_0/n9131 , \shifter_0/n9130 ,
         \shifter_0/n9129 , \shifter_0/n9128 , \shifter_0/n9127 ,
         \shifter_0/n9126 , \shifter_0/n9125 , \shifter_0/n9124 ,
         \shifter_0/n9123 , \shifter_0/n9122 , \shifter_0/n9121 ,
         \shifter_0/n9120 , \shifter_0/n9119 , \shifter_0/n9118 ,
         \shifter_0/n9117 , \shifter_0/n9116 , \shifter_0/n9115 ,
         \shifter_0/n9114 , \shifter_0/n9113 , \shifter_0/n9112 ,
         \shifter_0/n9111 , \shifter_0/n9110 , \shifter_0/n9109 ,
         \shifter_0/n9108 , \shifter_0/n9107 , \shifter_0/n9106 ,
         \shifter_0/n9105 , \shifter_0/n9104 , \shifter_0/n9103 ,
         \shifter_0/n9102 , \shifter_0/n9101 , \shifter_0/n9100 ,
         \shifter_0/n9099 , \shifter_0/n9098 , \shifter_0/n9097 ,
         \shifter_0/n9096 , \shifter_0/n9095 , \shifter_0/n9094 ,
         \shifter_0/n9093 , \shifter_0/n9092 , \shifter_0/n9091 ,
         \shifter_0/n9090 , \shifter_0/n9089 , \shifter_0/n9088 ,
         \shifter_0/n9087 , \shifter_0/n9086 , \shifter_0/n9085 ,
         \shifter_0/n9084 , \shifter_0/n9083 , \shifter_0/n9082 ,
         \shifter_0/n9081 , \shifter_0/n9080 , \shifter_0/n9079 ,
         \shifter_0/n9078 , \shifter_0/n9077 , \shifter_0/n9076 ,
         \shifter_0/n9075 , \shifter_0/n9074 , \shifter_0/n9073 ,
         \shifter_0/n9072 , \shifter_0/n9071 , \shifter_0/n9070 ,
         \shifter_0/n9069 , \shifter_0/n9068 , \shifter_0/n9067 ,
         \shifter_0/n9066 , \shifter_0/n9065 , \shifter_0/n9064 ,
         \shifter_0/n9063 , \shifter_0/n9062 , \shifter_0/n9061 ,
         \shifter_0/n9060 , \shifter_0/n9059 , \shifter_0/n9058 ,
         \shifter_0/n9057 , \shifter_0/n9056 , \shifter_0/n9055 ,
         \shifter_0/n9054 , \shifter_0/n9053 , \shifter_0/n9052 ,
         \shifter_0/n9051 , \shifter_0/n9050 , \shifter_0/n9049 ,
         \shifter_0/n9048 , \shifter_0/n9047 , \shifter_0/n9046 ,
         \shifter_0/n9045 , \shifter_0/n9044 , \shifter_0/n9043 ,
         \shifter_0/n9042 , \shifter_0/n9041 , \shifter_0/n9040 ,
         \shifter_0/n9039 , \shifter_0/n9038 , \shifter_0/n9037 ,
         \shifter_0/n9036 , \shifter_0/n9035 , \shifter_0/n9034 ,
         \shifter_0/n9033 , \shifter_0/n9032 , \shifter_0/n9031 ,
         \shifter_0/n9030 , \shifter_0/n9029 , \shifter_0/n9028 ,
         \shifter_0/n9027 , \shifter_0/n9026 , \shifter_0/n9025 ,
         \shifter_0/n9024 , \shifter_0/n9023 , \shifter_0/n9022 ,
         \shifter_0/n9021 , \shifter_0/n9020 , \shifter_0/n9019 ,
         \shifter_0/n9018 , \shifter_0/n9017 , \shifter_0/n9016 ,
         \shifter_0/n9015 , \shifter_0/n9014 , \shifter_0/n9013 ,
         \shifter_0/n9012 , \shifter_0/n9011 , \shifter_0/n9010 ,
         \shifter_0/n9009 , \shifter_0/n9008 , \shifter_0/n9007 ,
         \shifter_0/n9006 , \shifter_0/n9005 , \shifter_0/n9004 ,
         \shifter_0/n9003 , \shifter_0/n9002 , \shifter_0/n9001 ,
         \shifter_0/n9000 , \shifter_0/n8999 , \shifter_0/n8998 ,
         \shifter_0/n8997 , \shifter_0/n8996 , \shifter_0/n8995 ,
         \shifter_0/n8994 , \shifter_0/n8993 , \shifter_0/n8992 ,
         \shifter_0/n8991 , \shifter_0/n8990 , \shifter_0/n8989 ,
         \shifter_0/n8988 , \shifter_0/n8987 , \shifter_0/n8986 ,
         \shifter_0/n8985 , \shifter_0/n8984 , \shifter_0/n8983 ,
         \shifter_0/n8982 , \shifter_0/n8981 , \shifter_0/n8980 ,
         \shifter_0/n8979 , \shifter_0/n8978 , \shifter_0/n8977 ,
         \shifter_0/n8976 , \shifter_0/n8975 , \shifter_0/n8974 ,
         \shifter_0/n8973 , \shifter_0/n8972 , \shifter_0/n8971 ,
         \shifter_0/n8970 , \shifter_0/n8969 , \shifter_0/n8968 ,
         \shifter_0/n8967 , \shifter_0/n8966 , \shifter_0/n8965 ,
         \shifter_0/n8964 , \shifter_0/n8963 , \shifter_0/n8962 ,
         \shifter_0/n8961 , \shifter_0/n8960 , \shifter_0/n8959 ,
         \shifter_0/n8958 , \shifter_0/n8957 , \shifter_0/n8956 ,
         \shifter_0/n8955 , \shifter_0/n8954 , \shifter_0/n8953 ,
         \shifter_0/n8952 , \shifter_0/w_pointer[0] , \shifter_0/w_pointer[1] ,
         \shifter_0/w_pointer[2] , \shifter_0/w_pointer[3] ,
         \shifter_0/i_pointer[0] , \shifter_0/i_pointer[1] ,
         \shifter_0/i_pointer[2] , \shifter_0/i_pointer[3] ,
         \shifter_0/pointer[0] , \shifter_0/pointer[1] ,
         \shifter_0/pointer[2] , \shifter_0/pointer[3] ,
         \shifter_0/reg_w_15[0] , \shifter_0/reg_w_15[1] ,
         \shifter_0/reg_w_15[2] , \shifter_0/reg_w_15[3] ,
         \shifter_0/reg_w_15[4] , \shifter_0/reg_w_15[5] ,
         \shifter_0/reg_w_15[6] , \shifter_0/reg_w_15[7] ,
         \shifter_0/reg_w_15[8] , \shifter_0/reg_w_15[9] ,
         \shifter_0/reg_w_15[10] , \shifter_0/reg_w_15[11] ,
         \shifter_0/reg_w_15[12] , \shifter_0/reg_w_15[13] ,
         \shifter_0/reg_w_15[14] , \shifter_0/reg_w_15[15] ,
         \shifter_0/reg_w_15[16] , \shifter_0/reg_w_15[17] ,
         \shifter_0/reg_w_15[18] , \shifter_0/reg_w_15[19] ,
         \shifter_0/reg_w_14[0] , \shifter_0/reg_w_14[1] ,
         \shifter_0/reg_w_14[2] , \shifter_0/reg_w_14[3] ,
         \shifter_0/reg_w_14[4] , \shifter_0/reg_w_14[5] ,
         \shifter_0/reg_w_14[6] , \shifter_0/reg_w_14[7] ,
         \shifter_0/reg_w_14[8] , \shifter_0/reg_w_14[9] ,
         \shifter_0/reg_w_14[10] , \shifter_0/reg_w_14[11] ,
         \shifter_0/reg_w_14[12] , \shifter_0/reg_w_14[13] ,
         \shifter_0/reg_w_14[14] , \shifter_0/reg_w_14[15] ,
         \shifter_0/reg_w_14[16] , \shifter_0/reg_w_14[17] ,
         \shifter_0/reg_w_14[18] , \shifter_0/reg_w_14[19] ,
         \shifter_0/reg_w_13[0] , \shifter_0/reg_w_13[1] ,
         \shifter_0/reg_w_13[2] , \shifter_0/reg_w_13[3] ,
         \shifter_0/reg_w_13[4] , \shifter_0/reg_w_13[5] ,
         \shifter_0/reg_w_13[6] , \shifter_0/reg_w_13[7] ,
         \shifter_0/reg_w_13[8] , \shifter_0/reg_w_13[9] ,
         \shifter_0/reg_w_13[10] , \shifter_0/reg_w_13[11] ,
         \shifter_0/reg_w_13[12] , \shifter_0/reg_w_13[13] ,
         \shifter_0/reg_w_13[14] , \shifter_0/reg_w_13[15] ,
         \shifter_0/reg_w_13[16] , \shifter_0/reg_w_13[17] ,
         \shifter_0/reg_w_13[18] , \shifter_0/reg_w_13[19] ,
         \shifter_0/reg_w_12[0] , \shifter_0/reg_w_12[1] ,
         \shifter_0/reg_w_12[2] , \shifter_0/reg_w_12[3] ,
         \shifter_0/reg_w_12[4] , \shifter_0/reg_w_12[5] ,
         \shifter_0/reg_w_12[6] , \shifter_0/reg_w_12[7] ,
         \shifter_0/reg_w_12[8] , \shifter_0/reg_w_12[9] ,
         \shifter_0/reg_w_12[10] , \shifter_0/reg_w_12[11] ,
         \shifter_0/reg_w_12[12] , \shifter_0/reg_w_12[13] ,
         \shifter_0/reg_w_12[14] , \shifter_0/reg_w_12[15] ,
         \shifter_0/reg_w_12[16] , \shifter_0/reg_w_12[17] ,
         \shifter_0/reg_w_12[18] , \shifter_0/reg_w_12[19] ,
         \shifter_0/reg_w_11[0] , \shifter_0/reg_w_11[1] ,
         \shifter_0/reg_w_11[2] , \shifter_0/reg_w_11[3] ,
         \shifter_0/reg_w_11[4] , \shifter_0/reg_w_11[5] ,
         \shifter_0/reg_w_11[6] , \shifter_0/reg_w_11[7] ,
         \shifter_0/reg_w_11[8] , \shifter_0/reg_w_11[9] ,
         \shifter_0/reg_w_11[10] , \shifter_0/reg_w_11[11] ,
         \shifter_0/reg_w_11[12] , \shifter_0/reg_w_11[13] ,
         \shifter_0/reg_w_11[14] , \shifter_0/reg_w_11[15] ,
         \shifter_0/reg_w_11[16] , \shifter_0/reg_w_11[17] ,
         \shifter_0/reg_w_11[18] , \shifter_0/reg_w_11[19] ,
         \shifter_0/reg_w_10[0] , \shifter_0/reg_w_10[1] ,
         \shifter_0/reg_w_10[2] , \shifter_0/reg_w_10[3] ,
         \shifter_0/reg_w_10[4] , \shifter_0/reg_w_10[5] ,
         \shifter_0/reg_w_10[6] , \shifter_0/reg_w_10[7] ,
         \shifter_0/reg_w_10[8] , \shifter_0/reg_w_10[9] ,
         \shifter_0/reg_w_10[10] , \shifter_0/reg_w_10[11] ,
         \shifter_0/reg_w_10[12] , \shifter_0/reg_w_10[13] ,
         \shifter_0/reg_w_10[14] , \shifter_0/reg_w_10[15] ,
         \shifter_0/reg_w_10[16] , \shifter_0/reg_w_10[17] ,
         \shifter_0/reg_w_10[18] , \shifter_0/reg_w_10[19] ,
         \shifter_0/reg_w_9[0] , \shifter_0/reg_w_9[1] ,
         \shifter_0/reg_w_9[2] , \shifter_0/reg_w_9[3] ,
         \shifter_0/reg_w_9[4] , \shifter_0/reg_w_9[5] ,
         \shifter_0/reg_w_9[6] , \shifter_0/reg_w_9[7] ,
         \shifter_0/reg_w_9[8] , \shifter_0/reg_w_9[9] ,
         \shifter_0/reg_w_9[10] , \shifter_0/reg_w_9[11] ,
         \shifter_0/reg_w_9[12] , \shifter_0/reg_w_9[13] ,
         \shifter_0/reg_w_9[14] , \shifter_0/reg_w_9[15] ,
         \shifter_0/reg_w_9[16] , \shifter_0/reg_w_9[17] ,
         \shifter_0/reg_w_9[18] , \shifter_0/reg_w_9[19] ,
         \shifter_0/reg_w_8[0] , \shifter_0/reg_w_8[1] ,
         \shifter_0/reg_w_8[2] , \shifter_0/reg_w_8[3] ,
         \shifter_0/reg_w_8[4] , \shifter_0/reg_w_8[5] ,
         \shifter_0/reg_w_8[6] , \shifter_0/reg_w_8[7] ,
         \shifter_0/reg_w_8[8] , \shifter_0/reg_w_8[9] ,
         \shifter_0/reg_w_8[10] , \shifter_0/reg_w_8[11] ,
         \shifter_0/reg_w_8[12] , \shifter_0/reg_w_8[13] ,
         \shifter_0/reg_w_8[14] , \shifter_0/reg_w_8[15] ,
         \shifter_0/reg_w_8[16] , \shifter_0/reg_w_8[17] ,
         \shifter_0/reg_w_8[18] , \shifter_0/reg_w_8[19] ,
         \shifter_0/reg_w_7[0] , \shifter_0/reg_w_7[1] ,
         \shifter_0/reg_w_7[2] , \shifter_0/reg_w_7[3] ,
         \shifter_0/reg_w_7[4] , \shifter_0/reg_w_7[5] ,
         \shifter_0/reg_w_7[6] , \shifter_0/reg_w_7[7] ,
         \shifter_0/reg_w_7[8] , \shifter_0/reg_w_7[9] ,
         \shifter_0/reg_w_7[10] , \shifter_0/reg_w_7[11] ,
         \shifter_0/reg_w_7[12] , \shifter_0/reg_w_7[13] ,
         \shifter_0/reg_w_7[14] , \shifter_0/reg_w_7[15] ,
         \shifter_0/reg_w_7[16] , \shifter_0/reg_w_7[17] ,
         \shifter_0/reg_w_7[18] , \shifter_0/reg_w_7[19] ,
         \shifter_0/reg_w_6[0] , \shifter_0/reg_w_6[1] ,
         \shifter_0/reg_w_6[2] , \shifter_0/reg_w_6[3] ,
         \shifter_0/reg_w_6[4] , \shifter_0/reg_w_6[5] ,
         \shifter_0/reg_w_6[6] , \shifter_0/reg_w_6[7] ,
         \shifter_0/reg_w_6[8] , \shifter_0/reg_w_6[9] ,
         \shifter_0/reg_w_6[10] , \shifter_0/reg_w_6[11] ,
         \shifter_0/reg_w_6[12] , \shifter_0/reg_w_6[13] ,
         \shifter_0/reg_w_6[14] , \shifter_0/reg_w_6[15] ,
         \shifter_0/reg_w_6[16] , \shifter_0/reg_w_6[17] ,
         \shifter_0/reg_w_6[18] , \shifter_0/reg_w_6[19] ,
         \shifter_0/reg_w_5[0] , \shifter_0/reg_w_5[1] ,
         \shifter_0/reg_w_5[2] , \shifter_0/reg_w_5[3] ,
         \shifter_0/reg_w_5[4] , \shifter_0/reg_w_5[5] ,
         \shifter_0/reg_w_5[6] , \shifter_0/reg_w_5[7] ,
         \shifter_0/reg_w_5[8] , \shifter_0/reg_w_5[9] ,
         \shifter_0/reg_w_5[10] , \shifter_0/reg_w_5[11] ,
         \shifter_0/reg_w_5[12] , \shifter_0/reg_w_5[13] ,
         \shifter_0/reg_w_5[14] , \shifter_0/reg_w_5[15] ,
         \shifter_0/reg_w_5[16] , \shifter_0/reg_w_5[17] ,
         \shifter_0/reg_w_5[18] , \shifter_0/reg_w_5[19] ,
         \shifter_0/reg_w_4[0] , \shifter_0/reg_w_4[1] ,
         \shifter_0/reg_w_4[2] , \shifter_0/reg_w_4[3] ,
         \shifter_0/reg_w_4[4] , \shifter_0/reg_w_4[5] ,
         \shifter_0/reg_w_4[6] , \shifter_0/reg_w_4[7] ,
         \shifter_0/reg_w_4[8] , \shifter_0/reg_w_4[9] ,
         \shifter_0/reg_w_4[10] , \shifter_0/reg_w_4[11] ,
         \shifter_0/reg_w_4[12] , \shifter_0/reg_w_4[13] ,
         \shifter_0/reg_w_4[14] , \shifter_0/reg_w_4[15] ,
         \shifter_0/reg_w_4[16] , \shifter_0/reg_w_4[17] ,
         \shifter_0/reg_w_4[18] , \shifter_0/reg_w_4[19] ,
         \shifter_0/reg_w_3[0] , \shifter_0/reg_w_3[1] ,
         \shifter_0/reg_w_3[2] , \shifter_0/reg_w_3[3] ,
         \shifter_0/reg_w_3[4] , \shifter_0/reg_w_3[5] ,
         \shifter_0/reg_w_3[6] , \shifter_0/reg_w_3[7] ,
         \shifter_0/reg_w_3[8] , \shifter_0/reg_w_3[9] ,
         \shifter_0/reg_w_3[10] , \shifter_0/reg_w_3[11] ,
         \shifter_0/reg_w_3[12] , \shifter_0/reg_w_3[13] ,
         \shifter_0/reg_w_3[14] , \shifter_0/reg_w_3[15] ,
         \shifter_0/reg_w_3[16] , \shifter_0/reg_w_3[17] ,
         \shifter_0/reg_w_3[18] , \shifter_0/reg_w_3[19] ,
         \shifter_0/reg_w_2[0] , \shifter_0/reg_w_2[1] ,
         \shifter_0/reg_w_2[2] , \shifter_0/reg_w_2[3] ,
         \shifter_0/reg_w_2[4] , \shifter_0/reg_w_2[5] ,
         \shifter_0/reg_w_2[6] , \shifter_0/reg_w_2[7] ,
         \shifter_0/reg_w_2[8] , \shifter_0/reg_w_2[9] ,
         \shifter_0/reg_w_2[10] , \shifter_0/reg_w_2[11] ,
         \shifter_0/reg_w_2[12] , \shifter_0/reg_w_2[13] ,
         \shifter_0/reg_w_2[14] , \shifter_0/reg_w_2[15] ,
         \shifter_0/reg_w_2[16] , \shifter_0/reg_w_2[17] ,
         \shifter_0/reg_w_2[18] , \shifter_0/reg_w_2[19] ,
         \shifter_0/reg_w_1[0] , \shifter_0/reg_w_1[1] ,
         \shifter_0/reg_w_1[2] , \shifter_0/reg_w_1[3] ,
         \shifter_0/reg_w_1[4] , \shifter_0/reg_w_1[5] ,
         \shifter_0/reg_w_1[6] , \shifter_0/reg_w_1[7] ,
         \shifter_0/reg_w_1[8] , \shifter_0/reg_w_1[9] ,
         \shifter_0/reg_w_1[10] , \shifter_0/reg_w_1[11] ,
         \shifter_0/reg_w_1[12] , \shifter_0/reg_w_1[13] ,
         \shifter_0/reg_w_1[14] , \shifter_0/reg_w_1[15] ,
         \shifter_0/reg_w_1[16] , \shifter_0/reg_w_1[17] ,
         \shifter_0/reg_w_1[18] , \shifter_0/reg_w_1[19] ,
         \shifter_0/reg_w_0[0] , \shifter_0/reg_w_0[1] ,
         \shifter_0/reg_w_0[2] , \shifter_0/reg_w_0[3] ,
         \shifter_0/reg_w_0[4] , \shifter_0/reg_w_0[5] ,
         \shifter_0/reg_w_0[6] , \shifter_0/reg_w_0[7] ,
         \shifter_0/reg_w_0[8] , \shifter_0/reg_w_0[9] ,
         \shifter_0/reg_w_0[10] , \shifter_0/reg_w_0[11] ,
         \shifter_0/reg_w_0[12] , \shifter_0/reg_w_0[13] ,
         \shifter_0/reg_w_0[14] , \shifter_0/reg_w_0[15] ,
         \shifter_0/reg_w_0[16] , \shifter_0/reg_w_0[17] ,
         \shifter_0/reg_w_0[18] , \shifter_0/reg_w_0[19] ,
         \shifter_0/reg_i_15[0] , \shifter_0/reg_i_15[1] ,
         \shifter_0/reg_i_15[2] , \shifter_0/reg_i_15[3] ,
         \shifter_0/reg_i_15[4] , \shifter_0/reg_i_15[5] ,
         \shifter_0/reg_i_15[6] , \shifter_0/reg_i_15[7] ,
         \shifter_0/reg_i_15[8] , \shifter_0/reg_i_15[9] ,
         \shifter_0/reg_i_15[10] , \shifter_0/reg_i_15[11] ,
         \shifter_0/reg_i_15[12] , \shifter_0/reg_i_15[13] ,
         \shifter_0/reg_i_15[14] , \shifter_0/reg_i_15[15] ,
         \shifter_0/reg_i_15[16] , \shifter_0/reg_i_15[17] ,
         \shifter_0/reg_i_15[18] , \shifter_0/reg_i_15[19] ,
         \shifter_0/reg_i_14[0] , \shifter_0/reg_i_14[1] ,
         \shifter_0/reg_i_14[2] , \shifter_0/reg_i_14[3] ,
         \shifter_0/reg_i_14[4] , \shifter_0/reg_i_14[5] ,
         \shifter_0/reg_i_14[6] , \shifter_0/reg_i_14[7] ,
         \shifter_0/reg_i_14[8] , \shifter_0/reg_i_14[9] ,
         \shifter_0/reg_i_14[10] , \shifter_0/reg_i_14[11] ,
         \shifter_0/reg_i_14[12] , \shifter_0/reg_i_14[13] ,
         \shifter_0/reg_i_14[14] , \shifter_0/reg_i_14[15] ,
         \shifter_0/reg_i_14[16] , \shifter_0/reg_i_14[17] ,
         \shifter_0/reg_i_14[18] , \shifter_0/reg_i_14[19] ,
         \shifter_0/reg_i_13[0] , \shifter_0/reg_i_13[1] ,
         \shifter_0/reg_i_13[2] , \shifter_0/reg_i_13[3] ,
         \shifter_0/reg_i_13[4] , \shifter_0/reg_i_13[5] ,
         \shifter_0/reg_i_13[6] , \shifter_0/reg_i_13[7] ,
         \shifter_0/reg_i_13[8] , \shifter_0/reg_i_13[9] ,
         \shifter_0/reg_i_13[10] , \shifter_0/reg_i_13[11] ,
         \shifter_0/reg_i_13[12] , \shifter_0/reg_i_13[13] ,
         \shifter_0/reg_i_13[14] , \shifter_0/reg_i_13[15] ,
         \shifter_0/reg_i_13[16] , \shifter_0/reg_i_13[17] ,
         \shifter_0/reg_i_13[18] , \shifter_0/reg_i_13[19] ,
         \shifter_0/reg_i_12[0] , \shifter_0/reg_i_12[1] ,
         \shifter_0/reg_i_12[2] , \shifter_0/reg_i_12[3] ,
         \shifter_0/reg_i_12[4] , \shifter_0/reg_i_12[5] ,
         \shifter_0/reg_i_12[6] , \shifter_0/reg_i_12[7] ,
         \shifter_0/reg_i_12[8] , \shifter_0/reg_i_12[9] ,
         \shifter_0/reg_i_12[10] , \shifter_0/reg_i_12[11] ,
         \shifter_0/reg_i_12[12] , \shifter_0/reg_i_12[13] ,
         \shifter_0/reg_i_12[14] , \shifter_0/reg_i_12[15] ,
         \shifter_0/reg_i_12[16] , \shifter_0/reg_i_12[17] ,
         \shifter_0/reg_i_12[18] , \shifter_0/reg_i_12[19] ,
         \shifter_0/reg_i_11[0] , \shifter_0/reg_i_11[1] ,
         \shifter_0/reg_i_11[2] , \shifter_0/reg_i_11[3] ,
         \shifter_0/reg_i_11[4] , \shifter_0/reg_i_11[5] ,
         \shifter_0/reg_i_11[6] , \shifter_0/reg_i_11[7] ,
         \shifter_0/reg_i_11[8] , \shifter_0/reg_i_11[9] ,
         \shifter_0/reg_i_11[10] , \shifter_0/reg_i_11[11] ,
         \shifter_0/reg_i_11[12] , \shifter_0/reg_i_11[13] ,
         \shifter_0/reg_i_11[14] , \shifter_0/reg_i_11[15] ,
         \shifter_0/reg_i_11[16] , \shifter_0/reg_i_11[17] ,
         \shifter_0/reg_i_11[18] , \shifter_0/reg_i_11[19] ,
         \shifter_0/reg_i_10[0] , \shifter_0/reg_i_10[1] ,
         \shifter_0/reg_i_10[2] , \shifter_0/reg_i_10[3] ,
         \shifter_0/reg_i_10[4] , \shifter_0/reg_i_10[5] ,
         \shifter_0/reg_i_10[6] , \shifter_0/reg_i_10[7] ,
         \shifter_0/reg_i_10[8] , \shifter_0/reg_i_10[9] ,
         \shifter_0/reg_i_10[10] , \shifter_0/reg_i_10[11] ,
         \shifter_0/reg_i_10[12] , \shifter_0/reg_i_10[13] ,
         \shifter_0/reg_i_10[14] , \shifter_0/reg_i_10[15] ,
         \shifter_0/reg_i_10[16] , \shifter_0/reg_i_10[17] ,
         \shifter_0/reg_i_10[18] , \shifter_0/reg_i_10[19] ,
         \shifter_0/reg_i_9[0] , \shifter_0/reg_i_9[1] ,
         \shifter_0/reg_i_9[2] , \shifter_0/reg_i_9[3] ,
         \shifter_0/reg_i_9[4] , \shifter_0/reg_i_9[5] ,
         \shifter_0/reg_i_9[6] , \shifter_0/reg_i_9[7] ,
         \shifter_0/reg_i_9[8] , \shifter_0/reg_i_9[9] ,
         \shifter_0/reg_i_9[10] , \shifter_0/reg_i_9[11] ,
         \shifter_0/reg_i_9[12] , \shifter_0/reg_i_9[13] ,
         \shifter_0/reg_i_9[14] , \shifter_0/reg_i_9[15] ,
         \shifter_0/reg_i_9[16] , \shifter_0/reg_i_9[17] ,
         \shifter_0/reg_i_9[18] , \shifter_0/reg_i_9[19] ,
         \shifter_0/reg_i_8[0] , \shifter_0/reg_i_8[1] ,
         \shifter_0/reg_i_8[2] , \shifter_0/reg_i_8[3] ,
         \shifter_0/reg_i_8[4] , \shifter_0/reg_i_8[5] ,
         \shifter_0/reg_i_8[6] , \shifter_0/reg_i_8[7] ,
         \shifter_0/reg_i_8[8] , \shifter_0/reg_i_8[9] ,
         \shifter_0/reg_i_8[10] , \shifter_0/reg_i_8[11] ,
         \shifter_0/reg_i_8[12] , \shifter_0/reg_i_8[13] ,
         \shifter_0/reg_i_8[14] , \shifter_0/reg_i_8[15] ,
         \shifter_0/reg_i_8[16] , \shifter_0/reg_i_8[17] ,
         \shifter_0/reg_i_8[18] , \shifter_0/reg_i_8[19] ,
         \shifter_0/reg_i_7[0] , \shifter_0/reg_i_7[1] ,
         \shifter_0/reg_i_7[2] , \shifter_0/reg_i_7[3] ,
         \shifter_0/reg_i_7[4] , \shifter_0/reg_i_7[5] ,
         \shifter_0/reg_i_7[6] , \shifter_0/reg_i_7[7] ,
         \shifter_0/reg_i_7[8] , \shifter_0/reg_i_7[9] ,
         \shifter_0/reg_i_7[10] , \shifter_0/reg_i_7[11] ,
         \shifter_0/reg_i_7[12] , \shifter_0/reg_i_7[13] ,
         \shifter_0/reg_i_7[14] , \shifter_0/reg_i_7[15] ,
         \shifter_0/reg_i_7[16] , \shifter_0/reg_i_7[17] ,
         \shifter_0/reg_i_7[18] , \shifter_0/reg_i_7[19] ,
         \shifter_0/reg_i_6[0] , \shifter_0/reg_i_6[1] ,
         \shifter_0/reg_i_6[2] , \shifter_0/reg_i_6[3] ,
         \shifter_0/reg_i_6[4] , \shifter_0/reg_i_6[5] ,
         \shifter_0/reg_i_6[6] , \shifter_0/reg_i_6[7] ,
         \shifter_0/reg_i_6[8] , \shifter_0/reg_i_6[9] ,
         \shifter_0/reg_i_6[10] , \shifter_0/reg_i_6[11] ,
         \shifter_0/reg_i_6[12] , \shifter_0/reg_i_6[13] ,
         \shifter_0/reg_i_6[14] , \shifter_0/reg_i_6[15] ,
         \shifter_0/reg_i_6[16] , \shifter_0/reg_i_6[17] ,
         \shifter_0/reg_i_6[18] , \shifter_0/reg_i_6[19] ,
         \shifter_0/reg_i_5[0] , \shifter_0/reg_i_5[1] ,
         \shifter_0/reg_i_5[2] , \shifter_0/reg_i_5[3] ,
         \shifter_0/reg_i_5[4] , \shifter_0/reg_i_5[5] ,
         \shifter_0/reg_i_5[6] , \shifter_0/reg_i_5[7] ,
         \shifter_0/reg_i_5[8] , \shifter_0/reg_i_5[9] ,
         \shifter_0/reg_i_5[10] , \shifter_0/reg_i_5[11] ,
         \shifter_0/reg_i_5[12] , \shifter_0/reg_i_5[13] ,
         \shifter_0/reg_i_5[14] , \shifter_0/reg_i_5[15] ,
         \shifter_0/reg_i_5[16] , \shifter_0/reg_i_5[17] ,
         \shifter_0/reg_i_5[18] , \shifter_0/reg_i_5[19] ,
         \shifter_0/reg_i_4[0] , \shifter_0/reg_i_4[1] ,
         \shifter_0/reg_i_4[2] , \shifter_0/reg_i_4[3] ,
         \shifter_0/reg_i_4[4] , \shifter_0/reg_i_4[5] ,
         \shifter_0/reg_i_4[6] , \shifter_0/reg_i_4[7] ,
         \shifter_0/reg_i_4[8] , \shifter_0/reg_i_4[9] ,
         \shifter_0/reg_i_4[10] , \shifter_0/reg_i_4[11] ,
         \shifter_0/reg_i_4[12] , \shifter_0/reg_i_4[13] ,
         \shifter_0/reg_i_4[14] , \shifter_0/reg_i_4[15] ,
         \shifter_0/reg_i_4[16] , \shifter_0/reg_i_4[17] ,
         \shifter_0/reg_i_4[18] , \shifter_0/reg_i_4[19] ,
         \shifter_0/reg_i_3[0] , \shifter_0/reg_i_3[1] ,
         \shifter_0/reg_i_3[2] , \shifter_0/reg_i_3[3] ,
         \shifter_0/reg_i_3[4] , \shifter_0/reg_i_3[5] ,
         \shifter_0/reg_i_3[6] , \shifter_0/reg_i_3[7] ,
         \shifter_0/reg_i_3[8] , \shifter_0/reg_i_3[9] ,
         \shifter_0/reg_i_3[10] , \shifter_0/reg_i_3[11] ,
         \shifter_0/reg_i_3[12] , \shifter_0/reg_i_3[13] ,
         \shifter_0/reg_i_3[14] , \shifter_0/reg_i_3[15] ,
         \shifter_0/reg_i_3[16] , \shifter_0/reg_i_3[17] ,
         \shifter_0/reg_i_3[18] , \shifter_0/reg_i_3[19] ,
         \shifter_0/reg_i_2[0] , \shifter_0/reg_i_2[1] ,
         \shifter_0/reg_i_2[2] , \shifter_0/reg_i_2[3] ,
         \shifter_0/reg_i_2[4] , \shifter_0/reg_i_2[5] ,
         \shifter_0/reg_i_2[6] , \shifter_0/reg_i_2[7] ,
         \shifter_0/reg_i_2[8] , \shifter_0/reg_i_2[9] ,
         \shifter_0/reg_i_2[10] , \shifter_0/reg_i_2[11] ,
         \shifter_0/reg_i_2[12] , \shifter_0/reg_i_2[13] ,
         \shifter_0/reg_i_2[14] , \shifter_0/reg_i_2[15] ,
         \shifter_0/reg_i_2[16] , \shifter_0/reg_i_2[17] ,
         \shifter_0/reg_i_2[18] , \shifter_0/reg_i_2[19] ,
         \shifter_0/reg_i_1[0] , \shifter_0/reg_i_1[1] ,
         \shifter_0/reg_i_1[2] , \shifter_0/reg_i_1[3] ,
         \shifter_0/reg_i_1[4] , \shifter_0/reg_i_1[5] ,
         \shifter_0/reg_i_1[6] , \shifter_0/reg_i_1[7] ,
         \shifter_0/reg_i_1[8] , \shifter_0/reg_i_1[9] ,
         \shifter_0/reg_i_1[10] , \shifter_0/reg_i_1[11] ,
         \shifter_0/reg_i_1[12] , \shifter_0/reg_i_1[13] ,
         \shifter_0/reg_i_1[14] , \shifter_0/reg_i_1[15] ,
         \shifter_0/reg_i_1[16] , \shifter_0/reg_i_1[17] ,
         \shifter_0/reg_i_1[18] , \shifter_0/reg_i_1[19] ,
         \shifter_0/reg_i_0[0] , \shifter_0/reg_i_0[1] ,
         \shifter_0/reg_i_0[2] , \shifter_0/reg_i_0[3] ,
         \shifter_0/reg_i_0[4] , \shifter_0/reg_i_0[5] ,
         \shifter_0/reg_i_0[6] , \shifter_0/reg_i_0[7] ,
         \shifter_0/reg_i_0[8] , \shifter_0/reg_i_0[9] ,
         \shifter_0/reg_i_0[10] , \shifter_0/reg_i_0[11] ,
         \shifter_0/reg_i_0[12] , \shifter_0/reg_i_0[13] ,
         \shifter_0/reg_i_0[14] , \shifter_0/reg_i_0[15] ,
         \shifter_0/reg_i_0[16] , \shifter_0/reg_i_0[17] ,
         \shifter_0/reg_i_0[18] , \shifter_0/reg_i_0[19] , n18761, n18762,
         n18763, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,
         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,
         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
         n23633, n23634, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26214, n26215, n26216, n26217, n26218,
         n26219, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
         n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
         n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
         n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
         n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
         n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
         n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
         n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
         n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
         n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700,
         n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
         n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
         n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
         n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
         n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
         n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
         n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
         n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
         n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
         n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
         n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
         n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
         n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844,
         n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
         n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
         n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
         n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
         n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
         n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
         n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
         n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916,
         n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
         n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
         n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
         n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948,
         n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
         n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
         n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
         n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
         n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
         n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
         n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
         n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
         n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020,
         n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
         n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
         n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
         n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
         n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
         n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
         n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
         n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
         n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
         n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108,
         n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
         n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
         n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
         n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
         n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
         n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
         n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
         n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
         n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
         n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
         n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
         n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204,
         n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
         n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
         n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
         n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
         n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
         n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
         n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
         n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
         n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
         n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
         n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
         n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
         n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308,
         n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
         n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
         n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
         n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
         n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
         n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
         n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
         n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
         n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
         n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
         n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
         n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
         n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
         n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
         n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
         n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
         n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
         n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
         n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
         n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
         n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
         n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
         n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
         n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
         n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
         n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
         n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
         n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
         n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
         n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
         n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
         n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
         n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
         n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
         n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588,
         n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
         n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
         n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
         n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
         n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
         n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
         n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
         n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
         n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668,
         n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
         n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
         n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
         n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
         n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
         n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
         n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
         n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732,
         n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
         n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
         n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
         n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
         n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
         n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
         n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
         n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804,
         n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
         n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
         n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
         n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
         n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
         n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
         n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
         n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
         n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884,
         n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
         n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
         n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
         n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
         n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
         n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
         n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
         n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
         n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
         n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
         n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
         n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
         n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
         n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020,
         n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028,
         n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
         n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
         n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
         n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
         n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
         n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
         n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
         n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
         n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100,
         n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
         n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
         n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
         n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
         n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
         n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
         n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
         n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
         n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
         n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
         n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
         n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
         n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
         n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
         n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244,
         n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
         n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
         n28277, n28280, n28281, n28282, n28283, n28284, n28285, n28286,
         n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
         n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
         n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310,
         n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
         n28319, n28320, n28321, n28324, n28325, n28326, n28327, n28328,
         n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336,
         n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344,
         n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352,
         n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
         n28361, n28362, n28363, n28364, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28410, n28411, n28412,
         n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
         n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428,
         n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
         n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
         n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
         n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
         n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469,
         n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477,
         n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485,
         n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
         n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
         n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
         n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28623, n28624, n28625, n28626, n28627, n28628,
         n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
         n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644,
         n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28665, n28666, n28667, n28668, n28669, n28670,
         n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678,
         n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694,
         n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702,
         n28703, n28704, n28705, n28707, n28708, n28709, n28710, n28711,
         n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
         n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
         n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
         n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
         n28744, n28745, n28746, n28747, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28839, n28840, n28841, n28842, n28843, n28844, n28845,
         n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
         n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861,
         n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869,
         n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877,
         n28878, n28879, n28880, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
         n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
         n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
         n29061, n29062, n29063, n29064, n29066, n29067, n29068, n29069,
         n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077,
         n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085,
         n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093,
         n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101,
         n29102, n29103, n29104, n29105, n29106, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29237,
         n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245,
         n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253,
         n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261,
         n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
         n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29279,
         n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
         n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
         n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
         n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421,
         n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429,
         n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437,
         n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445,
         n29446, n29447, n29449, n29450, n29451, n29452, n29453, n29454,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
         n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478,
         n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
         n29487, n29488, n29489, n29490, n29491, n29492, n29494, n29495,
         n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
         n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511,
         n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
         n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527,
         n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29625, n29626, n29627, n29628,
         n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636,
         n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644,
         n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652,
         n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
         n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
         n29669, n29670, \shifter_0/n8950 , \shifter_0/n8949 ,
         \shifter_0/n8946 , \shifter_0/n8945 , \shifter_0/n8942 ,
         \shifter_0/n8941 , \shifter_0/n8938 , \shifter_0/n8937 ,
         \shifter_0/n8934 , \shifter_0/n8933 , \shifter_0/n8930 ,
         \shifter_0/n8929 , \shifter_0/n8926 , \shifter_0/n8925 ,
         \shifter_0/n8922 , \shifter_0/n8921 , \shifter_0/n8918 ,
         \shifter_0/n8917 , \shifter_0/n8914 , \shifter_0/n8913 ,
         \shifter_0/n8910 , \shifter_0/n8909 , \shifter_0/n8906 ,
         \shifter_0/n8905 , \shifter_0/n8902 , \shifter_0/n8901 ,
         \shifter_0/n8898 , \shifter_0/n8897 , \shifter_0/n8894 ,
         \shifter_0/n8893 , \shifter_0/n8890 , \shifter_0/n8889 ,
         \shifter_0/n8886 , \shifter_0/n8885 , \shifter_0/n8882 ,
         \shifter_0/n8881 , \shifter_0/n8878 , \shifter_0/n8877 ,
         \shifter_0/n8874 , \shifter_0/n8873 , \shifter_0/n8870 ,
         \shifter_0/n8869 , \shifter_0/n8866 , \shifter_0/n8865 ,
         \shifter_0/n8862 , \shifter_0/n8861 , \shifter_0/n8858 ,
         \shifter_0/n8857 , \shifter_0/n8854 , \shifter_0/n8853 ,
         \shifter_0/n8850 , \shifter_0/n8849 , \shifter_0/n8846 ,
         \shifter_0/n8845 , \shifter_0/n8842 , \shifter_0/n8841 ,
         \shifter_0/n8838 , \shifter_0/n8837 , \shifter_0/n8834 ,
         \shifter_0/n8833 , \shifter_0/n8830 , \shifter_0/n8829 ,
         \shifter_0/n8826 , \shifter_0/n8825 , \shifter_0/n8822 ,
         \shifter_0/n8821 , \shifter_0/n8818 , \shifter_0/n8817 ,
         \shifter_0/n8814 , \shifter_0/n8813 , \shifter_0/n8810 ,
         \shifter_0/n8809 , \shifter_0/n8806 , \shifter_0/n8805 ,
         \shifter_0/n8802 , \shifter_0/n8801 , \shifter_0/n8798 ,
         \shifter_0/n8797 , \shifter_0/n8794 , \shifter_0/n8793 ,
         \shifter_0/n8790 , \shifter_0/n8789 , \shifter_0/n8786 ,
         \shifter_0/n8785 , \shifter_0/n8782 , \shifter_0/n8781 ,
         \shifter_0/n8778 , \shifter_0/n8777 , \shifter_0/n8774 ,
         \shifter_0/n8773 , \shifter_0/n8770 , \shifter_0/n8769 ,
         \shifter_0/n8766 , \shifter_0/n8765 , \shifter_0/n8762 ,
         \shifter_0/n8761 , \shifter_0/n8758 , \shifter_0/n8757 ,
         \shifter_0/n8754 , \shifter_0/n8753 , \shifter_0/n8750 ,
         \shifter_0/n8749 , \shifter_0/n8746 , \shifter_0/n8745 ,
         \shifter_0/n8742 , \shifter_0/n8741 , \shifter_0/n8738 ,
         \shifter_0/n8737 , \shifter_0/n8734 , \shifter_0/n8733 ,
         \shifter_0/n8730 , \shifter_0/n8729 , \shifter_0/n8726 ,
         \shifter_0/n8725 , \shifter_0/n8722 , \shifter_0/n8721 ,
         \shifter_0/n8718 , \shifter_0/n8717 , \shifter_0/n8714 ,
         \shifter_0/n8713 , \shifter_0/n8710 , \shifter_0/n8709 ,
         \shifter_0/n8706 , \shifter_0/n8705 , \shifter_0/n8702 ,
         \shifter_0/n8701 , \shifter_0/n8698 , \shifter_0/n8697 ,
         \shifter_0/n8694 , \shifter_0/n8693 , \shifter_0/n8690 ,
         \shifter_0/n8689 , \shifter_0/n8686 , \shifter_0/n8685 ,
         \shifter_0/n8682 , \shifter_0/n8681 , \shifter_0/n8678 ,
         \shifter_0/n8677 , \shifter_0/n8674 , \shifter_0/n8673 ,
         \shifter_0/n8670 , \shifter_0/n8669 , \shifter_0/n8666 ,
         \shifter_0/n8665 , \shifter_0/n8662 , \shifter_0/n8661 ,
         \shifter_0/n8658 , \shifter_0/n8657 , \shifter_0/n8654 ,
         \shifter_0/n8653 , \shifter_0/n8650 , \shifter_0/n8649 ,
         \shifter_0/n8646 , \shifter_0/n8645 , \shifter_0/n8642 ,
         \shifter_0/n8641 , \shifter_0/n8638 , \shifter_0/n8637 ,
         \shifter_0/n8634 , \shifter_0/n8633 , \shifter_0/n8630 ,
         \shifter_0/n8629 , \shifter_0/n8626 , \shifter_0/n8625 ,
         \shifter_0/n8622 , \shifter_0/n8621 , \shifter_0/n8618 ,
         \shifter_0/n8617 , \shifter_0/n8614 , \shifter_0/n8613 ,
         \shifter_0/n8610 , \shifter_0/n8609 , \shifter_0/n8606 ,
         \shifter_0/n8605 , \shifter_0/n8602 , \shifter_0/n8601 ,
         \shifter_0/n8598 , \shifter_0/n8597 , \shifter_0/n8594 ,
         \shifter_0/n8593 , \shifter_0/n8590 , \shifter_0/n8589 ,
         \shifter_0/n8586 , \shifter_0/n8585 , \shifter_0/n8582 ,
         \shifter_0/n8581 , \shifter_0/n8578 , \shifter_0/n8577 ,
         \shifter_0/n8574 , \shifter_0/n8573 , \shifter_0/n8570 ,
         \shifter_0/n8569 , \shifter_0/n8566 , \shifter_0/n8565 ,
         \shifter_0/n8562 , \shifter_0/n8561 , \shifter_0/n8558 ,
         \shifter_0/n8557 , \shifter_0/n8554 , \shifter_0/n8553 ,
         \shifter_0/n8550 , \shifter_0/n8549 , \shifter_0/n8546 ,
         \shifter_0/n8545 , \shifter_0/n8542 , \shifter_0/n8541 ,
         \shifter_0/n8538 , \shifter_0/n8537 , \shifter_0/n8534 ,
         \shifter_0/n8533 , \shifter_0/n8530 , \shifter_0/n8529 ,
         \shifter_0/n8526 , \shifter_0/n8525 , \shifter_0/n8522 ,
         \shifter_0/n8521 , \shifter_0/n8518 , \shifter_0/n8517 ,
         \shifter_0/n8514 , \shifter_0/n8513 , \shifter_0/n8510 ,
         \shifter_0/n8509 , \shifter_0/n8506 , \shifter_0/n8505 ,
         \shifter_0/n8502 , \shifter_0/n8501 , \shifter_0/n8498 ,
         \shifter_0/n8497 , \shifter_0/n8494 , \shifter_0/n8493 ,
         \shifter_0/n8490 , \shifter_0/n8489 , \shifter_0/n8486 ,
         \shifter_0/n8485 , \shifter_0/n8482 , \shifter_0/n8481 ,
         \shifter_0/n8478 , \shifter_0/n8477 , \shifter_0/n8474 ,
         \shifter_0/n8473 , \shifter_0/n8470 , \shifter_0/n8469 ,
         \shifter_0/n8466 , \shifter_0/n8465 , \shifter_0/n8462 ,
         \shifter_0/n8461 , \shifter_0/n8458 , \shifter_0/n8457 ,
         \shifter_0/n8454 , \shifter_0/n8453 , \shifter_0/n8450 ,
         \shifter_0/n8449 , \shifter_0/n8446 , \shifter_0/n8445 ,
         \shifter_0/n8442 , \shifter_0/n8441 , \shifter_0/n8438 ,
         \shifter_0/n8437 , \shifter_0/n8434 , \shifter_0/n8433 ,
         \shifter_0/n8430 , \shifter_0/n8429 , \shifter_0/n8426 ,
         \shifter_0/n8425 , \shifter_0/n8422 , \shifter_0/n8421 ,
         \shifter_0/n8418 , \shifter_0/n8417 , \shifter_0/n8414 ,
         \shifter_0/n8413 , \shifter_0/n8410 , \shifter_0/n8409 ,
         \shifter_0/n8406 , \shifter_0/n8405 , \shifter_0/n8402 ,
         \shifter_0/n8401 , \shifter_0/n8398 , \shifter_0/n8397 ,
         \shifter_0/n8394 , \shifter_0/n8393 , \shifter_0/n8390 ,
         \shifter_0/n8389 , \shifter_0/n8386 , \shifter_0/n8385 ,
         \shifter_0/n8382 , \shifter_0/n8381 , \shifter_0/n8378 ,
         \shifter_0/n8377 , \shifter_0/n8374 , \shifter_0/n8373 ,
         \shifter_0/n8370 , \shifter_0/n8369 , \shifter_0/n8366 ,
         \shifter_0/n8365 , \shifter_0/n8362 , \shifter_0/n8361 ,
         \shifter_0/n8358 , \shifter_0/n8357 , \shifter_0/n8354 ,
         \shifter_0/n8353 , \shifter_0/n8350 , \shifter_0/n8349 ,
         \shifter_0/n8346 , \shifter_0/n8345 , \shifter_0/n8342 ,
         \shifter_0/n8341 , \shifter_0/n8338 , \shifter_0/n8337 ,
         \shifter_0/n8334 , \shifter_0/n8333 , \shifter_0/n8330 ,
         \shifter_0/n8329 , \shifter_0/n8326 , \shifter_0/n8325 ,
         \shifter_0/n8322 , \shifter_0/n8321 , \shifter_0/n8318 ,
         \shifter_0/n8317 , \shifter_0/n8314 , \shifter_0/n8313 ,
         \shifter_0/n8310 , \shifter_0/n8309 , \shifter_0/n8306 ,
         \shifter_0/n8305 , \shifter_0/n8302 , \shifter_0/n8301 ,
         \shifter_0/n8298 , \shifter_0/n8297 , \shifter_0/n8294 ,
         \shifter_0/n8293 , \shifter_0/n8290 , \shifter_0/n8289 ,
         \shifter_0/n8286 , \shifter_0/n8285 , \shifter_0/n8282 ,
         \shifter_0/n8281 , \shifter_0/n8278 , \shifter_0/n8277 ,
         \shifter_0/n8274 , \shifter_0/n8273 , \shifter_0/n8270 ,
         \shifter_0/n8269 , \shifter_0/n8266 , \shifter_0/n8265 ,
         \shifter_0/n8262 , \shifter_0/n8261 , \shifter_0/n8258 ,
         \shifter_0/n8257 , \shifter_0/n8254 , \shifter_0/n8253 ,
         \shifter_0/n8250 , \shifter_0/n8249 , \shifter_0/n8246 ,
         \shifter_0/n8245 , \shifter_0/n8242 , \shifter_0/n8241 ,
         \shifter_0/n8238 , \shifter_0/n8237 , \shifter_0/n8234 ,
         \shifter_0/n8233 , \shifter_0/n8230 , \shifter_0/n8229 ,
         \shifter_0/n8226 , \shifter_0/n8225 , \shifter_0/n8222 ,
         \shifter_0/n8221 , \shifter_0/n8218 , \shifter_0/n8217 ,
         \shifter_0/n8214 , \shifter_0/n8213 , \shifter_0/n8210 ,
         \shifter_0/n8209 , \shifter_0/n8206 , \shifter_0/n8205 ,
         \shifter_0/n8202 , \shifter_0/n8201 , \shifter_0/n8198 ,
         \shifter_0/n8197 , \shifter_0/n8194 , \shifter_0/n8193 ,
         \shifter_0/n8190 , \shifter_0/n8189 , \shifter_0/n8186 ,
         \shifter_0/n8185 , \shifter_0/n8182 , \shifter_0/n8181 ,
         \shifter_0/n8178 , \shifter_0/n8177 , \shifter_0/n8174 ,
         \shifter_0/n8173 , \shifter_0/n8170 , \shifter_0/n8169 ,
         \shifter_0/n8166 , \shifter_0/n8165 , \shifter_0/n8162 ,
         \shifter_0/n8161 , \shifter_0/n8158 , \shifter_0/n8157 ,
         \shifter_0/n8154 , \shifter_0/n8153 , \shifter_0/n8150 ,
         \shifter_0/n8149 , \shifter_0/n8146 , \shifter_0/n8145 ,
         \shifter_0/n8142 , \shifter_0/n8141 , \shifter_0/n8138 ,
         \shifter_0/n8137 , \shifter_0/n8134 , \shifter_0/n8133 ,
         \shifter_0/n8130 , \shifter_0/n8129 , \shifter_0/n8126 ,
         \shifter_0/n8125 , \shifter_0/n8122 , \shifter_0/n8121 ,
         \shifter_0/n8118 , \shifter_0/n8117 , \shifter_0/n8114 ,
         \shifter_0/n8113 , \shifter_0/n8110 , \shifter_0/n8109 ,
         \shifter_0/n8106 , \shifter_0/n8105 , \shifter_0/n8102 ,
         \shifter_0/n8101 , \shifter_0/n8098 , \shifter_0/n8097 ,
         \shifter_0/n8094 , \shifter_0/n8093 , \shifter_0/n8090 ,
         \shifter_0/n8089 , \shifter_0/n8086 , \shifter_0/n8085 ,
         \shifter_0/n8082 , \shifter_0/n8081 , \shifter_0/n8078 ,
         \shifter_0/n8077 , \shifter_0/n8073 , \shifter_0/n8069 ,
         \shifter_0/n8065 , \shifter_0/n8061 , \shifter_0/n8057 ,
         \shifter_0/n8053 , \shifter_0/n8049 , \shifter_0/n8045 ,
         \shifter_0/n8041 , \shifter_0/n8037 , \shifter_0/n8033 ,
         \shifter_0/n8029 , \shifter_0/n8025 , \shifter_0/n8021 ,
         \shifter_0/n8017 , \shifter_0/n8013 , \shifter_0/n8009 ,
         \shifter_0/n8005 , \shifter_0/n8001 , \shifter_0/n7997 ,
         \shifter_0/n7993 , \shifter_0/n7989 , \shifter_0/n7985 ,
         \shifter_0/n7981 , \shifter_0/n7977 , \shifter_0/n7973 ,
         \shifter_0/n7969 , \shifter_0/n7965 , \shifter_0/n7961 ,
         \shifter_0/n7957 , \shifter_0/n7953 , \shifter_0/n7949 ,
         \shifter_0/n7945 , \shifter_0/n7941 , \shifter_0/n7937 ,
         \shifter_0/n7933 , \shifter_0/n7929 , \shifter_0/n7925 ,
         \shifter_0/n7921 , \shifter_0/n7917 , \shifter_0/n7914 ,
         \shifter_0/n7913 , \shifter_0/n7910 , \shifter_0/n7909 ,
         \shifter_0/n7906 , \shifter_0/n7905 , \shifter_0/n7902 ,
         \shifter_0/n7901 , \shifter_0/n7898 , \shifter_0/n7897 ,
         \shifter_0/n7894 , \shifter_0/n7893 , \shifter_0/n7890 ,
         \shifter_0/n7889 , \shifter_0/n7886 , \shifter_0/n7885 ,
         \shifter_0/n7882 , \shifter_0/n7881 , \shifter_0/n7878 ,
         \shifter_0/n7877 , \shifter_0/n7874 , \shifter_0/n7873 ,
         \shifter_0/n7870 , \shifter_0/n7869 , \shifter_0/n7866 ,
         \shifter_0/n7865 , \shifter_0/n7862 , \shifter_0/n7861 ,
         \shifter_0/n7858 , \shifter_0/n7857 , \shifter_0/n7854 ,
         \shifter_0/n7853 , \shifter_0/n7850 , \shifter_0/n7849 ,
         \shifter_0/n7846 , \shifter_0/n7845 , \shifter_0/n7842 ,
         \shifter_0/n7841 , \shifter_0/n7838 , \shifter_0/n7837 ,
         \shifter_0/n7834 , \shifter_0/n7833 , \shifter_0/n7830 ,
         \shifter_0/n7829 , \shifter_0/n7826 , \shifter_0/n7825 ,
         \shifter_0/n7822 , \shifter_0/n7821 , \shifter_0/n7818 ,
         \shifter_0/n7817 , \shifter_0/n7814 , \shifter_0/n7813 ,
         \shifter_0/n7810 , \shifter_0/n7809 , \shifter_0/n7806 ,
         \shifter_0/n7805 , \shifter_0/n7802 , \shifter_0/n7801 ,
         \shifter_0/n7798 , \shifter_0/n7797 , \shifter_0/n7794 ,
         \shifter_0/n7793 , \shifter_0/n7790 , \shifter_0/n7789 ,
         \shifter_0/n7786 , \shifter_0/n7785 , \shifter_0/n7782 ,
         \shifter_0/n7781 , \shifter_0/n7778 , \shifter_0/n7777 ,
         \shifter_0/n7774 , \shifter_0/n7773 , \shifter_0/n7770 ,
         \shifter_0/n7769 , \shifter_0/n7766 , \shifter_0/n7765 ,
         \shifter_0/n7762 , \shifter_0/n7761 , \shifter_0/n7758 ,
         \shifter_0/n7757 , \shifter_0/n7754 , \shifter_0/n7753 ,
         \shifter_0/n7750 , \shifter_0/n7749 , \shifter_0/n7746 ,
         \shifter_0/n7745 , \shifter_0/n7742 , \shifter_0/n7741 ,
         \shifter_0/n7738 , \shifter_0/n7737 , \shifter_0/n7734 ,
         \shifter_0/n7733 , \shifter_0/n7730 , \shifter_0/n7729 ,
         \shifter_0/n7726 , \shifter_0/n7725 , \shifter_0/n7722 ,
         \shifter_0/n7721 , \shifter_0/n7718 , \shifter_0/n7717 ,
         \shifter_0/n7714 , \shifter_0/n7713 , \shifter_0/n7710 ,
         \shifter_0/n7709 , \shifter_0/n7706 , \shifter_0/n7705 ,
         \shifter_0/n7702 , \shifter_0/n7701 , \shifter_0/n7698 ,
         \shifter_0/n7697 , \shifter_0/n7694 , \shifter_0/n7693 ,
         \shifter_0/n7690 , \shifter_0/n7689 , \shifter_0/n7686 ,
         \shifter_0/n7685 , \shifter_0/n7682 , \shifter_0/n7681 ,
         \shifter_0/n7678 , \shifter_0/n7677 , \shifter_0/n7674 ,
         \shifter_0/n7673 , \shifter_0/n7670 , \shifter_0/n7669 ,
         \shifter_0/n7666 , \shifter_0/n7665 , \shifter_0/n7662 ,
         \shifter_0/n7661 , \shifter_0/n7658 , \shifter_0/n7657 ,
         \shifter_0/n7654 , \shifter_0/n7653 , \shifter_0/n7650 ,
         \shifter_0/n7649 , \shifter_0/n7646 , \shifter_0/n7645 ,
         \shifter_0/n7642 , \shifter_0/n7641 , \shifter_0/n7638 ,
         \shifter_0/n7637 , \shifter_0/n7634 , \shifter_0/n7633 ,
         \shifter_0/n7630 , \shifter_0/n7629 , \shifter_0/n7626 ,
         \shifter_0/n7625 , \shifter_0/n7622 , \shifter_0/n7621 ,
         \shifter_0/n7618 , \shifter_0/n7617 , \shifter_0/n7614 ,
         \shifter_0/n7613 , \shifter_0/n7610 , \shifter_0/n7609 ,
         \shifter_0/n7606 , \shifter_0/n7605 , \shifter_0/n7602 ,
         \shifter_0/n7601 , \shifter_0/n7598 , \shifter_0/n7597 ,
         \shifter_0/n7594 , \shifter_0/n7593 , \shifter_0/n7590 ,
         \shifter_0/n7589 , \shifter_0/n7586 , \shifter_0/n7585 ,
         \shifter_0/n7582 , \shifter_0/n7581 , \shifter_0/n7578 ,
         \shifter_0/n7577 , \shifter_0/n7574 , \shifter_0/n7573 ,
         \shifter_0/n7570 , \shifter_0/n7569 , \shifter_0/n7566 ,
         \shifter_0/n7565 , \shifter_0/n7562 , \shifter_0/n7561 ,
         \shifter_0/n7558 , \shifter_0/n7557 , \shifter_0/n7554 ,
         \shifter_0/n7553 , \shifter_0/n7550 , \shifter_0/n7549 ,
         \shifter_0/n7546 , \shifter_0/n7545 , \shifter_0/n7542 ,
         \shifter_0/n7541 , \shifter_0/n7538 , \shifter_0/n7537 ,
         \shifter_0/n7534 , \shifter_0/n7533 , \shifter_0/n7530 ,
         \shifter_0/n7529 , \shifter_0/n7526 , \shifter_0/n7525 ,
         \shifter_0/n7522 , \shifter_0/n7521 , \shifter_0/n7518 ,
         \shifter_0/n7517 , \shifter_0/n7514 , \shifter_0/n7513 ,
         \shifter_0/n7510 , \shifter_0/n7509 , \shifter_0/n7506 ,
         \shifter_0/n7505 , \shifter_0/n7502 , \shifter_0/n7501 ,
         \shifter_0/n7498 , \shifter_0/n7497 , \shifter_0/n7494 ,
         \shifter_0/n7493 , \shifter_0/n7490 , \shifter_0/n7489 ,
         \shifter_0/n7486 , \shifter_0/n7485 , \shifter_0/n7482 ,
         \shifter_0/n7481 , \shifter_0/n7478 , \shifter_0/n7477 ,
         \shifter_0/n7474 , \shifter_0/n7473 , \shifter_0/n7470 ,
         \shifter_0/n7469 , \shifter_0/n7466 , \shifter_0/n7465 ,
         \shifter_0/n7462 , \shifter_0/n7461 , \shifter_0/n7458 ,
         \shifter_0/n7457 , \shifter_0/n7454 , \shifter_0/n7453 ,
         \shifter_0/n7450 , \shifter_0/n7449 , \shifter_0/n7446 ,
         \shifter_0/n7445 , \shifter_0/n7442 , \shifter_0/n7441 ,
         \shifter_0/n7438 , \shifter_0/n7437 , \shifter_0/n7433 ,
         \shifter_0/n7429 , \shifter_0/n7425 , \shifter_0/n7421 ,
         \shifter_0/n7417 , \shifter_0/n7413 , \shifter_0/n7409 ,
         \shifter_0/n7405 , \shifter_0/n7401 , \shifter_0/n7397 ,
         \shifter_0/n7393 , \shifter_0/n7389 , \shifter_0/n7385 ,
         \shifter_0/n7381 , \shifter_0/n7377 , \shifter_0/n7373 ,
         \shifter_0/n7369 , \shifter_0/n7365 , \shifter_0/n7361 ,
         \shifter_0/n7357 , \shifter_0/n7353 , \shifter_0/n7349 ,
         \shifter_0/n7345 , \shifter_0/n7341 , \shifter_0/n7337 ,
         \shifter_0/n7333 , \shifter_0/n7329 , \shifter_0/n7325 ,
         \shifter_0/n7321 , \shifter_0/n7317 , \shifter_0/n7313 ,
         \shifter_0/n7309 , \shifter_0/n7305 , \shifter_0/n7301 ,
         \shifter_0/n7297 , \shifter_0/n7293 , \shifter_0/n7289 ,
         \shifter_0/n7285 , \shifter_0/n7281 , \shifter_0/n7277 ,
         \shifter_0/n7274 , \shifter_0/n7273 , \shifter_0/n7270 ,
         \shifter_0/n7269 , \shifter_0/n7266 , \shifter_0/n7265 ,
         \shifter_0/n7262 , \shifter_0/n7261 , \shifter_0/n7258 ,
         \shifter_0/n7257 , \shifter_0/n7254 , \shifter_0/n7253 ,
         \shifter_0/n7250 , \shifter_0/n7249 , \shifter_0/n7246 ,
         \shifter_0/n7245 , \shifter_0/n7242 , \shifter_0/n7241 ,
         \shifter_0/n7238 , \shifter_0/n7237 , \shifter_0/n7234 ,
         \shifter_0/n7233 , \shifter_0/n7230 , \shifter_0/n7229 ,
         \shifter_0/n7226 , \shifter_0/n7225 , \shifter_0/n7222 ,
         \shifter_0/n7221 , \shifter_0/n7218 , \shifter_0/n7217 ,
         \shifter_0/n7214 , \shifter_0/n7213 , \shifter_0/n7210 ,
         \shifter_0/n7209 , \shifter_0/n7206 , \shifter_0/n7205 ,
         \shifter_0/n7202 , \shifter_0/n7201 , \shifter_0/n7198 ,
         \shifter_0/n7197 , \shifter_0/n7194 , \shifter_0/n7193 ,
         \shifter_0/n7190 , \shifter_0/n7189 , \shifter_0/n7186 ,
         \shifter_0/n7185 , \shifter_0/n7182 , \shifter_0/n7181 ,
         \shifter_0/n7178 , \shifter_0/n7177 , \shifter_0/n7174 ,
         \shifter_0/n7173 , \shifter_0/n7170 , \shifter_0/n7169 ,
         \shifter_0/n7166 , \shifter_0/n7165 , \shifter_0/n7162 ,
         \shifter_0/n7161 , \shifter_0/n7158 , \shifter_0/n7157 ,
         \shifter_0/n7154 , \shifter_0/n7153 , \shifter_0/n7150 ,
         \shifter_0/n7149 , \shifter_0/n7146 , \shifter_0/n7145 ,
         \shifter_0/n7142 , \shifter_0/n7141 , \shifter_0/n7138 ,
         \shifter_0/n7137 , \shifter_0/n7134 , \shifter_0/n7133 ,
         \shifter_0/n7130 , \shifter_0/n7129 , \shifter_0/n7126 ,
         \shifter_0/n7125 , \shifter_0/n7122 , \shifter_0/n7121 ,
         \shifter_0/n7118 , \shifter_0/n7117 , \shifter_0/n7113 ,
         \shifter_0/n7109 , \shifter_0/n7105 , \shifter_0/n7101 ,
         \shifter_0/n7097 , \shifter_0/n7093 , \shifter_0/n7089 ,
         \shifter_0/n7085 , \shifter_0/n7081 , \shifter_0/n7077 ,
         \shifter_0/n7073 , \shifter_0/n7069 , \shifter_0/n7065 ,
         \shifter_0/n7061 , \shifter_0/n7057 , \shifter_0/n7053 ,
         \shifter_0/n7049 , \shifter_0/n7045 , \shifter_0/n7041 ,
         \shifter_0/n7037 , \shifter_0/n7033 , \shifter_0/n7029 ,
         \shifter_0/n7025 , \shifter_0/n7021 , \shifter_0/n7017 ,
         \shifter_0/n7013 , \shifter_0/n7009 , \shifter_0/n7005 ,
         \shifter_0/n7001 , \shifter_0/n6997 , \shifter_0/n6993 ,
         \shifter_0/n6989 , \shifter_0/n6985 , \shifter_0/n6981 ,
         \shifter_0/n6977 , \shifter_0/n6973 , \shifter_0/n6969 ,
         \shifter_0/n6965 , \shifter_0/n6961 , \shifter_0/n6957 ,
         \shifter_0/n6953 , \shifter_0/n6949 , \shifter_0/n6945 ,
         \shifter_0/n6941 , \shifter_0/n6937 , \shifter_0/n6933 ,
         \shifter_0/n6929 , \shifter_0/n6925 , \shifter_0/n6921 ,
         \shifter_0/n6917 , \shifter_0/n6913 , \shifter_0/n6909 ,
         \shifter_0/n6905 , \shifter_0/n6901 , \shifter_0/n6897 ,
         \shifter_0/n6893 , \shifter_0/n6889 , \shifter_0/n6885 ,
         \shifter_0/n6881 , \shifter_0/n6877 , \shifter_0/n6873 ,
         \shifter_0/n6869 , \shifter_0/n6865 , \shifter_0/n6861 ,
         \shifter_0/n6857 , \shifter_0/n6853 , \shifter_0/n6849 ,
         \shifter_0/n6845 , \shifter_0/n6841 , \shifter_0/n6837 ,
         \shifter_0/n6833 , \shifter_0/n6829 , \shifter_0/n6825 ,
         \shifter_0/n6821 , \shifter_0/n6817 , \shifter_0/n6813 ,
         \shifter_0/n6809 , \shifter_0/n6805 , \shifter_0/n6801 ,
         \shifter_0/n6797 , \shifter_0/n6793 , \shifter_0/n6789 ,
         \shifter_0/n6785 , \shifter_0/n6781 , \shifter_0/n6777 ,
         \shifter_0/n6773 , \shifter_0/n6769 , \shifter_0/n6765 ,
         \shifter_0/n6761 , \shifter_0/n6757 , \shifter_0/n6753 ,
         \shifter_0/n6749 , \shifter_0/n6745 , \shifter_0/n6741 ,
         \shifter_0/n6737 , \shifter_0/n6733 , \shifter_0/n6729 ,
         \shifter_0/n6725 , \shifter_0/n6721 , \shifter_0/n6717 ,
         \shifter_0/n6713 , \shifter_0/n6709 , \shifter_0/n6705 ,
         \shifter_0/n6701 , \shifter_0/n6697 , \shifter_0/n6693 ,
         \shifter_0/n6689 , \shifter_0/n6685 , \shifter_0/n6681 ,
         \shifter_0/n6677 , \shifter_0/n6673 , \shifter_0/n6669 ,
         \shifter_0/n6665 , \shifter_0/n6661 , \shifter_0/n6657 ,
         \shifter_0/n6653 , \shifter_0/n6649 , \shifter_0/n6645 ,
         \shifter_0/n6641 , \shifter_0/n6637 , \shifter_0/n6633 ,
         \shifter_0/n6629 , \shifter_0/n6625 , \shifter_0/n6621 ,
         \shifter_0/n6617 , \shifter_0/n6613 , \shifter_0/n6609 ,
         \shifter_0/n6605 , \shifter_0/n6601 , \shifter_0/n6597 ,
         \shifter_0/n6593 , \shifter_0/n6589 , \shifter_0/n6585 ,
         \shifter_0/n6581 , \shifter_0/n6577 , \shifter_0/n6573 ,
         \shifter_0/n6569 , \shifter_0/n6565 , \shifter_0/n6561 ,
         \shifter_0/n6557 , \shifter_0/n6553 , \shifter_0/n6549 ,
         \shifter_0/n6545 , \shifter_0/n6541 , \shifter_0/n6537 ,
         \shifter_0/n6533 , \shifter_0/n6529 , \shifter_0/n6525 ,
         \shifter_0/n6521 , \shifter_0/n6517 , \shifter_0/n6513 ,
         \shifter_0/n6509 , \shifter_0/n6505 , \shifter_0/n6501 ,
         \shifter_0/n6497 , \shifter_0/n6493 , \shifter_0/n6489 ,
         \shifter_0/n6485 , \shifter_0/n6481 , \shifter_0/n6477 ,
         \shifter_0/n6474 , \shifter_0/n6473 , \shifter_0/n6470 ,
         \shifter_0/n6469 , \shifter_0/n6466 , \shifter_0/n6465 ,
         \shifter_0/n6462 , \shifter_0/n6461 , \shifter_0/n6458 ,
         \shifter_0/n6457 , \shifter_0/n6454 , \shifter_0/n6453 ,
         \shifter_0/n6450 , \shifter_0/n6449 , \shifter_0/n6446 ,
         \shifter_0/n6445 , \shifter_0/n6442 , \shifter_0/n6441 ,
         \shifter_0/n6438 , \shifter_0/n6437 , \shifter_0/n6434 ,
         \shifter_0/n6433 , \shifter_0/n6430 , \shifter_0/n6429 ,
         \shifter_0/n6426 , \shifter_0/n6425 , \shifter_0/n6422 ,
         \shifter_0/n6421 , \shifter_0/n6418 , \shifter_0/n6417 ,
         \shifter_0/n6414 , \shifter_0/n6413 , \shifter_0/n6410 ,
         \shifter_0/n6409 , \shifter_0/n6406 , \shifter_0/n6405 ,
         \shifter_0/n6402 , \shifter_0/n6401 , \shifter_0/n6398 ,
         \shifter_0/n6397 , \shifter_0/n6394 , \shifter_0/n6393 , n15356,
         n15355, n15354, n15353, n15352, n15351, n15350, n15349, n15348,
         n15347, n15346, n15345, n15344, n15343, n15342, n15341, n15340,
         n15339, n15338, n15337, n15336, n15335, n15334, n15333, n15332,
         n15331, n15330, n15329, n15328, n15327, n15326, n15325, n15324,
         n15323, n15322, n15321, n15320, n15319, n15318, n15317, n15316,
         n15315, n15314, n15313, n15312, n15311, n15310, n15309, n15308,
         n15307, n15306, n15305, n15304, n15303, n15302, n15301, n15300,
         n15299, n15298, n15297, n15296, n15295, n15294, n15293, n15292,
         n15291, n15290, n15289, n15288, n15287, n15286, n15285, n15284,
         n15283, n15282, n15281, n15280, n15279, n15278, n15277, n15276,
         n15275, n15274, n15273, n15272, n15271, n15270, n15269, n15268,
         n15267, n15266, n15265, n15264, n15263, n15262, n15261, n15260,
         n15259, n15258, n15257, n15256, n15255, n15254, n15253, n15252,
         n15251, n15250, n15249, n15248, n15247, n15246, n15245, n15244,
         n15243, n15242, n15241, n15240, n15239, n15238, n15237, n15236,
         n15235, n15234, n15233, n15232, n15231, n15230, n15229, n15228,
         n15227, n15226, n15225, n15224, n15223, n15222, n15221, n15220,
         n15219, n15218, n15217, n15216, n15215, n15214, n15213, n15212,
         n15211, n15210, n15209, n15208, n15207, n15206, n15205, n15204,
         n15203, n15202, n15201, n15200, n15199, n15198, n15197, n15195,
         n15194, n15193, n15192, n15191, n15190, n15189, n15188, n15187,
         n15186, n15185, n15184, n15183, n15182, n15181, n15180, n15179,
         n15178, n15177, n15172, n15171, n15170, n15168, n15167, n15166,
         n15165, n15164, n15163, n15162, n15161, n15160, n15159, n15158,
         n15157, n15156, n15155, n15154, n15153, n15152, n15151, n15150,
         n15149, n15148, n15147, n15146, n15145, n15144, n15143, n15142,
         n15141, n15140, n15139, n15138, n15137, n15136, n15135, n15134,
         n15133, n15132, n15131, n15130, n15129, n15128, n15127, n15126,
         n15125, n15124, n15123, n15122, n15121, n15120, n15119, n15118,
         n15117, n15116, n15115, n15114, n15113, n15112, n15111, n15110,
         n15109, n15108, n15107, n15106, n15105, n15104, n15103, n15102,
         n15101, n15100, n15099, n15098, n15097, n15096, n15095, n15094,
         n15093, n15092, n15091, n15090, n15089, n15088, n15087, n15086,
         n15085, n15084, n15083, n15082, n15081, n15080, n15079, n15078,
         n15077, n15076, n15075, n15074, n15073, n15072, n15071, n15070,
         n15069, n15068, n15067, n15066, n15065, n15064, n15063, n15062,
         n15061, n15059, n15058, n15057, n15056, n15055, n15054, n15053,
         n15052, n15051, n15050, n15049, n15048, n15047, n15046, n15045,
         n15044, n15039, n15038, n15037, n15035, n15034, n15032, n15031,
         n15030, n15029, n15028, n15027, n15026, n15025, n15024, n15023,
         n15022, n15021, n15020, n15019, n15018, n15017, n15016, n15015,
         n15014, n15013, n15012, n15011, n15010, n15009, n15008, n15007,
         n15006, n15005, n15004, n15003, n15002, n15001, n15000, n14999,
         n14998, n14997, n14996, n14995, n14994, n14993, n14992, n14991,
         n14990, n14989, n14988, n14987, n14986, n14985, n14984, n14983,
         n14982, n14981, n14980, n14979, n14978, n14977, n14976, n14975,
         n14974, n14973, n14972, n14971, n14970, n14969, n14968, n14967,
         n14966, n14965, n14964, n14963, n14962, n14961, n14960, n14959,
         n14958, n14957, n14956, n14955, n14954, n14953, n14952, n14951,
         n14950, n14949, n14948, n14947, n14946, n14945, n14944, n14943,
         n14942, n14941, n14940, n14939, n14938, n14937, n14936, n14935,
         n14934, n14933, n14932, n14931, n14930, n14929, n14928, n14927,
         n14926, n14925, n14924, n14923, n14922, n14921, n14920, n14919,
         n14918, n14917, n14916, n14915, n14914, n14913, n14912, n14911,
         n14910, n14909, n14908, n14907, n14906, n14905, n14904, n14903,
         n14902, n14901, n14900, n14899, n14898, n14897, n14896, n14895,
         n14894, n14893, n14892, n14891, n14890, n14889, n14888, n14887,
         n14886, n14885, n14884, n14883, n14882, n14881, n14880, n14879,
         n14878, n14877, n14876, n14875, n14874, n14873, n14872, n14871,
         n14870, n14869, n14868, n14867, n14866, n14865, n14864, n14863,
         n14862, n14861, n14860, n14859, n14858, n14857, n14856, n14855,
         n14854, n14853, n14852, n14851, n14850, n14849, n14848, n14847,
         n14846, n14845, n14844, n14843, n14842, n14841, n14840, n14839,
         n14838, n14837, n14836, n14835, n14834, n14833, n14832, n14831,
         n14830, n14829, n14828, n14827, n14826, n14825, n14824, n14823,
         n14822, n14821, n14820, n14819, n14818, n14817, n14816, n14815,
         n14814, n14813, n14812, n14811, n14810, n14809, n14808, n14807,
         n14806, n14805, n14804, n14803, n14802, n14801, n14800, n14799,
         n14798, n14797, n14796, n14795, n14794, n14793, n14792, n14791,
         n14790, n14789, n14788, n14787, n14786, n14785, n14784, n14783,
         n14782, n14781, n14780, n14779, n14778, n14777, n14776, n14775,
         n14774, n14773, n14772, n14771, n14770, n14769, n14768, n14767,
         n14766, n14765, n14764, n14763, n14762, n14761, n14760, n14759,
         n14758, n14757, n14756, n14755, n14754, n14753, n14752, n14751,
         n14750, n14749, n14748, n14747, n14746, n14745, n14744, n14743,
         n14742, n14741, n14740, n14739, n14738, n14737, n14736, n14735,
         n14734, n14733, n14732, n14731, n14730, n14729, n14728, n14727,
         n14726, n14725, n14724, n14723, n14722, n14721, n14720, n14719,
         n14718, n14717, n14716, n14715, n14714, n14713, n14712, n14711,
         n14710, n14709, n14708, n14707, n14706, n14705, n14704, n14703,
         n14702, n14701, n14700, n14699, n14698, n14697, n14696, n14695,
         n14694, n14693, n14692, n14691, n14690, n14689, n14688, n14687,
         n14686, n14685, n14684, n14683, n14682, n14681, n14680, n14679,
         n14678, n14677, n14676, n14675, n14674, n14673, n14672, n14671,
         n14670, n14669, n14668, n14667, n14666, n14665, n14664, n14663,
         n14662, n14661, n14660, n14659, n14658, n14657, n14656, n14655,
         n14654, n14653, n14652, n14651, n14650, n14649, n14648, n14647,
         n14646, n14645, n14644, n14643, n14642, n14641, n14640, n14639,
         n14638, n14637, n14636, n14635, n14634, n14633, n14632, n14631,
         n14630, n14629, n14628, n14627, n14626, n14625, n14624, n14623,
         n14622, n14621, n14620, n14619, n14618, n14617, n14616, n14615,
         n14614, n14613, n14612, n14611, n14610, n14609, n14608, n14607,
         n14606, n14605, n14604, n14603, n14602, n14601, n14600, n14599,
         n14598, n14597, n14596, n14595, n14594, n14593, n14592, n14591,
         n14590, n14589, n14588, n14587, n14586, n14585, n14584, n14583,
         n14582, n14581, n14580, n14579, n14578, n14577, n14576, n14575,
         n14574, n14573, n14572, n14571, n14570, n14569, n14568, n14567,
         n14566, n14565, n14564, n14563, n14562, n14561, n14560, n14559,
         n14558, n14557, n14556, n14555, n14554, n14553, n14552, n14551,
         n14550, n14549, n14548, n14547, n14546, n14545, n14544, n14543,
         n14542, n14541, n14540, n14539, n14538, n14537, n14536, n14535,
         n14534, n14533, n14532, n14531, n14530, n14529, n14528, n14527,
         n14526, n14525, n14524, n14523, n14522, n14521, n14520, n14519,
         n14518, n14517, n14516, n14515, n14514, n14513, n14512, n14511,
         n14510, n14509, n14508, n14507, n14506, n14505, n14504, n14503,
         n14502, n14501, n14500, n14499, n14498, n14497, n14496, n14495,
         n14494, n14493, n14492, n14491, n14490, n14489, n14488, n14487,
         n14486, n14485, n14484, n14483, n14482, n14481, n14480, n14479,
         n14478, n14477, n14476, n14475, n14474, n14473, n14472, n14471,
         n14470, n14469, n14468, n14467, n14466, n14465, n14464, n14463,
         n14462, n14461, n14460, n14459, n14458, n14457, n14456, n14455,
         n14454, n14453, n14452, n14451, n14450, n14449, n14448, n14447,
         n14446, n14445, n14444, n14443, n14442, n14441, n14440, n14439,
         n14438, n14437, n14436, n14435, n14434, n14433, n14432, n14431,
         n14430, n14429, n14428, n14427, n14426, n14425, n14424, n14423,
         n14422, n14421, n14420, n14419, n14418, n14417, n14416, n14415,
         n14414, n14413, n14412, n14411, n14410, n14409, n14408, n14407,
         n14406, n14405, n14404, n14403, n14402, n14401, n14400, n14399,
         n14398, n14397, n14396, n14395, n14394, n14393, n14392, n14391,
         n14390, n14389, n14388, n14387, n14386, n14385, n14384, n14383,
         n14382, n14381, n14380, n14379, n14378, n14377, n14376, n14375,
         n14374, n14373, n14372, n14371, n14370, n14369, n14368, n14367,
         n14366, n14365, n14364, n14363, n14362, n14361, n14360, n14359,
         n14358, n14357, n14356, n14355, n14354, n14353, n14352, n14351,
         n14350, n14349, n14348, n14347, n14346, n14345, n14344, n14343,
         n14342, n14341, n14340, n14339, n14338, n14337, n14336, n14335,
         n14334, n14333, n14332, n14331, n14330, n14329, n14328, n14327,
         n14326, n14325, n14324, n14323, n14322, n14321, n14320, n14319,
         n14318, n14317, n14316, n14315, n14314, n14313, n14312, n14311,
         n14310, n14309, n14308, n14307, n14306, n14305, n14304, n14303,
         n14302, n14301, n14300, n14299, n14298, n14297, n14296, n14295,
         n14294, n14293, n14292, n14291, n14290, n14289, n14288, n14287,
         n14286, n14285, n14284, n14283, n14282, n14281, n14280, n14279,
         n14278, n14277, n14276, n14275, n14274, n14273, n14272, n14271,
         n14270, n14269, n14268, n14267, n14266, n14265, n14264, n14263,
         n14262, n14261, n14260, n14259, n14258, n14257, n14256, n14255,
         n14254, n14253, n14252, n14251, n14250, n14249, n14248, n14247,
         n14246, n14245, n14244, n14243, n14242, n14241, n14240, n14239,
         n14238, n14237, n14236, n14235, n14234, n14233, n14232, n14231,
         n14230, n14229, n14228, n14227, n14226, n14225, n14224, n14223,
         n14222, n14221, n14220, n14219, n14218, n14217, n14216, n14215,
         n14214, n14213, n14212, n14211, n14210, n14209, n14208, n14207,
         n14206, n14205, n14204, n14203, n14202, n14201, n14200, n14199,
         n14198, n14197, n14196, n14195, n14194, n14193, n14192, n14191,
         n14190, n14189, n14188, n14187, n14186, n14185, n14184, n14183,
         n14182, n14181, n14180, n14179, n14178, n14177, n14176, n14175,
         n14174, n14173, n14172, n14171, n14170, n14169, n14168, n14167,
         n14166, n14165, n14164, n14163, n14162, n14161, n14160, n14159,
         n14158, n14157, n14156, n14155, n14154, n14153, n14152, n14151,
         n14150, n14149, n14148, n14147, n14146, n14145, n14144, n14143,
         n14142, n14141, n14140, n14139, n14138, n14137, n14136, n14135,
         n14134, n14133, n14132, n14131, n14130, n14129, n14128, n14127,
         n14126, n14125, n14124, n14123, n14122, n14121, n14120, n14119,
         n14118, n14117, n14116, n14115, n14114, n14113, n14112, n14111,
         n14110, n14109, n14108, n14107, n14106, n14105, n14104, n14103,
         n14102, n14101, n14100, n14099, n14098, n14097, n14096, n14095,
         n14094, n14093, n14092, n14091, n14090, n14089, n14088, n14087,
         n14086, n14085, n14084, n14083, n14082, n14081, n14080, n14079,
         n14078, n14077, n14076, n14075, n14074, n14073, n14072, n14071,
         n14070, n14069, n14068, n14067, n14066, n14065, n14064, n14063,
         n14062, n14061, n14060, n14059, n14058, n14057, n14056, n14055,
         n14054, n14053, n14052, n14051, n14050, n14049, n14048, n14047,
         n14046, n14045, n14044, n14043, n14042, n14041, n14040, n14039,
         n14038, n14037, n14036, n14035, n14034, n14033, n14032, n14031,
         n14030, n14029, n14028, n14027, n14026, n14025, n14024, n14023,
         n14022, n14021, n14020, n14019, n14018, n14017, n14016, n14015,
         n14014, n14013, n14012, n14011, n14010, n14009, n14008, n14007,
         n14006, n14005, n14004, n14003, n14002, n14001, n14000, n13999,
         n13998, n13997, n13996, n13995, n13994, n13993, n13992, n13991,
         n13990, n13989, n13988, n13987, n13986, n13985, n13984, n13983,
         n13982, n13981, n13980, n13979, n13978, n13977, n13976, n13975,
         n13974, n13973, n13972, n13971, n13970, n13969, n13968, n13967,
         n13966, n13965, n13964, n13963, n13962, n13961, n13960, n13959,
         n13958, n13957, n13956, n13955, n13954, n13953, n13952, n13951,
         n13950, n13949, n13948, n13947, n13946, n13945, n13944, n13943,
         n13942, n13941, n13940, n13939, n13938, n13937, n13936, n13935,
         n13934, n13933, n13932, n13931, n13930, n13929, n13928, n13927,
         n13926, n13925, n13924, n13923, n13922, n13921, n13920, n13919,
         n13918, n13917, n13916, n13915, n13914, n13913, n13912, n13911,
         n13910, n13909, n13908, n13907, n13906, n13905, n13904, n13903,
         n13902, n13901, n13900, n13899, n13898, n13897, n13896, n13895,
         n13894, n13893, n13892, n13891, n13890, n13889, n13888, n13887,
         n13886, n13885, n13884, n13883, n13882, n13881, n13880, n13879,
         n13878, n13877, n13876, n13875, n13874, n13873, n13872, n13871,
         n13870, n13869, n13868, n13867, n13866, n13865, n13864, n13863,
         n13862, n13861, n13860, n13859, n13858, n13857, n13856, n13855,
         n13854, n13853, n13852, n13851, n13850, n13849, n13848, n13847,
         n13846, n13845, n13844, n13843, n13842, n13841, n13840, n13839,
         n13838, n13837, n13836, n13835, n13834, n13833, n13832, n13831,
         n13830, n13829, n13828, n13827, n13826, n13825, n13824, n13823,
         n13822, n13821, n13819, n13818, n13816, n13815, n13814, n13813,
         n13812, n13811, n13810, n13809, n13808, n13807, n13806, n13805,
         n13804, n13803, n13802, n13801, n13800, n13799, n13798, n13797,
         n13796, n13795, n13794, n13793, n13792, n13791, n13790, n13789,
         n13788, n13787, n13786, n13785, n13784, n13782, n13781, n13780,
         n13779, n13778, n13777, n13776, n13775, n13774, n13773, n13772,
         n13771, n13770, n13769, n13768, n13767, n13766, n13765, n13764,
         n13763, n13762, n13761, n13760, n13759, n13758, n13757, n13756,
         n13755, n13754, n13753, n13752, n13751, n13750, n13749, n13748,
         n13747, n13746, n13745, n13744, n13743, n13742, n13741, n13740,
         n13739, n13738, n13737, n13736, n13735, n13734, n13733, n13732,
         n13731, n13730, n13729, n13728, n13727, n13726, n13725, n13724,
         n13723, n13722, n13721, n13720, n13719, n13718, n13717, n13716,
         n13715, n13714, n13713, n13712, n13711, n13710, n13709, n13708,
         n13707, n13706, n13705, n13704, n13703, n13701, n13700, n13699,
         n13698, n13697, n13696, n13695, n13694, n13693, n13692, n13691,
         n13690, n13689, n13688, n13687, n13686, n13685, n13684, n13683,
         n13682, n13681, n13680, n13679, n13678, n13677, n13676, n13675,
         n13674, n13673, n13672, n13671, n13670, n13669, n13668, n13667,
         n13666, n13665, n13664, n13663, n13662, n13661, n13660, n13659,
         n13658, n13657, n13656, n13655, n13654, n13653, n13652, n13651,
         n13650, n13649, n13648, n13647, n13646, n13645, n13644, n13643,
         n13642, n13641, n13640, n13639, n13638, n13637, n13636, n13635,
         n13634, n13633, n13632, n13631, n13630, n13629, n13628, n13627,
         n13626, n13625, n13624, n13623, n13622, n13621, n13620, n13619,
         n13618, n13617, n13616, n13614, n13613, n13612, n13611, n13610,
         n13609, n13608, n13607, n13606, n13605, n13604, n13603, n13602,
         n13601, n13600, n13599, n13598, n13597, n13596, n13595, n13594,
         n13593, n13592, n13591, n13590, n13589, n13588, n13587, n13586,
         n13585, n13584, n13583, n13582, n13581, n13580, n13579, n13578,
         n13577, n13576, n13575, n13574, n13573, n13572, n13571, n13570,
         n13569, n13568, n13567, n13566, n13565, n13564, n13563, n13562,
         n13561, n13560, n13559, n13558, n13557, n13556, n13555, n13554,
         n13553, n13552, n13551, n13550, n13549, n13548, n13547, n13546,
         n13545, n13544, n13543, n13542, n13541, n13540, n13539, n13538,
         n13537, n13536, n13535, n13534, n13533, n13532, n13531, n13530,
         n13529, n13528, n13527, n13526, n13525, n13524, n13523, n13522,
         n13521, n13520, n13519, n13518, n13517, n13516, n13515, n13514,
         n13513, n13512, n13511, n13510, n13509, n13508, n13507, n13506,
         n13505, n13504, n13503, n13502, n13501, n13500, n13499, n13498,
         n13497, n13496, n13495, n13494, n13493, n13492, n13491, n13489,
         n13488, n13487, n13486, n13485, n13484, n13483, n13482, n13481,
         n13480, n13479, n13478, n13477, n13476, n13475, n13474, n13473,
         n13472, n13471, n13470, n13469, n13468, n13467, n13466, n13465,
         n13464, n13463, n13462, n13461, n13460, n13459, n13458, n13457,
         n13456, n13455, n13454, n13453, n13452, n13451, n13450, n13449,
         n13448, n13447, n13446, n13445, n13444, n13443, n13442, n13441,
         n13440, n13439, n13438, n13437, n13436, n13435, n13434, n13433,
         n13432, n13431, n13430, n13429, n13428, n13427, n13426, n13425,
         n13424, n13423, n13422, n13421, n13420, n13419, n13418, n13417,
         n13416, n13415, n13414, n13413, n13412, n13411, n13410, n13409,
         n13408, n13407, n13406, n13405, n13404, n13403, n13402, n13401,
         n13400, n13399, n13398, n13397, n13396, n13395, n13394, n13393,
         n13392, n13391, n13390, n13389, n13388, n13387, n13386, n13385,
         n13384, n13383, n13382, n13381, n13380, n13379, n13378, n13377,
         n13376, n13375, n13374, n13373, n13372, n13371, n13370, n13369,
         n13368, n13367, n13366, n13365, n13364, n13363, n13362, n13360,
         n13359, n13358, n13357, n13356, n13355, n13354, n13353, n13352,
         n13351, n13350, n13349, n13348, n13347, n13346, n13345, n13344,
         n13343, n13342, n13341, n13340, n13339, n13338, n13337, n13336,
         n13335, n13334, n13333, n13332, n13331, n13330, n13329, n13328,
         n13327, n13326, n13325, n13324, n13323, n13322, n13321, n13320,
         n13319, n13318, n13317, n13316, n13315, n13314, n13313, n13312,
         n13311, n13310, n13309, n13308, n13307, n13306, n13305, n13304,
         n13303, n13302, n13301, n13300, n13299, n13298, n13297, n13296,
         n13295, n13294, n13292, n13291, n13290, n13289, n13288, n13287,
         n13286, n13285, n13284, n13283, n13282, n13281, n13280, n13279,
         n13278, n13277, n13276, n13275, n13274, n13273, n13272, n13271,
         n13270, n13269, n13268, n13267, n13266, n13265, n13264, n13263,
         n13262, n13261, n13260, n13259, n13258, n13257, n13256, n13255,
         n13254, n13253, n13252, n13251, n13250, n13249, n13248, n13247,
         n13246, n13245, n13244, n13243, n13242, n13241, n13240, n13239,
         n13238, n13237, n13236, n13235, n13234, n13233, n13232, n13231,
         n13230, n13229, n13228, n13226, n13225, n13224, n13223, n13222,
         n13221, n13220, n13219, n13218, n13217, n13216, n13215, n13214,
         n13213, n13212, n13211, n13210, n13209, n13208, n13207, n13206,
         n13205, n13204, n13203, n13202, n13201, n13200, n13199, n13198,
         n13197, n13196, n13195, n13194, n13193, n13192, n13191, n13190,
         n13189, n13188, n13187, n13186, n13185, n13184, n13183, n13182,
         n13181, n13180, n13179, n13178, n13177, n13176, n13175, n13174,
         n13173, n13172, n13171, n13170, n13169, n13168, n13167, n13166,
         n13165, n13164, n13163, n13162, n13161, n13160, n13159, n13158,
         n13157, n13156, n13155, n13154, n13153, n13152, n13151, n13150,
         n13149, n13148, n13147, n13146, n13145, n13144, n13143, n13142,
         n13141, n13140, n13139, n13138, n13137, n13136, n13135, n13134,
         n13133, n13132, n13131, n13130, n13129, n13127, n13126, n13125,
         n13124, n13123, n13122, n13121, n13120, n13119, n13118, n13117,
         n13116, n13115, n13114, n13113, n13112, n13111, n13110, n13109,
         n13108, n13106, n13105, n13104, n13103, n13101, n13100, n13099,
         n13098, n13097, n13096, n13095, n13094, n13093, n13092, n13091,
         n13090, n13089, n13088, n13087, n13086, n13085, n13084, n13083,
         n13082, n13081, n13080, n13079, n13078, n13077, n13076, n13075,
         n13074, n13073, n13072, n13071, n13070, n13069, n13068, n13067,
         n13066, n13065, n13064, n13063, n13062, n13061, n13060, n13059,
         n13058, n13057, n13056, n13055, n13054, n13053, n13052, n13051,
         n13050, n13049, n13048, n13047, n13046, n13045, n13044, n13043,
         n13042, n13041, n13040, n13039, n13038, n13037, n13036, n13035,
         n13034, n13033, n13032, n13031, n13030, n13029, n13028, n13027,
         n13026, n13025, n13024, n13023, n13022, n13021, n13020, n13019,
         n13018, n13017, n13016, n13015, n13014, n13013, n13012, n13011,
         n13010, n13009, n13008, n13007, n13006, n13005, n13004, n13003,
         n13002, n13001, n13000, n12999, n12998, n12997, n12996, n12995,
         n12994, n12993, n12992, n12991, n12990, n12989, n12988, n12987,
         n12986, n12985, n12984, n12983, n12982, n12981, n12980, n12979,
         n12978, n12977, n12976, n12975, n12974, n12972, n12970, n12969,
         n12968, n12967, n12966, n12965, n12964, n12963, n12962, n12961,
         n12960, n12959, n12958, n12956, n12955, n12954, n12953, n12952,
         n12950, n12949, n12948, n12947, n12946, n12944, n12943, n12942,
         n12941, n12940, n12938, n12937, n12936, n12935, n12934, n12932,
         n12931, n12930, n12929, n12928, n12926, n12925, n12924, n12923,
         n12922, n12920, n12919, n12918, n12917, n12916, n12914, n12913,
         n12912, n12911, n12910, n12908, n12907, n12906, n12905, n12904,
         n12902, n12901, n12900, n12899, n12898, n12896, n12895, n12894,
         n12893, n12892, n12890, n12889, n12888, n12887, n12886, n12884,
         n12883, n12882, n12881, n12880, n12878, n12877, n12876, n12875,
         n12874, n12872, n12871, n12870, n12869, n12868, n12866, n12865,
         n12864, n12863, n12862, n12861, n12860, n12859, n12858, n12857,
         n12856, n12854, n12853, n12852, n12851, n12850, n12848, n12847,
         n12846, n12845, n12844, n12842, n12841, n12840, n12839, n12838,
         n12837, n12836, n12835, n12834, n12832, n12831, n12830, n12829,
         n12828, n12826, n12825, n12824, n12823, n12822, n12820, n12819,
         n12818, n12817, n12816, n12814, n12813, n12812, n12811, n12810,
         n12808, n12807, n12806, n12805, n12804, n12802, n12801, n12800,
         n12799, n12798, n12797, n12796, n12795, n12794, n12793, n12792,
         n12790, n12789, n12788, n12787, n12786, n12785, n12784, n12783,
         n12782, n12781, n12780, n12778, n12777, n12776, n12775, n12774,
         n12772, n12771, n12770, n12769, n12768, n12766, n12765, n12764,
         n12763, n12762, n12760, n12759, n12758, n12757, n12756, n12755,
         n12754, n12753, n12752, n12751, n12750, n12748, n12747, n12746,
         n12745, n12744, n12742, n12741, n12740, n12739, n12738, n12737,
         n12736, n12735, n12734, n12733, n12732, n12731, n12730, n12729,
         n12728, n12727, n12726, n12724, n12723, n12722, n12721, n12720,
         n12719, n12718, n12717, n12716, n12715, n12714, n12713, n12710,
         n12709, n12708, n12707, n12706, n12705, n12704, n12703, n12702,
         n12701, n12700, n12699, n12698, n12697, n12696, n12695, n12694,
         n12693, n12692, n12691, n12690, n12689, n12688, n12687, n12686,
         n12685, n12684, n12683, n12682, n12681, n12680, n12679, n12678,
         n12677, n12676, n12675, n12674, n12673, n12672, n12671, n12670,
         n12669, n12668, n12667, n12666, n12665, n12664, n12663, n12662,
         n12661, n12660, n12659, n12658, n12657, n12656, n12655, n12654,
         n12653, n12652, n12651, n12650, n12649, n12648, n12647, n12646,
         n12645, n12644, n12643, n12642, n12641, n12640, n12639, n12638,
         n12637, n12636, n12635, n12634, n12633, n12632, n12631, n12630,
         n12629, n12628, n12627, n12626, n12625, n12624, n12623, n12622,
         n12621, n12620, n12619, n12617, n12616, n12615, n12614, n12613,
         n12612, n12611, n12610, n12609, n12608, n12607, n12606, n12605,
         n12604, n12603, n12602, n12601, n12600, n12599, n12598, n12597,
         n12596, n12595, n12594, n12593, n12592, n12591, n12590, n12589,
         n12588, n12587, n12586, n12585, n12584, n12583, n12582, n12581,
         n12580, n12579, n12578, n12577, n12576, n12575, n12574, n12573,
         n12572, n12571, n12570, n12569, n12568, n12567, n12566, n12565,
         n12564, n12563, n12562, n12561, n12560, n12559, n12558, n12557,
         n12556, n12555, n12554, n12553, n12552, n12551, n12550, n12549,
         n12548, n12547, n12546, n12545, n12544, n12543, n12542, n12541,
         n12540, n12539, n12538, n12537, n12536, n12535, n12534, n12533,
         n12532, n12531, n12530, n12529, n12528, n12526, n12525, n12524,
         n12523, n12522, n12521, n12520, n12519, n12518, n12517, n12516,
         n12515, n12514, n12513, n12512, n12511, n12510, n12509, n12508,
         n12507, n12506, n12505, n12504, n12503, n12502, n12501, n12500,
         n12499, n12498, n12497, n12496, n12495, n12494, n12493, n12492,
         n12491, n12490, n12489, n12488, n12487, n12486, n12485, n12484,
         n12483, n12482, n12481, n12480, n12479, n12478, n12477, n12476,
         n12475, n12474, n12473, n12472, n12471, n12470, n12469, n12468,
         n12467, n12466, n12465, n12464, n12463, n12462, n12461, n12460,
         n12459, n12458, n12457, n12456, n12455, n12454, n12453, n12452,
         n12451, n12450, n12449, n12448, n12447, n12446, n12445, n12444,
         n12443, n12442, n12440, n12439, n12438, n12436, n12435, n12434,
         n12433, n12432, n12431, n12430, n12429, n12428, n12427, n12426,
         n12425, n12424, n12423, n12422, n12421, n12420, n12419, n12418,
         n12417, n12416, n12415, n12414, n12413, n12412, n12411, n12410,
         n12409, n12408, n12407, n12406, n12405, n12404, n12403, n12402,
         n12401, n12400, n12399, n12398, n12397, n12396, n12395, n12394,
         n12393, n12392, n12391, n12390, n12389, n12388, n12387, n12386,
         n12385, n12384, n12383, n12382, n12381, n12380, n12379, n12378,
         n12377, n12376, n12375, n12374, n12373, n12372, n12371, n12370,
         n12369, n12368, n12367, n12366, n12365, n12364, n12363, n12362,
         n12361, n12360, n12359, n12358, n12357, n12356, n12355, n12354,
         n12353, n12352, n12351, n12348, n12347, n12346, n12345, n12344,
         n12343, n12342, n12341, n12340, n12339, n12338, n12337, n12336,
         n12335, n12334, n12333, n12332, n12331, n12330, n12329, n12328,
         n12327, n12326, n12325, n12324, n12323, n12322, n12321, n12320,
         n12319, n12318, n12317, n12316, n12315, n12314, n12313, n12312,
         n12311, n12310, n12309, n12308, n12307, n12306, n12305, n12304,
         n12303, n12302, n12301, n12300, n12299, n12298, n12297, n12296,
         n12295, n12294, n12293, n12292, n12291, n12290, n12289, n12288,
         n12287, n12286, n12285, n12284, n12283, n12282, n12281, n12280,
         n12279, n12278, n12277, n12276, n12275, n12274, n12273, n12272,
         n12271, n12270, n12269, n12268, n12267, n12266, n12265, n12264,
         n12263, n12262, n12261, n12260, n12259, n12258, n12257, n12256,
         n12255, n12254, n12253, n12252, n12251, n12250, n12249, n12248,
         n12247, n12246, n12245, n12244, n12243, n12242, n12241, n12240,
         n12239, n12238, n12237, n12236, n12235, n12234, n12233, n12232,
         n12231, n12230, n12229, n12228, n12227, n12226, n12225, n12224,
         n12223, n12222, n12221, n12220, n12219, n12218, n12217, n12216,
         n12215, n12214, n12213, n12212, n12211, n12210, n12209, n12208,
         n12207, n12206, n12205, n12204, n12203, n12202, n12201, n12200,
         n12199, n12198, n12197, n12196, n12195, n12194, n12193, n12192,
         n12191, n12190, n12189, n12188, n12187, n12186, n12185, n12184,
         n12183, n12182, n12181, n12180, n12179, n12178, n12177, n12176,
         n12175, n12174, n12173, n12172, n12171, n12170, n12169, n12168,
         n12167, n12166, n12165, n12164, n12163, n12162, n12161, n12160,
         n12159, n12158, n12157, n12156, n12155, n12154, n12153, n12152,
         n12151, n12150, n12149, n12148, n12147, n12146, n12145, n12144,
         n12143, n12142, n12141, n12140, n12139, n12138, n12137, n12136,
         n12135, n12134, n12133, n12132, n12131, n12130, n12129, n12128,
         n12127, n12126, n12125, n12122, n12121, n12120, n12119, n12117,
         n12116, n12115, n12114, n12113, n12112, n12111, n12110, n12109,
         n12108, n12107, n12106, n12105, n12104, n12103, n12102, n12101,
         n12100, n12099, n12098, n12097, n12096, n12095, n12094, n12093,
         n12092, n12091, n12090, n12089, n12088, n12087, n12086, n12085,
         n12084, n12083, n12082, n12081, n12080, n12079, n12078, n12077,
         n12076, n12075, n12074, n12073, n12072, n12071, n12070, n12069,
         n12068, n12067, n12066, n12065, n12064, n12063, n12062, n12061,
         n12060, n12059, n12058, n12057, n12056, n12055, n12054, n12053,
         n12052, n12051, n12050, n12049, n12048, n12047, n12046, n12045,
         n12044, n12043, n12042, n12041, n12040, n12039, n12038, n12037,
         n12036, n12035, n12034, n12033, n12032, n12031, n12030, n12029,
         n12028, n12027, n12026, n12025, n12024, n12023, n12022, n12021,
         n12020, n12019, n12018, n12017, n12016, n12015, n12014, n12013,
         n12012, n12011, n12010, n12009, n12008, n12007, n12006, n12005,
         n12004, n12003, n12002, n12001, n12000, n11999, n11998, n11997,
         n11996, n11995, n11994, n11993, n11992, n11991, n11990, n11989,
         n11988, n11987, n11986, n11985, n11984, n11983, n11982, n11981,
         n11980, n11979, n11978, n11977, n11976, n11975, n11974, n11973,
         n11972, n11971, n11970, n11969, n11968, n11967, n11966, n11965,
         n11964, n11963, n11962, n11961, n11960, n11959, n11958, n11957,
         n11956, n11955, n11954, n11953, n11952, n11951, n11950, n11949,
         n11948, n11947, n11946, n11945, n11944, n11943, n11942, n11941,
         n11940, n11939, n11938, n11937, n11936, n11935, n11934, n11933,
         n11932, n11931, n11930, n11929, n11928, n11927, n11926, n11925,
         n11924, n11923, n11922, n11921, n11920, n11919, n11918, n11917,
         n11916, n11915, n11914, n11913, n11912, n11911, n11910, n11909,
         n11908, n11907, n11906, n11905, n11904, n11903, n11902, n11901,
         n11900, n11899, n11898, n11897, n11895, n11894, n11893, n11892,
         n11891, n11890, n11889, n11888, n11887, n11886, n11885, n11884,
         n11883, n11882, n11881, n11880, n11879, n11878, n11877, n11876,
         n11875, n11874, n11873, n11872, n11871, n11870, n11869, n11868,
         n11867, n11866, n11865, n11864, n11863, n11862, n11861, n11860,
         n11859, n11858, n11857, n11856, n11855, n11854, n11853, n11852,
         n11851, n11850, n11848, n11847, n11846, n11845, n11843, n11842,
         n11841, n11840, n11839, n11838, n11837, n11836, n11835, n11834,
         n11833, n11832, n11831, n11830, n11829, n11828, n11827, n11826,
         n11825, n11824, n11823, n11822, n11821, n11820, n11819, n11818,
         n11817, n11816, n11815, n11814, n11813, n11812, n11811, n11810,
         n11809, n11808, n11807, n11806, n11805, n11804, n11803, n11802,
         n11800, n11799, n11798, n11797, n11796, n11795, n11794, n11793,
         n11792, n11791, n11790, n11789, n11788, n11787, n11786, n11785,
         n11784, n11783, n11782, n11781, n11780, n11779, n11778, n11777,
         n11776, n11775, n11774, n11773, n11772, n11771, n11770, n11768,
         n11767, n11766, n11765, n11764, n11762, n11761, n11760, n11759,
         n11758, n11757, n11756, n11755, n11754, n11753, n11752, n11751,
         n11750, n11749, n11748, n11747, n11746, n11745, n11744, n11743,
         n11742, n11741, n11740, n11739, n11738, n11737, n11736, n11735,
         n11734, n11733, n11732, n11731, n11730, n11729, n11728, n11727,
         n11726, n11725, n11724, n11723, n11722, n11721, n11720, n11719,
         n11718, n11717, n11716, n11715, n11714, n11713, n11712, n11711,
         n11710, n11709, n11708, n11707, n11706, n11705, n11704, n11703,
         n11702, n11701, n11700, n11699, n11698, n11697, n11696, n11695,
         n11694, n11693, n11692, n11691, n11690, n11689, n11688, n11687,
         n11686, n11685, n11684, n11683, n11682, n11681, n11680, n11679,
         n11678, n11677, n11676, n11675, n11674, n11673, n11672, n11671,
         n11670, n11669, n11668, n11667, n11665, n11664, n11663, n11662,
         n11661, n11660, n11659, n11658, n11657, n11656, n11655, n11654,
         n11653, n11652, n11651, n11650, n11649, n11648, n11647, n11646,
         n11645, n11644, n11643, n11642, n11641, n11640, n11639, n11638,
         n11637, n11636, n11635, n11634, n11633, n11632, n11631, n11630,
         n11629, n11628, n11627, n11626, n11625, n11624, n11623, n11622,
         n11621, n11620, n11619, n11618, n11617, n11616, n11615, n11614,
         n11612, n11611, n11610, n11609, n11608, n11607, n11606, n11605,
         n11604, n11603, n11602, n11601, n11600, n11599, n11598, n11597,
         n11596, n11595, n11594, n11593, n11592, n11591, n11590, n11589,
         n11588, n11587, n11586, n11585, n11584, n11583, n11582, n11581,
         n11580, n11579, n11578, n11577, n11576, n11575, n11574, n11573,
         n11572, n11571, n11570, n11569, n11568, n11567, n11566, n11565,
         n11564, n11563, n11562, n11561, n11560, n11559, n11558, n11557,
         n11556, n11555, n11554, n11553, n11552, n11551, n11550, n11549,
         n11548, n11547, n11546, n11545, n11544, n11543, n11542, n11541,
         n11540, n11539, n11538, n11537, n11536, n11535, \filter_0/n7589 ,
         \filter_0/n7588 , \filter_0/n7585 , \filter_0/n7584 ,
         \filter_0/n7581 , \filter_0/n7580 , \filter_0/n7577 ,
         \filter_0/n7576 , \filter_0/n7573 , \filter_0/n7572 ,
         \filter_0/n7569 , \filter_0/n7568 , \filter_0/n7565 ,
         \filter_0/n7564 , \filter_0/n7561 , \filter_0/n7560 ,
         \filter_0/n7557 , \filter_0/n7556 , \filter_0/n7553 ,
         \filter_0/n7552 , \filter_0/n7549 , \filter_0/n7548 ,
         \filter_0/n7545 , \filter_0/n7544 , \filter_0/n7541 ,
         \filter_0/n7540 , \filter_0/n7537 , \filter_0/n7536 ,
         \filter_0/n7533 , \filter_0/n7532 , \filter_0/n7529 ,
         \filter_0/n7528 , \filter_0/n7525 , \filter_0/n7524 ,
         \filter_0/n7521 , \filter_0/n7520 , \filter_0/n7517 ,
         \filter_0/n7516 , \filter_0/n7513 , \filter_0/n7512 ,
         \filter_0/n7509 , \filter_0/n7508 , \filter_0/n7505 ,
         \filter_0/n7504 , \filter_0/n7501 , \filter_0/n7500 ,
         \filter_0/n7497 , \filter_0/n7496 , \filter_0/n7493 ,
         \filter_0/n7492 , \filter_0/n7489 , \filter_0/n7488 ,
         \filter_0/n7485 , \filter_0/n7484 , \filter_0/n7481 ,
         \filter_0/n7480 , \filter_0/n7477 , \filter_0/n7476 ,
         \filter_0/n7473 , \filter_0/n7472 , \filter_0/n7469 ,
         \filter_0/n7468 , \filter_0/n7465 , \filter_0/n7464 ,
         \filter_0/n7461 , \filter_0/n7460 , \filter_0/n7457 ,
         \filter_0/n7456 , \filter_0/n7453 , \filter_0/n7452 ,
         \filter_0/n7449 , \filter_0/n7448 , \filter_0/n7445 ,
         \filter_0/n7444 , \filter_0/n7441 , \filter_0/n7440 ,
         \filter_0/n7437 , \filter_0/n7436 , \filter_0/n7433 ,
         \filter_0/n7432 , \filter_0/n7429 , \filter_0/n7428 ,
         \filter_0/n7425 , \filter_0/n7424 , \filter_0/n7421 ,
         \filter_0/n7420 , \filter_0/n7417 , \filter_0/n7416 ,
         \filter_0/n7413 , \filter_0/n7412 , \filter_0/n7409 ,
         \filter_0/n7408 , \filter_0/n7405 , \filter_0/n7404 ,
         \filter_0/n7401 , \filter_0/n7400 , \filter_0/n7397 ,
         \filter_0/n7396 , \filter_0/n7393 , \filter_0/n7392 ,
         \filter_0/n7389 , \filter_0/n7388 , \filter_0/n7385 ,
         \filter_0/n7384 , \filter_0/n7381 , \filter_0/n7380 ,
         \filter_0/n7377 , \filter_0/n7376 , \filter_0/n7373 ,
         \filter_0/n7372 , \filter_0/n7369 , \filter_0/n7368 ,
         \filter_0/n7365 , \filter_0/n7364 , \filter_0/n7361 ,
         \filter_0/n7360 , \filter_0/n7357 , \filter_0/n7356 ,
         \filter_0/n7353 , \filter_0/n7352 , \filter_0/n7349 ,
         \filter_0/n7348 , \filter_0/n7345 , \filter_0/n7344 ,
         \filter_0/n7341 , \filter_0/n7340 , \filter_0/n7337 ,
         \filter_0/n7336 , \filter_0/n7333 , \filter_0/n7332 ,
         \filter_0/n7329 , \filter_0/n7328 , \filter_0/n7325 ,
         \filter_0/n7324 , \filter_0/n7321 , \filter_0/n7320 ,
         \filter_0/n7317 , \filter_0/n7316 , \filter_0/n7313 ,
         \filter_0/n7312 , \filter_0/n7309 , \filter_0/n7308 ,
         \filter_0/n7305 , \filter_0/n7304 , \filter_0/n7301 ,
         \filter_0/n7300 , \filter_0/n7297 , \filter_0/n7296 ,
         \filter_0/n7293 , \filter_0/n7292 , \filter_0/n7289 ,
         \filter_0/n7288 , \filter_0/n7285 , \filter_0/n7284 ,
         \filter_0/n7281 , \filter_0/n7280 , \filter_0/n7277 ,
         \filter_0/n7276 , \filter_0/n7273 , \filter_0/n7272 ,
         \filter_0/n7269 , \filter_0/n7268 , \filter_0/n7265 ,
         \filter_0/n7264 , \filter_0/n7261 , \filter_0/n7260 ,
         \filter_0/n7257 , \filter_0/n7256 , \filter_0/n7253 ,
         \filter_0/n7252 , \filter_0/n7249 , \filter_0/n7248 ,
         \filter_0/n7245 , \filter_0/n7244 , \filter_0/n7241 ,
         \filter_0/n7240 , \filter_0/n7237 , \filter_0/n7236 ,
         \filter_0/n7233 , \filter_0/n7232 , \filter_0/n7229 ,
         \filter_0/n7228 , \filter_0/n7225 , \filter_0/n7224 ,
         \filter_0/n7221 , \filter_0/n7220 , \filter_0/n7217 ,
         \filter_0/n7216 , \filter_0/n7213 , \filter_0/n7212 ,
         \filter_0/n7209 , \filter_0/n7208 , \filter_0/n7205 ,
         \filter_0/n7204 , \filter_0/n7201 , \filter_0/n7200 ,
         \filter_0/n7197 , \filter_0/n7196 , \filter_0/n7193 ,
         \filter_0/n7192 , \filter_0/n7189 , \filter_0/n7188 ,
         \filter_0/n7185 , \filter_0/n7184 , \filter_0/n7181 ,
         \filter_0/n7180 , \filter_0/n7177 , \filter_0/n7176 ,
         \filter_0/n7173 , \filter_0/n7172 , \filter_0/n7169 ,
         \filter_0/n7168 , \filter_0/n7165 , \filter_0/n7164 ,
         \filter_0/n7161 , \filter_0/n7160 , \filter_0/n7157 ,
         \filter_0/n7156 , \filter_0/n7153 , \filter_0/n7152 ,
         \filter_0/n7149 , \filter_0/n7148 , \filter_0/n7145 ,
         \filter_0/n7144 , \filter_0/n7141 , \filter_0/n7140 ,
         \filter_0/n7137 , \filter_0/n7136 , \filter_0/n7133 ,
         \filter_0/n7132 , \filter_0/n7129 , \filter_0/n7128 ,
         \filter_0/n7125 , \filter_0/n7124 , \filter_0/n7121 ,
         \filter_0/n7120 , \filter_0/n7117 , \filter_0/n7116 ,
         \filter_0/n7113 , \filter_0/n7112 , \filter_0/n7109 ,
         \filter_0/n7108 , \filter_0/n7105 , \filter_0/n7104 ,
         \filter_0/n7101 , \filter_0/n7100 , \filter_0/n7097 ,
         \filter_0/n7096 , \filter_0/n7093 , \filter_0/n7092 ,
         \filter_0/n7089 , \filter_0/n7088 , \filter_0/n7085 ,
         \filter_0/n7084 , \filter_0/n7081 , \filter_0/n7080 ,
         \filter_0/n7077 , \filter_0/n7076 , \filter_0/n7073 ,
         \filter_0/n7072 , \filter_0/n7069 , \filter_0/n7068 ,
         \filter_0/n7065 , \filter_0/n7064 , \filter_0/n7061 ,
         \filter_0/n7060 , \filter_0/n7057 , \filter_0/n7056 ,
         \filter_0/n7053 , \filter_0/n7052 , \filter_0/n7049 ,
         \filter_0/n7048 , \filter_0/n7045 , \filter_0/n7044 ,
         \filter_0/n7041 , \filter_0/n7040 , \filter_0/n7037 ,
         \filter_0/n7036 , \filter_0/n7033 , \filter_0/n7032 ,
         \filter_0/n7029 , \filter_0/n7028 , \filter_0/n7025 ,
         \filter_0/n7024 , \filter_0/n7021 , \filter_0/n7020 ,
         \filter_0/n7017 , \filter_0/n7016 , \filter_0/n7013 ,
         \filter_0/n7012 , \filter_0/n7009 , \filter_0/n7008 ,
         \filter_0/n7005 , \filter_0/n7004 , \filter_0/n7001 ,
         \filter_0/n7000 , \filter_0/n6997 , \filter_0/n6996 ,
         \filter_0/n6993 , \filter_0/n6992 , \filter_0/n6989 ,
         \filter_0/n6988 , \filter_0/n6985 , \filter_0/n6984 ,
         \filter_0/n6981 , \filter_0/n6980 , \filter_0/n6977 ,
         \filter_0/n6976 , \filter_0/n6973 , \filter_0/n6972 ,
         \filter_0/n6969 , \filter_0/n6968 , \filter_0/n6965 ,
         \filter_0/n6964 , \filter_0/n6961 , \filter_0/n6960 ,
         \filter_0/n6957 , \filter_0/n6956 , \filter_0/n6953 ,
         \filter_0/n6952 , \filter_0/n6949 , \filter_0/n6948 ,
         \filter_0/n6945 , \filter_0/n6944 , \filter_0/n6941 ,
         \filter_0/n6940 , \filter_0/n6937 , \filter_0/n6936 ,
         \filter_0/n6933 , \filter_0/n6932 , \filter_0/n6929 ,
         \filter_0/n6928 , \filter_0/n6925 , \filter_0/n6924 ,
         \filter_0/n6921 , \filter_0/n6920 , \filter_0/n6917 ,
         \filter_0/n6916 , \filter_0/n6913 , \filter_0/n6912 ,
         \filter_0/n6909 , \filter_0/n6908 , \filter_0/n6905 ,
         \filter_0/n6904 , \filter_0/n6901 , \filter_0/n6900 ,
         \filter_0/n6897 , \filter_0/n6896 , \filter_0/n6893 ,
         \filter_0/n6892 , \filter_0/n6889 , \filter_0/n6888 ,
         \filter_0/n6885 , \filter_0/n6884 , \filter_0/n6881 ,
         \filter_0/n6880 , \filter_0/n6877 , \filter_0/n6876 ,
         \filter_0/n6873 , \filter_0/n6872 , \filter_0/n6869 ,
         \filter_0/n6868 , \filter_0/n6865 , \filter_0/n6864 ,
         \filter_0/n6861 , \filter_0/n6860 , \filter_0/n6857 ,
         \filter_0/n6856 , \filter_0/n6853 , \filter_0/n6852 ,
         \filter_0/n6849 , \filter_0/n6848 , \filter_0/n6845 ,
         \filter_0/n6844 , \filter_0/n6841 , \filter_0/n6840 ,
         \filter_0/n6837 , \filter_0/n6836 , \filter_0/n6833 ,
         \filter_0/n6832 , \filter_0/n6829 , \filter_0/n6828 ,
         \filter_0/n6825 , \filter_0/n6824 , \filter_0/n6821 ,
         \filter_0/n6820 , \filter_0/n6817 , \filter_0/n6816 ,
         \filter_0/n6813 , \filter_0/n6812 , \filter_0/n6809 ,
         \filter_0/n6808 , \filter_0/n6805 , \filter_0/n6804 ,
         \filter_0/n6801 , \filter_0/n6800 , \filter_0/n6797 ,
         \filter_0/n6796 , \filter_0/n6793 , \filter_0/n6792 ,
         \filter_0/n6789 , \filter_0/n6788 , \filter_0/n6785 ,
         \filter_0/n6784 , \filter_0/n6781 , \filter_0/n6780 ,
         \filter_0/n6777 , \filter_0/n6776 , \filter_0/n6773 ,
         \filter_0/n6772 , \filter_0/n6769 , \filter_0/n6768 ,
         \filter_0/n6765 , \filter_0/n6764 , \filter_0/n6761 ,
         \filter_0/n6760 , \filter_0/n6757 , \filter_0/n6756 ,
         \filter_0/n6753 , \filter_0/n6752 , \filter_0/n6749 ,
         \filter_0/n6748 , \filter_0/n6745 , \filter_0/n6744 ,
         \filter_0/n6741 , \filter_0/n6740 , \filter_0/n6737 ,
         \filter_0/n6736 , \filter_0/n6733 , \filter_0/n6732 ,
         \filter_0/n6729 , \filter_0/n6728 , \filter_0/n6725 ,
         \filter_0/n6724 , \filter_0/n6721 , \filter_0/n6720 ,
         \filter_0/n6717 , \filter_0/n6716 , \filter_0/n6713 ,
         \filter_0/n6712 , \filter_0/n6709 , \filter_0/n6708 ,
         \filter_0/n6705 , \filter_0/n6704 , \filter_0/n6701 ,
         \filter_0/n6700 , \filter_0/n6697 , \filter_0/n6696 ,
         \filter_0/n6693 , \filter_0/n6692 , \filter_0/n6689 ,
         \filter_0/n6688 , \filter_0/n6685 , \filter_0/n6684 ,
         \filter_0/n6681 , \filter_0/n6680 , \filter_0/n6677 ,
         \filter_0/n6676 , \filter_0/n6673 , \filter_0/n6672 ,
         \filter_0/n6669 , \filter_0/n6668 , \filter_0/n6665 ,
         \filter_0/n6664 , \filter_0/n6661 , \filter_0/n6660 ,
         \filter_0/n6657 , \filter_0/n6656 , \filter_0/n6653 ,
         \filter_0/n6652 , \filter_0/n6649 , \filter_0/n6648 ,
         \filter_0/n6645 , \filter_0/n6644 , \filter_0/n6641 ,
         \filter_0/n6640 , \filter_0/n6637 , \filter_0/n6636 ,
         \filter_0/n6633 , \filter_0/n6632 , \filter_0/n6629 ,
         \filter_0/n6628 , \filter_0/n6625 , \filter_0/n6624 ,
         \filter_0/n6621 , \filter_0/n6620 , \filter_0/n6617 ,
         \filter_0/n6616 , \filter_0/n6613 , \filter_0/n6612 ,
         \filter_0/n6609 , \filter_0/n6608 , \filter_0/n6605 ,
         \filter_0/n6604 , \filter_0/n6601 , \filter_0/n6600 ,
         \filter_0/n6597 , \filter_0/n6596 , \filter_0/n6593 ,
         \filter_0/n6592 , \filter_0/n6589 , \filter_0/n6588 ,
         \filter_0/n6585 , \filter_0/n6584 , \filter_0/n6581 ,
         \filter_0/n6580 , \filter_0/n6577 , \filter_0/n6576 ,
         \filter_0/n6573 , \filter_0/n6572 , \filter_0/n6569 ,
         \filter_0/n6568 , \filter_0/n6565 , \filter_0/n6564 ,
         \filter_0/n6561 , \filter_0/n6560 , \filter_0/n6557 ,
         \filter_0/n6556 , \filter_0/n6553 , \filter_0/n6552 ,
         \filter_0/n6549 , \filter_0/n6548 , \filter_0/n6545 ,
         \filter_0/n6544 , \filter_0/n6541 , \filter_0/n6540 ,
         \filter_0/n6537 , \filter_0/n6536 , \filter_0/n6533 ,
         \filter_0/n6532 , \filter_0/n6529 , \filter_0/n6528 ,
         \filter_0/n6525 , \filter_0/n6524 , \filter_0/n6521 ,
         \filter_0/n6520 , \filter_0/n6517 , \filter_0/n6516 ,
         \filter_0/n6513 , \filter_0/n6512 , \filter_0/n6509 ,
         \filter_0/n6508 , \filter_0/n6505 , \filter_0/n6504 ,
         \filter_0/n6501 , \filter_0/n6500 , \filter_0/n6497 ,
         \filter_0/n6496 , \filter_0/n6493 , \filter_0/n6492 ,
         \filter_0/n6489 , \filter_0/n6488 , \filter_0/n6485 ,
         \filter_0/n6484 , \filter_0/n6481 , \filter_0/n6480 ,
         \filter_0/n6477 , \filter_0/n6476 , \filter_0/n6473 ,
         \filter_0/n6472 , \filter_0/n6469 , \filter_0/n6468 ,
         \filter_0/n6465 , \filter_0/n6464 , \filter_0/n6461 ,
         \filter_0/n6460 , \filter_0/n6457 , \filter_0/n6456 ,
         \filter_0/n6453 , \filter_0/n6452 , \filter_0/n6449 ,
         \filter_0/n6448 , \filter_0/n6445 , \filter_0/n6444 ,
         \filter_0/n6441 , \filter_0/n6440 , \filter_0/n6437 ,
         \filter_0/n6436 , \filter_0/n6433 , \filter_0/n6432 ,
         \filter_0/n6429 , \filter_0/n6428 , \filter_0/n6425 ,
         \filter_0/n6424 , \filter_0/n6421 , \filter_0/n6420 ,
         \filter_0/n6417 , \filter_0/n6416 , \filter_0/n6413 ,
         \filter_0/n6412 , \filter_0/n6409 , \filter_0/n6408 ,
         \filter_0/n6405 , \filter_0/n6404 , \filter_0/n6401 ,
         \filter_0/n6400 , \filter_0/n6397 , \filter_0/n6396 ,
         \filter_0/n6393 , \filter_0/n6392 , \filter_0/n6389 ,
         \filter_0/n6388 , \filter_0/n6385 , \filter_0/n6384 ,
         \filter_0/n6381 , \filter_0/n6380 , \filter_0/n6377 ,
         \filter_0/n6376 , \filter_0/n6373 , \filter_0/n6372 ,
         \filter_0/n6369 , \filter_0/n6368 , \filter_0/n6365 ,
         \filter_0/n6364 , \filter_0/n6361 , \filter_0/n6360 ,
         \filter_0/n6357 , \filter_0/n6356 , \filter_0/n6353 ,
         \filter_0/n6352 , \filter_0/n6349 , \filter_0/n6348 ,
         \filter_0/n6345 , \filter_0/n6344 , \filter_0/n6341 ,
         \filter_0/n6340 , \filter_0/n6337 , \filter_0/n6336 ,
         \filter_0/n6333 , \filter_0/n6332 , \filter_0/n6329 ,
         \filter_0/n6328 , \filter_0/n6325 , \filter_0/n6324 ,
         \filter_0/n6321 , \filter_0/n6320 , \filter_0/n6317 ,
         \filter_0/n6316 , \filter_0/n6313 , \filter_0/n6312 ,
         \filter_0/n6309 , \filter_0/n6308 , \filter_0/n6305 ,
         \filter_0/n6304 , \filter_0/n6301 , \filter_0/n6300 ,
         \filter_0/n6297 , \filter_0/n6296 , \filter_0/n6293 ,
         \filter_0/n6292 , \filter_0/n6289 , \filter_0/n6288 ,
         \filter_0/n6285 , \filter_0/n6284 , \filter_0/n6281 ,
         \filter_0/n6280 , \filter_0/n6277 , \filter_0/n6276 ,
         \filter_0/n6273 , \filter_0/n6272 , \filter_0/n6269 ,
         \filter_0/n6268 , \filter_0/n6265 , \filter_0/n6264 ,
         \filter_0/n6261 , \filter_0/n6260 , \filter_0/n6257 ,
         \filter_0/n6256 , \filter_0/n6253 , \filter_0/n6252 ,
         \filter_0/n6249 , \filter_0/n6248 , \filter_0/n6245 ,
         \filter_0/n6244 , \filter_0/n6241 , \filter_0/n6240 ,
         \filter_0/n6237 , \filter_0/n6236 , \filter_0/n6233 ,
         \filter_0/n6232 , \filter_0/n6229 , \filter_0/n6228 ,
         \filter_0/n6225 , \filter_0/n6224 , \filter_0/n6221 ,
         \filter_0/n6220 , \filter_0/n6217 , \filter_0/n6216 ,
         \filter_0/n6213 , \filter_0/n6212 , \filter_0/n6209 ,
         \filter_0/n6208 , \filter_0/n6205 , \filter_0/n6204 ,
         \filter_0/n6201 , \filter_0/n6200 , \filter_0/n6197 ,
         \filter_0/n6196 , \filter_0/n6193 , \filter_0/n6192 ,
         \filter_0/n6189 , \filter_0/n6188 , \filter_0/n6185 ,
         \filter_0/n6184 , \filter_0/n6181 , \filter_0/n6180 ,
         \filter_0/n6177 , \filter_0/n6176 , \filter_0/n6173 ,
         \filter_0/n6172 , \filter_0/n6169 , \filter_0/n6168 ,
         \filter_0/n6165 , \filter_0/n6164 , \filter_0/n6161 ,
         \filter_0/n6160 , \filter_0/n6157 , \filter_0/n6156 ,
         \filter_0/n6153 , \filter_0/n6152 , \filter_0/n6149 ,
         \filter_0/n6148 , \filter_0/n6145 , \filter_0/n6144 ,
         \filter_0/n6141 , \filter_0/n6140 , \filter_0/n6137 ,
         \filter_0/n6136 , \filter_0/n6133 , \filter_0/n6132 ,
         \filter_0/n6129 , \filter_0/n6128 , \filter_0/n6125 ,
         \filter_0/n6124 , \filter_0/n6121 , \filter_0/n6120 ,
         \filter_0/n6117 , \filter_0/n6116 , \filter_0/n6113 ,
         \filter_0/n6112 , \filter_0/n6109 , \filter_0/n6108 ,
         \filter_0/n6105 , \filter_0/n6104 , \filter_0/n6101 ,
         \filter_0/n6100 , \filter_0/n6097 , \filter_0/n6096 ,
         \filter_0/n6093 , \filter_0/n6092 , \filter_0/n6089 ,
         \filter_0/n6088 , \filter_0/n6085 , \filter_0/n6084 ,
         \filter_0/n6081 , \filter_0/n6080 , \filter_0/n6077 ,
         \filter_0/n6076 , \filter_0/n6073 , \filter_0/n6072 ,
         \filter_0/n6069 , \filter_0/n6068 , \filter_0/n6065 ,
         \filter_0/n6064 , \filter_0/n6061 , \filter_0/n6060 ,
         \filter_0/n6057 , \filter_0/n6056 , \filter_0/n6053 ,
         \filter_0/n6052 , \filter_0/n6049 , \filter_0/n6048 ,
         \filter_0/n6045 , \filter_0/n6044 , \filter_0/n6041 ,
         \filter_0/n6040 , \filter_0/n6037 , \filter_0/n6036 ,
         \filter_0/n6033 , \filter_0/n6032 , \filter_0/n6029 ,
         \filter_0/n6028 , \filter_0/n6025 , \filter_0/n6024 ,
         \filter_0/n6021 , \filter_0/n6020 , \filter_0/n6017 ,
         \filter_0/n6016 , \filter_0/n6013 , \filter_0/n6012 ,
         \filter_0/n6009 , \filter_0/n6008 , \filter_0/n6005 ,
         \filter_0/n6004 , \filter_0/n6001 , \filter_0/n6000 ,
         \filter_0/n5997 , \filter_0/n5996 , \filter_0/n5993 ,
         \filter_0/n5992 , \filter_0/n5989 , \filter_0/n5988 ,
         \filter_0/n5985 , \filter_0/n5984 , \filter_0/n5981 ,
         \filter_0/n5980 , \filter_0/n5977 , \filter_0/n5976 ,
         \filter_0/n5973 , \filter_0/n5972 , \filter_0/n5969 ,
         \filter_0/n5968 , \filter_0/n5965 , \filter_0/n5964 ,
         \filter_0/n5961 , \filter_0/n5960 , \filter_0/n5957 ,
         \filter_0/n5956 , \filter_0/n5953 , \filter_0/n5952 ,
         \filter_0/n5949 , \filter_0/n5948 , \filter_0/n5945 ,
         \filter_0/n5944 , \filter_0/n5941 , \filter_0/n5940 ,
         \filter_0/n5937 , \filter_0/n5936 , \filter_0/n5933 ,
         \filter_0/n5932 , \filter_0/n5929 , \filter_0/n5928 ,
         \filter_0/n5925 , \filter_0/n5924 , \filter_0/n5921 ,
         \filter_0/n5920 , \filter_0/n5917 , \filter_0/n5916 ,
         \filter_0/n5913 , \filter_0/n5912 , \filter_0/n5909 ,
         \filter_0/n5908 , \filter_0/n5905 , \filter_0/n5904 ,
         \filter_0/n5901 , \filter_0/n5900 , \filter_0/n5897 ,
         \filter_0/n5896 , \filter_0/n5893 , \filter_0/n5892 ,
         \filter_0/n5889 , \filter_0/n5888 , \filter_0/n5885 ,
         \filter_0/n5884 , \filter_0/n5881 , \filter_0/n5880 ,
         \filter_0/n5877 , \filter_0/n5876 , \filter_0/n5873 ,
         \filter_0/n5872 , \filter_0/n5869 , \filter_0/n5868 ,
         \filter_0/n5865 , \filter_0/n5864 , \filter_0/n5861 ,
         \filter_0/n5860 , \filter_0/n5857 , \filter_0/n5856 ,
         \filter_0/n5853 , \filter_0/n5852 , \filter_0/n5849 ,
         \filter_0/n5848 , \filter_0/n5845 , \filter_0/n5844 ,
         \filter_0/n5841 , \filter_0/n5840 , \filter_0/n5837 ,
         \filter_0/n5836 , \filter_0/n5833 , \filter_0/n5832 ,
         \filter_0/n5829 , \filter_0/n5828 , \filter_0/n5825 ,
         \filter_0/n5824 , \filter_0/n5821 , \filter_0/n5820 ,
         \filter_0/n5817 , \filter_0/n5816 , \filter_0/n5813 ,
         \filter_0/n5812 , \filter_0/n5809 , \filter_0/n5808 ,
         \filter_0/n5805 , \filter_0/n5804 , \filter_0/n5801 ,
         \filter_0/n5800 , \filter_0/n5797 , \filter_0/n5796 ,
         \filter_0/n5793 , \filter_0/n5792 , \filter_0/n5789 ,
         \filter_0/n5788 , \filter_0/n5785 , \filter_0/n5784 ,
         \filter_0/n5781 , \filter_0/n5780 , \filter_0/n5777 ,
         \filter_0/n5776 , \filter_0/n5773 , \filter_0/n5772 ,
         \filter_0/n5769 , \filter_0/n5768 , \filter_0/n5765 ,
         \filter_0/n5764 , \filter_0/n5761 , \filter_0/n5760 ,
         \filter_0/n5757 , \filter_0/n5756 , \filter_0/n5753 ,
         \filter_0/n5752 , \filter_0/n5749 , \filter_0/n5748 ,
         \filter_0/n5745 , \filter_0/n5744 , \filter_0/n5741 ,
         \filter_0/n5740 , \filter_0/n5737 , \filter_0/n5736 ,
         \filter_0/n5733 , \filter_0/n5732 , \filter_0/n5729 ,
         \filter_0/n5728 , \filter_0/n5725 , \filter_0/n5724 ,
         \filter_0/n5721 , \filter_0/n5720 , \filter_0/n5717 ,
         \filter_0/n5716 , \filter_0/n5713 , \filter_0/n5712 ,
         \filter_0/n5709 , \filter_0/n5708 , \filter_0/n5705 ,
         \filter_0/n5704 , \filter_0/n5701 , \filter_0/n5700 ,
         \filter_0/n5697 , \filter_0/n5696 , \filter_0/n5693 ,
         \filter_0/n5692 , \filter_0/n5689 , \filter_0/n5688 ,
         \filter_0/n5685 , \filter_0/n5684 , \filter_0/n5681 ,
         \filter_0/n5680 , \filter_0/n5677 , \filter_0/n5676 ,
         \filter_0/n5673 , \filter_0/n5672 , \filter_0/n5669 ,
         \filter_0/n5668 , \filter_0/n5665 , \filter_0/n5664 ,
         \filter_0/n5661 , \filter_0/n5660 , \filter_0/n5657 ,
         \filter_0/n5656 , \filter_0/n5653 , \filter_0/n5652 ,
         \filter_0/n5649 , \filter_0/n5648 , \filter_0/n5645 ,
         \filter_0/n5644 , \filter_0/n5641 , \filter_0/n5640 ,
         \filter_0/n5637 , \filter_0/n5636 , \filter_0/n5633 ,
         \filter_0/n5632 , \filter_0/n5629 , \filter_0/n5628 ,
         \filter_0/n5625 , \filter_0/n5624 , \filter_0/n5621 ,
         \filter_0/n5620 , \filter_0/n5617 , \filter_0/n5616 ,
         \filter_0/n5613 , \filter_0/n5612 , \filter_0/n5609 ,
         \filter_0/n5608 , \filter_0/n5605 , \filter_0/n5604 ,
         \filter_0/n5601 , \filter_0/n5600 , \filter_0/n5597 ,
         \filter_0/n5596 , \filter_0/n5593 , \filter_0/n5592 ,
         \filter_0/n5589 , \filter_0/n5588 , \filter_0/n5585 ,
         \filter_0/n5584 , \filter_0/n5581 , \filter_0/n5580 ,
         \filter_0/n5577 , \filter_0/n5576 , \filter_0/n5573 ,
         \filter_0/n5572 , \filter_0/n5569 , \filter_0/n5568 ,
         \filter_0/n5565 , \filter_0/n5564 , \filter_0/n5561 ,
         \filter_0/n5560 , \filter_0/n5557 , \filter_0/n5556 ,
         \filter_0/n5553 , \filter_0/n5552 , \filter_0/n5549 ,
         \filter_0/n5548 , \filter_0/n5545 , \filter_0/n5544 ,
         \filter_0/n5541 , \filter_0/n5540 , \filter_0/n5537 ,
         \filter_0/n5536 , \filter_0/n5533 , \filter_0/n5532 ,
         \filter_0/n5529 , \filter_0/n5528 , \filter_0/n5525 ,
         \filter_0/n5524 , \filter_0/n5521 , \filter_0/n5520 ,
         \filter_0/n5517 , \filter_0/n5516 , \filter_0/n5513 ,
         \filter_0/n5512 , \filter_0/n5509 , \filter_0/n5508 ,
         \filter_0/n5505 , \filter_0/n5504 , \filter_0/n5501 ,
         \filter_0/n5500 , \filter_0/n5497 , \filter_0/n5496 ,
         \filter_0/n5493 , \filter_0/n5492 , \filter_0/n5489 ,
         \filter_0/n5488 , \filter_0/n5485 , \filter_0/n5484 ,
         \filter_0/n5481 , \filter_0/n5480 , \filter_0/n5477 ,
         \filter_0/n5476 , \filter_0/n5473 , \filter_0/n5472 ,
         \filter_0/n5469 , \filter_0/n5468 , \filter_0/n5465 ,
         \filter_0/n5464 , \filter_0/n5461 , \filter_0/n5460 ,
         \filter_0/n5457 , \filter_0/n5456 , \filter_0/n5453 ,
         \filter_0/n5452 , \filter_0/n5449 , \filter_0/n5448 ,
         \filter_0/n5445 , \filter_0/n5444 , \filter_0/n5441 ,
         \filter_0/n5440 , \filter_0/n5437 , \filter_0/n5436 ,
         \filter_0/n5433 , \filter_0/n5432 , \filter_0/n5429 ,
         \filter_0/n5428 , \filter_0/n5425 , \filter_0/n5424 ,
         \filter_0/n5421 , \filter_0/n5420 , \filter_0/n5417 ,
         \filter_0/n5416 , \filter_0/n5413 , \filter_0/n5412 ,
         \filter_0/n5409 , \filter_0/n5408 , \filter_0/n5405 ,
         \filter_0/n5404 , \filter_0/n5401 , \filter_0/n5400 ,
         \filter_0/n5397 , \filter_0/n5396 , \filter_0/n5393 ,
         \filter_0/n5392 , \filter_0/n5389 , \filter_0/n5388 ,
         \filter_0/n5385 , \filter_0/n5384 , \filter_0/n5381 ,
         \filter_0/n5380 , \filter_0/n5377 , \filter_0/n5376 ,
         \filter_0/n5373 , \filter_0/n5372 , \filter_0/n5369 ,
         \filter_0/n5368 , \filter_0/n5365 , \filter_0/n5364 ,
         \filter_0/n5361 , \filter_0/n5360 , \filter_0/n5357 ,
         \filter_0/n5356 , \filter_0/n5353 , \filter_0/n5352 ,
         \filter_0/n5349 , \filter_0/n5348 , \filter_0/n5345 ,
         \filter_0/n5344 , \filter_0/n5341 , \filter_0/n5340 ,
         \filter_0/n5337 , \filter_0/n5336 , \filter_0/n5333 ,
         \filter_0/n5332 , \filter_0/n5329 , \filter_0/n5328 ,
         \filter_0/n5325 , \filter_0/n5324 , \filter_0/n5321 ,
         \filter_0/n5320 , \filter_0/n5317 , \filter_0/n5316 ,
         \filter_0/n5313 , \filter_0/n5312 , \filter_0/n5309 ,
         \filter_0/n5308 , \filter_0/n5305 , \filter_0/n5304 ,
         \filter_0/n5301 , \filter_0/n5300 , \filter_0/n5297 ,
         \filter_0/n5296 , \filter_0/n5293 , \filter_0/n5292 ,
         \filter_0/n5289 , \filter_0/n5288 , \filter_0/n5285 ,
         \filter_0/n5284 , \filter_0/n5281 , \filter_0/n5280 ,
         \filter_0/n5277 , \filter_0/n5276 , \filter_0/n5273 ,
         \filter_0/n5272 , \filter_0/n5269 , \filter_0/n5268 ,
         \filter_0/n5265 , \filter_0/n5264 , \filter_0/n5261 ,
         \filter_0/n5260 , \filter_0/n5257 , \filter_0/n5256 ,
         \filter_0/n5253 , \filter_0/n5252 , \filter_0/n5249 ,
         \filter_0/n5248 , \filter_0/n5245 , \filter_0/n5244 ,
         \filter_0/n5241 , \filter_0/n5240 , \filter_0/n5237 ,
         \filter_0/n5236 , \filter_0/n5233 , \filter_0/n5232 ,
         \filter_0/n5229 , \filter_0/n5228 , \filter_0/n5225 ,
         \filter_0/n5224 , \filter_0/n5221 , \filter_0/n5220 ,
         \filter_0/n5217 , \filter_0/n5216 , \filter_0/n5213 ,
         \filter_0/n5212 , \filter_0/n5209 , \filter_0/n5208 ,
         \filter_0/n5205 , \filter_0/n5204 , \filter_0/n5201 ,
         \filter_0/n5200 , \filter_0/n5197 , \filter_0/n5196 ,
         \filter_0/n5193 , \filter_0/n5192 , \filter_0/n5189 ,
         \filter_0/n5188 , \filter_0/n5185 , \filter_0/n5184 ,
         \filter_0/n5181 , \filter_0/n5180 , \filter_0/n5177 ,
         \filter_0/n5176 , \filter_0/n5173 , \filter_0/n5172 ,
         \filter_0/n5169 , \filter_0/n5168 , \filter_0/n5165 ,
         \filter_0/n5164 , \filter_0/n5161 , \filter_0/n5160 ,
         \filter_0/n5157 , \filter_0/n5156 , \filter_0/n5153 ,
         \filter_0/n5152 , \filter_0/n5149 , \filter_0/n5148 ,
         \filter_0/n5145 , \filter_0/n5144 , \filter_0/n5141 ,
         \filter_0/n5140 , \filter_0/n5137 , \filter_0/n5136 ,
         \filter_0/n5133 , \filter_0/n5132 , \filter_0/n5129 ,
         \filter_0/n5128 , \filter_0/n5125 , \filter_0/n5124 ,
         \filter_0/n5121 , \filter_0/n5120 , \filter_0/n5117 ,
         \filter_0/n5116 , \filter_0/n5113 , \filter_0/n5112 ,
         \filter_0/n5109 , \filter_0/n5108 , \filter_0/n5105 ,
         \filter_0/n5104 , \filter_0/n5101 , \filter_0/n5100 ,
         \filter_0/n5097 , \filter_0/n5096 , \filter_0/n5093 ,
         \filter_0/n5092 , \filter_0/n5089 , \filter_0/n5088 ,
         \filter_0/n5085 , \filter_0/n5084 , \filter_0/n5081 ,
         \filter_0/n5080 , \filter_0/n5077 , \filter_0/n5076 ,
         \filter_0/n5073 , \filter_0/n5072 , \filter_0/n5069 ,
         \filter_0/n5068 , \filter_0/n5065 , \filter_0/n5064 ,
         \filter_0/n5061 , \filter_0/n5060 , \filter_0/n5057 ,
         \filter_0/n5056 , \filter_0/n5053 , \filter_0/n5052 ,
         \filter_0/n5049 , \filter_0/n5048 , \filter_0/n5045 ,
         \filter_0/n5044 , \filter_0/n5041 , \filter_0/n5040 ,
         \filter_0/n5037 , \filter_0/n5036 , \filter_0/n5033 ,
         \filter_0/n5032 , \filter_0/n5029 , \filter_0/n5028 ,
         \filter_0/n5025 , \filter_0/n5024 , \filter_0/n5021 ,
         \filter_0/n5020 , \filter_0/n5017 , \filter_0/n5016 ,
         \filter_0/n5013 , \filter_0/n5012 , \filter_0/n5009 ,
         \filter_0/n5008 , \filter_0/n5005 , \filter_0/n5004 ,
         \filter_0/n5001 , \filter_0/n5000 , \filter_0/n4997 ,
         \filter_0/n4996 , \filter_0/n4993 , \filter_0/n4992 ,
         \filter_0/n4989 , \filter_0/n4988 , \filter_0/n4985 ,
         \filter_0/n4984 , \filter_0/n4981 , \filter_0/n4980 , n29671, n29672,
         n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
         n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688,
         n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696,
         n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
         n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712,
         n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720,
         n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
         n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736,
         n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
         n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752,
         n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760,
         n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
         n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
         n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784,
         n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792,
         n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
         n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
         n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
         n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
         n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832,
         n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840,
         n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
         n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856,
         n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
         n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
         n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880,
         n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
         n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
         n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904,
         n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912,
         n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
         n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
         n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936,
         n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
         n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952,
         n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
         n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968,
         n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976,
         n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
         n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
         n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000,
         n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
         n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
         n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
         n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
         n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
         n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048,
         n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
         n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
         n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
         n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080,
         n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
         n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
         n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
         n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
         n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120,
         n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
         n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
         n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144,
         n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152,
         n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
         n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168,
         n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
         n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184,
         n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192,
         n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
         n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
         n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216,
         n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
         n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
         n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240,
         n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
         n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256,
         n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264,
         n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272,
         n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
         n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288,
         n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
         n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
         n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312,
         n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
         n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
         n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336,
         n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344,
         n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
         n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360,
         n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368,
         n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
         n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384,
         n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
         n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
         n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408,
         n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
         n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424,
         n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432,
         n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440,
         n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
         n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456,
         n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
         n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472,
         n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480,
         n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
         n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496,
         n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
         n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
         n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
         n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528,
         n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
         n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
         n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552,
         n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
         n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
         n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
         n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584,
         n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
         n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600,
         n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
         n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616,
         n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624,
         n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
         n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
         n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648,
         n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656,
         n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
         n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672,
         n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
         n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
         n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696,
         n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
         n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
         n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
         n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728,
         n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
         n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744,
         n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
         n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
         n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768,
         n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
         n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784,
         n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792,
         n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800,
         n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
         n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816,
         n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
         n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832,
         n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840,
         n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
         n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
         n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864,
         n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872,
         n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
         n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888,
         n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
         n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904,
         n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
         n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920,
         n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
         n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936,
         n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944,
         n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
         n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960,
         n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
         n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
         n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
         n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992,
         n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
         n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008,
         n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016,
         n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
         n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032,
         n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
         n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
         n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056,
         n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064,
         n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
         n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
         n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088,
         n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
         n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104,
         n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
         n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
         n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128,
         n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136,
         n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
         n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
         n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160,
         n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
         n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176,
         n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
         n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
         n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200,
         n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
         n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
         n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224,
         n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232,
         n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
         n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248,
         n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
         n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
         n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272,
         n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280,
         n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
         n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
         n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304,
         n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
         n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320,
         n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
         n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
         n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344,
         n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
         n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360,
         n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368,
         n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376,
         n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
         n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392,
         n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
         n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
         n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416,
         n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
         n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432,
         n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440,
         n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
         n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
         n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464,
         n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
         n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480,
         n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488,
         n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
         n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
         n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512,
         n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520,
         n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
         n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536,
         n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
         n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552,
         n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
         n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
         n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
         n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584,
         n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
         n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
         n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608,
         n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
         n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
         n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632,
         n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
         n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
         n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
         n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
         n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
         n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680,
         n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
         n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
         n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704,
         n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
         n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720,
         n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
         n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
         n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
         n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752,
         n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
         n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768,
         n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776,
         n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784,
         n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
         n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800,
         n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808,
         n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816,
         n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824,
         n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832,
         n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840,
         n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848,
         n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856,
         n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864,
         n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872,
         n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880,
         n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888,
         n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896,
         n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904,
         n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912,
         n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920,
         n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928,
         n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
         n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944,
         n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952,
         n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960,
         n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968,
         n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976,
         n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984,
         n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992,
         n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000,
         n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008,
         n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016,
         n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024,
         n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
         n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040,
         n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048,
         n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056,
         n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064,
         n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072,
         n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080,
         n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088,
         n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096,
         n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
         n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112,
         n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
         n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
         n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136,
         n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
         n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152,
         n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160,
         n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168,
         n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176,
         n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184,
         n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192,
         n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200,
         n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208,
         n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216,
         n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224,
         n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232,
         n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240,
         n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248,
         n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256,
         n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264,
         n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272,
         n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280,
         n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288,
         n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296,
         n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304,
         n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312,
         n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320,
         n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328,
         n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336,
         n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344,
         n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352,
         n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360,
         n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368,
         n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376,
         n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384,
         n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
         n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400,
         n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
         n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
         n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424,
         n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432,
         n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440,
         n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448,
         n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
         n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
         n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472,
         n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480,
         n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488,
         n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496,
         n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504,
         n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512,
         n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520,
         n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528,
         n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
         n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544,
         n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552,
         n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560,
         n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568,
         n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576,
         n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
         n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592,
         n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600,
         n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608,
         n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616,
         n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624,
         n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632,
         n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640,
         n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648,
         n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656,
         n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664,
         n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672,
         n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680,
         n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688,
         n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696,
         n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
         n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712,
         n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720,
         n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728,
         n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736,
         n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744,
         n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752,
         n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760,
         n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
         n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776,
         n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784,
         n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792,
         n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800,
         n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808,
         n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816,
         n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824,
         n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832,
         n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
         n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848,
         n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856,
         n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864,
         n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872,
         n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880,
         n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888,
         n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
         n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904,
         n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
         n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
         n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928,
         n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936,
         n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944,
         n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952,
         n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960,
         n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968,
         n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976,
         n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
         n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992,
         n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000,
         n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008,
         n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016,
         n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024,
         n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032,
         n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040,
         n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048,
         n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
         n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064,
         n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072,
         n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
         n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
         n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096,
         n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104,
         n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
         n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120,
         n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
         n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136,
         n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144,
         n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152,
         n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160,
         n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168,
         n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176,
         n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184,
         n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192,
         n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
         n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208,
         n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216,
         n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224,
         n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232,
         n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240,
         n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248,
         n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
         n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264,
         n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
         n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280,
         n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288,
         n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296,
         n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304,
         n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312,
         n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320,
         n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328,
         n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336,
         n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344,
         n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352,
         n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360,
         n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368,
         n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
         n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384,
         n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392,
         n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400,
         n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408,
         n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416,
         n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424,
         n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432,
         n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440,
         n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448,
         n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456,
         n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464,
         n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472,
         n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480,
         n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488,
         n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496,
         n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504,
         n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512,
         n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520,
         n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528,
         n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536,
         n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544,
         n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552,
         n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
         n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568,
         n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576,
         n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584,
         n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592,
         n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600,
         n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608,
         n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616,
         n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624,
         n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632,
         n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640,
         n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648,
         n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656,
         n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664,
         n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672,
         n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680,
         n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688,
         n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696,
         n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
         n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712,
         n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720,
         n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728,
         n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736,
         n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744,
         n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752,
         n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
         n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768,
         n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776,
         n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784,
         n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792,
         n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800,
         n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808,
         n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
         n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824,
         n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832,
         n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840,
         n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848,
         n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856,
         n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864,
         n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
         n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880,
         n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888,
         n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896,
         n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904,
         n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912,
         n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
         n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928,
         n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936,
         n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944,
         n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952,
         n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960,
         n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968,
         n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976,
         n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984,
         n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
         n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000,
         n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008,
         n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
         n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
         n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032,
         n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040,
         n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048,
         n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056,
         n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064,
         n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072,
         n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080,
         n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
         n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096,
         n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104,
         n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112,
         n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120,
         n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128,
         n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136,
         n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
         n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152,
         n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
         n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
         n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176,
         n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184,
         n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192,
         n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200,
         n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
         n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216,
         n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224,
         n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232,
         n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
         n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248,
         n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256,
         n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264,
         n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272,
         n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280,
         n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288,
         n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296,
         n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304,
         n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312,
         n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320,
         n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328,
         n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
         n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344,
         n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352,
         n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360,
         n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368,
         n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
         n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384,
         n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392,
         n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400,
         n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
         n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416,
         n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424,
         n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432,
         n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440,
         n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448,
         n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456,
         n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464,
         n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472,
         n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
         n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488,
         n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
         n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504,
         n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512,
         n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520,
         n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528,
         n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536,
         n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544,
         n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552,
         n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560,
         n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568,
         n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576,
         n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584,
         n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592,
         n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600,
         n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608,
         n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616,
         n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624,
         n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632,
         n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
         n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648,
         n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656,
         n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664,
         n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672,
         n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680,
         n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688,
         n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696,
         n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704,
         n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712,
         n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720,
         n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728,
         n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736,
         n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744,
         n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752,
         n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760,
         n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
         n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776,
         n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
         n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792,
         n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800,
         n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808,
         n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816,
         n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824,
         n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832,
         n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840,
         n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848,
         n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856,
         n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864,
         n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872,
         n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880,
         n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888,
         n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896,
         n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904,
         n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912,
         n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920,
         n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928,
         n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936,
         n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944,
         n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952,
         n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960,
         n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968,
         n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976,
         n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984,
         n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992,
         n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000,
         n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008,
         n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016,
         n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024,
         n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032,
         n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040,
         n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048,
         n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056,
         n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064,
         n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072,
         n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080,
         n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088,
         n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096,
         n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104,
         n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112,
         n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120,
         n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128,
         n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136,
         n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144,
         n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152,
         n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160,
         n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168,
         n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176,
         n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184,
         n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192,
         n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200,
         n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208,
         n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216,
         n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224,
         n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232,
         n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
         n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
         n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256,
         n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264,
         n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
         n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280,
         n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288,
         n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296,
         n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304,
         n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312,
         n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320,
         n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328,
         n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336,
         n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
         n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352,
         n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360,
         n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368,
         n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376,
         n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384,
         n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392,
         n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400,
         n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408,
         n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
         n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424,
         n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
         n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
         n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448,
         n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456,
         n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
         n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472,
         n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480,
         n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
         n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496,
         n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
         n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512,
         n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520,
         n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528,
         n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536,
         n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544,
         n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552,
         n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
         n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568,
         n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
         n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584,
         n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592,
         n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600,
         n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608,
         n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616,
         n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624,
         n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632,
         n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640,
         n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
         n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656,
         n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664,
         n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672,
         n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680,
         n35681, n35682, n35683, n35684, n35685, n40858, n40859, n40860,
         n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868,
         n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876,
         n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884,
         n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892,
         n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900,
         n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908,
         n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916,
         n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924,
         n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932,
         n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940,
         n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948,
         n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956,
         n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964,
         n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972,
         n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980,
         n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988,
         n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996,
         n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004,
         n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012,
         n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020,
         n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028,
         n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036,
         n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044,
         n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052,
         n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060,
         n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068,
         n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076,
         n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084,
         n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092,
         n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100,
         n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108,
         n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116,
         n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124,
         n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132,
         n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
         n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148,
         n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156,
         n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164,
         n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172,
         n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180,
         n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188,
         n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196,
         n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204,
         n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212,
         n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220,
         n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228,
         n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236,
         n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244,
         n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252,
         n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260,
         n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268,
         n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276,
         n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284,
         n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292,
         n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300,
         n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308,
         n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316,
         n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324,
         n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332,
         n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340,
         n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348,
         n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356,
         n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364,
         n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372,
         n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380,
         n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388,
         n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396,
         n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404,
         n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412,
         n41413, n41414, n41415, n41416, n41417, n41418, n41419, n41420,
         n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428,
         n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436,
         n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444,
         n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452,
         n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460,
         n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468,
         n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476,
         n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484,
         n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492,
         n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500,
         n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508,
         n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516,
         n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524,
         n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532,
         n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540,
         n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548,
         n41549, n41550, n41551, n41552, n41553, n41554, n41555, n41556,
         n41557, n41558, n41559, n41560, n41561, n41562, n41563, n41564,
         n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572,
         n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580,
         n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588,
         n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596,
         n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604,
         n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612,
         n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620,
         n41621, n41622, n41623, n41624, n41625, n41626, n41627, n41628,
         n41629, n41630, n41631, n41632, n41633, n41634, n41635, n41636,
         n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644,
         n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652,
         n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660,
         n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668,
         n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676,
         n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684,
         n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692,
         n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700,
         n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708,
         n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716,
         n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724,
         n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732,
         n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740,
         n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748,
         n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756,
         n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764,
         n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772,
         n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780,
         n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788,
         n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796,
         n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804,
         n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812,
         n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820,
         n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828,
         n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836,
         n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844,
         n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852,
         n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860,
         n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868,
         n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876,
         n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884,
         n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892,
         n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900,
         n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908,
         n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916,
         n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924,
         n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932,
         n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940,
         n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948,
         n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956,
         n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964,
         n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972,
         n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980,
         n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988,
         n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996,
         n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004,
         n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012,
         n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020,
         n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028,
         n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036,
         n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044,
         n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052,
         n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060,
         n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068,
         n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076,
         n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084,
         n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092,
         n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100,
         n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108,
         n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116,
         n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124,
         n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132,
         n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140,
         n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148,
         n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156,
         n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
         n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172,
         n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180,
         n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188,
         n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196,
         n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204,
         n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212,
         n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220,
         n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228,
         n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236,
         n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244,
         n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252,
         n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260,
         n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268,
         n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276,
         n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284,
         n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292,
         n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300,
         n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
         n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316,
         n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324,
         n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332,
         n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340,
         n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348,
         n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356,
         n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364,
         n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372,
         n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380,
         n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388,
         n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396,
         n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404,
         n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412,
         n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420,
         n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428,
         n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436,
         n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444,
         n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452,
         n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460,
         n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468,
         n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476,
         n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484,
         n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492,
         n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500,
         n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508,
         n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516,
         n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524,
         n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532,
         n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540,
         n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548,
         n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556,
         n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564,
         n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572,
         n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580,
         n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588,
         n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596,
         n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604,
         n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612,
         n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620,
         n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628,
         n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636,
         n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644,
         n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652,
         n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660,
         n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668,
         n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676,
         n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684,
         n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692,
         n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700,
         n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708,
         n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716,
         n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724,
         n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732,
         n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740,
         n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748,
         n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756,
         n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764,
         n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772,
         n42773, n42774, n42775;
  wire   [19:0] reg_i_0;
  wire   [19:0] reg_i_1;
  wire   [19:0] reg_i_2;
  wire   [19:0] reg_i_3;
  wire   [19:0] reg_i_4;
  wire   [19:0] reg_i_5;
  wire   [19:0] reg_i_6;
  wire   [19:0] reg_i_7;
  wire   [19:0] reg_i_8;
  wire   [19:0] reg_i_9;
  wire   [19:0] reg_i_10;
  wire   [19:0] reg_i_11;
  wire   [19:0] reg_i_12;
  wire   [19:0] reg_i_13;
  wire   [19:0] reg_i_14;
  wire   [19:0] reg_i_15;
  wire   [19:0] reg_w_0;
  wire   [19:0] reg_w_1;
  wire   [19:0] reg_w_2;
  wire   [19:0] reg_w_3;
  wire   [19:0] reg_w_4;
  wire   [19:0] reg_w_5;
  wire   [19:0] reg_w_6;
  wire   [19:0] reg_w_7;
  wire   [19:0] reg_w_8;
  wire   [19:0] reg_w_9;
  wire   [19:0] reg_w_10;
  wire   [19:0] reg_w_11;
  wire   [19:0] reg_w_12;
  wire   [19:0] reg_w_13;
  wire   [19:0] reg_w_14;
  wire   [19:0] reg_w_15;
  wire   [19:0] reg_ii_0;
  wire   [19:0] reg_ii_1;
  wire   [19:0] reg_ii_2;
  wire   [19:0] reg_ii_3;
  wire   [19:0] reg_ii_4;
  wire   [19:0] reg_ii_5;
  wire   [19:0] reg_ii_6;
  wire   [19:0] reg_ii_7;
  wire   [19:0] reg_ii_8;
  wire   [19:0] reg_ii_9;
  wire   [19:0] reg_ii_10;
  wire   [19:0] reg_ii_11;
  wire   [19:0] reg_ii_12;
  wire   [19:0] reg_ii_13;
  wire   [19:0] reg_ii_14;
  wire   [19:0] reg_ii_15;
  wire   [19:0] reg_ww_0;
  wire   [19:0] reg_ww_1;
  wire   [19:0] reg_ww_2;
  wire   [19:0] reg_ww_3;
  wire   [19:0] reg_ww_4;
  wire   [19:0] reg_ww_5;
  wire   [19:0] reg_ww_6;
  wire   [19:0] reg_ww_7;
  wire   [19:0] reg_ww_8;
  wire   [19:0] reg_ww_9;
  wire   [19:0] reg_ww_10;
  wire   [19:0] reg_ww_11;
  wire   [19:0] reg_ww_12;
  wire   [19:0] reg_ww_13;
  wire   [19:0] reg_ww_14;
  wire   [19:0] reg_ww_15;
  wire   [19:0] reg_iii_0;
  wire   [19:0] reg_iii_1;
  wire   [19:0] reg_iii_2;
  wire   [19:0] reg_iii_3;
  wire   [19:0] reg_iii_4;
  wire   [19:0] reg_iii_5;
  wire   [19:0] reg_iii_6;
  wire   [19:0] reg_iii_7;
  wire   [19:0] reg_iii_8;
  wire   [19:0] reg_iii_9;
  wire   [19:0] reg_iii_10;
  wire   [19:0] reg_iii_11;
  wire   [19:0] reg_iii_12;
  wire   [19:0] reg_iii_13;
  wire   [19:0] reg_iii_14;
  wire   [19:0] reg_iii_15;
  wire   [19:0] reg_www_0;
  wire   [19:0] reg_www_1;
  wire   [19:0] reg_www_2;
  wire   [19:0] reg_www_3;
  wire   [19:0] reg_www_4;
  wire   [19:0] reg_www_5;
  wire   [19:0] reg_www_6;
  wire   [19:0] reg_www_7;
  wire   [19:0] reg_www_8;
  wire   [19:0] reg_www_9;
  wire   [19:0] reg_www_10;
  wire   [19:0] reg_www_11;
  wire   [19:0] reg_www_12;
  wire   [19:0] reg_www_13;
  wire   [19:0] reg_www_14;
  wire   [19:0] reg_www_15;
  wire   [31:0] reg_i_mask;
  wire   [31:0] reg_w_mask;
  wire   [19:0] reg_oi_0;
  wire   [19:0] reg_oi_1;
  wire   [19:0] reg_oi_2;
  wire   [19:0] reg_oi_3;
  wire   [19:0] reg_oi_4;
  wire   [19:0] reg_oi_5;
  wire   [19:0] reg_oi_6;
  wire   [19:0] reg_oi_7;
  wire   [19:0] reg_oi_8;
  wire   [19:0] reg_oi_9;
  wire   [19:0] reg_oi_10;
  wire   [19:0] reg_oi_11;
  wire   [19:0] reg_oi_12;
  wire   [19:0] reg_oi_13;
  wire   [19:0] reg_oi_14;
  wire   [19:0] reg_oi_15;
  wire   [19:0] reg_ow_0;
  wire   [19:0] reg_ow_1;
  wire   [19:0] reg_ow_2;
  wire   [19:0] reg_ow_3;
  wire   [19:0] reg_ow_4;
  wire   [19:0] reg_ow_5;
  wire   [19:0] reg_ow_6;
  wire   [19:0] reg_ow_7;
  wire   [19:0] reg_ow_8;
  wire   [19:0] reg_ow_9;
  wire   [19:0] reg_ow_10;
  wire   [19:0] reg_ow_11;
  wire   [19:0] reg_ow_12;
  wire   [19:0] reg_ow_13;
  wire   [19:0] reg_ow_14;
  wire   [19:0] reg_ow_15;
  wire   [1:0] filter_state;
  wire   [1:0] shifter_state;

  dff_sg mask_input_ready_reg ( .D(input_ready), .CP(clk), .Q(mask_input_ready) );
  dff_sg delayed_input_ready_reg ( .D(mask_input_ready), .CP(clk), .Q(
        delayed_input_ready) );
  dff_sg filter_input_ready_reg ( .D(delayed_input_ready), .CP(clk), .Q(
        filter_input_ready) );
  dff_sg \state_reg[1]  ( .D(n5982), .CP(clk), .Q(state[1]) );
  dff_sg \state_reg[0]  ( .D(n5981), .CP(clk), .Q(state[0]) );
  dff_sg \reg_w_mask_reg[31]  ( .D(n5277), .CP(clk), .Q(reg_w_mask[31]) );
  dff_sg \reg_w_mask_reg[30]  ( .D(n5278), .CP(clk), .Q(reg_w_mask[30]) );
  dff_sg \reg_w_mask_reg[29]  ( .D(n5279), .CP(clk), .Q(reg_w_mask[29]) );
  dff_sg \reg_w_mask_reg[28]  ( .D(n5280), .CP(clk), .Q(reg_w_mask[28]) );
  dff_sg \reg_w_mask_reg[27]  ( .D(n5281), .CP(clk), .Q(reg_w_mask[27]) );
  dff_sg \reg_w_mask_reg[26]  ( .D(n5282), .CP(clk), .Q(reg_w_mask[26]) );
  dff_sg \reg_w_mask_reg[25]  ( .D(n5283), .CP(clk), .Q(reg_w_mask[25]) );
  dff_sg \reg_w_mask_reg[24]  ( .D(n5284), .CP(clk), .Q(reg_w_mask[24]) );
  dff_sg \reg_w_mask_reg[23]  ( .D(n5285), .CP(clk), .Q(reg_w_mask[23]) );
  dff_sg \reg_w_mask_reg[22]  ( .D(n5286), .CP(clk), .Q(reg_w_mask[22]) );
  dff_sg \reg_w_mask_reg[21]  ( .D(n5287), .CP(clk), .Q(reg_w_mask[21]) );
  dff_sg \reg_w_mask_reg[20]  ( .D(n5288), .CP(clk), .Q(reg_w_mask[20]) );
  dff_sg \reg_w_mask_reg[19]  ( .D(n5289), .CP(clk), .Q(reg_w_mask[19]) );
  dff_sg \reg_w_mask_reg[18]  ( .D(n5290), .CP(clk), .Q(reg_w_mask[18]) );
  dff_sg \reg_w_mask_reg[17]  ( .D(n5291), .CP(clk), .Q(reg_w_mask[17]) );
  dff_sg \reg_w_mask_reg[16]  ( .D(n5292), .CP(clk), .Q(reg_w_mask[16]) );
  dff_sg \reg_w_mask_reg[15]  ( .D(n5293), .CP(clk), .Q(reg_w_mask[15]) );
  dff_sg \reg_w_mask_reg[14]  ( .D(n5294), .CP(clk), .Q(reg_w_mask[14]) );
  dff_sg \reg_w_mask_reg[13]  ( .D(n5295), .CP(clk), .Q(reg_w_mask[13]) );
  dff_sg \reg_w_mask_reg[12]  ( .D(n5296), .CP(clk), .Q(reg_w_mask[12]) );
  dff_sg \reg_w_mask_reg[11]  ( .D(n5297), .CP(clk), .Q(reg_w_mask[11]) );
  dff_sg \reg_w_mask_reg[10]  ( .D(n5298), .CP(clk), .Q(reg_w_mask[10]) );
  dff_sg \reg_w_mask_reg[9]  ( .D(n5299), .CP(clk), .Q(reg_w_mask[9]) );
  dff_sg \reg_w_mask_reg[8]  ( .D(n5300), .CP(clk), .Q(reg_w_mask[8]) );
  dff_sg \reg_w_mask_reg[7]  ( .D(n5301), .CP(clk), .Q(reg_w_mask[7]) );
  dff_sg \reg_w_mask_reg[6]  ( .D(n5302), .CP(clk), .Q(reg_w_mask[6]) );
  dff_sg \reg_w_mask_reg[5]  ( .D(n5303), .CP(clk), .Q(reg_w_mask[5]) );
  dff_sg \reg_w_mask_reg[4]  ( .D(n5304), .CP(clk), .Q(reg_w_mask[4]) );
  dff_sg \reg_w_mask_reg[3]  ( .D(n5305), .CP(clk), .Q(reg_w_mask[3]) );
  dff_sg \reg_w_mask_reg[2]  ( .D(n5306), .CP(clk), .Q(reg_w_mask[2]) );
  dff_sg \reg_w_mask_reg[1]  ( .D(n5307), .CP(clk), .Q(reg_w_mask[1]) );
  dff_sg \reg_w_mask_reg[0]  ( .D(n5308), .CP(clk), .Q(reg_w_mask[0]) );
  dff_sg \reg_i_mask_reg[31]  ( .D(n5309), .CP(clk), .Q(reg_i_mask[31]) );
  dff_sg \reg_i_mask_reg[30]  ( .D(n5310), .CP(clk), .Q(reg_i_mask[30]) );
  dff_sg \reg_i_mask_reg[29]  ( .D(n5311), .CP(clk), .Q(reg_i_mask[29]) );
  dff_sg \reg_i_mask_reg[28]  ( .D(n5312), .CP(clk), .Q(reg_i_mask[28]) );
  dff_sg \reg_i_mask_reg[27]  ( .D(n5313), .CP(clk), .Q(reg_i_mask[27]) );
  dff_sg \reg_i_mask_reg[26]  ( .D(n5314), .CP(clk), .Q(reg_i_mask[26]) );
  dff_sg \reg_i_mask_reg[25]  ( .D(n5315), .CP(clk), .Q(reg_i_mask[25]) );
  dff_sg \reg_i_mask_reg[24]  ( .D(n5316), .CP(clk), .Q(reg_i_mask[24]) );
  dff_sg \reg_i_mask_reg[23]  ( .D(n5317), .CP(clk), .Q(reg_i_mask[23]) );
  dff_sg \reg_i_mask_reg[22]  ( .D(n5318), .CP(clk), .Q(reg_i_mask[22]) );
  dff_sg \reg_i_mask_reg[21]  ( .D(n5319), .CP(clk), .Q(reg_i_mask[21]) );
  dff_sg \reg_i_mask_reg[20]  ( .D(n5320), .CP(clk), .Q(reg_i_mask[20]) );
  dff_sg \reg_i_mask_reg[19]  ( .D(n5321), .CP(clk), .Q(reg_i_mask[19]) );
  dff_sg \reg_i_mask_reg[18]  ( .D(n5322), .CP(clk), .Q(reg_i_mask[18]) );
  dff_sg \reg_i_mask_reg[17]  ( .D(n5323), .CP(clk), .Q(reg_i_mask[17]) );
  dff_sg \reg_i_mask_reg[16]  ( .D(n5324), .CP(clk), .Q(reg_i_mask[16]) );
  dff_sg \reg_i_mask_reg[15]  ( .D(n5325), .CP(clk), .Q(reg_i_mask[15]) );
  dff_sg \reg_i_mask_reg[14]  ( .D(n5326), .CP(clk), .Q(reg_i_mask[14]) );
  dff_sg \reg_i_mask_reg[13]  ( .D(n5327), .CP(clk), .Q(reg_i_mask[13]) );
  dff_sg \reg_i_mask_reg[12]  ( .D(n5328), .CP(clk), .Q(reg_i_mask[12]) );
  dff_sg \reg_i_mask_reg[11]  ( .D(n5329), .CP(clk), .Q(reg_i_mask[11]) );
  dff_sg \reg_i_mask_reg[10]  ( .D(n5330), .CP(clk), .Q(reg_i_mask[10]) );
  dff_sg \reg_i_mask_reg[9]  ( .D(n5331), .CP(clk), .Q(reg_i_mask[9]) );
  dff_sg \reg_i_mask_reg[8]  ( .D(n5332), .CP(clk), .Q(reg_i_mask[8]) );
  dff_sg \reg_i_mask_reg[7]  ( .D(n5333), .CP(clk), .Q(reg_i_mask[7]) );
  dff_sg \reg_i_mask_reg[6]  ( .D(n5334), .CP(clk), .Q(reg_i_mask[6]) );
  dff_sg \reg_i_mask_reg[5]  ( .D(n5335), .CP(clk), .Q(reg_i_mask[5]) );
  dff_sg \reg_i_mask_reg[4]  ( .D(n5336), .CP(clk), .Q(reg_i_mask[4]) );
  dff_sg \reg_i_mask_reg[3]  ( .D(n5337), .CP(clk), .Q(reg_i_mask[3]) );
  dff_sg \reg_i_mask_reg[2]  ( .D(n5338), .CP(clk), .Q(reg_i_mask[2]) );
  dff_sg \reg_i_mask_reg[1]  ( .D(n5339), .CP(clk), .Q(reg_i_mask[1]) );
  dff_sg \reg_i_mask_reg[0]  ( .D(n5340), .CP(clk), .Q(reg_i_mask[0]) );
  dff_sg \reg_w_15_reg[19]  ( .D(n5341), .CP(clk), .Q(reg_w_15[19]) );
  dff_sg \reg_ww_15_reg[19]  ( .D(n5210), .CP(clk), .Q(reg_ww_15[19]) );
  dff_sg \reg_www_15_reg[19]  ( .D(n5190), .CP(clk), .Q(reg_www_15[19]) );
  dff_sg \reg_w_15_reg[18]  ( .D(n5342), .CP(clk), .Q(reg_w_15[18]) );
  dff_sg \reg_ww_15_reg[18]  ( .D(n5211), .CP(clk), .Q(reg_ww_15[18]) );
  dff_sg \reg_www_15_reg[18]  ( .D(n5191), .CP(clk), .Q(reg_www_15[18]) );
  dff_sg \reg_w_15_reg[17]  ( .D(n5343), .CP(clk), .Q(reg_w_15[17]) );
  dff_sg \reg_ww_15_reg[17]  ( .D(n5212), .CP(clk), .Q(reg_ww_15[17]) );
  dff_sg \reg_www_15_reg[17]  ( .D(n5192), .CP(clk), .Q(reg_www_15[17]) );
  dff_sg \reg_w_15_reg[16]  ( .D(n5344), .CP(clk), .Q(reg_w_15[16]) );
  dff_sg \reg_ww_15_reg[16]  ( .D(n5213), .CP(clk), .Q(reg_ww_15[16]) );
  dff_sg \reg_www_15_reg[16]  ( .D(n5193), .CP(clk), .Q(reg_www_15[16]) );
  dff_sg \reg_w_15_reg[15]  ( .D(n5345), .CP(clk), .Q(reg_w_15[15]) );
  dff_sg \reg_ww_15_reg[15]  ( .D(n5214), .CP(clk), .Q(reg_ww_15[15]) );
  dff_sg \reg_www_15_reg[15]  ( .D(n5194), .CP(clk), .Q(reg_www_15[15]) );
  dff_sg \reg_w_15_reg[14]  ( .D(n5346), .CP(clk), .Q(reg_w_15[14]) );
  dff_sg \reg_ww_15_reg[14]  ( .D(n5215), .CP(clk), .Q(reg_ww_15[14]) );
  dff_sg \reg_www_15_reg[14]  ( .D(n5195), .CP(clk), .Q(reg_www_15[14]) );
  dff_sg \reg_w_15_reg[13]  ( .D(n5347), .CP(clk), .Q(reg_w_15[13]) );
  dff_sg \reg_ww_15_reg[13]  ( .D(n5216), .CP(clk), .Q(reg_ww_15[13]) );
  dff_sg \reg_www_15_reg[13]  ( .D(n5196), .CP(clk), .Q(reg_www_15[13]) );
  dff_sg \reg_w_15_reg[12]  ( .D(n5348), .CP(clk), .Q(reg_w_15[12]) );
  dff_sg \reg_ww_15_reg[12]  ( .D(n5217), .CP(clk), .Q(reg_ww_15[12]) );
  dff_sg \reg_www_15_reg[12]  ( .D(n5197), .CP(clk), .Q(reg_www_15[12]) );
  dff_sg \reg_w_15_reg[11]  ( .D(n5349), .CP(clk), .Q(reg_w_15[11]) );
  dff_sg \reg_ww_15_reg[11]  ( .D(n5218), .CP(clk), .Q(reg_ww_15[11]) );
  dff_sg \reg_www_15_reg[11]  ( .D(n5198), .CP(clk), .Q(reg_www_15[11]) );
  dff_sg \reg_w_15_reg[10]  ( .D(n5350), .CP(clk), .Q(reg_w_15[10]) );
  dff_sg \reg_ww_15_reg[10]  ( .D(n5219), .CP(clk), .Q(reg_ww_15[10]) );
  dff_sg \reg_www_15_reg[10]  ( .D(n5199), .CP(clk), .Q(reg_www_15[10]) );
  dff_sg \reg_w_15_reg[9]  ( .D(n5351), .CP(clk), .Q(reg_w_15[9]) );
  dff_sg \reg_ww_15_reg[9]  ( .D(n5220), .CP(clk), .Q(reg_ww_15[9]) );
  dff_sg \reg_www_15_reg[9]  ( .D(n5200), .CP(clk), .Q(reg_www_15[9]) );
  dff_sg \reg_w_15_reg[8]  ( .D(n5352), .CP(clk), .Q(reg_w_15[8]) );
  dff_sg \reg_ww_15_reg[8]  ( .D(n5221), .CP(clk), .Q(reg_ww_15[8]) );
  dff_sg \reg_www_15_reg[8]  ( .D(n5201), .CP(clk), .Q(reg_www_15[8]) );
  dff_sg \reg_w_15_reg[7]  ( .D(n5353), .CP(clk), .Q(reg_w_15[7]) );
  dff_sg \reg_ww_15_reg[7]  ( .D(n5222), .CP(clk), .Q(reg_ww_15[7]) );
  dff_sg \reg_www_15_reg[7]  ( .D(n5202), .CP(clk), .Q(reg_www_15[7]) );
  dff_sg \reg_w_15_reg[6]  ( .D(n5354), .CP(clk), .Q(reg_w_15[6]) );
  dff_sg \reg_ww_15_reg[6]  ( .D(n5223), .CP(clk), .Q(reg_ww_15[6]) );
  dff_sg \reg_www_15_reg[6]  ( .D(n5203), .CP(clk), .Q(reg_www_15[6]) );
  dff_sg \reg_w_15_reg[5]  ( .D(n5355), .CP(clk), .Q(reg_w_15[5]) );
  dff_sg \reg_ww_15_reg[5]  ( .D(n5224), .CP(clk), .Q(reg_ww_15[5]) );
  dff_sg \reg_www_15_reg[5]  ( .D(n5204), .CP(clk), .Q(reg_www_15[5]) );
  dff_sg \reg_w_15_reg[4]  ( .D(n5356), .CP(clk), .Q(reg_w_15[4]) );
  dff_sg \reg_ww_15_reg[4]  ( .D(n5225), .CP(clk), .Q(reg_ww_15[4]) );
  dff_sg \reg_www_15_reg[4]  ( .D(n5205), .CP(clk), .Q(reg_www_15[4]) );
  dff_sg \reg_w_15_reg[3]  ( .D(n5357), .CP(clk), .Q(reg_w_15[3]) );
  dff_sg \reg_ww_15_reg[3]  ( .D(n5226), .CP(clk), .Q(reg_ww_15[3]) );
  dff_sg \reg_www_15_reg[3]  ( .D(n5206), .CP(clk), .Q(reg_www_15[3]) );
  dff_sg \reg_w_15_reg[2]  ( .D(n5358), .CP(clk), .Q(reg_w_15[2]) );
  dff_sg \reg_ww_15_reg[2]  ( .D(n5227), .CP(clk), .Q(reg_ww_15[2]) );
  dff_sg \reg_www_15_reg[2]  ( .D(n5207), .CP(clk), .Q(reg_www_15[2]) );
  dff_sg \reg_w_15_reg[1]  ( .D(n5359), .CP(clk), .Q(reg_w_15[1]) );
  dff_sg \reg_ww_15_reg[1]  ( .D(n5228), .CP(clk), .Q(reg_ww_15[1]) );
  dff_sg \reg_www_15_reg[1]  ( .D(n5208), .CP(clk), .Q(reg_www_15[1]) );
  dff_sg \reg_w_15_reg[0]  ( .D(n5360), .CP(clk), .Q(reg_w_15[0]) );
  dff_sg \reg_ww_15_reg[0]  ( .D(n5229), .CP(clk), .Q(reg_ww_15[0]) );
  dff_sg \reg_www_15_reg[0]  ( .D(n5209), .CP(clk), .Q(reg_www_15[0]) );
  dff_sg \reg_w_14_reg[19]  ( .D(n5361), .CP(clk), .Q(reg_w_14[19]) );
  dff_sg \reg_ww_14_reg[19]  ( .D(n5250), .CP(clk), .Q(reg_ww_14[19]) );
  dff_sg \reg_www_14_reg[19]  ( .D(n5230), .CP(clk), .Q(reg_www_14[19]) );
  dff_sg \reg_w_14_reg[18]  ( .D(n5362), .CP(clk), .Q(reg_w_14[18]) );
  dff_sg \reg_ww_14_reg[18]  ( .D(n5251), .CP(clk), .Q(reg_ww_14[18]) );
  dff_sg \reg_www_14_reg[18]  ( .D(n5231), .CP(clk), .Q(reg_www_14[18]) );
  dff_sg \reg_w_14_reg[17]  ( .D(n5363), .CP(clk), .Q(reg_w_14[17]) );
  dff_sg \reg_ww_14_reg[17]  ( .D(n5252), .CP(clk), .Q(reg_ww_14[17]) );
  dff_sg \reg_www_14_reg[17]  ( .D(n5232), .CP(clk), .Q(reg_www_14[17]) );
  dff_sg \reg_w_14_reg[16]  ( .D(n5364), .CP(clk), .Q(reg_w_14[16]) );
  dff_sg \reg_ww_14_reg[16]  ( .D(n5253), .CP(clk), .Q(reg_ww_14[16]) );
  dff_sg \reg_www_14_reg[16]  ( .D(n5233), .CP(clk), .Q(reg_www_14[16]) );
  dff_sg \reg_w_14_reg[15]  ( .D(n5365), .CP(clk), .Q(reg_w_14[15]) );
  dff_sg \reg_ww_14_reg[15]  ( .D(n5254), .CP(clk), .Q(reg_ww_14[15]) );
  dff_sg \reg_www_14_reg[15]  ( .D(n5234), .CP(clk), .Q(reg_www_14[15]) );
  dff_sg \reg_w_14_reg[14]  ( .D(n5366), .CP(clk), .Q(reg_w_14[14]) );
  dff_sg \reg_ww_14_reg[14]  ( .D(n5255), .CP(clk), .Q(reg_ww_14[14]) );
  dff_sg \reg_www_14_reg[14]  ( .D(n5235), .CP(clk), .Q(reg_www_14[14]) );
  dff_sg \reg_w_14_reg[13]  ( .D(n5367), .CP(clk), .Q(reg_w_14[13]) );
  dff_sg \reg_ww_14_reg[13]  ( .D(n5256), .CP(clk), .Q(reg_ww_14[13]) );
  dff_sg \reg_www_14_reg[13]  ( .D(n5236), .CP(clk), .Q(reg_www_14[13]) );
  dff_sg \reg_w_14_reg[12]  ( .D(n5368), .CP(clk), .Q(reg_w_14[12]) );
  dff_sg \reg_ww_14_reg[12]  ( .D(n5257), .CP(clk), .Q(reg_ww_14[12]) );
  dff_sg \reg_www_14_reg[12]  ( .D(n5237), .CP(clk), .Q(reg_www_14[12]) );
  dff_sg \reg_w_14_reg[11]  ( .D(n5369), .CP(clk), .Q(reg_w_14[11]) );
  dff_sg \reg_ww_14_reg[11]  ( .D(n5258), .CP(clk), .Q(reg_ww_14[11]) );
  dff_sg \reg_www_14_reg[11]  ( .D(n5238), .CP(clk), .Q(reg_www_14[11]) );
  dff_sg \reg_w_14_reg[10]  ( .D(n5370), .CP(clk), .Q(reg_w_14[10]) );
  dff_sg \reg_ww_14_reg[10]  ( .D(n5259), .CP(clk), .Q(reg_ww_14[10]) );
  dff_sg \reg_www_14_reg[10]  ( .D(n5239), .CP(clk), .Q(reg_www_14[10]) );
  dff_sg \reg_w_14_reg[9]  ( .D(n5371), .CP(clk), .Q(reg_w_14[9]) );
  dff_sg \reg_ww_14_reg[9]  ( .D(n5260), .CP(clk), .Q(reg_ww_14[9]) );
  dff_sg \reg_www_14_reg[9]  ( .D(n5240), .CP(clk), .Q(reg_www_14[9]) );
  dff_sg \reg_w_14_reg[8]  ( .D(n5372), .CP(clk), .Q(reg_w_14[8]) );
  dff_sg \reg_ww_14_reg[8]  ( .D(n5261), .CP(clk), .Q(reg_ww_14[8]) );
  dff_sg \reg_www_14_reg[8]  ( .D(n5241), .CP(clk), .Q(reg_www_14[8]) );
  dff_sg \reg_w_14_reg[7]  ( .D(n5373), .CP(clk), .Q(reg_w_14[7]) );
  dff_sg \reg_ww_14_reg[7]  ( .D(n5262), .CP(clk), .Q(reg_ww_14[7]) );
  dff_sg \reg_www_14_reg[7]  ( .D(n5242), .CP(clk), .Q(reg_www_14[7]) );
  dff_sg \reg_w_14_reg[6]  ( .D(n5374), .CP(clk), .Q(reg_w_14[6]) );
  dff_sg \reg_ww_14_reg[6]  ( .D(n5263), .CP(clk), .Q(reg_ww_14[6]) );
  dff_sg \reg_www_14_reg[6]  ( .D(n5243), .CP(clk), .Q(reg_www_14[6]) );
  dff_sg \reg_w_14_reg[5]  ( .D(n5375), .CP(clk), .Q(reg_w_14[5]) );
  dff_sg \reg_ww_14_reg[5]  ( .D(n5264), .CP(clk), .Q(reg_ww_14[5]) );
  dff_sg \reg_www_14_reg[5]  ( .D(n5244), .CP(clk), .Q(reg_www_14[5]) );
  dff_sg \reg_w_14_reg[4]  ( .D(n5376), .CP(clk), .Q(reg_w_14[4]) );
  dff_sg \reg_ww_14_reg[4]  ( .D(n5265), .CP(clk), .Q(reg_ww_14[4]) );
  dff_sg \reg_www_14_reg[4]  ( .D(n5245), .CP(clk), .Q(reg_www_14[4]) );
  dff_sg \reg_w_14_reg[3]  ( .D(n5377), .CP(clk), .Q(reg_w_14[3]) );
  dff_sg \reg_ww_14_reg[3]  ( .D(n5266), .CP(clk), .Q(reg_ww_14[3]) );
  dff_sg \reg_www_14_reg[3]  ( .D(n5246), .CP(clk), .Q(reg_www_14[3]) );
  dff_sg \reg_w_14_reg[2]  ( .D(n5378), .CP(clk), .Q(reg_w_14[2]) );
  dff_sg \reg_ww_14_reg[2]  ( .D(n5267), .CP(clk), .Q(reg_ww_14[2]) );
  dff_sg \reg_www_14_reg[2]  ( .D(n5247), .CP(clk), .Q(reg_www_14[2]) );
  dff_sg \reg_w_14_reg[1]  ( .D(n5379), .CP(clk), .Q(reg_w_14[1]) );
  dff_sg \reg_ww_14_reg[1]  ( .D(n5268), .CP(clk), .Q(reg_ww_14[1]) );
  dff_sg \reg_www_14_reg[1]  ( .D(n5248), .CP(clk), .Q(reg_www_14[1]) );
  dff_sg \reg_w_14_reg[0]  ( .D(n5380), .CP(clk), .Q(reg_w_14[0]) );
  dff_sg \reg_ww_14_reg[0]  ( .D(n5269), .CP(clk), .Q(reg_ww_14[0]) );
  dff_sg \reg_www_14_reg[0]  ( .D(n5249), .CP(clk), .Q(reg_www_14[0]) );
  dff_sg \reg_w_13_reg[19]  ( .D(n5381), .CP(clk), .Q(reg_w_13[19]) );
  dff_sg \reg_ww_13_reg[19]  ( .D(n5270), .CP(clk), .Q(reg_ww_13[19]) );
  dff_sg \reg_www_13_reg[19]  ( .D(n4991), .CP(clk), .Q(reg_www_13[19]) );
  dff_sg \reg_w_13_reg[18]  ( .D(n5382), .CP(clk), .Q(reg_w_13[18]) );
  dff_sg \reg_ww_13_reg[18]  ( .D(n5271), .CP(clk), .Q(reg_ww_13[18]) );
  dff_sg \reg_www_13_reg[18]  ( .D(n4992), .CP(clk), .Q(reg_www_13[18]) );
  dff_sg \reg_w_13_reg[17]  ( .D(n5383), .CP(clk), .Q(reg_w_13[17]) );
  dff_sg \reg_ww_13_reg[17]  ( .D(n5272), .CP(clk), .Q(reg_ww_13[17]) );
  dff_sg \reg_www_13_reg[17]  ( .D(n4993), .CP(clk), .Q(reg_www_13[17]) );
  dff_sg \reg_w_13_reg[16]  ( .D(n5384), .CP(clk), .Q(reg_w_13[16]) );
  dff_sg \reg_ww_13_reg[16]  ( .D(n5273), .CP(clk), .Q(reg_ww_13[16]) );
  dff_sg \reg_www_13_reg[16]  ( .D(n4994), .CP(clk), .Q(reg_www_13[16]) );
  dff_sg \reg_w_13_reg[15]  ( .D(n5385), .CP(clk), .Q(reg_w_13[15]) );
  dff_sg \reg_ww_13_reg[15]  ( .D(n5274), .CP(clk), .Q(reg_ww_13[15]) );
  dff_sg \reg_www_13_reg[15]  ( .D(n4995), .CP(clk), .Q(reg_www_13[15]) );
  dff_sg \reg_w_13_reg[14]  ( .D(n5386), .CP(clk), .Q(reg_w_13[14]) );
  dff_sg \reg_ww_13_reg[14]  ( .D(n5275), .CP(clk), .Q(reg_ww_13[14]) );
  dff_sg \reg_www_13_reg[14]  ( .D(n4996), .CP(clk), .Q(reg_www_13[14]) );
  dff_sg \reg_w_13_reg[13]  ( .D(n5387), .CP(clk), .Q(reg_w_13[13]) );
  dff_sg \reg_ww_13_reg[13]  ( .D(n5011), .CP(clk), .Q(reg_ww_13[13]) );
  dff_sg \reg_www_13_reg[13]  ( .D(n4997), .CP(clk), .Q(reg_www_13[13]) );
  dff_sg \reg_w_13_reg[12]  ( .D(n5388), .CP(clk), .Q(reg_w_13[12]) );
  dff_sg \reg_ww_13_reg[12]  ( .D(n5012), .CP(clk), .Q(reg_ww_13[12]) );
  dff_sg \reg_www_13_reg[12]  ( .D(n4998), .CP(clk), .Q(reg_www_13[12]) );
  dff_sg \reg_w_13_reg[11]  ( .D(n5389), .CP(clk), .Q(reg_w_13[11]) );
  dff_sg \reg_ww_13_reg[11]  ( .D(n5013), .CP(clk), .Q(reg_ww_13[11]) );
  dff_sg \reg_www_13_reg[11]  ( .D(n4999), .CP(clk), .Q(reg_www_13[11]) );
  dff_sg \reg_w_13_reg[10]  ( .D(n5390), .CP(clk), .Q(reg_w_13[10]) );
  dff_sg \reg_ww_13_reg[10]  ( .D(n5014), .CP(clk), .Q(reg_ww_13[10]) );
  dff_sg \reg_www_13_reg[10]  ( .D(n5000), .CP(clk), .Q(reg_www_13[10]) );
  dff_sg \reg_w_13_reg[9]  ( .D(n5391), .CP(clk), .Q(reg_w_13[9]) );
  dff_sg \reg_ww_13_reg[9]  ( .D(n5015), .CP(clk), .Q(reg_ww_13[9]) );
  dff_sg \reg_www_13_reg[9]  ( .D(n5001), .CP(clk), .Q(reg_www_13[9]) );
  dff_sg \reg_w_13_reg[8]  ( .D(n5392), .CP(clk), .Q(reg_w_13[8]) );
  dff_sg \reg_ww_13_reg[8]  ( .D(n5016), .CP(clk), .Q(reg_ww_13[8]) );
  dff_sg \reg_www_13_reg[8]  ( .D(n5002), .CP(clk), .Q(reg_www_13[8]) );
  dff_sg \reg_w_13_reg[7]  ( .D(n5393), .CP(clk), .Q(reg_w_13[7]) );
  dff_sg \reg_ww_13_reg[7]  ( .D(n5017), .CP(clk), .Q(reg_ww_13[7]) );
  dff_sg \reg_www_13_reg[7]  ( .D(n5003), .CP(clk), .Q(reg_www_13[7]) );
  dff_sg \reg_w_13_reg[6]  ( .D(n5394), .CP(clk), .Q(reg_w_13[6]) );
  dff_sg \reg_ww_13_reg[6]  ( .D(n5018), .CP(clk), .Q(reg_ww_13[6]) );
  dff_sg \reg_www_13_reg[6]  ( .D(n5004), .CP(clk), .Q(reg_www_13[6]) );
  dff_sg \reg_w_13_reg[5]  ( .D(n5395), .CP(clk), .Q(reg_w_13[5]) );
  dff_sg \reg_ww_13_reg[5]  ( .D(n5019), .CP(clk), .Q(reg_ww_13[5]) );
  dff_sg \reg_www_13_reg[5]  ( .D(n5005), .CP(clk), .Q(reg_www_13[5]) );
  dff_sg \reg_w_13_reg[4]  ( .D(n5396), .CP(clk), .Q(reg_w_13[4]) );
  dff_sg \reg_ww_13_reg[4]  ( .D(n5020), .CP(clk), .Q(reg_ww_13[4]) );
  dff_sg \reg_www_13_reg[4]  ( .D(n5006), .CP(clk), .Q(reg_www_13[4]) );
  dff_sg \reg_w_13_reg[3]  ( .D(n5397), .CP(clk), .Q(reg_w_13[3]) );
  dff_sg \reg_ww_13_reg[3]  ( .D(n5021), .CP(clk), .Q(reg_ww_13[3]) );
  dff_sg \reg_www_13_reg[3]  ( .D(n5007), .CP(clk), .Q(reg_www_13[3]) );
  dff_sg \reg_w_13_reg[2]  ( .D(n5398), .CP(clk), .Q(reg_w_13[2]) );
  dff_sg \reg_ww_13_reg[2]  ( .D(n5022), .CP(clk), .Q(reg_ww_13[2]) );
  dff_sg \reg_www_13_reg[2]  ( .D(n5008), .CP(clk), .Q(reg_www_13[2]) );
  dff_sg \reg_w_13_reg[1]  ( .D(n5399), .CP(clk), .Q(reg_w_13[1]) );
  dff_sg \reg_ww_13_reg[1]  ( .D(n5023), .CP(clk), .Q(reg_ww_13[1]) );
  dff_sg \reg_www_13_reg[1]  ( .D(n5009), .CP(clk), .Q(reg_www_13[1]) );
  dff_sg \reg_w_13_reg[0]  ( .D(n5400), .CP(clk), .Q(reg_w_13[0]) );
  dff_sg \reg_ww_13_reg[0]  ( .D(n5024), .CP(clk), .Q(reg_ww_13[0]) );
  dff_sg \reg_www_13_reg[0]  ( .D(n5010), .CP(clk), .Q(reg_www_13[0]) );
  dff_sg \reg_w_12_reg[19]  ( .D(n5401), .CP(clk), .Q(reg_w_12[19]) );
  dff_sg \reg_ww_12_reg[19]  ( .D(n5045), .CP(clk), .Q(reg_ww_12[19]) );
  dff_sg \reg_www_12_reg[19]  ( .D(n5025), .CP(clk), .Q(reg_www_12[19]) );
  dff_sg \reg_w_12_reg[18]  ( .D(n5402), .CP(clk), .Q(reg_w_12[18]) );
  dff_sg \reg_ww_12_reg[18]  ( .D(n5046), .CP(clk), .Q(reg_ww_12[18]) );
  dff_sg \reg_www_12_reg[18]  ( .D(n5026), .CP(clk), .Q(reg_www_12[18]) );
  dff_sg \reg_w_12_reg[17]  ( .D(n5403), .CP(clk), .Q(reg_w_12[17]) );
  dff_sg \reg_ww_12_reg[17]  ( .D(n5047), .CP(clk), .Q(reg_ww_12[17]) );
  dff_sg \reg_www_12_reg[17]  ( .D(n5027), .CP(clk), .Q(reg_www_12[17]) );
  dff_sg \reg_w_12_reg[16]  ( .D(n5404), .CP(clk), .Q(reg_w_12[16]) );
  dff_sg \reg_ww_12_reg[16]  ( .D(n5048), .CP(clk), .Q(reg_ww_12[16]) );
  dff_sg \reg_www_12_reg[16]  ( .D(n5028), .CP(clk), .Q(reg_www_12[16]) );
  dff_sg \reg_w_12_reg[15]  ( .D(n5405), .CP(clk), .Q(reg_w_12[15]) );
  dff_sg \reg_ww_12_reg[15]  ( .D(n5049), .CP(clk), .Q(reg_ww_12[15]) );
  dff_sg \reg_www_12_reg[15]  ( .D(n5029), .CP(clk), .Q(reg_www_12[15]) );
  dff_sg \reg_w_12_reg[14]  ( .D(n5406), .CP(clk), .Q(reg_w_12[14]) );
  dff_sg \reg_ww_12_reg[14]  ( .D(n5050), .CP(clk), .Q(reg_ww_12[14]) );
  dff_sg \reg_www_12_reg[14]  ( .D(n5030), .CP(clk), .Q(reg_www_12[14]) );
  dff_sg \reg_w_12_reg[13]  ( .D(n5407), .CP(clk), .Q(reg_w_12[13]) );
  dff_sg \reg_ww_12_reg[13]  ( .D(n5051), .CP(clk), .Q(reg_ww_12[13]) );
  dff_sg \reg_www_12_reg[13]  ( .D(n5031), .CP(clk), .Q(reg_www_12[13]) );
  dff_sg \reg_w_12_reg[12]  ( .D(n5408), .CP(clk), .Q(reg_w_12[12]) );
  dff_sg \reg_ww_12_reg[12]  ( .D(n5052), .CP(clk), .Q(reg_ww_12[12]) );
  dff_sg \reg_www_12_reg[12]  ( .D(n5032), .CP(clk), .Q(reg_www_12[12]) );
  dff_sg \reg_w_12_reg[11]  ( .D(n5409), .CP(clk), .Q(reg_w_12[11]) );
  dff_sg \reg_ww_12_reg[11]  ( .D(n5053), .CP(clk), .Q(reg_ww_12[11]) );
  dff_sg \reg_www_12_reg[11]  ( .D(n5033), .CP(clk), .Q(reg_www_12[11]) );
  dff_sg \reg_w_12_reg[10]  ( .D(n5410), .CP(clk), .Q(reg_w_12[10]) );
  dff_sg \reg_ww_12_reg[10]  ( .D(n5054), .CP(clk), .Q(reg_ww_12[10]) );
  dff_sg \reg_www_12_reg[10]  ( .D(n5034), .CP(clk), .Q(reg_www_12[10]) );
  dff_sg \reg_w_12_reg[9]  ( .D(n5411), .CP(clk), .Q(reg_w_12[9]) );
  dff_sg \reg_ww_12_reg[9]  ( .D(n5055), .CP(clk), .Q(reg_ww_12[9]) );
  dff_sg \reg_www_12_reg[9]  ( .D(n5035), .CP(clk), .Q(reg_www_12[9]) );
  dff_sg \reg_w_12_reg[8]  ( .D(n5412), .CP(clk), .Q(reg_w_12[8]) );
  dff_sg \reg_ww_12_reg[8]  ( .D(n5056), .CP(clk), .Q(reg_ww_12[8]) );
  dff_sg \reg_www_12_reg[8]  ( .D(n5036), .CP(clk), .Q(reg_www_12[8]) );
  dff_sg \reg_w_12_reg[7]  ( .D(n5413), .CP(clk), .Q(reg_w_12[7]) );
  dff_sg \reg_ww_12_reg[7]  ( .D(n5057), .CP(clk), .Q(reg_ww_12[7]) );
  dff_sg \reg_www_12_reg[7]  ( .D(n5037), .CP(clk), .Q(reg_www_12[7]) );
  dff_sg \reg_w_12_reg[6]  ( .D(n5414), .CP(clk), .Q(reg_w_12[6]) );
  dff_sg \reg_ww_12_reg[6]  ( .D(n5058), .CP(clk), .Q(reg_ww_12[6]) );
  dff_sg \reg_www_12_reg[6]  ( .D(n5038), .CP(clk), .Q(reg_www_12[6]) );
  dff_sg \reg_w_12_reg[5]  ( .D(n5415), .CP(clk), .Q(reg_w_12[5]) );
  dff_sg \reg_ww_12_reg[5]  ( .D(n5059), .CP(clk), .Q(reg_ww_12[5]) );
  dff_sg \reg_www_12_reg[5]  ( .D(n5039), .CP(clk), .Q(reg_www_12[5]) );
  dff_sg \reg_w_12_reg[4]  ( .D(n5416), .CP(clk), .Q(reg_w_12[4]) );
  dff_sg \reg_ww_12_reg[4]  ( .D(n5060), .CP(clk), .Q(reg_ww_12[4]) );
  dff_sg \reg_www_12_reg[4]  ( .D(n5040), .CP(clk), .Q(reg_www_12[4]) );
  dff_sg \reg_w_12_reg[3]  ( .D(n5417), .CP(clk), .Q(reg_w_12[3]) );
  dff_sg \reg_ww_12_reg[3]  ( .D(n5061), .CP(clk), .Q(reg_ww_12[3]) );
  dff_sg \reg_www_12_reg[3]  ( .D(n5041), .CP(clk), .Q(reg_www_12[3]) );
  dff_sg \reg_w_12_reg[2]  ( .D(n5418), .CP(clk), .Q(reg_w_12[2]) );
  dff_sg \reg_ww_12_reg[2]  ( .D(n5062), .CP(clk), .Q(reg_ww_12[2]) );
  dff_sg \reg_www_12_reg[2]  ( .D(n5042), .CP(clk), .Q(reg_www_12[2]) );
  dff_sg \reg_w_12_reg[1]  ( .D(n5419), .CP(clk), .Q(reg_w_12[1]) );
  dff_sg \reg_ww_12_reg[1]  ( .D(n5063), .CP(clk), .Q(reg_ww_12[1]) );
  dff_sg \reg_www_12_reg[1]  ( .D(n5043), .CP(clk), .Q(reg_www_12[1]) );
  dff_sg \reg_w_12_reg[0]  ( .D(n5420), .CP(clk), .Q(reg_w_12[0]) );
  dff_sg \reg_ww_12_reg[0]  ( .D(n5064), .CP(clk), .Q(reg_ww_12[0]) );
  dff_sg \reg_www_12_reg[0]  ( .D(n5044), .CP(clk), .Q(reg_www_12[0]) );
  dff_sg \reg_w_11_reg[19]  ( .D(n5421), .CP(clk), .Q(reg_w_11[19]) );
  dff_sg \reg_ww_11_reg[19]  ( .D(n5085), .CP(clk), .Q(reg_ww_11[19]) );
  dff_sg \reg_www_11_reg[19]  ( .D(n5065), .CP(clk), .Q(reg_www_11[19]) );
  dff_sg \reg_w_11_reg[18]  ( .D(n5422), .CP(clk), .Q(reg_w_11[18]) );
  dff_sg \reg_ww_11_reg[18]  ( .D(n5086), .CP(clk), .Q(reg_ww_11[18]) );
  dff_sg \reg_www_11_reg[18]  ( .D(n5066), .CP(clk), .Q(reg_www_11[18]) );
  dff_sg \reg_w_11_reg[17]  ( .D(n5423), .CP(clk), .Q(reg_w_11[17]) );
  dff_sg \reg_ww_11_reg[17]  ( .D(n5087), .CP(clk), .Q(reg_ww_11[17]) );
  dff_sg \reg_www_11_reg[17]  ( .D(n5067), .CP(clk), .Q(reg_www_11[17]) );
  dff_sg \reg_w_11_reg[16]  ( .D(n5424), .CP(clk), .Q(reg_w_11[16]) );
  dff_sg \reg_ww_11_reg[16]  ( .D(n5088), .CP(clk), .Q(reg_ww_11[16]) );
  dff_sg \reg_www_11_reg[16]  ( .D(n5068), .CP(clk), .Q(reg_www_11[16]) );
  dff_sg \reg_w_11_reg[15]  ( .D(n5425), .CP(clk), .Q(reg_w_11[15]) );
  dff_sg \reg_ww_11_reg[15]  ( .D(n5089), .CP(clk), .Q(reg_ww_11[15]) );
  dff_sg \reg_www_11_reg[15]  ( .D(n5069), .CP(clk), .Q(reg_www_11[15]) );
  dff_sg \reg_w_11_reg[14]  ( .D(n5426), .CP(clk), .Q(reg_w_11[14]) );
  dff_sg \reg_ww_11_reg[14]  ( .D(n5090), .CP(clk), .Q(reg_ww_11[14]) );
  dff_sg \reg_www_11_reg[14]  ( .D(n5070), .CP(clk), .Q(reg_www_11[14]) );
  dff_sg \reg_w_11_reg[13]  ( .D(n5427), .CP(clk), .Q(reg_w_11[13]) );
  dff_sg \reg_ww_11_reg[13]  ( .D(n5091), .CP(clk), .Q(reg_ww_11[13]) );
  dff_sg \reg_www_11_reg[13]  ( .D(n5071), .CP(clk), .Q(reg_www_11[13]) );
  dff_sg \reg_w_11_reg[12]  ( .D(n5428), .CP(clk), .Q(reg_w_11[12]) );
  dff_sg \reg_ww_11_reg[12]  ( .D(n5092), .CP(clk), .Q(reg_ww_11[12]) );
  dff_sg \reg_www_11_reg[12]  ( .D(n5072), .CP(clk), .Q(reg_www_11[12]) );
  dff_sg \reg_w_11_reg[11]  ( .D(n5429), .CP(clk), .Q(reg_w_11[11]) );
  dff_sg \reg_ww_11_reg[11]  ( .D(n5093), .CP(clk), .Q(reg_ww_11[11]) );
  dff_sg \reg_www_11_reg[11]  ( .D(n5073), .CP(clk), .Q(reg_www_11[11]) );
  dff_sg \reg_w_11_reg[10]  ( .D(n5430), .CP(clk), .Q(reg_w_11[10]) );
  dff_sg \reg_ww_11_reg[10]  ( .D(n5094), .CP(clk), .Q(reg_ww_11[10]) );
  dff_sg \reg_www_11_reg[10]  ( .D(n5074), .CP(clk), .Q(reg_www_11[10]) );
  dff_sg \reg_w_11_reg[9]  ( .D(n5431), .CP(clk), .Q(reg_w_11[9]) );
  dff_sg \reg_ww_11_reg[9]  ( .D(n5095), .CP(clk), .Q(reg_ww_11[9]) );
  dff_sg \reg_www_11_reg[9]  ( .D(n5075), .CP(clk), .Q(reg_www_11[9]) );
  dff_sg \reg_w_11_reg[8]  ( .D(n5432), .CP(clk), .Q(reg_w_11[8]) );
  dff_sg \reg_ww_11_reg[8]  ( .D(n5096), .CP(clk), .Q(reg_ww_11[8]) );
  dff_sg \reg_www_11_reg[8]  ( .D(n5076), .CP(clk), .Q(reg_www_11[8]) );
  dff_sg \reg_w_11_reg[7]  ( .D(n5433), .CP(clk), .Q(reg_w_11[7]) );
  dff_sg \reg_ww_11_reg[7]  ( .D(n5097), .CP(clk), .Q(reg_ww_11[7]) );
  dff_sg \reg_www_11_reg[7]  ( .D(n5077), .CP(clk), .Q(reg_www_11[7]) );
  dff_sg \reg_w_11_reg[6]  ( .D(n5434), .CP(clk), .Q(reg_w_11[6]) );
  dff_sg \reg_ww_11_reg[6]  ( .D(n5098), .CP(clk), .Q(reg_ww_11[6]) );
  dff_sg \reg_www_11_reg[6]  ( .D(n5078), .CP(clk), .Q(reg_www_11[6]) );
  dff_sg \reg_w_11_reg[5]  ( .D(n5435), .CP(clk), .Q(reg_w_11[5]) );
  dff_sg \reg_ww_11_reg[5]  ( .D(n5099), .CP(clk), .Q(reg_ww_11[5]) );
  dff_sg \reg_www_11_reg[5]  ( .D(n5079), .CP(clk), .Q(reg_www_11[5]) );
  dff_sg \reg_w_11_reg[4]  ( .D(n5436), .CP(clk), .Q(reg_w_11[4]) );
  dff_sg \reg_ww_11_reg[4]  ( .D(n5100), .CP(clk), .Q(reg_ww_11[4]) );
  dff_sg \reg_www_11_reg[4]  ( .D(n5080), .CP(clk), .Q(reg_www_11[4]) );
  dff_sg \reg_w_11_reg[3]  ( .D(n5437), .CP(clk), .Q(reg_w_11[3]) );
  dff_sg \reg_ww_11_reg[3]  ( .D(n5101), .CP(clk), .Q(reg_ww_11[3]) );
  dff_sg \reg_www_11_reg[3]  ( .D(n5081), .CP(clk), .Q(reg_www_11[3]) );
  dff_sg \reg_w_11_reg[2]  ( .D(n5438), .CP(clk), .Q(reg_w_11[2]) );
  dff_sg \reg_ww_11_reg[2]  ( .D(n5102), .CP(clk), .Q(reg_ww_11[2]) );
  dff_sg \reg_www_11_reg[2]  ( .D(n5082), .CP(clk), .Q(reg_www_11[2]) );
  dff_sg \reg_w_11_reg[1]  ( .D(n5439), .CP(clk), .Q(reg_w_11[1]) );
  dff_sg \reg_ww_11_reg[1]  ( .D(n5103), .CP(clk), .Q(reg_ww_11[1]) );
  dff_sg \reg_www_11_reg[1]  ( .D(n5083), .CP(clk), .Q(reg_www_11[1]) );
  dff_sg \reg_w_11_reg[0]  ( .D(n5440), .CP(clk), .Q(reg_w_11[0]) );
  dff_sg \reg_ww_11_reg[0]  ( .D(n5104), .CP(clk), .Q(reg_ww_11[0]) );
  dff_sg \reg_www_11_reg[0]  ( .D(n5084), .CP(clk), .Q(reg_www_11[0]) );
  dff_sg \reg_w_10_reg[19]  ( .D(n5441), .CP(clk), .Q(reg_w_10[19]) );
  dff_sg \reg_ww_10_reg[19]  ( .D(n5125), .CP(clk), .Q(reg_ww_10[19]) );
  dff_sg \reg_www_10_reg[19]  ( .D(n5105), .CP(clk), .Q(reg_www_10[19]) );
  dff_sg \reg_w_10_reg[18]  ( .D(n5442), .CP(clk), .Q(reg_w_10[18]) );
  dff_sg \reg_ww_10_reg[18]  ( .D(n5126), .CP(clk), .Q(reg_ww_10[18]) );
  dff_sg \reg_www_10_reg[18]  ( .D(n5106), .CP(clk), .Q(reg_www_10[18]) );
  dff_sg \reg_w_10_reg[17]  ( .D(n5443), .CP(clk), .Q(reg_w_10[17]) );
  dff_sg \reg_ww_10_reg[17]  ( .D(n5127), .CP(clk), .Q(reg_ww_10[17]) );
  dff_sg \reg_www_10_reg[17]  ( .D(n5107), .CP(clk), .Q(reg_www_10[17]) );
  dff_sg \reg_w_10_reg[16]  ( .D(n5444), .CP(clk), .Q(reg_w_10[16]) );
  dff_sg \reg_ww_10_reg[16]  ( .D(n5128), .CP(clk), .Q(reg_ww_10[16]) );
  dff_sg \reg_www_10_reg[16]  ( .D(n5108), .CP(clk), .Q(reg_www_10[16]) );
  dff_sg \reg_w_10_reg[15]  ( .D(n5445), .CP(clk), .Q(reg_w_10[15]) );
  dff_sg \reg_ww_10_reg[15]  ( .D(n5129), .CP(clk), .Q(reg_ww_10[15]) );
  dff_sg \reg_www_10_reg[15]  ( .D(n5109), .CP(clk), .Q(reg_www_10[15]) );
  dff_sg \reg_w_10_reg[14]  ( .D(n5446), .CP(clk), .Q(reg_w_10[14]) );
  dff_sg \reg_ww_10_reg[14]  ( .D(n5130), .CP(clk), .Q(reg_ww_10[14]) );
  dff_sg \reg_www_10_reg[14]  ( .D(n5110), .CP(clk), .Q(reg_www_10[14]) );
  dff_sg \reg_w_10_reg[13]  ( .D(n5447), .CP(clk), .Q(reg_w_10[13]) );
  dff_sg \reg_ww_10_reg[13]  ( .D(n5131), .CP(clk), .Q(reg_ww_10[13]) );
  dff_sg \reg_www_10_reg[13]  ( .D(n5111), .CP(clk), .Q(reg_www_10[13]) );
  dff_sg \reg_w_10_reg[12]  ( .D(n5448), .CP(clk), .Q(reg_w_10[12]) );
  dff_sg \reg_ww_10_reg[12]  ( .D(n5132), .CP(clk), .Q(reg_ww_10[12]) );
  dff_sg \reg_www_10_reg[12]  ( .D(n5112), .CP(clk), .Q(reg_www_10[12]) );
  dff_sg \reg_w_10_reg[11]  ( .D(n5449), .CP(clk), .Q(reg_w_10[11]) );
  dff_sg \reg_ww_10_reg[11]  ( .D(n5133), .CP(clk), .Q(reg_ww_10[11]) );
  dff_sg \reg_www_10_reg[11]  ( .D(n5113), .CP(clk), .Q(reg_www_10[11]) );
  dff_sg \reg_w_10_reg[10]  ( .D(n5450), .CP(clk), .Q(reg_w_10[10]) );
  dff_sg \reg_ww_10_reg[10]  ( .D(n5134), .CP(clk), .Q(reg_ww_10[10]) );
  dff_sg \reg_www_10_reg[10]  ( .D(n5114), .CP(clk), .Q(reg_www_10[10]) );
  dff_sg \reg_w_10_reg[9]  ( .D(n5451), .CP(clk), .Q(reg_w_10[9]) );
  dff_sg \reg_ww_10_reg[9]  ( .D(n5135), .CP(clk), .Q(reg_ww_10[9]) );
  dff_sg \reg_www_10_reg[9]  ( .D(n5115), .CP(clk), .Q(reg_www_10[9]) );
  dff_sg \reg_w_10_reg[8]  ( .D(n5452), .CP(clk), .Q(reg_w_10[8]) );
  dff_sg \reg_ww_10_reg[8]  ( .D(n5136), .CP(clk), .Q(reg_ww_10[8]) );
  dff_sg \reg_www_10_reg[8]  ( .D(n5116), .CP(clk), .Q(reg_www_10[8]) );
  dff_sg \reg_w_10_reg[7]  ( .D(n5453), .CP(clk), .Q(reg_w_10[7]) );
  dff_sg \reg_ww_10_reg[7]  ( .D(n5137), .CP(clk), .Q(reg_ww_10[7]) );
  dff_sg \reg_www_10_reg[7]  ( .D(n5117), .CP(clk), .Q(reg_www_10[7]) );
  dff_sg \reg_w_10_reg[6]  ( .D(n5454), .CP(clk), .Q(reg_w_10[6]) );
  dff_sg \reg_ww_10_reg[6]  ( .D(n5138), .CP(clk), .Q(reg_ww_10[6]) );
  dff_sg \reg_www_10_reg[6]  ( .D(n5118), .CP(clk), .Q(reg_www_10[6]) );
  dff_sg \reg_w_10_reg[5]  ( .D(n5455), .CP(clk), .Q(reg_w_10[5]) );
  dff_sg \reg_ww_10_reg[5]  ( .D(n5139), .CP(clk), .Q(reg_ww_10[5]) );
  dff_sg \reg_www_10_reg[5]  ( .D(n5119), .CP(clk), .Q(reg_www_10[5]) );
  dff_sg \reg_w_10_reg[4]  ( .D(n5456), .CP(clk), .Q(reg_w_10[4]) );
  dff_sg \reg_ww_10_reg[4]  ( .D(n5140), .CP(clk), .Q(reg_ww_10[4]) );
  dff_sg \reg_www_10_reg[4]  ( .D(n5120), .CP(clk), .Q(reg_www_10[4]) );
  dff_sg \reg_w_10_reg[3]  ( .D(n5457), .CP(clk), .Q(reg_w_10[3]) );
  dff_sg \reg_ww_10_reg[3]  ( .D(n5141), .CP(clk), .Q(reg_ww_10[3]) );
  dff_sg \reg_www_10_reg[3]  ( .D(n5121), .CP(clk), .Q(reg_www_10[3]) );
  dff_sg \reg_w_10_reg[2]  ( .D(n5458), .CP(clk), .Q(reg_w_10[2]) );
  dff_sg \reg_ww_10_reg[2]  ( .D(n5142), .CP(clk), .Q(reg_ww_10[2]) );
  dff_sg \reg_www_10_reg[2]  ( .D(n5122), .CP(clk), .Q(reg_www_10[2]) );
  dff_sg \reg_w_10_reg[1]  ( .D(n5459), .CP(clk), .Q(reg_w_10[1]) );
  dff_sg \reg_ww_10_reg[1]  ( .D(n5143), .CP(clk), .Q(reg_ww_10[1]) );
  dff_sg \reg_www_10_reg[1]  ( .D(n5123), .CP(clk), .Q(reg_www_10[1]) );
  dff_sg \reg_w_10_reg[0]  ( .D(n5460), .CP(clk), .Q(reg_w_10[0]) );
  dff_sg \reg_ww_10_reg[0]  ( .D(n5144), .CP(clk), .Q(reg_ww_10[0]) );
  dff_sg \reg_www_10_reg[0]  ( .D(n5124), .CP(clk), .Q(reg_www_10[0]) );
  dff_sg \reg_w_9_reg[19]  ( .D(n5461), .CP(clk), .Q(reg_w_9[19]) );
  dff_sg \reg_ww_9_reg[19]  ( .D(n5165), .CP(clk), .Q(reg_ww_9[19]) );
  dff_sg \reg_www_9_reg[19]  ( .D(n5145), .CP(clk), .Q(reg_www_9[19]) );
  dff_sg \reg_w_9_reg[18]  ( .D(n5462), .CP(clk), .Q(reg_w_9[18]) );
  dff_sg \reg_ww_9_reg[18]  ( .D(n5166), .CP(clk), .Q(reg_ww_9[18]) );
  dff_sg \reg_www_9_reg[18]  ( .D(n5146), .CP(clk), .Q(reg_www_9[18]) );
  dff_sg \reg_w_9_reg[17]  ( .D(n5463), .CP(clk), .Q(reg_w_9[17]) );
  dff_sg \reg_ww_9_reg[17]  ( .D(n5167), .CP(clk), .Q(reg_ww_9[17]) );
  dff_sg \reg_www_9_reg[17]  ( .D(n5147), .CP(clk), .Q(reg_www_9[17]) );
  dff_sg \reg_w_9_reg[16]  ( .D(n5464), .CP(clk), .Q(reg_w_9[16]) );
  dff_sg \reg_ww_9_reg[16]  ( .D(n5168), .CP(clk), .Q(reg_ww_9[16]) );
  dff_sg \reg_www_9_reg[16]  ( .D(n5148), .CP(clk), .Q(reg_www_9[16]) );
  dff_sg \reg_w_9_reg[15]  ( .D(n5465), .CP(clk), .Q(reg_w_9[15]) );
  dff_sg \reg_ww_9_reg[15]  ( .D(n5169), .CP(clk), .Q(reg_ww_9[15]) );
  dff_sg \reg_www_9_reg[15]  ( .D(n5149), .CP(clk), .Q(reg_www_9[15]) );
  dff_sg \reg_w_9_reg[14]  ( .D(n5466), .CP(clk), .Q(reg_w_9[14]) );
  dff_sg \reg_ww_9_reg[14]  ( .D(n5170), .CP(clk), .Q(reg_ww_9[14]) );
  dff_sg \reg_www_9_reg[14]  ( .D(n5150), .CP(clk), .Q(reg_www_9[14]) );
  dff_sg \reg_w_9_reg[13]  ( .D(n5467), .CP(clk), .Q(reg_w_9[13]) );
  dff_sg \reg_ww_9_reg[13]  ( .D(n5171), .CP(clk), .Q(reg_ww_9[13]) );
  dff_sg \reg_www_9_reg[13]  ( .D(n5151), .CP(clk), .Q(reg_www_9[13]) );
  dff_sg \reg_w_9_reg[12]  ( .D(n5468), .CP(clk), .Q(reg_w_9[12]) );
  dff_sg \reg_ww_9_reg[12]  ( .D(n5172), .CP(clk), .Q(reg_ww_9[12]) );
  dff_sg \reg_www_9_reg[12]  ( .D(n5152), .CP(clk), .Q(reg_www_9[12]) );
  dff_sg \reg_w_9_reg[11]  ( .D(n5469), .CP(clk), .Q(reg_w_9[11]) );
  dff_sg \reg_ww_9_reg[11]  ( .D(n5173), .CP(clk), .Q(reg_ww_9[11]) );
  dff_sg \reg_www_9_reg[11]  ( .D(n5153), .CP(clk), .Q(reg_www_9[11]) );
  dff_sg \reg_w_9_reg[10]  ( .D(n5470), .CP(clk), .Q(reg_w_9[10]) );
  dff_sg \reg_ww_9_reg[10]  ( .D(n5174), .CP(clk), .Q(reg_ww_9[10]) );
  dff_sg \reg_www_9_reg[10]  ( .D(n5154), .CP(clk), .Q(reg_www_9[10]) );
  dff_sg \reg_w_9_reg[9]  ( .D(n5471), .CP(clk), .Q(reg_w_9[9]) );
  dff_sg \reg_ww_9_reg[9]  ( .D(n5175), .CP(clk), .Q(reg_ww_9[9]) );
  dff_sg \reg_www_9_reg[9]  ( .D(n5155), .CP(clk), .Q(reg_www_9[9]) );
  dff_sg \reg_w_9_reg[8]  ( .D(n5472), .CP(clk), .Q(reg_w_9[8]) );
  dff_sg \reg_ww_9_reg[8]  ( .D(n5176), .CP(clk), .Q(reg_ww_9[8]) );
  dff_sg \reg_www_9_reg[8]  ( .D(n5156), .CP(clk), .Q(reg_www_9[8]) );
  dff_sg \reg_w_9_reg[7]  ( .D(n5473), .CP(clk), .Q(reg_w_9[7]) );
  dff_sg \reg_ww_9_reg[7]  ( .D(n5177), .CP(clk), .Q(reg_ww_9[7]) );
  dff_sg \reg_www_9_reg[7]  ( .D(n5157), .CP(clk), .Q(reg_www_9[7]) );
  dff_sg \reg_w_9_reg[6]  ( .D(n5474), .CP(clk), .Q(reg_w_9[6]) );
  dff_sg \reg_ww_9_reg[6]  ( .D(n5178), .CP(clk), .Q(reg_ww_9[6]) );
  dff_sg \reg_www_9_reg[6]  ( .D(n5158), .CP(clk), .Q(reg_www_9[6]) );
  dff_sg \reg_w_9_reg[5]  ( .D(n5475), .CP(clk), .Q(reg_w_9[5]) );
  dff_sg \reg_ww_9_reg[5]  ( .D(n5179), .CP(clk), .Q(reg_ww_9[5]) );
  dff_sg \reg_www_9_reg[5]  ( .D(n5159), .CP(clk), .Q(reg_www_9[5]) );
  dff_sg \reg_w_9_reg[4]  ( .D(n5476), .CP(clk), .Q(reg_w_9[4]) );
  dff_sg \reg_ww_9_reg[4]  ( .D(n5180), .CP(clk), .Q(reg_ww_9[4]) );
  dff_sg \reg_www_9_reg[4]  ( .D(n5160), .CP(clk), .Q(reg_www_9[4]) );
  dff_sg \reg_w_9_reg[3]  ( .D(n5477), .CP(clk), .Q(reg_w_9[3]) );
  dff_sg \reg_ww_9_reg[3]  ( .D(n5181), .CP(clk), .Q(reg_ww_9[3]) );
  dff_sg \reg_www_9_reg[3]  ( .D(n5161), .CP(clk), .Q(reg_www_9[3]) );
  dff_sg \reg_w_9_reg[2]  ( .D(n5478), .CP(clk), .Q(reg_w_9[2]) );
  dff_sg \reg_ww_9_reg[2]  ( .D(n5182), .CP(clk), .Q(reg_ww_9[2]) );
  dff_sg \reg_www_9_reg[2]  ( .D(n5162), .CP(clk), .Q(reg_www_9[2]) );
  dff_sg \reg_w_9_reg[1]  ( .D(n5479), .CP(clk), .Q(reg_w_9[1]) );
  dff_sg \reg_ww_9_reg[1]  ( .D(n5183), .CP(clk), .Q(reg_ww_9[1]) );
  dff_sg \reg_www_9_reg[1]  ( .D(n5163), .CP(clk), .Q(reg_www_9[1]) );
  dff_sg \reg_w_9_reg[0]  ( .D(n5480), .CP(clk), .Q(reg_w_9[0]) );
  dff_sg \reg_ww_9_reg[0]  ( .D(n5184), .CP(clk), .Q(reg_ww_9[0]) );
  dff_sg \reg_www_9_reg[0]  ( .D(n5164), .CP(clk), .Q(reg_www_9[0]) );
  dff_sg \reg_w_8_reg[19]  ( .D(n5481), .CP(clk), .Q(reg_w_8[19]) );
  dff_sg \reg_ww_8_reg[19]  ( .D(n5185), .CP(clk), .Q(reg_ww_8[19]) );
  dff_sg \reg_www_8_reg[19]  ( .D(n4792), .CP(clk), .Q(reg_www_8[19]) );
  dff_sg \reg_w_8_reg[18]  ( .D(n5482), .CP(clk), .Q(reg_w_8[18]) );
  dff_sg \reg_ww_8_reg[18]  ( .D(n5186), .CP(clk), .Q(reg_ww_8[18]) );
  dff_sg \reg_www_8_reg[18]  ( .D(n4793), .CP(clk), .Q(reg_www_8[18]) );
  dff_sg \reg_w_8_reg[17]  ( .D(n5483), .CP(clk), .Q(reg_w_8[17]) );
  dff_sg \reg_ww_8_reg[17]  ( .D(n5187), .CP(clk), .Q(reg_ww_8[17]) );
  dff_sg \reg_www_8_reg[17]  ( .D(n4794), .CP(clk), .Q(reg_www_8[17]) );
  dff_sg \reg_w_8_reg[16]  ( .D(n5484), .CP(clk), .Q(reg_w_8[16]) );
  dff_sg \reg_ww_8_reg[16]  ( .D(n5188), .CP(clk), .Q(reg_ww_8[16]) );
  dff_sg \reg_www_8_reg[16]  ( .D(n4795), .CP(clk), .Q(reg_www_8[16]) );
  dff_sg \reg_w_8_reg[15]  ( .D(n5485), .CP(clk), .Q(reg_w_8[15]) );
  dff_sg \reg_ww_8_reg[15]  ( .D(n5189), .CP(clk), .Q(reg_ww_8[15]) );
  dff_sg \reg_www_8_reg[15]  ( .D(n4796), .CP(clk), .Q(reg_www_8[15]) );
  dff_sg \reg_w_8_reg[14]  ( .D(n5486), .CP(clk), .Q(reg_w_8[14]) );
  dff_sg \reg_ww_8_reg[14]  ( .D(n4812), .CP(clk), .Q(reg_ww_8[14]) );
  dff_sg \reg_www_8_reg[14]  ( .D(n4797), .CP(clk), .Q(reg_www_8[14]) );
  dff_sg \reg_w_8_reg[13]  ( .D(n5487), .CP(clk), .Q(reg_w_8[13]) );
  dff_sg \reg_ww_8_reg[13]  ( .D(n4813), .CP(clk), .Q(reg_ww_8[13]) );
  dff_sg \reg_www_8_reg[13]  ( .D(n4798), .CP(clk), .Q(reg_www_8[13]) );
  dff_sg \reg_w_8_reg[12]  ( .D(n5488), .CP(clk), .Q(reg_w_8[12]) );
  dff_sg \reg_ww_8_reg[12]  ( .D(n4814), .CP(clk), .Q(reg_ww_8[12]) );
  dff_sg \reg_www_8_reg[12]  ( .D(n4799), .CP(clk), .Q(reg_www_8[12]) );
  dff_sg \reg_w_8_reg[11]  ( .D(n5489), .CP(clk), .Q(reg_w_8[11]) );
  dff_sg \reg_ww_8_reg[11]  ( .D(n4815), .CP(clk), .Q(reg_ww_8[11]) );
  dff_sg \reg_www_8_reg[11]  ( .D(n4800), .CP(clk), .Q(reg_www_8[11]) );
  dff_sg \reg_w_8_reg[10]  ( .D(n5490), .CP(clk), .Q(reg_w_8[10]) );
  dff_sg \reg_ww_8_reg[10]  ( .D(n4816), .CP(clk), .Q(reg_ww_8[10]) );
  dff_sg \reg_www_8_reg[10]  ( .D(n4801), .CP(clk), .Q(reg_www_8[10]) );
  dff_sg \reg_w_8_reg[9]  ( .D(n5491), .CP(clk), .Q(reg_w_8[9]) );
  dff_sg \reg_ww_8_reg[9]  ( .D(n4817), .CP(clk), .Q(reg_ww_8[9]) );
  dff_sg \reg_www_8_reg[9]  ( .D(n4802), .CP(clk), .Q(reg_www_8[9]) );
  dff_sg \reg_w_8_reg[8]  ( .D(n5492), .CP(clk), .Q(reg_w_8[8]) );
  dff_sg \reg_ww_8_reg[8]  ( .D(n4818), .CP(clk), .Q(reg_ww_8[8]) );
  dff_sg \reg_www_8_reg[8]  ( .D(n4803), .CP(clk), .Q(reg_www_8[8]) );
  dff_sg \reg_w_8_reg[7]  ( .D(n5493), .CP(clk), .Q(reg_w_8[7]) );
  dff_sg \reg_ww_8_reg[7]  ( .D(n4819), .CP(clk), .Q(reg_ww_8[7]) );
  dff_sg \reg_www_8_reg[7]  ( .D(n4804), .CP(clk), .Q(reg_www_8[7]) );
  dff_sg \reg_w_8_reg[6]  ( .D(n5494), .CP(clk), .Q(reg_w_8[6]) );
  dff_sg \reg_ww_8_reg[6]  ( .D(n4820), .CP(clk), .Q(reg_ww_8[6]) );
  dff_sg \reg_www_8_reg[6]  ( .D(n4805), .CP(clk), .Q(reg_www_8[6]) );
  dff_sg \reg_w_8_reg[5]  ( .D(n5495), .CP(clk), .Q(reg_w_8[5]) );
  dff_sg \reg_ww_8_reg[5]  ( .D(n4821), .CP(clk), .Q(reg_ww_8[5]) );
  dff_sg \reg_www_8_reg[5]  ( .D(n4806), .CP(clk), .Q(reg_www_8[5]) );
  dff_sg \reg_w_8_reg[4]  ( .D(n5496), .CP(clk), .Q(reg_w_8[4]) );
  dff_sg \reg_ww_8_reg[4]  ( .D(n4822), .CP(clk), .Q(reg_ww_8[4]) );
  dff_sg \reg_www_8_reg[4]  ( .D(n4807), .CP(clk), .Q(reg_www_8[4]) );
  dff_sg \reg_w_8_reg[3]  ( .D(n5497), .CP(clk), .Q(reg_w_8[3]) );
  dff_sg \reg_ww_8_reg[3]  ( .D(n4823), .CP(clk), .Q(reg_ww_8[3]) );
  dff_sg \reg_www_8_reg[3]  ( .D(n4808), .CP(clk), .Q(reg_www_8[3]) );
  dff_sg \reg_w_8_reg[2]  ( .D(n5498), .CP(clk), .Q(reg_w_8[2]) );
  dff_sg \reg_ww_8_reg[2]  ( .D(n4824), .CP(clk), .Q(reg_ww_8[2]) );
  dff_sg \reg_www_8_reg[2]  ( .D(n4809), .CP(clk), .Q(reg_www_8[2]) );
  dff_sg \reg_w_8_reg[1]  ( .D(n5499), .CP(clk), .Q(reg_w_8[1]) );
  dff_sg \reg_ww_8_reg[1]  ( .D(n4825), .CP(clk), .Q(reg_ww_8[1]) );
  dff_sg \reg_www_8_reg[1]  ( .D(n4810), .CP(clk), .Q(reg_www_8[1]) );
  dff_sg \reg_w_8_reg[0]  ( .D(n5500), .CP(clk), .Q(reg_w_8[0]) );
  dff_sg \reg_ww_8_reg[0]  ( .D(n4826), .CP(clk), .Q(reg_ww_8[0]) );
  dff_sg \reg_www_8_reg[0]  ( .D(n4811), .CP(clk), .Q(reg_www_8[0]) );
  dff_sg \reg_w_7_reg[19]  ( .D(n5501), .CP(clk), .Q(reg_w_7[19]) );
  dff_sg \reg_ww_7_reg[19]  ( .D(n4847), .CP(clk), .Q(reg_ww_7[19]) );
  dff_sg \reg_www_7_reg[19]  ( .D(n4827), .CP(clk), .Q(reg_www_7[19]) );
  dff_sg \reg_w_7_reg[18]  ( .D(n5502), .CP(clk), .Q(reg_w_7[18]) );
  dff_sg \reg_ww_7_reg[18]  ( .D(n4848), .CP(clk), .Q(reg_ww_7[18]) );
  dff_sg \reg_www_7_reg[18]  ( .D(n4828), .CP(clk), .Q(reg_www_7[18]) );
  dff_sg \reg_w_7_reg[17]  ( .D(n5503), .CP(clk), .Q(reg_w_7[17]) );
  dff_sg \reg_ww_7_reg[17]  ( .D(n4849), .CP(clk), .Q(reg_ww_7[17]) );
  dff_sg \reg_www_7_reg[17]  ( .D(n4829), .CP(clk), .Q(reg_www_7[17]) );
  dff_sg \reg_w_7_reg[16]  ( .D(n5504), .CP(clk), .Q(reg_w_7[16]) );
  dff_sg \reg_ww_7_reg[16]  ( .D(n4850), .CP(clk), .Q(reg_ww_7[16]) );
  dff_sg \reg_www_7_reg[16]  ( .D(n4830), .CP(clk), .Q(reg_www_7[16]) );
  dff_sg \reg_w_7_reg[15]  ( .D(n5505), .CP(clk), .Q(reg_w_7[15]) );
  dff_sg \reg_ww_7_reg[15]  ( .D(n4851), .CP(clk), .Q(reg_ww_7[15]) );
  dff_sg \reg_www_7_reg[15]  ( .D(n4831), .CP(clk), .Q(reg_www_7[15]) );
  dff_sg \reg_w_7_reg[14]  ( .D(n5506), .CP(clk), .Q(reg_w_7[14]) );
  dff_sg \reg_ww_7_reg[14]  ( .D(n4852), .CP(clk), .Q(reg_ww_7[14]) );
  dff_sg \reg_www_7_reg[14]  ( .D(n4832), .CP(clk), .Q(reg_www_7[14]) );
  dff_sg \reg_w_7_reg[13]  ( .D(n5507), .CP(clk), .Q(reg_w_7[13]) );
  dff_sg \reg_ww_7_reg[13]  ( .D(n4853), .CP(clk), .Q(reg_ww_7[13]) );
  dff_sg \reg_www_7_reg[13]  ( .D(n4833), .CP(clk), .Q(reg_www_7[13]) );
  dff_sg \reg_w_7_reg[12]  ( .D(n5508), .CP(clk), .Q(reg_w_7[12]) );
  dff_sg \reg_ww_7_reg[12]  ( .D(n4854), .CP(clk), .Q(reg_ww_7[12]) );
  dff_sg \reg_www_7_reg[12]  ( .D(n4834), .CP(clk), .Q(reg_www_7[12]) );
  dff_sg \reg_w_7_reg[11]  ( .D(n5509), .CP(clk), .Q(reg_w_7[11]) );
  dff_sg \reg_ww_7_reg[11]  ( .D(n4855), .CP(clk), .Q(reg_ww_7[11]) );
  dff_sg \reg_www_7_reg[11]  ( .D(n4835), .CP(clk), .Q(reg_www_7[11]) );
  dff_sg \reg_w_7_reg[10]  ( .D(n5510), .CP(clk), .Q(reg_w_7[10]) );
  dff_sg \reg_ww_7_reg[10]  ( .D(n4856), .CP(clk), .Q(reg_ww_7[10]) );
  dff_sg \reg_www_7_reg[10]  ( .D(n4836), .CP(clk), .Q(reg_www_7[10]) );
  dff_sg \reg_w_7_reg[9]  ( .D(n5511), .CP(clk), .Q(reg_w_7[9]) );
  dff_sg \reg_ww_7_reg[9]  ( .D(n4857), .CP(clk), .Q(reg_ww_7[9]) );
  dff_sg \reg_www_7_reg[9]  ( .D(n4837), .CP(clk), .Q(reg_www_7[9]) );
  dff_sg \reg_w_7_reg[8]  ( .D(n5512), .CP(clk), .Q(reg_w_7[8]) );
  dff_sg \reg_ww_7_reg[8]  ( .D(n4858), .CP(clk), .Q(reg_ww_7[8]) );
  dff_sg \reg_www_7_reg[8]  ( .D(n4838), .CP(clk), .Q(reg_www_7[8]) );
  dff_sg \reg_w_7_reg[7]  ( .D(n5513), .CP(clk), .Q(reg_w_7[7]) );
  dff_sg \reg_ww_7_reg[7]  ( .D(n4859), .CP(clk), .Q(reg_ww_7[7]) );
  dff_sg \reg_www_7_reg[7]  ( .D(n4839), .CP(clk), .Q(reg_www_7[7]) );
  dff_sg \reg_w_7_reg[6]  ( .D(n5514), .CP(clk), .Q(reg_w_7[6]) );
  dff_sg \reg_ww_7_reg[6]  ( .D(n4860), .CP(clk), .Q(reg_ww_7[6]) );
  dff_sg \reg_www_7_reg[6]  ( .D(n4840), .CP(clk), .Q(reg_www_7[6]) );
  dff_sg \reg_w_7_reg[5]  ( .D(n5515), .CP(clk), .Q(reg_w_7[5]) );
  dff_sg \reg_ww_7_reg[5]  ( .D(n4861), .CP(clk), .Q(reg_ww_7[5]) );
  dff_sg \reg_www_7_reg[5]  ( .D(n4841), .CP(clk), .Q(reg_www_7[5]) );
  dff_sg \reg_w_7_reg[4]  ( .D(n5516), .CP(clk), .Q(reg_w_7[4]) );
  dff_sg \reg_ww_7_reg[4]  ( .D(n4862), .CP(clk), .Q(reg_ww_7[4]) );
  dff_sg \reg_www_7_reg[4]  ( .D(n4842), .CP(clk), .Q(reg_www_7[4]) );
  dff_sg \reg_w_7_reg[3]  ( .D(n5517), .CP(clk), .Q(reg_w_7[3]) );
  dff_sg \reg_ww_7_reg[3]  ( .D(n4863), .CP(clk), .Q(reg_ww_7[3]) );
  dff_sg \reg_www_7_reg[3]  ( .D(n4843), .CP(clk), .Q(reg_www_7[3]) );
  dff_sg \reg_w_7_reg[2]  ( .D(n5518), .CP(clk), .Q(reg_w_7[2]) );
  dff_sg \reg_ww_7_reg[2]  ( .D(n4864), .CP(clk), .Q(reg_ww_7[2]) );
  dff_sg \reg_www_7_reg[2]  ( .D(n4844), .CP(clk), .Q(reg_www_7[2]) );
  dff_sg \reg_w_7_reg[1]  ( .D(n5519), .CP(clk), .Q(reg_w_7[1]) );
  dff_sg \reg_ww_7_reg[1]  ( .D(n4865), .CP(clk), .Q(reg_ww_7[1]) );
  dff_sg \reg_www_7_reg[1]  ( .D(n4845), .CP(clk), .Q(reg_www_7[1]) );
  dff_sg \reg_w_7_reg[0]  ( .D(n5520), .CP(clk), .Q(reg_w_7[0]) );
  dff_sg \reg_ww_7_reg[0]  ( .D(n4866), .CP(clk), .Q(reg_ww_7[0]) );
  dff_sg \reg_www_7_reg[0]  ( .D(n4846), .CP(clk), .Q(reg_www_7[0]) );
  dff_sg \reg_w_6_reg[19]  ( .D(n5521), .CP(clk), .Q(reg_w_6[19]) );
  dff_sg \reg_ww_6_reg[19]  ( .D(n4887), .CP(clk), .Q(reg_ww_6[19]) );
  dff_sg \reg_www_6_reg[19]  ( .D(n4867), .CP(clk), .Q(reg_www_6[19]) );
  dff_sg \reg_w_6_reg[18]  ( .D(n5522), .CP(clk), .Q(reg_w_6[18]) );
  dff_sg \reg_ww_6_reg[18]  ( .D(n4888), .CP(clk), .Q(reg_ww_6[18]) );
  dff_sg \reg_www_6_reg[18]  ( .D(n4868), .CP(clk), .Q(reg_www_6[18]) );
  dff_sg \reg_w_6_reg[17]  ( .D(n5523), .CP(clk), .Q(reg_w_6[17]) );
  dff_sg \reg_ww_6_reg[17]  ( .D(n4889), .CP(clk), .Q(reg_ww_6[17]) );
  dff_sg \reg_www_6_reg[17]  ( .D(n4869), .CP(clk), .Q(reg_www_6[17]) );
  dff_sg \reg_w_6_reg[16]  ( .D(n5524), .CP(clk), .Q(reg_w_6[16]) );
  dff_sg \reg_ww_6_reg[16]  ( .D(n4890), .CP(clk), .Q(reg_ww_6[16]) );
  dff_sg \reg_www_6_reg[16]  ( .D(n4870), .CP(clk), .Q(reg_www_6[16]) );
  dff_sg \reg_w_6_reg[15]  ( .D(n5525), .CP(clk), .Q(reg_w_6[15]) );
  dff_sg \reg_ww_6_reg[15]  ( .D(n4891), .CP(clk), .Q(reg_ww_6[15]) );
  dff_sg \reg_www_6_reg[15]  ( .D(n4871), .CP(clk), .Q(reg_www_6[15]) );
  dff_sg \reg_w_6_reg[14]  ( .D(n5526), .CP(clk), .Q(reg_w_6[14]) );
  dff_sg \reg_ww_6_reg[14]  ( .D(n4892), .CP(clk), .Q(reg_ww_6[14]) );
  dff_sg \reg_www_6_reg[14]  ( .D(n4872), .CP(clk), .Q(reg_www_6[14]) );
  dff_sg \reg_w_6_reg[13]  ( .D(n5527), .CP(clk), .Q(reg_w_6[13]) );
  dff_sg \reg_ww_6_reg[13]  ( .D(n4893), .CP(clk), .Q(reg_ww_6[13]) );
  dff_sg \reg_www_6_reg[13]  ( .D(n4873), .CP(clk), .Q(reg_www_6[13]) );
  dff_sg \reg_w_6_reg[12]  ( .D(n5528), .CP(clk), .Q(reg_w_6[12]) );
  dff_sg \reg_ww_6_reg[12]  ( .D(n4894), .CP(clk), .Q(reg_ww_6[12]) );
  dff_sg \reg_www_6_reg[12]  ( .D(n4874), .CP(clk), .Q(reg_www_6[12]) );
  dff_sg \reg_w_6_reg[11]  ( .D(n5529), .CP(clk), .Q(reg_w_6[11]) );
  dff_sg \reg_ww_6_reg[11]  ( .D(n4895), .CP(clk), .Q(reg_ww_6[11]) );
  dff_sg \reg_www_6_reg[11]  ( .D(n4875), .CP(clk), .Q(reg_www_6[11]) );
  dff_sg \reg_w_6_reg[10]  ( .D(n5530), .CP(clk), .Q(reg_w_6[10]) );
  dff_sg \reg_ww_6_reg[10]  ( .D(n4896), .CP(clk), .Q(reg_ww_6[10]) );
  dff_sg \reg_www_6_reg[10]  ( .D(n4876), .CP(clk), .Q(reg_www_6[10]) );
  dff_sg \reg_w_6_reg[9]  ( .D(n5531), .CP(clk), .Q(reg_w_6[9]) );
  dff_sg \reg_ww_6_reg[9]  ( .D(n4897), .CP(clk), .Q(reg_ww_6[9]) );
  dff_sg \reg_www_6_reg[9]  ( .D(n4877), .CP(clk), .Q(reg_www_6[9]) );
  dff_sg \reg_w_6_reg[8]  ( .D(n5532), .CP(clk), .Q(reg_w_6[8]) );
  dff_sg \reg_ww_6_reg[8]  ( .D(n4898), .CP(clk), .Q(reg_ww_6[8]) );
  dff_sg \reg_www_6_reg[8]  ( .D(n4878), .CP(clk), .Q(reg_www_6[8]) );
  dff_sg \reg_w_6_reg[7]  ( .D(n5533), .CP(clk), .Q(reg_w_6[7]) );
  dff_sg \reg_ww_6_reg[7]  ( .D(n4899), .CP(clk), .Q(reg_ww_6[7]) );
  dff_sg \reg_www_6_reg[7]  ( .D(n4879), .CP(clk), .Q(reg_www_6[7]) );
  dff_sg \reg_w_6_reg[6]  ( .D(n5534), .CP(clk), .Q(reg_w_6[6]) );
  dff_sg \reg_ww_6_reg[6]  ( .D(n4900), .CP(clk), .Q(reg_ww_6[6]) );
  dff_sg \reg_www_6_reg[6]  ( .D(n4880), .CP(clk), .Q(reg_www_6[6]) );
  dff_sg \reg_w_6_reg[5]  ( .D(n5535), .CP(clk), .Q(reg_w_6[5]) );
  dff_sg \reg_ww_6_reg[5]  ( .D(n4901), .CP(clk), .Q(reg_ww_6[5]) );
  dff_sg \reg_www_6_reg[5]  ( .D(n4881), .CP(clk), .Q(reg_www_6[5]) );
  dff_sg \reg_w_6_reg[4]  ( .D(n5536), .CP(clk), .Q(reg_w_6[4]) );
  dff_sg \reg_ww_6_reg[4]  ( .D(n4902), .CP(clk), .Q(reg_ww_6[4]) );
  dff_sg \reg_www_6_reg[4]  ( .D(n4882), .CP(clk), .Q(reg_www_6[4]) );
  dff_sg \reg_w_6_reg[3]  ( .D(n5537), .CP(clk), .Q(reg_w_6[3]) );
  dff_sg \reg_ww_6_reg[3]  ( .D(n4903), .CP(clk), .Q(reg_ww_6[3]) );
  dff_sg \reg_www_6_reg[3]  ( .D(n4883), .CP(clk), .Q(reg_www_6[3]) );
  dff_sg \reg_w_6_reg[2]  ( .D(n5538), .CP(clk), .Q(reg_w_6[2]) );
  dff_sg \reg_ww_6_reg[2]  ( .D(n4904), .CP(clk), .Q(reg_ww_6[2]) );
  dff_sg \reg_www_6_reg[2]  ( .D(n4884), .CP(clk), .Q(reg_www_6[2]) );
  dff_sg \reg_w_6_reg[1]  ( .D(n5539), .CP(clk), .Q(reg_w_6[1]) );
  dff_sg \reg_ww_6_reg[1]  ( .D(n4905), .CP(clk), .Q(reg_ww_6[1]) );
  dff_sg \reg_www_6_reg[1]  ( .D(n4885), .CP(clk), .Q(reg_www_6[1]) );
  dff_sg \reg_w_6_reg[0]  ( .D(n5540), .CP(clk), .Q(reg_w_6[0]) );
  dff_sg \reg_ww_6_reg[0]  ( .D(n4906), .CP(clk), .Q(reg_ww_6[0]) );
  dff_sg \reg_www_6_reg[0]  ( .D(n4886), .CP(clk), .Q(reg_www_6[0]) );
  dff_sg \reg_w_5_reg[19]  ( .D(n5541), .CP(clk), .Q(reg_w_5[19]) );
  dff_sg \reg_ww_5_reg[19]  ( .D(n4927), .CP(clk), .Q(reg_ww_5[19]) );
  dff_sg \reg_www_5_reg[19]  ( .D(n4907), .CP(clk), .Q(reg_www_5[19]) );
  dff_sg \reg_w_5_reg[18]  ( .D(n5542), .CP(clk), .Q(reg_w_5[18]) );
  dff_sg \reg_ww_5_reg[18]  ( .D(n4928), .CP(clk), .Q(reg_ww_5[18]) );
  dff_sg \reg_www_5_reg[18]  ( .D(n4908), .CP(clk), .Q(reg_www_5[18]) );
  dff_sg \reg_w_5_reg[17]  ( .D(n5543), .CP(clk), .Q(reg_w_5[17]) );
  dff_sg \reg_ww_5_reg[17]  ( .D(n4929), .CP(clk), .Q(reg_ww_5[17]) );
  dff_sg \reg_www_5_reg[17]  ( .D(n4909), .CP(clk), .Q(reg_www_5[17]) );
  dff_sg \reg_w_5_reg[16]  ( .D(n5544), .CP(clk), .Q(reg_w_5[16]) );
  dff_sg \reg_ww_5_reg[16]  ( .D(n4930), .CP(clk), .Q(reg_ww_5[16]) );
  dff_sg \reg_www_5_reg[16]  ( .D(n4910), .CP(clk), .Q(reg_www_5[16]) );
  dff_sg \reg_w_5_reg[15]  ( .D(n5545), .CP(clk), .Q(reg_w_5[15]) );
  dff_sg \reg_ww_5_reg[15]  ( .D(n4931), .CP(clk), .Q(reg_ww_5[15]) );
  dff_sg \reg_www_5_reg[15]  ( .D(n4911), .CP(clk), .Q(reg_www_5[15]) );
  dff_sg \reg_w_5_reg[14]  ( .D(n5546), .CP(clk), .Q(reg_w_5[14]) );
  dff_sg \reg_ww_5_reg[14]  ( .D(n4932), .CP(clk), .Q(reg_ww_5[14]) );
  dff_sg \reg_www_5_reg[14]  ( .D(n4912), .CP(clk), .Q(reg_www_5[14]) );
  dff_sg \reg_w_5_reg[13]  ( .D(n5547), .CP(clk), .Q(reg_w_5[13]) );
  dff_sg \reg_ww_5_reg[13]  ( .D(n4933), .CP(clk), .Q(reg_ww_5[13]) );
  dff_sg \reg_www_5_reg[13]  ( .D(n4913), .CP(clk), .Q(reg_www_5[13]) );
  dff_sg \reg_w_5_reg[12]  ( .D(n5548), .CP(clk), .Q(reg_w_5[12]) );
  dff_sg \reg_ww_5_reg[12]  ( .D(n4934), .CP(clk), .Q(reg_ww_5[12]) );
  dff_sg \reg_www_5_reg[12]  ( .D(n4914), .CP(clk), .Q(reg_www_5[12]) );
  dff_sg \reg_w_5_reg[11]  ( .D(n5549), .CP(clk), .Q(reg_w_5[11]) );
  dff_sg \reg_ww_5_reg[11]  ( .D(n4935), .CP(clk), .Q(reg_ww_5[11]) );
  dff_sg \reg_www_5_reg[11]  ( .D(n4915), .CP(clk), .Q(reg_www_5[11]) );
  dff_sg \reg_w_5_reg[10]  ( .D(n5550), .CP(clk), .Q(reg_w_5[10]) );
  dff_sg \reg_ww_5_reg[10]  ( .D(n4936), .CP(clk), .Q(reg_ww_5[10]) );
  dff_sg \reg_www_5_reg[10]  ( .D(n4916), .CP(clk), .Q(reg_www_5[10]) );
  dff_sg \reg_w_5_reg[9]  ( .D(n5551), .CP(clk), .Q(reg_w_5[9]) );
  dff_sg \reg_ww_5_reg[9]  ( .D(n4937), .CP(clk), .Q(reg_ww_5[9]) );
  dff_sg \reg_www_5_reg[9]  ( .D(n4917), .CP(clk), .Q(reg_www_5[9]) );
  dff_sg \reg_w_5_reg[8]  ( .D(n5552), .CP(clk), .Q(reg_w_5[8]) );
  dff_sg \reg_ww_5_reg[8]  ( .D(n4938), .CP(clk), .Q(reg_ww_5[8]) );
  dff_sg \reg_www_5_reg[8]  ( .D(n4918), .CP(clk), .Q(reg_www_5[8]) );
  dff_sg \reg_w_5_reg[7]  ( .D(n5553), .CP(clk), .Q(reg_w_5[7]) );
  dff_sg \reg_ww_5_reg[7]  ( .D(n4939), .CP(clk), .Q(reg_ww_5[7]) );
  dff_sg \reg_www_5_reg[7]  ( .D(n4919), .CP(clk), .Q(reg_www_5[7]) );
  dff_sg \reg_w_5_reg[6]  ( .D(n5554), .CP(clk), .Q(reg_w_5[6]) );
  dff_sg \reg_ww_5_reg[6]  ( .D(n4940), .CP(clk), .Q(reg_ww_5[6]) );
  dff_sg \reg_www_5_reg[6]  ( .D(n4920), .CP(clk), .Q(reg_www_5[6]) );
  dff_sg \reg_w_5_reg[5]  ( .D(n5555), .CP(clk), .Q(reg_w_5[5]) );
  dff_sg \reg_ww_5_reg[5]  ( .D(n4941), .CP(clk), .Q(reg_ww_5[5]) );
  dff_sg \reg_www_5_reg[5]  ( .D(n4921), .CP(clk), .Q(reg_www_5[5]) );
  dff_sg \reg_w_5_reg[4]  ( .D(n5556), .CP(clk), .Q(reg_w_5[4]) );
  dff_sg \reg_ww_5_reg[4]  ( .D(n4942), .CP(clk), .Q(reg_ww_5[4]) );
  dff_sg \reg_www_5_reg[4]  ( .D(n4922), .CP(clk), .Q(reg_www_5[4]) );
  dff_sg \reg_w_5_reg[3]  ( .D(n5557), .CP(clk), .Q(reg_w_5[3]) );
  dff_sg \reg_ww_5_reg[3]  ( .D(n4943), .CP(clk), .Q(reg_ww_5[3]) );
  dff_sg \reg_www_5_reg[3]  ( .D(n4923), .CP(clk), .Q(reg_www_5[3]) );
  dff_sg \reg_w_5_reg[2]  ( .D(n5558), .CP(clk), .Q(reg_w_5[2]) );
  dff_sg \reg_ww_5_reg[2]  ( .D(n4944), .CP(clk), .Q(reg_ww_5[2]) );
  dff_sg \reg_www_5_reg[2]  ( .D(n4924), .CP(clk), .Q(reg_www_5[2]) );
  dff_sg \reg_w_5_reg[1]  ( .D(n5559), .CP(clk), .Q(reg_w_5[1]) );
  dff_sg \reg_ww_5_reg[1]  ( .D(n4945), .CP(clk), .Q(reg_ww_5[1]) );
  dff_sg \reg_www_5_reg[1]  ( .D(n4925), .CP(clk), .Q(reg_www_5[1]) );
  dff_sg \reg_w_5_reg[0]  ( .D(n5560), .CP(clk), .Q(reg_w_5[0]) );
  dff_sg \reg_ww_5_reg[0]  ( .D(n4946), .CP(clk), .Q(reg_ww_5[0]) );
  dff_sg \reg_www_5_reg[0]  ( .D(n4926), .CP(clk), .Q(reg_www_5[0]) );
  dff_sg \reg_w_4_reg[19]  ( .D(n5561), .CP(clk), .Q(reg_w_4[19]) );
  dff_sg \reg_ww_4_reg[19]  ( .D(n4967), .CP(clk), .Q(reg_ww_4[19]) );
  dff_sg \reg_www_4_reg[19]  ( .D(n4947), .CP(clk), .Q(reg_www_4[19]) );
  dff_sg \reg_w_4_reg[18]  ( .D(n5562), .CP(clk), .Q(reg_w_4[18]) );
  dff_sg \reg_ww_4_reg[18]  ( .D(n4968), .CP(clk), .Q(reg_ww_4[18]) );
  dff_sg \reg_www_4_reg[18]  ( .D(n4948), .CP(clk), .Q(reg_www_4[18]) );
  dff_sg \reg_w_4_reg[17]  ( .D(n5563), .CP(clk), .Q(reg_w_4[17]) );
  dff_sg \reg_ww_4_reg[17]  ( .D(n4969), .CP(clk), .Q(reg_ww_4[17]) );
  dff_sg \reg_www_4_reg[17]  ( .D(n4949), .CP(clk), .Q(reg_www_4[17]) );
  dff_sg \reg_w_4_reg[16]  ( .D(n5564), .CP(clk), .Q(reg_w_4[16]) );
  dff_sg \reg_ww_4_reg[16]  ( .D(n4970), .CP(clk), .Q(reg_ww_4[16]) );
  dff_sg \reg_www_4_reg[16]  ( .D(n4950), .CP(clk), .Q(reg_www_4[16]) );
  dff_sg \reg_w_4_reg[15]  ( .D(n5565), .CP(clk), .Q(reg_w_4[15]) );
  dff_sg \reg_ww_4_reg[15]  ( .D(n4971), .CP(clk), .Q(reg_ww_4[15]) );
  dff_sg \reg_www_4_reg[15]  ( .D(n4951), .CP(clk), .Q(reg_www_4[15]) );
  dff_sg \reg_w_4_reg[14]  ( .D(n5566), .CP(clk), .Q(reg_w_4[14]) );
  dff_sg \reg_ww_4_reg[14]  ( .D(n4972), .CP(clk), .Q(reg_ww_4[14]) );
  dff_sg \reg_www_4_reg[14]  ( .D(n4952), .CP(clk), .Q(reg_www_4[14]) );
  dff_sg \reg_w_4_reg[13]  ( .D(n5567), .CP(clk), .Q(reg_w_4[13]) );
  dff_sg \reg_ww_4_reg[13]  ( .D(n4973), .CP(clk), .Q(reg_ww_4[13]) );
  dff_sg \reg_www_4_reg[13]  ( .D(n4953), .CP(clk), .Q(reg_www_4[13]) );
  dff_sg \reg_w_4_reg[12]  ( .D(n5568), .CP(clk), .Q(reg_w_4[12]) );
  dff_sg \reg_ww_4_reg[12]  ( .D(n4974), .CP(clk), .Q(reg_ww_4[12]) );
  dff_sg \reg_www_4_reg[12]  ( .D(n4954), .CP(clk), .Q(reg_www_4[12]) );
  dff_sg \reg_w_4_reg[11]  ( .D(n5569), .CP(clk), .Q(reg_w_4[11]) );
  dff_sg \reg_ww_4_reg[11]  ( .D(n4975), .CP(clk), .Q(reg_ww_4[11]) );
  dff_sg \reg_www_4_reg[11]  ( .D(n4955), .CP(clk), .Q(reg_www_4[11]) );
  dff_sg \reg_w_4_reg[10]  ( .D(n5570), .CP(clk), .Q(reg_w_4[10]) );
  dff_sg \reg_ww_4_reg[10]  ( .D(n4976), .CP(clk), .Q(reg_ww_4[10]) );
  dff_sg \reg_www_4_reg[10]  ( .D(n4956), .CP(clk), .Q(reg_www_4[10]) );
  dff_sg \reg_w_4_reg[9]  ( .D(n5571), .CP(clk), .Q(reg_w_4[9]) );
  dff_sg \reg_ww_4_reg[9]  ( .D(n4977), .CP(clk), .Q(reg_ww_4[9]) );
  dff_sg \reg_www_4_reg[9]  ( .D(n4957), .CP(clk), .Q(reg_www_4[9]) );
  dff_sg \reg_w_4_reg[8]  ( .D(n5572), .CP(clk), .Q(reg_w_4[8]) );
  dff_sg \reg_ww_4_reg[8]  ( .D(n4978), .CP(clk), .Q(reg_ww_4[8]) );
  dff_sg \reg_www_4_reg[8]  ( .D(n4958), .CP(clk), .Q(reg_www_4[8]) );
  dff_sg \reg_w_4_reg[7]  ( .D(n5573), .CP(clk), .Q(reg_w_4[7]) );
  dff_sg \reg_ww_4_reg[7]  ( .D(n4979), .CP(clk), .Q(reg_ww_4[7]) );
  dff_sg \reg_www_4_reg[7]  ( .D(n4959), .CP(clk), .Q(reg_www_4[7]) );
  dff_sg \reg_w_4_reg[6]  ( .D(n5574), .CP(clk), .Q(reg_w_4[6]) );
  dff_sg \reg_ww_4_reg[6]  ( .D(n4980), .CP(clk), .Q(reg_ww_4[6]) );
  dff_sg \reg_www_4_reg[6]  ( .D(n4960), .CP(clk), .Q(reg_www_4[6]) );
  dff_sg \reg_w_4_reg[5]  ( .D(n5575), .CP(clk), .Q(reg_w_4[5]) );
  dff_sg \reg_ww_4_reg[5]  ( .D(n4981), .CP(clk), .Q(reg_ww_4[5]) );
  dff_sg \reg_www_4_reg[5]  ( .D(n4961), .CP(clk), .Q(reg_www_4[5]) );
  dff_sg \reg_w_4_reg[4]  ( .D(n5576), .CP(clk), .Q(reg_w_4[4]) );
  dff_sg \reg_ww_4_reg[4]  ( .D(n4982), .CP(clk), .Q(reg_ww_4[4]) );
  dff_sg \reg_www_4_reg[4]  ( .D(n4962), .CP(clk), .Q(reg_www_4[4]) );
  dff_sg \reg_w_4_reg[3]  ( .D(n5577), .CP(clk), .Q(reg_w_4[3]) );
  dff_sg \reg_ww_4_reg[3]  ( .D(n4983), .CP(clk), .Q(reg_ww_4[3]) );
  dff_sg \reg_www_4_reg[3]  ( .D(n4963), .CP(clk), .Q(reg_www_4[3]) );
  dff_sg \reg_w_4_reg[2]  ( .D(n5578), .CP(clk), .Q(reg_w_4[2]) );
  dff_sg \reg_ww_4_reg[2]  ( .D(n4984), .CP(clk), .Q(reg_ww_4[2]) );
  dff_sg \reg_www_4_reg[2]  ( .D(n4964), .CP(clk), .Q(reg_www_4[2]) );
  dff_sg \reg_w_4_reg[1]  ( .D(n5579), .CP(clk), .Q(reg_w_4[1]) );
  dff_sg \reg_ww_4_reg[1]  ( .D(n4985), .CP(clk), .Q(reg_ww_4[1]) );
  dff_sg \reg_www_4_reg[1]  ( .D(n4965), .CP(clk), .Q(reg_www_4[1]) );
  dff_sg \reg_w_4_reg[0]  ( .D(n5580), .CP(clk), .Q(reg_w_4[0]) );
  dff_sg \reg_ww_4_reg[0]  ( .D(n4986), .CP(clk), .Q(reg_ww_4[0]) );
  dff_sg \reg_www_4_reg[0]  ( .D(n4966), .CP(clk), .Q(reg_www_4[0]) );
  dff_sg \reg_w_3_reg[19]  ( .D(n5581), .CP(clk), .Q(reg_w_3[19]) );
  dff_sg \reg_ww_3_reg[19]  ( .D(n4987), .CP(clk), .Q(reg_ww_3[19]) );
  dff_sg \reg_www_3_reg[19]  ( .D(n4593), .CP(clk), .Q(reg_www_3[19]) );
  dff_sg \reg_w_3_reg[18]  ( .D(n5582), .CP(clk), .Q(reg_w_3[18]) );
  dff_sg \reg_ww_3_reg[18]  ( .D(n4988), .CP(clk), .Q(reg_ww_3[18]) );
  dff_sg \reg_www_3_reg[18]  ( .D(n4594), .CP(clk), .Q(reg_www_3[18]) );
  dff_sg \reg_w_3_reg[17]  ( .D(n5583), .CP(clk), .Q(reg_w_3[17]) );
  dff_sg \reg_ww_3_reg[17]  ( .D(n4989), .CP(clk), .Q(reg_ww_3[17]) );
  dff_sg \reg_www_3_reg[17]  ( .D(n4595), .CP(clk), .Q(reg_www_3[17]) );
  dff_sg \reg_w_3_reg[16]  ( .D(n5584), .CP(clk), .Q(reg_w_3[16]) );
  dff_sg \reg_ww_3_reg[16]  ( .D(n4990), .CP(clk), .Q(reg_ww_3[16]) );
  dff_sg \reg_www_3_reg[16]  ( .D(n4596), .CP(clk), .Q(reg_www_3[16]) );
  dff_sg \reg_w_3_reg[15]  ( .D(n5585), .CP(clk), .Q(reg_w_3[15]) );
  dff_sg \reg_ww_3_reg[15]  ( .D(n4613), .CP(clk), .Q(reg_ww_3[15]) );
  dff_sg \reg_www_3_reg[15]  ( .D(n4597), .CP(clk), .Q(reg_www_3[15]) );
  dff_sg \reg_w_3_reg[14]  ( .D(n5586), .CP(clk), .Q(reg_w_3[14]) );
  dff_sg \reg_ww_3_reg[14]  ( .D(n4614), .CP(clk), .Q(reg_ww_3[14]) );
  dff_sg \reg_www_3_reg[14]  ( .D(n4598), .CP(clk), .Q(reg_www_3[14]) );
  dff_sg \reg_w_3_reg[13]  ( .D(n5587), .CP(clk), .Q(reg_w_3[13]) );
  dff_sg \reg_ww_3_reg[13]  ( .D(n4615), .CP(clk), .Q(reg_ww_3[13]) );
  dff_sg \reg_www_3_reg[13]  ( .D(n4599), .CP(clk), .Q(reg_www_3[13]) );
  dff_sg \reg_w_3_reg[12]  ( .D(n5588), .CP(clk), .Q(reg_w_3[12]) );
  dff_sg \reg_ww_3_reg[12]  ( .D(n4616), .CP(clk), .Q(reg_ww_3[12]) );
  dff_sg \reg_www_3_reg[12]  ( .D(n4600), .CP(clk), .Q(reg_www_3[12]) );
  dff_sg \reg_w_3_reg[11]  ( .D(n5589), .CP(clk), .Q(reg_w_3[11]) );
  dff_sg \reg_ww_3_reg[11]  ( .D(n4617), .CP(clk), .Q(reg_ww_3[11]) );
  dff_sg \reg_www_3_reg[11]  ( .D(n4601), .CP(clk), .Q(reg_www_3[11]) );
  dff_sg \reg_w_3_reg[10]  ( .D(n5590), .CP(clk), .Q(reg_w_3[10]) );
  dff_sg \reg_ww_3_reg[10]  ( .D(n4618), .CP(clk), .Q(reg_ww_3[10]) );
  dff_sg \reg_www_3_reg[10]  ( .D(n4602), .CP(clk), .Q(reg_www_3[10]) );
  dff_sg \reg_w_3_reg[9]  ( .D(n5591), .CP(clk), .Q(reg_w_3[9]) );
  dff_sg \reg_ww_3_reg[9]  ( .D(n4619), .CP(clk), .Q(reg_ww_3[9]) );
  dff_sg \reg_www_3_reg[9]  ( .D(n4603), .CP(clk), .Q(reg_www_3[9]) );
  dff_sg \reg_w_3_reg[8]  ( .D(n5592), .CP(clk), .Q(reg_w_3[8]) );
  dff_sg \reg_ww_3_reg[8]  ( .D(n4620), .CP(clk), .Q(reg_ww_3[8]) );
  dff_sg \reg_www_3_reg[8]  ( .D(n4604), .CP(clk), .Q(reg_www_3[8]) );
  dff_sg \reg_w_3_reg[7]  ( .D(n5593), .CP(clk), .Q(reg_w_3[7]) );
  dff_sg \reg_ww_3_reg[7]  ( .D(n4621), .CP(clk), .Q(reg_ww_3[7]) );
  dff_sg \reg_www_3_reg[7]  ( .D(n4605), .CP(clk), .Q(reg_www_3[7]) );
  dff_sg \reg_w_3_reg[6]  ( .D(n5594), .CP(clk), .Q(reg_w_3[6]) );
  dff_sg \reg_ww_3_reg[6]  ( .D(n4622), .CP(clk), .Q(reg_ww_3[6]) );
  dff_sg \reg_www_3_reg[6]  ( .D(n4606), .CP(clk), .Q(reg_www_3[6]) );
  dff_sg \reg_w_3_reg[5]  ( .D(n5595), .CP(clk), .Q(reg_w_3[5]) );
  dff_sg \reg_ww_3_reg[5]  ( .D(n4623), .CP(clk), .Q(reg_ww_3[5]) );
  dff_sg \reg_www_3_reg[5]  ( .D(n4607), .CP(clk), .Q(reg_www_3[5]) );
  dff_sg \reg_w_3_reg[4]  ( .D(n5596), .CP(clk), .Q(reg_w_3[4]) );
  dff_sg \reg_ww_3_reg[4]  ( .D(n4624), .CP(clk), .Q(reg_ww_3[4]) );
  dff_sg \reg_www_3_reg[4]  ( .D(n4608), .CP(clk), .Q(reg_www_3[4]) );
  dff_sg \reg_w_3_reg[3]  ( .D(n5597), .CP(clk), .Q(reg_w_3[3]) );
  dff_sg \reg_ww_3_reg[3]  ( .D(n4625), .CP(clk), .Q(reg_ww_3[3]) );
  dff_sg \reg_www_3_reg[3]  ( .D(n4609), .CP(clk), .Q(reg_www_3[3]) );
  dff_sg \reg_w_3_reg[2]  ( .D(n5598), .CP(clk), .Q(reg_w_3[2]) );
  dff_sg \reg_ww_3_reg[2]  ( .D(n4626), .CP(clk), .Q(reg_ww_3[2]) );
  dff_sg \reg_www_3_reg[2]  ( .D(n4610), .CP(clk), .Q(reg_www_3[2]) );
  dff_sg \reg_w_3_reg[1]  ( .D(n5599), .CP(clk), .Q(reg_w_3[1]) );
  dff_sg \reg_ww_3_reg[1]  ( .D(n4627), .CP(clk), .Q(reg_ww_3[1]) );
  dff_sg \reg_www_3_reg[1]  ( .D(n4611), .CP(clk), .Q(reg_www_3[1]) );
  dff_sg \reg_w_3_reg[0]  ( .D(n5600), .CP(clk), .Q(reg_w_3[0]) );
  dff_sg \reg_ww_3_reg[0]  ( .D(n4628), .CP(clk), .Q(reg_ww_3[0]) );
  dff_sg \reg_www_3_reg[0]  ( .D(n4612), .CP(clk), .Q(reg_www_3[0]) );
  dff_sg \reg_w_2_reg[19]  ( .D(n5601), .CP(clk), .Q(reg_w_2[19]) );
  dff_sg \reg_ww_2_reg[19]  ( .D(n4649), .CP(clk), .Q(reg_ww_2[19]) );
  dff_sg \reg_www_2_reg[19]  ( .D(n4629), .CP(clk), .Q(reg_www_2[19]) );
  dff_sg \reg_w_2_reg[18]  ( .D(n5602), .CP(clk), .Q(reg_w_2[18]) );
  dff_sg \reg_ww_2_reg[18]  ( .D(n4650), .CP(clk), .Q(reg_ww_2[18]) );
  dff_sg \reg_www_2_reg[18]  ( .D(n4630), .CP(clk), .Q(reg_www_2[18]) );
  dff_sg \reg_w_2_reg[17]  ( .D(n5603), .CP(clk), .Q(reg_w_2[17]) );
  dff_sg \reg_ww_2_reg[17]  ( .D(n4651), .CP(clk), .Q(reg_ww_2[17]) );
  dff_sg \reg_www_2_reg[17]  ( .D(n4631), .CP(clk), .Q(reg_www_2[17]) );
  dff_sg \reg_w_2_reg[16]  ( .D(n5604), .CP(clk), .Q(reg_w_2[16]) );
  dff_sg \reg_ww_2_reg[16]  ( .D(n4652), .CP(clk), .Q(reg_ww_2[16]) );
  dff_sg \reg_www_2_reg[16]  ( .D(n4632), .CP(clk), .Q(reg_www_2[16]) );
  dff_sg \reg_w_2_reg[15]  ( .D(n5605), .CP(clk), .Q(reg_w_2[15]) );
  dff_sg \reg_ww_2_reg[15]  ( .D(n4653), .CP(clk), .Q(reg_ww_2[15]) );
  dff_sg \reg_www_2_reg[15]  ( .D(n4633), .CP(clk), .Q(reg_www_2[15]) );
  dff_sg \reg_w_2_reg[14]  ( .D(n5606), .CP(clk), .Q(reg_w_2[14]) );
  dff_sg \reg_ww_2_reg[14]  ( .D(n4654), .CP(clk), .Q(reg_ww_2[14]) );
  dff_sg \reg_www_2_reg[14]  ( .D(n4634), .CP(clk), .Q(reg_www_2[14]) );
  dff_sg \reg_w_2_reg[13]  ( .D(n5607), .CP(clk), .Q(reg_w_2[13]) );
  dff_sg \reg_ww_2_reg[13]  ( .D(n4655), .CP(clk), .Q(reg_ww_2[13]) );
  dff_sg \reg_www_2_reg[13]  ( .D(n4635), .CP(clk), .Q(reg_www_2[13]) );
  dff_sg \reg_w_2_reg[12]  ( .D(n5608), .CP(clk), .Q(reg_w_2[12]) );
  dff_sg \reg_ww_2_reg[12]  ( .D(n4656), .CP(clk), .Q(reg_ww_2[12]) );
  dff_sg \reg_www_2_reg[12]  ( .D(n4636), .CP(clk), .Q(reg_www_2[12]) );
  dff_sg \reg_w_2_reg[11]  ( .D(n5609), .CP(clk), .Q(reg_w_2[11]) );
  dff_sg \reg_ww_2_reg[11]  ( .D(n4657), .CP(clk), .Q(reg_ww_2[11]) );
  dff_sg \reg_www_2_reg[11]  ( .D(n4637), .CP(clk), .Q(reg_www_2[11]) );
  dff_sg \reg_w_2_reg[10]  ( .D(n5610), .CP(clk), .Q(reg_w_2[10]) );
  dff_sg \reg_ww_2_reg[10]  ( .D(n4658), .CP(clk), .Q(reg_ww_2[10]) );
  dff_sg \reg_www_2_reg[10]  ( .D(n4638), .CP(clk), .Q(reg_www_2[10]) );
  dff_sg \reg_w_2_reg[9]  ( .D(n5611), .CP(clk), .Q(reg_w_2[9]) );
  dff_sg \reg_ww_2_reg[9]  ( .D(n4659), .CP(clk), .Q(reg_ww_2[9]) );
  dff_sg \reg_www_2_reg[9]  ( .D(n4639), .CP(clk), .Q(reg_www_2[9]) );
  dff_sg \reg_w_2_reg[8]  ( .D(n5612), .CP(clk), .Q(reg_w_2[8]) );
  dff_sg \reg_ww_2_reg[8]  ( .D(n4660), .CP(clk), .Q(reg_ww_2[8]) );
  dff_sg \reg_www_2_reg[8]  ( .D(n4640), .CP(clk), .Q(reg_www_2[8]) );
  dff_sg \reg_w_2_reg[7]  ( .D(n5613), .CP(clk), .Q(reg_w_2[7]) );
  dff_sg \reg_ww_2_reg[7]  ( .D(n4661), .CP(clk), .Q(reg_ww_2[7]) );
  dff_sg \reg_www_2_reg[7]  ( .D(n4641), .CP(clk), .Q(reg_www_2[7]) );
  dff_sg \reg_w_2_reg[6]  ( .D(n5614), .CP(clk), .Q(reg_w_2[6]) );
  dff_sg \reg_ww_2_reg[6]  ( .D(n4662), .CP(clk), .Q(reg_ww_2[6]) );
  dff_sg \reg_www_2_reg[6]  ( .D(n4642), .CP(clk), .Q(reg_www_2[6]) );
  dff_sg \reg_w_2_reg[5]  ( .D(n5615), .CP(clk), .Q(reg_w_2[5]) );
  dff_sg \reg_ww_2_reg[5]  ( .D(n4663), .CP(clk), .Q(reg_ww_2[5]) );
  dff_sg \reg_www_2_reg[5]  ( .D(n4643), .CP(clk), .Q(reg_www_2[5]) );
  dff_sg \reg_w_2_reg[4]  ( .D(n5616), .CP(clk), .Q(reg_w_2[4]) );
  dff_sg \reg_ww_2_reg[4]  ( .D(n4664), .CP(clk), .Q(reg_ww_2[4]) );
  dff_sg \reg_www_2_reg[4]  ( .D(n4644), .CP(clk), .Q(reg_www_2[4]) );
  dff_sg \reg_w_2_reg[3]  ( .D(n5617), .CP(clk), .Q(reg_w_2[3]) );
  dff_sg \reg_ww_2_reg[3]  ( .D(n4665), .CP(clk), .Q(reg_ww_2[3]) );
  dff_sg \reg_www_2_reg[3]  ( .D(n4645), .CP(clk), .Q(reg_www_2[3]) );
  dff_sg \reg_w_2_reg[2]  ( .D(n5618), .CP(clk), .Q(reg_w_2[2]) );
  dff_sg \reg_ww_2_reg[2]  ( .D(n4666), .CP(clk), .Q(reg_ww_2[2]) );
  dff_sg \reg_www_2_reg[2]  ( .D(n4646), .CP(clk), .Q(reg_www_2[2]) );
  dff_sg \reg_w_2_reg[1]  ( .D(n5619), .CP(clk), .Q(reg_w_2[1]) );
  dff_sg \reg_ww_2_reg[1]  ( .D(n4667), .CP(clk), .Q(reg_ww_2[1]) );
  dff_sg \reg_www_2_reg[1]  ( .D(n4647), .CP(clk), .Q(reg_www_2[1]) );
  dff_sg \reg_w_2_reg[0]  ( .D(n5620), .CP(clk), .Q(reg_w_2[0]) );
  dff_sg \reg_ww_2_reg[0]  ( .D(n4668), .CP(clk), .Q(reg_ww_2[0]) );
  dff_sg \reg_www_2_reg[0]  ( .D(n4648), .CP(clk), .Q(reg_www_2[0]) );
  dff_sg \reg_w_1_reg[19]  ( .D(n5621), .CP(clk), .Q(reg_w_1[19]) );
  dff_sg \reg_ww_1_reg[19]  ( .D(n4689), .CP(clk), .Q(reg_ww_1[19]) );
  dff_sg \reg_www_1_reg[19]  ( .D(n4669), .CP(clk), .Q(reg_www_1[19]) );
  dff_sg \reg_w_1_reg[18]  ( .D(n5622), .CP(clk), .Q(reg_w_1[18]) );
  dff_sg \reg_ww_1_reg[18]  ( .D(n4690), .CP(clk), .Q(reg_ww_1[18]) );
  dff_sg \reg_www_1_reg[18]  ( .D(n4670), .CP(clk), .Q(reg_www_1[18]) );
  dff_sg \reg_w_1_reg[17]  ( .D(n5623), .CP(clk), .Q(reg_w_1[17]) );
  dff_sg \reg_ww_1_reg[17]  ( .D(n4691), .CP(clk), .Q(reg_ww_1[17]) );
  dff_sg \reg_www_1_reg[17]  ( .D(n4671), .CP(clk), .Q(reg_www_1[17]) );
  dff_sg \reg_w_1_reg[16]  ( .D(n5624), .CP(clk), .Q(reg_w_1[16]) );
  dff_sg \reg_ww_1_reg[16]  ( .D(n4692), .CP(clk), .Q(reg_ww_1[16]) );
  dff_sg \reg_www_1_reg[16]  ( .D(n4672), .CP(clk), .Q(reg_www_1[16]) );
  dff_sg \reg_w_1_reg[15]  ( .D(n5625), .CP(clk), .Q(reg_w_1[15]) );
  dff_sg \reg_ww_1_reg[15]  ( .D(n4693), .CP(clk), .Q(reg_ww_1[15]) );
  dff_sg \reg_www_1_reg[15]  ( .D(n4673), .CP(clk), .Q(reg_www_1[15]) );
  dff_sg \reg_w_1_reg[14]  ( .D(n5626), .CP(clk), .Q(reg_w_1[14]) );
  dff_sg \reg_ww_1_reg[14]  ( .D(n4694), .CP(clk), .Q(reg_ww_1[14]) );
  dff_sg \reg_www_1_reg[14]  ( .D(n4674), .CP(clk), .Q(reg_www_1[14]) );
  dff_sg \reg_w_1_reg[13]  ( .D(n5627), .CP(clk), .Q(reg_w_1[13]) );
  dff_sg \reg_ww_1_reg[13]  ( .D(n4695), .CP(clk), .Q(reg_ww_1[13]) );
  dff_sg \reg_www_1_reg[13]  ( .D(n4675), .CP(clk), .Q(reg_www_1[13]) );
  dff_sg \reg_w_1_reg[12]  ( .D(n5628), .CP(clk), .Q(reg_w_1[12]) );
  dff_sg \reg_ww_1_reg[12]  ( .D(n4696), .CP(clk), .Q(reg_ww_1[12]) );
  dff_sg \reg_www_1_reg[12]  ( .D(n4676), .CP(clk), .Q(reg_www_1[12]) );
  dff_sg \reg_w_1_reg[11]  ( .D(n5629), .CP(clk), .Q(reg_w_1[11]) );
  dff_sg \reg_ww_1_reg[11]  ( .D(n4697), .CP(clk), .Q(reg_ww_1[11]) );
  dff_sg \reg_www_1_reg[11]  ( .D(n4677), .CP(clk), .Q(reg_www_1[11]) );
  dff_sg \reg_w_1_reg[10]  ( .D(n5630), .CP(clk), .Q(reg_w_1[10]) );
  dff_sg \reg_ww_1_reg[10]  ( .D(n4698), .CP(clk), .Q(reg_ww_1[10]) );
  dff_sg \reg_www_1_reg[10]  ( .D(n4678), .CP(clk), .Q(reg_www_1[10]) );
  dff_sg \reg_w_1_reg[9]  ( .D(n5631), .CP(clk), .Q(reg_w_1[9]) );
  dff_sg \reg_ww_1_reg[9]  ( .D(n4699), .CP(clk), .Q(reg_ww_1[9]) );
  dff_sg \reg_www_1_reg[9]  ( .D(n4679), .CP(clk), .Q(reg_www_1[9]) );
  dff_sg \reg_w_1_reg[8]  ( .D(n5632), .CP(clk), .Q(reg_w_1[8]) );
  dff_sg \reg_ww_1_reg[8]  ( .D(n4700), .CP(clk), .Q(reg_ww_1[8]) );
  dff_sg \reg_www_1_reg[8]  ( .D(n4680), .CP(clk), .Q(reg_www_1[8]) );
  dff_sg \reg_w_1_reg[7]  ( .D(n5633), .CP(clk), .Q(reg_w_1[7]) );
  dff_sg \reg_ww_1_reg[7]  ( .D(n4701), .CP(clk), .Q(reg_ww_1[7]) );
  dff_sg \reg_www_1_reg[7]  ( .D(n4681), .CP(clk), .Q(reg_www_1[7]) );
  dff_sg \reg_w_1_reg[6]  ( .D(n5634), .CP(clk), .Q(reg_w_1[6]) );
  dff_sg \reg_ww_1_reg[6]  ( .D(n4702), .CP(clk), .Q(reg_ww_1[6]) );
  dff_sg \reg_www_1_reg[6]  ( .D(n4682), .CP(clk), .Q(reg_www_1[6]) );
  dff_sg \reg_w_1_reg[5]  ( .D(n5635), .CP(clk), .Q(reg_w_1[5]) );
  dff_sg \reg_ww_1_reg[5]  ( .D(n4703), .CP(clk), .Q(reg_ww_1[5]) );
  dff_sg \reg_www_1_reg[5]  ( .D(n4683), .CP(clk), .Q(reg_www_1[5]) );
  dff_sg \reg_w_1_reg[4]  ( .D(n5636), .CP(clk), .Q(reg_w_1[4]) );
  dff_sg \reg_ww_1_reg[4]  ( .D(n4704), .CP(clk), .Q(reg_ww_1[4]) );
  dff_sg \reg_www_1_reg[4]  ( .D(n4684), .CP(clk), .Q(reg_www_1[4]) );
  dff_sg \reg_w_1_reg[3]  ( .D(n5637), .CP(clk), .Q(reg_w_1[3]) );
  dff_sg \reg_ww_1_reg[3]  ( .D(n4705), .CP(clk), .Q(reg_ww_1[3]) );
  dff_sg \reg_www_1_reg[3]  ( .D(n4685), .CP(clk), .Q(reg_www_1[3]) );
  dff_sg \reg_w_1_reg[2]  ( .D(n5638), .CP(clk), .Q(reg_w_1[2]) );
  dff_sg \reg_ww_1_reg[2]  ( .D(n4706), .CP(clk), .Q(reg_ww_1[2]) );
  dff_sg \reg_www_1_reg[2]  ( .D(n4686), .CP(clk), .Q(reg_www_1[2]) );
  dff_sg \reg_w_1_reg[1]  ( .D(n5639), .CP(clk), .Q(reg_w_1[1]) );
  dff_sg \reg_ww_1_reg[1]  ( .D(n4707), .CP(clk), .Q(reg_ww_1[1]) );
  dff_sg \reg_www_1_reg[1]  ( .D(n4687), .CP(clk), .Q(reg_www_1[1]) );
  dff_sg \reg_w_1_reg[0]  ( .D(n5640), .CP(clk), .Q(reg_w_1[0]) );
  dff_sg \reg_ww_1_reg[0]  ( .D(n4708), .CP(clk), .Q(reg_ww_1[0]) );
  dff_sg \reg_www_1_reg[0]  ( .D(n4688), .CP(clk), .Q(reg_www_1[0]) );
  dff_sg \reg_w_0_reg[19]  ( .D(n5641), .CP(clk), .Q(reg_w_0[19]) );
  dff_sg \reg_ww_0_reg[19]  ( .D(n4729), .CP(clk), .Q(reg_ww_0[19]) );
  dff_sg \reg_www_0_reg[19]  ( .D(n4709), .CP(clk), .Q(reg_www_0[19]) );
  dff_sg \reg_w_0_reg[18]  ( .D(n5642), .CP(clk), .Q(reg_w_0[18]) );
  dff_sg \reg_ww_0_reg[18]  ( .D(n4730), .CP(clk), .Q(reg_ww_0[18]) );
  dff_sg \reg_www_0_reg[18]  ( .D(n4710), .CP(clk), .Q(reg_www_0[18]) );
  dff_sg \reg_w_0_reg[17]  ( .D(n5643), .CP(clk), .Q(reg_w_0[17]) );
  dff_sg \reg_ww_0_reg[17]  ( .D(n4731), .CP(clk), .Q(reg_ww_0[17]) );
  dff_sg \reg_www_0_reg[17]  ( .D(n4711), .CP(clk), .Q(reg_www_0[17]) );
  dff_sg \reg_w_0_reg[16]  ( .D(n5644), .CP(clk), .Q(reg_w_0[16]) );
  dff_sg \reg_ww_0_reg[16]  ( .D(n4732), .CP(clk), .Q(reg_ww_0[16]) );
  dff_sg \reg_www_0_reg[16]  ( .D(n4712), .CP(clk), .Q(reg_www_0[16]) );
  dff_sg \reg_w_0_reg[15]  ( .D(n5645), .CP(clk), .Q(reg_w_0[15]) );
  dff_sg \reg_ww_0_reg[15]  ( .D(n4733), .CP(clk), .Q(reg_ww_0[15]) );
  dff_sg \reg_www_0_reg[15]  ( .D(n4713), .CP(clk), .Q(reg_www_0[15]) );
  dff_sg \reg_w_0_reg[14]  ( .D(n5646), .CP(clk), .Q(reg_w_0[14]) );
  dff_sg \reg_ww_0_reg[14]  ( .D(n4734), .CP(clk), .Q(reg_ww_0[14]) );
  dff_sg \reg_www_0_reg[14]  ( .D(n4714), .CP(clk), .Q(reg_www_0[14]) );
  dff_sg \reg_w_0_reg[13]  ( .D(n5647), .CP(clk), .Q(reg_w_0[13]) );
  dff_sg \reg_ww_0_reg[13]  ( .D(n4735), .CP(clk), .Q(reg_ww_0[13]) );
  dff_sg \reg_www_0_reg[13]  ( .D(n4715), .CP(clk), .Q(reg_www_0[13]) );
  dff_sg \reg_w_0_reg[12]  ( .D(n5648), .CP(clk), .Q(reg_w_0[12]) );
  dff_sg \reg_ww_0_reg[12]  ( .D(n4736), .CP(clk), .Q(reg_ww_0[12]) );
  dff_sg \reg_www_0_reg[12]  ( .D(n4716), .CP(clk), .Q(reg_www_0[12]) );
  dff_sg \reg_w_0_reg[11]  ( .D(n5649), .CP(clk), .Q(reg_w_0[11]) );
  dff_sg \reg_ww_0_reg[11]  ( .D(n4737), .CP(clk), .Q(reg_ww_0[11]) );
  dff_sg \reg_www_0_reg[11]  ( .D(n4717), .CP(clk), .Q(reg_www_0[11]) );
  dff_sg \reg_w_0_reg[10]  ( .D(n5650), .CP(clk), .Q(reg_w_0[10]) );
  dff_sg \reg_ww_0_reg[10]  ( .D(n4738), .CP(clk), .Q(reg_ww_0[10]) );
  dff_sg \reg_www_0_reg[10]  ( .D(n4718), .CP(clk), .Q(reg_www_0[10]) );
  dff_sg \reg_w_0_reg[9]  ( .D(n5651), .CP(clk), .Q(reg_w_0[9]) );
  dff_sg \reg_ww_0_reg[9]  ( .D(n4739), .CP(clk), .Q(reg_ww_0[9]) );
  dff_sg \reg_www_0_reg[9]  ( .D(n4719), .CP(clk), .Q(reg_www_0[9]) );
  dff_sg \reg_w_0_reg[8]  ( .D(n5652), .CP(clk), .Q(reg_w_0[8]) );
  dff_sg \reg_ww_0_reg[8]  ( .D(n4740), .CP(clk), .Q(reg_ww_0[8]) );
  dff_sg \reg_www_0_reg[8]  ( .D(n4720), .CP(clk), .Q(reg_www_0[8]) );
  dff_sg \reg_w_0_reg[7]  ( .D(n5653), .CP(clk), .Q(reg_w_0[7]) );
  dff_sg \reg_ww_0_reg[7]  ( .D(n4741), .CP(clk), .Q(reg_ww_0[7]) );
  dff_sg \reg_www_0_reg[7]  ( .D(n4721), .CP(clk), .Q(reg_www_0[7]) );
  dff_sg \reg_w_0_reg[6]  ( .D(n5654), .CP(clk), .Q(reg_w_0[6]) );
  dff_sg \reg_ww_0_reg[6]  ( .D(n4742), .CP(clk), .Q(reg_ww_0[6]) );
  dff_sg \reg_www_0_reg[6]  ( .D(n4722), .CP(clk), .Q(reg_www_0[6]) );
  dff_sg \reg_w_0_reg[5]  ( .D(n5655), .CP(clk), .Q(reg_w_0[5]) );
  dff_sg \reg_ww_0_reg[5]  ( .D(n4743), .CP(clk), .Q(reg_ww_0[5]) );
  dff_sg \reg_www_0_reg[5]  ( .D(n4723), .CP(clk), .Q(reg_www_0[5]) );
  dff_sg \reg_w_0_reg[4]  ( .D(n5656), .CP(clk), .Q(reg_w_0[4]) );
  dff_sg \reg_ww_0_reg[4]  ( .D(n4744), .CP(clk), .Q(reg_ww_0[4]) );
  dff_sg \reg_www_0_reg[4]  ( .D(n4724), .CP(clk), .Q(reg_www_0[4]) );
  dff_sg \reg_w_0_reg[3]  ( .D(n5657), .CP(clk), .Q(reg_w_0[3]) );
  dff_sg \reg_ww_0_reg[3]  ( .D(n4745), .CP(clk), .Q(reg_ww_0[3]) );
  dff_sg \reg_www_0_reg[3]  ( .D(n4725), .CP(clk), .Q(reg_www_0[3]) );
  dff_sg \reg_w_0_reg[2]  ( .D(n5658), .CP(clk), .Q(reg_w_0[2]) );
  dff_sg \reg_ww_0_reg[2]  ( .D(n4746), .CP(clk), .Q(reg_ww_0[2]) );
  dff_sg \reg_www_0_reg[2]  ( .D(n4726), .CP(clk), .Q(reg_www_0[2]) );
  dff_sg \reg_w_0_reg[1]  ( .D(n5659), .CP(clk), .Q(reg_w_0[1]) );
  dff_sg \reg_ww_0_reg[1]  ( .D(n4747), .CP(clk), .Q(reg_ww_0[1]) );
  dff_sg \reg_www_0_reg[1]  ( .D(n4727), .CP(clk), .Q(reg_www_0[1]) );
  dff_sg \reg_w_0_reg[0]  ( .D(n5660), .CP(clk), .Q(reg_w_0[0]) );
  dff_sg \reg_ww_0_reg[0]  ( .D(n4748), .CP(clk), .Q(reg_ww_0[0]) );
  dff_sg \reg_www_0_reg[0]  ( .D(n4728), .CP(clk), .Q(reg_www_0[0]) );
  dff_sg \reg_i_15_reg[19]  ( .D(n5661), .CP(clk), .Q(reg_i_15[19]) );
  dff_sg \reg_ii_15_reg[19]  ( .D(n4769), .CP(clk), .Q(reg_ii_15[19]) );
  dff_sg \reg_iii_15_reg[19]  ( .D(n4749), .CP(clk), .Q(reg_iii_15[19]) );
  dff_sg \reg_i_15_reg[18]  ( .D(n5662), .CP(clk), .Q(reg_i_15[18]) );
  dff_sg \reg_ii_15_reg[18]  ( .D(n4770), .CP(clk), .Q(reg_ii_15[18]) );
  dff_sg \reg_iii_15_reg[18]  ( .D(n4750), .CP(clk), .Q(reg_iii_15[18]) );
  dff_sg \reg_i_15_reg[17]  ( .D(n5663), .CP(clk), .Q(reg_i_15[17]) );
  dff_sg \reg_ii_15_reg[17]  ( .D(n4771), .CP(clk), .Q(reg_ii_15[17]) );
  dff_sg \reg_iii_15_reg[17]  ( .D(n4751), .CP(clk), .Q(reg_iii_15[17]) );
  dff_sg \reg_i_15_reg[16]  ( .D(n5664), .CP(clk), .Q(reg_i_15[16]) );
  dff_sg \reg_ii_15_reg[16]  ( .D(n4772), .CP(clk), .Q(reg_ii_15[16]) );
  dff_sg \reg_iii_15_reg[16]  ( .D(n4752), .CP(clk), .Q(reg_iii_15[16]) );
  dff_sg \reg_i_15_reg[15]  ( .D(n5665), .CP(clk), .Q(reg_i_15[15]) );
  dff_sg \reg_ii_15_reg[15]  ( .D(n4773), .CP(clk), .Q(reg_ii_15[15]) );
  dff_sg \reg_iii_15_reg[15]  ( .D(n4753), .CP(clk), .Q(reg_iii_15[15]) );
  dff_sg \reg_i_15_reg[14]  ( .D(n5666), .CP(clk), .Q(reg_i_15[14]) );
  dff_sg \reg_ii_15_reg[14]  ( .D(n4774), .CP(clk), .Q(reg_ii_15[14]) );
  dff_sg \reg_iii_15_reg[14]  ( .D(n4754), .CP(clk), .Q(reg_iii_15[14]) );
  dff_sg \reg_i_15_reg[13]  ( .D(n5667), .CP(clk), .Q(reg_i_15[13]) );
  dff_sg \reg_ii_15_reg[13]  ( .D(n4775), .CP(clk), .Q(reg_ii_15[13]) );
  dff_sg \reg_iii_15_reg[13]  ( .D(n4755), .CP(clk), .Q(reg_iii_15[13]) );
  dff_sg \reg_i_15_reg[12]  ( .D(n5668), .CP(clk), .Q(reg_i_15[12]) );
  dff_sg \reg_ii_15_reg[12]  ( .D(n4776), .CP(clk), .Q(reg_ii_15[12]) );
  dff_sg \reg_iii_15_reg[12]  ( .D(n4756), .CP(clk), .Q(reg_iii_15[12]) );
  dff_sg \reg_i_15_reg[11]  ( .D(n5669), .CP(clk), .Q(reg_i_15[11]) );
  dff_sg \reg_ii_15_reg[11]  ( .D(n4777), .CP(clk), .Q(reg_ii_15[11]) );
  dff_sg \reg_iii_15_reg[11]  ( .D(n4757), .CP(clk), .Q(reg_iii_15[11]) );
  dff_sg \reg_i_15_reg[10]  ( .D(n5670), .CP(clk), .Q(reg_i_15[10]) );
  dff_sg \reg_ii_15_reg[10]  ( .D(n4778), .CP(clk), .Q(reg_ii_15[10]) );
  dff_sg \reg_iii_15_reg[10]  ( .D(n4758), .CP(clk), .Q(reg_iii_15[10]) );
  dff_sg \reg_i_15_reg[9]  ( .D(n5671), .CP(clk), .Q(reg_i_15[9]) );
  dff_sg \reg_ii_15_reg[9]  ( .D(n4779), .CP(clk), .Q(reg_ii_15[9]) );
  dff_sg \reg_iii_15_reg[9]  ( .D(n4759), .CP(clk), .Q(reg_iii_15[9]) );
  dff_sg \reg_i_15_reg[8]  ( .D(n5672), .CP(clk), .Q(reg_i_15[8]) );
  dff_sg \reg_ii_15_reg[8]  ( .D(n4780), .CP(clk), .Q(reg_ii_15[8]) );
  dff_sg \reg_iii_15_reg[8]  ( .D(n4760), .CP(clk), .Q(reg_iii_15[8]) );
  dff_sg \reg_i_15_reg[7]  ( .D(n5673), .CP(clk), .Q(reg_i_15[7]) );
  dff_sg \reg_ii_15_reg[7]  ( .D(n4781), .CP(clk), .Q(reg_ii_15[7]) );
  dff_sg \reg_iii_15_reg[7]  ( .D(n4761), .CP(clk), .Q(reg_iii_15[7]) );
  dff_sg \reg_i_15_reg[6]  ( .D(n5674), .CP(clk), .Q(reg_i_15[6]) );
  dff_sg \reg_ii_15_reg[6]  ( .D(n4782), .CP(clk), .Q(reg_ii_15[6]) );
  dff_sg \reg_iii_15_reg[6]  ( .D(n4762), .CP(clk), .Q(reg_iii_15[6]) );
  dff_sg \reg_i_15_reg[5]  ( .D(n5675), .CP(clk), .Q(reg_i_15[5]) );
  dff_sg \reg_ii_15_reg[5]  ( .D(n4783), .CP(clk), .Q(reg_ii_15[5]) );
  dff_sg \reg_iii_15_reg[5]  ( .D(n4763), .CP(clk), .Q(reg_iii_15[5]) );
  dff_sg \reg_i_15_reg[4]  ( .D(n5676), .CP(clk), .Q(reg_i_15[4]) );
  dff_sg \reg_ii_15_reg[4]  ( .D(n4784), .CP(clk), .Q(reg_ii_15[4]) );
  dff_sg \reg_iii_15_reg[4]  ( .D(n4764), .CP(clk), .Q(reg_iii_15[4]) );
  dff_sg \reg_i_15_reg[3]  ( .D(n5677), .CP(clk), .Q(reg_i_15[3]) );
  dff_sg \reg_ii_15_reg[3]  ( .D(n4785), .CP(clk), .Q(reg_ii_15[3]) );
  dff_sg \reg_iii_15_reg[3]  ( .D(n4765), .CP(clk), .Q(reg_iii_15[3]) );
  dff_sg \reg_i_15_reg[2]  ( .D(n5678), .CP(clk), .Q(reg_i_15[2]) );
  dff_sg \reg_ii_15_reg[2]  ( .D(n4786), .CP(clk), .Q(reg_ii_15[2]) );
  dff_sg \reg_iii_15_reg[2]  ( .D(n4766), .CP(clk), .Q(reg_iii_15[2]) );
  dff_sg \reg_i_15_reg[1]  ( .D(n5679), .CP(clk), .Q(reg_i_15[1]) );
  dff_sg \reg_ii_15_reg[1]  ( .D(n4787), .CP(clk), .Q(reg_ii_15[1]) );
  dff_sg \reg_iii_15_reg[1]  ( .D(n4767), .CP(clk), .Q(reg_iii_15[1]) );
  dff_sg \reg_i_15_reg[0]  ( .D(n5680), .CP(clk), .Q(reg_i_15[0]) );
  dff_sg \reg_ii_15_reg[0]  ( .D(n4788), .CP(clk), .Q(reg_ii_15[0]) );
  dff_sg \reg_iii_15_reg[0]  ( .D(n4768), .CP(clk), .Q(reg_iii_15[0]) );
  dff_sg \reg_i_14_reg[19]  ( .D(n5681), .CP(clk), .Q(reg_i_14[19]) );
  dff_sg \reg_ii_14_reg[19]  ( .D(n4789), .CP(clk), .Q(reg_ii_14[19]) );
  dff_sg \reg_iii_14_reg[19]  ( .D(n4394), .CP(clk), .Q(reg_iii_14[19]) );
  dff_sg \reg_i_14_reg[18]  ( .D(n5682), .CP(clk), .Q(reg_i_14[18]) );
  dff_sg \reg_ii_14_reg[18]  ( .D(n4790), .CP(clk), .Q(reg_ii_14[18]) );
  dff_sg \reg_iii_14_reg[18]  ( .D(n4395), .CP(clk), .Q(reg_iii_14[18]) );
  dff_sg \reg_i_14_reg[17]  ( .D(n5683), .CP(clk), .Q(reg_i_14[17]) );
  dff_sg \reg_ii_14_reg[17]  ( .D(n4791), .CP(clk), .Q(reg_ii_14[17]) );
  dff_sg \reg_iii_14_reg[17]  ( .D(n4396), .CP(clk), .Q(reg_iii_14[17]) );
  dff_sg \reg_i_14_reg[16]  ( .D(n5684), .CP(clk), .Q(reg_i_14[16]) );
  dff_sg \reg_ii_14_reg[16]  ( .D(n4414), .CP(clk), .Q(reg_ii_14[16]) );
  dff_sg \reg_iii_14_reg[16]  ( .D(n4397), .CP(clk), .Q(reg_iii_14[16]) );
  dff_sg \reg_i_14_reg[15]  ( .D(n5685), .CP(clk), .Q(reg_i_14[15]) );
  dff_sg \reg_ii_14_reg[15]  ( .D(n4415), .CP(clk), .Q(reg_ii_14[15]) );
  dff_sg \reg_iii_14_reg[15]  ( .D(n4398), .CP(clk), .Q(reg_iii_14[15]) );
  dff_sg \reg_i_14_reg[14]  ( .D(n5686), .CP(clk), .Q(reg_i_14[14]) );
  dff_sg \reg_ii_14_reg[14]  ( .D(n4416), .CP(clk), .Q(reg_ii_14[14]) );
  dff_sg \reg_iii_14_reg[14]  ( .D(n4399), .CP(clk), .Q(reg_iii_14[14]) );
  dff_sg \reg_i_14_reg[13]  ( .D(n5687), .CP(clk), .Q(reg_i_14[13]) );
  dff_sg \reg_ii_14_reg[13]  ( .D(n4417), .CP(clk), .Q(reg_ii_14[13]) );
  dff_sg \reg_iii_14_reg[13]  ( .D(n4400), .CP(clk), .Q(reg_iii_14[13]) );
  dff_sg \reg_i_14_reg[12]  ( .D(n5688), .CP(clk), .Q(reg_i_14[12]) );
  dff_sg \reg_ii_14_reg[12]  ( .D(n4418), .CP(clk), .Q(reg_ii_14[12]) );
  dff_sg \reg_iii_14_reg[12]  ( .D(n4401), .CP(clk), .Q(reg_iii_14[12]) );
  dff_sg \reg_i_14_reg[11]  ( .D(n5689), .CP(clk), .Q(reg_i_14[11]) );
  dff_sg \reg_ii_14_reg[11]  ( .D(n4419), .CP(clk), .Q(reg_ii_14[11]) );
  dff_sg \reg_iii_14_reg[11]  ( .D(n4402), .CP(clk), .Q(reg_iii_14[11]) );
  dff_sg \reg_i_14_reg[10]  ( .D(n5690), .CP(clk), .Q(reg_i_14[10]) );
  dff_sg \reg_ii_14_reg[10]  ( .D(n4420), .CP(clk), .Q(reg_ii_14[10]) );
  dff_sg \reg_iii_14_reg[10]  ( .D(n4403), .CP(clk), .Q(reg_iii_14[10]) );
  dff_sg \reg_i_14_reg[9]  ( .D(n5691), .CP(clk), .Q(reg_i_14[9]) );
  dff_sg \reg_ii_14_reg[9]  ( .D(n4421), .CP(clk), .Q(reg_ii_14[9]) );
  dff_sg \reg_iii_14_reg[9]  ( .D(n4404), .CP(clk), .Q(reg_iii_14[9]) );
  dff_sg \reg_i_14_reg[8]  ( .D(n5692), .CP(clk), .Q(reg_i_14[8]) );
  dff_sg \reg_ii_14_reg[8]  ( .D(n4422), .CP(clk), .Q(reg_ii_14[8]) );
  dff_sg \reg_iii_14_reg[8]  ( .D(n4405), .CP(clk), .Q(reg_iii_14[8]) );
  dff_sg \reg_i_14_reg[7]  ( .D(n5693), .CP(clk), .Q(reg_i_14[7]) );
  dff_sg \reg_ii_14_reg[7]  ( .D(n4423), .CP(clk), .Q(reg_ii_14[7]) );
  dff_sg \reg_iii_14_reg[7]  ( .D(n4406), .CP(clk), .Q(reg_iii_14[7]) );
  dff_sg \reg_i_14_reg[6]  ( .D(n5694), .CP(clk), .Q(reg_i_14[6]) );
  dff_sg \reg_ii_14_reg[6]  ( .D(n4424), .CP(clk), .Q(reg_ii_14[6]) );
  dff_sg \reg_iii_14_reg[6]  ( .D(n4407), .CP(clk), .Q(reg_iii_14[6]) );
  dff_sg \reg_i_14_reg[5]  ( .D(n5695), .CP(clk), .Q(reg_i_14[5]) );
  dff_sg \reg_ii_14_reg[5]  ( .D(n4425), .CP(clk), .Q(reg_ii_14[5]) );
  dff_sg \reg_iii_14_reg[5]  ( .D(n4408), .CP(clk), .Q(reg_iii_14[5]) );
  dff_sg \reg_i_14_reg[4]  ( .D(n5696), .CP(clk), .Q(reg_i_14[4]) );
  dff_sg \reg_ii_14_reg[4]  ( .D(n4426), .CP(clk), .Q(reg_ii_14[4]) );
  dff_sg \reg_iii_14_reg[4]  ( .D(n4409), .CP(clk), .Q(reg_iii_14[4]) );
  dff_sg \reg_i_14_reg[3]  ( .D(n5697), .CP(clk), .Q(reg_i_14[3]) );
  dff_sg \reg_ii_14_reg[3]  ( .D(n4427), .CP(clk), .Q(reg_ii_14[3]) );
  dff_sg \reg_iii_14_reg[3]  ( .D(n4410), .CP(clk), .Q(reg_iii_14[3]) );
  dff_sg \reg_i_14_reg[2]  ( .D(n5698), .CP(clk), .Q(reg_i_14[2]) );
  dff_sg \reg_ii_14_reg[2]  ( .D(n4428), .CP(clk), .Q(reg_ii_14[2]) );
  dff_sg \reg_iii_14_reg[2]  ( .D(n4411), .CP(clk), .Q(reg_iii_14[2]) );
  dff_sg \reg_i_14_reg[1]  ( .D(n5699), .CP(clk), .Q(reg_i_14[1]) );
  dff_sg \reg_ii_14_reg[1]  ( .D(n4429), .CP(clk), .Q(reg_ii_14[1]) );
  dff_sg \reg_iii_14_reg[1]  ( .D(n4412), .CP(clk), .Q(reg_iii_14[1]) );
  dff_sg \reg_i_14_reg[0]  ( .D(n5700), .CP(clk), .Q(reg_i_14[0]) );
  dff_sg \reg_ii_14_reg[0]  ( .D(n4430), .CP(clk), .Q(reg_ii_14[0]) );
  dff_sg \reg_iii_14_reg[0]  ( .D(n4413), .CP(clk), .Q(reg_iii_14[0]) );
  dff_sg \reg_i_13_reg[19]  ( .D(n5701), .CP(clk), .Q(reg_i_13[19]) );
  dff_sg \reg_ii_13_reg[19]  ( .D(n4451), .CP(clk), .Q(reg_ii_13[19]) );
  dff_sg \reg_iii_13_reg[19]  ( .D(n4431), .CP(clk), .Q(reg_iii_13[19]) );
  dff_sg \reg_i_13_reg[18]  ( .D(n5702), .CP(clk), .Q(reg_i_13[18]) );
  dff_sg \reg_ii_13_reg[18]  ( .D(n4452), .CP(clk), .Q(reg_ii_13[18]) );
  dff_sg \reg_iii_13_reg[18]  ( .D(n4432), .CP(clk), .Q(reg_iii_13[18]) );
  dff_sg \reg_i_13_reg[17]  ( .D(n5703), .CP(clk), .Q(reg_i_13[17]) );
  dff_sg \reg_ii_13_reg[17]  ( .D(n4453), .CP(clk), .Q(reg_ii_13[17]) );
  dff_sg \reg_iii_13_reg[17]  ( .D(n4433), .CP(clk), .Q(reg_iii_13[17]) );
  dff_sg \reg_i_13_reg[16]  ( .D(n5704), .CP(clk), .Q(reg_i_13[16]) );
  dff_sg \reg_ii_13_reg[16]  ( .D(n4454), .CP(clk), .Q(reg_ii_13[16]) );
  dff_sg \reg_iii_13_reg[16]  ( .D(n4434), .CP(clk), .Q(reg_iii_13[16]) );
  dff_sg \reg_i_13_reg[15]  ( .D(n5705), .CP(clk), .Q(reg_i_13[15]) );
  dff_sg \reg_ii_13_reg[15]  ( .D(n4455), .CP(clk), .Q(reg_ii_13[15]) );
  dff_sg \reg_iii_13_reg[15]  ( .D(n4435), .CP(clk), .Q(reg_iii_13[15]) );
  dff_sg \reg_i_13_reg[14]  ( .D(n5706), .CP(clk), .Q(reg_i_13[14]) );
  dff_sg \reg_ii_13_reg[14]  ( .D(n4456), .CP(clk), .Q(reg_ii_13[14]) );
  dff_sg \reg_iii_13_reg[14]  ( .D(n4436), .CP(clk), .Q(reg_iii_13[14]) );
  dff_sg \reg_i_13_reg[13]  ( .D(n5707), .CP(clk), .Q(reg_i_13[13]) );
  dff_sg \reg_ii_13_reg[13]  ( .D(n4457), .CP(clk), .Q(reg_ii_13[13]) );
  dff_sg \reg_iii_13_reg[13]  ( .D(n4437), .CP(clk), .Q(reg_iii_13[13]) );
  dff_sg \reg_i_13_reg[12]  ( .D(n5708), .CP(clk), .Q(reg_i_13[12]) );
  dff_sg \reg_ii_13_reg[12]  ( .D(n4458), .CP(clk), .Q(reg_ii_13[12]) );
  dff_sg \reg_iii_13_reg[12]  ( .D(n4438), .CP(clk), .Q(reg_iii_13[12]) );
  dff_sg \reg_i_13_reg[11]  ( .D(n5709), .CP(clk), .Q(reg_i_13[11]) );
  dff_sg \reg_ii_13_reg[11]  ( .D(n4459), .CP(clk), .Q(reg_ii_13[11]) );
  dff_sg \reg_iii_13_reg[11]  ( .D(n4439), .CP(clk), .Q(reg_iii_13[11]) );
  dff_sg \reg_i_13_reg[10]  ( .D(n5710), .CP(clk), .Q(reg_i_13[10]) );
  dff_sg \reg_ii_13_reg[10]  ( .D(n4460), .CP(clk), .Q(reg_ii_13[10]) );
  dff_sg \reg_iii_13_reg[10]  ( .D(n4440), .CP(clk), .Q(reg_iii_13[10]) );
  dff_sg \reg_i_13_reg[9]  ( .D(n5711), .CP(clk), .Q(reg_i_13[9]) );
  dff_sg \reg_ii_13_reg[9]  ( .D(n4461), .CP(clk), .Q(reg_ii_13[9]) );
  dff_sg \reg_iii_13_reg[9]  ( .D(n4441), .CP(clk), .Q(reg_iii_13[9]) );
  dff_sg \reg_i_13_reg[8]  ( .D(n5712), .CP(clk), .Q(reg_i_13[8]) );
  dff_sg \reg_ii_13_reg[8]  ( .D(n4462), .CP(clk), .Q(reg_ii_13[8]) );
  dff_sg \reg_iii_13_reg[8]  ( .D(n4442), .CP(clk), .Q(reg_iii_13[8]) );
  dff_sg \reg_i_13_reg[7]  ( .D(n5713), .CP(clk), .Q(reg_i_13[7]) );
  dff_sg \reg_ii_13_reg[7]  ( .D(n4463), .CP(clk), .Q(reg_ii_13[7]) );
  dff_sg \reg_iii_13_reg[7]  ( .D(n4443), .CP(clk), .Q(reg_iii_13[7]) );
  dff_sg \reg_i_13_reg[6]  ( .D(n5714), .CP(clk), .Q(reg_i_13[6]) );
  dff_sg \reg_ii_13_reg[6]  ( .D(n4464), .CP(clk), .Q(reg_ii_13[6]) );
  dff_sg \reg_iii_13_reg[6]  ( .D(n4444), .CP(clk), .Q(reg_iii_13[6]) );
  dff_sg \reg_i_13_reg[5]  ( .D(n5715), .CP(clk), .Q(reg_i_13[5]) );
  dff_sg \reg_ii_13_reg[5]  ( .D(n4465), .CP(clk), .Q(reg_ii_13[5]) );
  dff_sg \reg_iii_13_reg[5]  ( .D(n4445), .CP(clk), .Q(reg_iii_13[5]) );
  dff_sg \reg_i_13_reg[4]  ( .D(n5716), .CP(clk), .Q(reg_i_13[4]) );
  dff_sg \reg_ii_13_reg[4]  ( .D(n4466), .CP(clk), .Q(reg_ii_13[4]) );
  dff_sg \reg_iii_13_reg[4]  ( .D(n4446), .CP(clk), .Q(reg_iii_13[4]) );
  dff_sg \reg_i_13_reg[3]  ( .D(n5717), .CP(clk), .Q(reg_i_13[3]) );
  dff_sg \reg_ii_13_reg[3]  ( .D(n4467), .CP(clk), .Q(reg_ii_13[3]) );
  dff_sg \reg_iii_13_reg[3]  ( .D(n4447), .CP(clk), .Q(reg_iii_13[3]) );
  dff_sg \reg_i_13_reg[2]  ( .D(n5718), .CP(clk), .Q(reg_i_13[2]) );
  dff_sg \reg_ii_13_reg[2]  ( .D(n4468), .CP(clk), .Q(reg_ii_13[2]) );
  dff_sg \reg_iii_13_reg[2]  ( .D(n4448), .CP(clk), .Q(reg_iii_13[2]) );
  dff_sg \reg_i_13_reg[1]  ( .D(n5719), .CP(clk), .Q(reg_i_13[1]) );
  dff_sg \reg_ii_13_reg[1]  ( .D(n4469), .CP(clk), .Q(reg_ii_13[1]) );
  dff_sg \reg_iii_13_reg[1]  ( .D(n4449), .CP(clk), .Q(reg_iii_13[1]) );
  dff_sg \reg_i_13_reg[0]  ( .D(n5720), .CP(clk), .Q(reg_i_13[0]) );
  dff_sg \reg_ii_13_reg[0]  ( .D(n4470), .CP(clk), .Q(reg_ii_13[0]) );
  dff_sg \reg_iii_13_reg[0]  ( .D(n4450), .CP(clk), .Q(reg_iii_13[0]) );
  dff_sg \reg_i_12_reg[19]  ( .D(n5721), .CP(clk), .Q(reg_i_12[19]) );
  dff_sg \reg_ii_12_reg[19]  ( .D(n4491), .CP(clk), .Q(reg_ii_12[19]) );
  dff_sg \reg_iii_12_reg[19]  ( .D(n4471), .CP(clk), .Q(reg_iii_12[19]) );
  dff_sg \reg_i_12_reg[18]  ( .D(n5722), .CP(clk), .Q(reg_i_12[18]) );
  dff_sg \reg_ii_12_reg[18]  ( .D(n4492), .CP(clk), .Q(reg_ii_12[18]) );
  dff_sg \reg_iii_12_reg[18]  ( .D(n4472), .CP(clk), .Q(reg_iii_12[18]) );
  dff_sg \reg_i_12_reg[17]  ( .D(n5723), .CP(clk), .Q(reg_i_12[17]) );
  dff_sg \reg_ii_12_reg[17]  ( .D(n4493), .CP(clk), .Q(reg_ii_12[17]) );
  dff_sg \reg_iii_12_reg[17]  ( .D(n4473), .CP(clk), .Q(reg_iii_12[17]) );
  dff_sg \reg_i_12_reg[16]  ( .D(n5724), .CP(clk), .Q(reg_i_12[16]) );
  dff_sg \reg_ii_12_reg[16]  ( .D(n4494), .CP(clk), .Q(reg_ii_12[16]) );
  dff_sg \reg_iii_12_reg[16]  ( .D(n4474), .CP(clk), .Q(reg_iii_12[16]) );
  dff_sg \reg_i_12_reg[15]  ( .D(n5725), .CP(clk), .Q(reg_i_12[15]) );
  dff_sg \reg_ii_12_reg[15]  ( .D(n4495), .CP(clk), .Q(reg_ii_12[15]) );
  dff_sg \reg_iii_12_reg[15]  ( .D(n4475), .CP(clk), .Q(reg_iii_12[15]) );
  dff_sg \reg_i_12_reg[14]  ( .D(n5726), .CP(clk), .Q(reg_i_12[14]) );
  dff_sg \reg_ii_12_reg[14]  ( .D(n4496), .CP(clk), .Q(reg_ii_12[14]) );
  dff_sg \reg_iii_12_reg[14]  ( .D(n4476), .CP(clk), .Q(reg_iii_12[14]) );
  dff_sg \reg_i_12_reg[13]  ( .D(n5727), .CP(clk), .Q(reg_i_12[13]) );
  dff_sg \reg_ii_12_reg[13]  ( .D(n4497), .CP(clk), .Q(reg_ii_12[13]) );
  dff_sg \reg_iii_12_reg[13]  ( .D(n4477), .CP(clk), .Q(reg_iii_12[13]) );
  dff_sg \reg_i_12_reg[12]  ( .D(n5728), .CP(clk), .Q(reg_i_12[12]) );
  dff_sg \reg_ii_12_reg[12]  ( .D(n4498), .CP(clk), .Q(reg_ii_12[12]) );
  dff_sg \reg_iii_12_reg[12]  ( .D(n4478), .CP(clk), .Q(reg_iii_12[12]) );
  dff_sg \reg_i_12_reg[11]  ( .D(n5729), .CP(clk), .Q(reg_i_12[11]) );
  dff_sg \reg_ii_12_reg[11]  ( .D(n4499), .CP(clk), .Q(reg_ii_12[11]) );
  dff_sg \reg_iii_12_reg[11]  ( .D(n4479), .CP(clk), .Q(reg_iii_12[11]) );
  dff_sg \reg_i_12_reg[10]  ( .D(n5730), .CP(clk), .Q(reg_i_12[10]) );
  dff_sg \reg_ii_12_reg[10]  ( .D(n4500), .CP(clk), .Q(reg_ii_12[10]) );
  dff_sg \reg_iii_12_reg[10]  ( .D(n4480), .CP(clk), .Q(reg_iii_12[10]) );
  dff_sg \reg_i_12_reg[9]  ( .D(n5731), .CP(clk), .Q(reg_i_12[9]) );
  dff_sg \reg_ii_12_reg[9]  ( .D(n4501), .CP(clk), .Q(reg_ii_12[9]) );
  dff_sg \reg_iii_12_reg[9]  ( .D(n4481), .CP(clk), .Q(reg_iii_12[9]) );
  dff_sg \reg_i_12_reg[8]  ( .D(n5732), .CP(clk), .Q(reg_i_12[8]) );
  dff_sg \reg_ii_12_reg[8]  ( .D(n4502), .CP(clk), .Q(reg_ii_12[8]) );
  dff_sg \reg_iii_12_reg[8]  ( .D(n4482), .CP(clk), .Q(reg_iii_12[8]) );
  dff_sg \reg_i_12_reg[7]  ( .D(n5733), .CP(clk), .Q(reg_i_12[7]) );
  dff_sg \reg_ii_12_reg[7]  ( .D(n4503), .CP(clk), .Q(reg_ii_12[7]) );
  dff_sg \reg_iii_12_reg[7]  ( .D(n4483), .CP(clk), .Q(reg_iii_12[7]) );
  dff_sg \reg_i_12_reg[6]  ( .D(n5734), .CP(clk), .Q(reg_i_12[6]) );
  dff_sg \reg_ii_12_reg[6]  ( .D(n4504), .CP(clk), .Q(reg_ii_12[6]) );
  dff_sg \reg_iii_12_reg[6]  ( .D(n4484), .CP(clk), .Q(reg_iii_12[6]) );
  dff_sg \reg_i_12_reg[5]  ( .D(n5735), .CP(clk), .Q(reg_i_12[5]) );
  dff_sg \reg_ii_12_reg[5]  ( .D(n4505), .CP(clk), .Q(reg_ii_12[5]) );
  dff_sg \reg_iii_12_reg[5]  ( .D(n4485), .CP(clk), .Q(reg_iii_12[5]) );
  dff_sg \reg_i_12_reg[4]  ( .D(n5736), .CP(clk), .Q(reg_i_12[4]) );
  dff_sg \reg_ii_12_reg[4]  ( .D(n4506), .CP(clk), .Q(reg_ii_12[4]) );
  dff_sg \reg_iii_12_reg[4]  ( .D(n4486), .CP(clk), .Q(reg_iii_12[4]) );
  dff_sg \reg_i_12_reg[3]  ( .D(n5737), .CP(clk), .Q(reg_i_12[3]) );
  dff_sg \reg_ii_12_reg[3]  ( .D(n4507), .CP(clk), .Q(reg_ii_12[3]) );
  dff_sg \reg_iii_12_reg[3]  ( .D(n4487), .CP(clk), .Q(reg_iii_12[3]) );
  dff_sg \reg_i_12_reg[2]  ( .D(n5738), .CP(clk), .Q(reg_i_12[2]) );
  dff_sg \reg_ii_12_reg[2]  ( .D(n4508), .CP(clk), .Q(reg_ii_12[2]) );
  dff_sg \reg_iii_12_reg[2]  ( .D(n4488), .CP(clk), .Q(reg_iii_12[2]) );
  dff_sg \reg_i_12_reg[1]  ( .D(n5739), .CP(clk), .Q(reg_i_12[1]) );
  dff_sg \reg_ii_12_reg[1]  ( .D(n4509), .CP(clk), .Q(reg_ii_12[1]) );
  dff_sg \reg_iii_12_reg[1]  ( .D(n4489), .CP(clk), .Q(reg_iii_12[1]) );
  dff_sg \reg_i_12_reg[0]  ( .D(n5740), .CP(clk), .Q(reg_i_12[0]) );
  dff_sg \reg_ii_12_reg[0]  ( .D(n4510), .CP(clk), .Q(reg_ii_12[0]) );
  dff_sg \reg_iii_12_reg[0]  ( .D(n4490), .CP(clk), .Q(reg_iii_12[0]) );
  dff_sg \reg_i_11_reg[19]  ( .D(n5741), .CP(clk), .Q(reg_i_11[19]) );
  dff_sg \reg_ii_11_reg[19]  ( .D(n4531), .CP(clk), .Q(reg_ii_11[19]) );
  dff_sg \reg_iii_11_reg[19]  ( .D(n4511), .CP(clk), .Q(reg_iii_11[19]) );
  dff_sg \reg_i_11_reg[18]  ( .D(n5742), .CP(clk), .Q(reg_i_11[18]) );
  dff_sg \reg_ii_11_reg[18]  ( .D(n4532), .CP(clk), .Q(reg_ii_11[18]) );
  dff_sg \reg_iii_11_reg[18]  ( .D(n4512), .CP(clk), .Q(reg_iii_11[18]) );
  dff_sg \reg_i_11_reg[17]  ( .D(n5743), .CP(clk), .Q(reg_i_11[17]) );
  dff_sg \reg_ii_11_reg[17]  ( .D(n4533), .CP(clk), .Q(reg_ii_11[17]) );
  dff_sg \reg_iii_11_reg[17]  ( .D(n4513), .CP(clk), .Q(reg_iii_11[17]) );
  dff_sg \reg_i_11_reg[16]  ( .D(n5744), .CP(clk), .Q(reg_i_11[16]) );
  dff_sg \reg_ii_11_reg[16]  ( .D(n4534), .CP(clk), .Q(reg_ii_11[16]) );
  dff_sg \reg_iii_11_reg[16]  ( .D(n4514), .CP(clk), .Q(reg_iii_11[16]) );
  dff_sg \reg_i_11_reg[15]  ( .D(n5745), .CP(clk), .Q(reg_i_11[15]) );
  dff_sg \reg_ii_11_reg[15]  ( .D(n4535), .CP(clk), .Q(reg_ii_11[15]) );
  dff_sg \reg_iii_11_reg[15]  ( .D(n4515), .CP(clk), .Q(reg_iii_11[15]) );
  dff_sg \reg_i_11_reg[14]  ( .D(n5746), .CP(clk), .Q(reg_i_11[14]) );
  dff_sg \reg_ii_11_reg[14]  ( .D(n4536), .CP(clk), .Q(reg_ii_11[14]) );
  dff_sg \reg_iii_11_reg[14]  ( .D(n4516), .CP(clk), .Q(reg_iii_11[14]) );
  dff_sg \reg_i_11_reg[13]  ( .D(n5747), .CP(clk), .Q(reg_i_11[13]) );
  dff_sg \reg_ii_11_reg[13]  ( .D(n4537), .CP(clk), .Q(reg_ii_11[13]) );
  dff_sg \reg_iii_11_reg[13]  ( .D(n4517), .CP(clk), .Q(reg_iii_11[13]) );
  dff_sg \reg_i_11_reg[12]  ( .D(n5748), .CP(clk), .Q(reg_i_11[12]) );
  dff_sg \reg_ii_11_reg[12]  ( .D(n4538), .CP(clk), .Q(reg_ii_11[12]) );
  dff_sg \reg_iii_11_reg[12]  ( .D(n4518), .CP(clk), .Q(reg_iii_11[12]) );
  dff_sg \reg_i_11_reg[11]  ( .D(n5749), .CP(clk), .Q(reg_i_11[11]) );
  dff_sg \reg_ii_11_reg[11]  ( .D(n4539), .CP(clk), .Q(reg_ii_11[11]) );
  dff_sg \reg_iii_11_reg[11]  ( .D(n4519), .CP(clk), .Q(reg_iii_11[11]) );
  dff_sg \reg_i_11_reg[10]  ( .D(n5750), .CP(clk), .Q(reg_i_11[10]) );
  dff_sg \reg_ii_11_reg[10]  ( .D(n4540), .CP(clk), .Q(reg_ii_11[10]) );
  dff_sg \reg_iii_11_reg[10]  ( .D(n4520), .CP(clk), .Q(reg_iii_11[10]) );
  dff_sg \reg_i_11_reg[9]  ( .D(n5751), .CP(clk), .Q(reg_i_11[9]) );
  dff_sg \reg_ii_11_reg[9]  ( .D(n4541), .CP(clk), .Q(reg_ii_11[9]) );
  dff_sg \reg_iii_11_reg[9]  ( .D(n4521), .CP(clk), .Q(reg_iii_11[9]) );
  dff_sg \reg_i_11_reg[8]  ( .D(n5752), .CP(clk), .Q(reg_i_11[8]) );
  dff_sg \reg_ii_11_reg[8]  ( .D(n4542), .CP(clk), .Q(reg_ii_11[8]) );
  dff_sg \reg_iii_11_reg[8]  ( .D(n4522), .CP(clk), .Q(reg_iii_11[8]) );
  dff_sg \reg_i_11_reg[7]  ( .D(n5753), .CP(clk), .Q(reg_i_11[7]) );
  dff_sg \reg_ii_11_reg[7]  ( .D(n4543), .CP(clk), .Q(reg_ii_11[7]) );
  dff_sg \reg_iii_11_reg[7]  ( .D(n4523), .CP(clk), .Q(reg_iii_11[7]) );
  dff_sg \reg_i_11_reg[6]  ( .D(n5754), .CP(clk), .Q(reg_i_11[6]) );
  dff_sg \reg_ii_11_reg[6]  ( .D(n4544), .CP(clk), .Q(reg_ii_11[6]) );
  dff_sg \reg_iii_11_reg[6]  ( .D(n4524), .CP(clk), .Q(reg_iii_11[6]) );
  dff_sg \reg_i_11_reg[5]  ( .D(n5755), .CP(clk), .Q(reg_i_11[5]) );
  dff_sg \reg_ii_11_reg[5]  ( .D(n4545), .CP(clk), .Q(reg_ii_11[5]) );
  dff_sg \reg_iii_11_reg[5]  ( .D(n4525), .CP(clk), .Q(reg_iii_11[5]) );
  dff_sg \reg_i_11_reg[4]  ( .D(n5756), .CP(clk), .Q(reg_i_11[4]) );
  dff_sg \reg_ii_11_reg[4]  ( .D(n4546), .CP(clk), .Q(reg_ii_11[4]) );
  dff_sg \reg_iii_11_reg[4]  ( .D(n4526), .CP(clk), .Q(reg_iii_11[4]) );
  dff_sg \reg_i_11_reg[3]  ( .D(n5757), .CP(clk), .Q(reg_i_11[3]) );
  dff_sg \reg_ii_11_reg[3]  ( .D(n4547), .CP(clk), .Q(reg_ii_11[3]) );
  dff_sg \reg_iii_11_reg[3]  ( .D(n4527), .CP(clk), .Q(reg_iii_11[3]) );
  dff_sg \reg_i_11_reg[2]  ( .D(n5758), .CP(clk), .Q(reg_i_11[2]) );
  dff_sg \reg_ii_11_reg[2]  ( .D(n4548), .CP(clk), .Q(reg_ii_11[2]) );
  dff_sg \reg_iii_11_reg[2]  ( .D(n4528), .CP(clk), .Q(reg_iii_11[2]) );
  dff_sg \reg_i_11_reg[1]  ( .D(n5759), .CP(clk), .Q(reg_i_11[1]) );
  dff_sg \reg_ii_11_reg[1]  ( .D(n4549), .CP(clk), .Q(reg_ii_11[1]) );
  dff_sg \reg_iii_11_reg[1]  ( .D(n4529), .CP(clk), .Q(reg_iii_11[1]) );
  dff_sg \reg_i_11_reg[0]  ( .D(n5760), .CP(clk), .Q(reg_i_11[0]) );
  dff_sg \reg_ii_11_reg[0]  ( .D(n4550), .CP(clk), .Q(reg_ii_11[0]) );
  dff_sg \reg_iii_11_reg[0]  ( .D(n4530), .CP(clk), .Q(reg_iii_11[0]) );
  dff_sg \reg_i_10_reg[19]  ( .D(n5761), .CP(clk), .Q(reg_i_10[19]) );
  dff_sg \reg_ii_10_reg[19]  ( .D(n4571), .CP(clk), .Q(reg_ii_10[19]) );
  dff_sg \reg_iii_10_reg[19]  ( .D(n4551), .CP(clk), .Q(reg_iii_10[19]) );
  dff_sg \reg_i_10_reg[18]  ( .D(n5762), .CP(clk), .Q(reg_i_10[18]) );
  dff_sg \reg_ii_10_reg[18]  ( .D(n4572), .CP(clk), .Q(reg_ii_10[18]) );
  dff_sg \reg_iii_10_reg[18]  ( .D(n4552), .CP(clk), .Q(reg_iii_10[18]) );
  dff_sg \reg_i_10_reg[17]  ( .D(n5763), .CP(clk), .Q(reg_i_10[17]) );
  dff_sg \reg_ii_10_reg[17]  ( .D(n4573), .CP(clk), .Q(reg_ii_10[17]) );
  dff_sg \reg_iii_10_reg[17]  ( .D(n4553), .CP(clk), .Q(reg_iii_10[17]) );
  dff_sg \reg_i_10_reg[16]  ( .D(n5764), .CP(clk), .Q(reg_i_10[16]) );
  dff_sg \reg_ii_10_reg[16]  ( .D(n4574), .CP(clk), .Q(reg_ii_10[16]) );
  dff_sg \reg_iii_10_reg[16]  ( .D(n4554), .CP(clk), .Q(reg_iii_10[16]) );
  dff_sg \reg_i_10_reg[15]  ( .D(n5765), .CP(clk), .Q(reg_i_10[15]) );
  dff_sg \reg_ii_10_reg[15]  ( .D(n4575), .CP(clk), .Q(reg_ii_10[15]) );
  dff_sg \reg_iii_10_reg[15]  ( .D(n4555), .CP(clk), .Q(reg_iii_10[15]) );
  dff_sg \reg_i_10_reg[14]  ( .D(n5766), .CP(clk), .Q(reg_i_10[14]) );
  dff_sg \reg_ii_10_reg[14]  ( .D(n4576), .CP(clk), .Q(reg_ii_10[14]) );
  dff_sg \reg_iii_10_reg[14]  ( .D(n4556), .CP(clk), .Q(reg_iii_10[14]) );
  dff_sg \reg_i_10_reg[13]  ( .D(n5767), .CP(clk), .Q(reg_i_10[13]) );
  dff_sg \reg_ii_10_reg[13]  ( .D(n4577), .CP(clk), .Q(reg_ii_10[13]) );
  dff_sg \reg_iii_10_reg[13]  ( .D(n4557), .CP(clk), .Q(reg_iii_10[13]) );
  dff_sg \reg_i_10_reg[12]  ( .D(n5768), .CP(clk), .Q(reg_i_10[12]) );
  dff_sg \reg_ii_10_reg[12]  ( .D(n4578), .CP(clk), .Q(reg_ii_10[12]) );
  dff_sg \reg_iii_10_reg[12]  ( .D(n4558), .CP(clk), .Q(reg_iii_10[12]) );
  dff_sg \reg_i_10_reg[11]  ( .D(n5769), .CP(clk), .Q(reg_i_10[11]) );
  dff_sg \reg_ii_10_reg[11]  ( .D(n4579), .CP(clk), .Q(reg_ii_10[11]) );
  dff_sg \reg_iii_10_reg[11]  ( .D(n4559), .CP(clk), .Q(reg_iii_10[11]) );
  dff_sg \reg_i_10_reg[10]  ( .D(n5770), .CP(clk), .Q(reg_i_10[10]) );
  dff_sg \reg_ii_10_reg[10]  ( .D(n4580), .CP(clk), .Q(reg_ii_10[10]) );
  dff_sg \reg_iii_10_reg[10]  ( .D(n4560), .CP(clk), .Q(reg_iii_10[10]) );
  dff_sg \reg_i_10_reg[9]  ( .D(n5771), .CP(clk), .Q(reg_i_10[9]) );
  dff_sg \reg_ii_10_reg[9]  ( .D(n4581), .CP(clk), .Q(reg_ii_10[9]) );
  dff_sg \reg_iii_10_reg[9]  ( .D(n4561), .CP(clk), .Q(reg_iii_10[9]) );
  dff_sg \reg_i_10_reg[8]  ( .D(n5772), .CP(clk), .Q(reg_i_10[8]) );
  dff_sg \reg_ii_10_reg[8]  ( .D(n4582), .CP(clk), .Q(reg_ii_10[8]) );
  dff_sg \reg_iii_10_reg[8]  ( .D(n4562), .CP(clk), .Q(reg_iii_10[8]) );
  dff_sg \reg_i_10_reg[7]  ( .D(n5773), .CP(clk), .Q(reg_i_10[7]) );
  dff_sg \reg_ii_10_reg[7]  ( .D(n4583), .CP(clk), .Q(reg_ii_10[7]) );
  dff_sg \reg_iii_10_reg[7]  ( .D(n4563), .CP(clk), .Q(reg_iii_10[7]) );
  dff_sg \reg_i_10_reg[6]  ( .D(n5774), .CP(clk), .Q(reg_i_10[6]) );
  dff_sg \reg_ii_10_reg[6]  ( .D(n4584), .CP(clk), .Q(reg_ii_10[6]) );
  dff_sg \reg_iii_10_reg[6]  ( .D(n4564), .CP(clk), .Q(reg_iii_10[6]) );
  dff_sg \reg_i_10_reg[5]  ( .D(n5775), .CP(clk), .Q(reg_i_10[5]) );
  dff_sg \reg_ii_10_reg[5]  ( .D(n4585), .CP(clk), .Q(reg_ii_10[5]) );
  dff_sg \reg_iii_10_reg[5]  ( .D(n4565), .CP(clk), .Q(reg_iii_10[5]) );
  dff_sg \reg_i_10_reg[4]  ( .D(n5776), .CP(clk), .Q(reg_i_10[4]) );
  dff_sg \reg_ii_10_reg[4]  ( .D(n4586), .CP(clk), .Q(reg_ii_10[4]) );
  dff_sg \reg_iii_10_reg[4]  ( .D(n4566), .CP(clk), .Q(reg_iii_10[4]) );
  dff_sg \reg_i_10_reg[3]  ( .D(n5777), .CP(clk), .Q(reg_i_10[3]) );
  dff_sg \reg_ii_10_reg[3]  ( .D(n4587), .CP(clk), .Q(reg_ii_10[3]) );
  dff_sg \reg_iii_10_reg[3]  ( .D(n4567), .CP(clk), .Q(reg_iii_10[3]) );
  dff_sg \reg_i_10_reg[2]  ( .D(n5778), .CP(clk), .Q(reg_i_10[2]) );
  dff_sg \reg_ii_10_reg[2]  ( .D(n4588), .CP(clk), .Q(reg_ii_10[2]) );
  dff_sg \reg_iii_10_reg[2]  ( .D(n4568), .CP(clk), .Q(reg_iii_10[2]) );
  dff_sg \reg_i_10_reg[1]  ( .D(n5779), .CP(clk), .Q(reg_i_10[1]) );
  dff_sg \reg_ii_10_reg[1]  ( .D(n4589), .CP(clk), .Q(reg_ii_10[1]) );
  dff_sg \reg_iii_10_reg[1]  ( .D(n4569), .CP(clk), .Q(reg_iii_10[1]) );
  dff_sg \reg_i_10_reg[0]  ( .D(n5780), .CP(clk), .Q(reg_i_10[0]) );
  dff_sg \reg_ii_10_reg[0]  ( .D(n4590), .CP(clk), .Q(reg_ii_10[0]) );
  dff_sg \reg_iii_10_reg[0]  ( .D(n4570), .CP(clk), .Q(reg_iii_10[0]) );
  dff_sg \reg_i_9_reg[19]  ( .D(n5781), .CP(clk), .Q(reg_i_9[19]) );
  dff_sg \reg_ii_9_reg[19]  ( .D(n4591), .CP(clk), .Q(reg_ii_9[19]) );
  dff_sg \reg_iii_9_reg[19]  ( .D(n4195), .CP(clk), .Q(reg_iii_9[19]) );
  dff_sg \reg_i_9_reg[18]  ( .D(n5782), .CP(clk), .Q(reg_i_9[18]) );
  dff_sg \reg_ii_9_reg[18]  ( .D(n4592), .CP(clk), .Q(reg_ii_9[18]) );
  dff_sg \reg_iii_9_reg[18]  ( .D(n4196), .CP(clk), .Q(reg_iii_9[18]) );
  dff_sg \reg_i_9_reg[17]  ( .D(n5783), .CP(clk), .Q(reg_i_9[17]) );
  dff_sg \reg_ii_9_reg[17]  ( .D(n4215), .CP(clk), .Q(reg_ii_9[17]) );
  dff_sg \reg_iii_9_reg[17]  ( .D(n4197), .CP(clk), .Q(reg_iii_9[17]) );
  dff_sg \reg_i_9_reg[16]  ( .D(n5784), .CP(clk), .Q(reg_i_9[16]) );
  dff_sg \reg_ii_9_reg[16]  ( .D(n4216), .CP(clk), .Q(reg_ii_9[16]) );
  dff_sg \reg_iii_9_reg[16]  ( .D(n4198), .CP(clk), .Q(reg_iii_9[16]) );
  dff_sg \reg_i_9_reg[15]  ( .D(n5785), .CP(clk), .Q(reg_i_9[15]) );
  dff_sg \reg_ii_9_reg[15]  ( .D(n4217), .CP(clk), .Q(reg_ii_9[15]) );
  dff_sg \reg_iii_9_reg[15]  ( .D(n4199), .CP(clk), .Q(reg_iii_9[15]) );
  dff_sg \reg_i_9_reg[14]  ( .D(n5786), .CP(clk), .Q(reg_i_9[14]) );
  dff_sg \reg_ii_9_reg[14]  ( .D(n4218), .CP(clk), .Q(reg_ii_9[14]) );
  dff_sg \reg_iii_9_reg[14]  ( .D(n4200), .CP(clk), .Q(reg_iii_9[14]) );
  dff_sg \reg_i_9_reg[13]  ( .D(n5787), .CP(clk), .Q(reg_i_9[13]) );
  dff_sg \reg_ii_9_reg[13]  ( .D(n4219), .CP(clk), .Q(reg_ii_9[13]) );
  dff_sg \reg_iii_9_reg[13]  ( .D(n4201), .CP(clk), .Q(reg_iii_9[13]) );
  dff_sg \reg_i_9_reg[12]  ( .D(n5788), .CP(clk), .Q(reg_i_9[12]) );
  dff_sg \reg_ii_9_reg[12]  ( .D(n4220), .CP(clk), .Q(reg_ii_9[12]) );
  dff_sg \reg_iii_9_reg[12]  ( .D(n4202), .CP(clk), .Q(reg_iii_9[12]) );
  dff_sg \reg_i_9_reg[11]  ( .D(n5789), .CP(clk), .Q(reg_i_9[11]) );
  dff_sg \reg_ii_9_reg[11]  ( .D(n4221), .CP(clk), .Q(reg_ii_9[11]) );
  dff_sg \reg_iii_9_reg[11]  ( .D(n4203), .CP(clk), .Q(reg_iii_9[11]) );
  dff_sg \reg_i_9_reg[10]  ( .D(n5790), .CP(clk), .Q(reg_i_9[10]) );
  dff_sg \reg_ii_9_reg[10]  ( .D(n4222), .CP(clk), .Q(reg_ii_9[10]) );
  dff_sg \reg_iii_9_reg[10]  ( .D(n4204), .CP(clk), .Q(reg_iii_9[10]) );
  dff_sg \reg_i_9_reg[9]  ( .D(n5791), .CP(clk), .Q(reg_i_9[9]) );
  dff_sg \reg_ii_9_reg[9]  ( .D(n4223), .CP(clk), .Q(reg_ii_9[9]) );
  dff_sg \reg_iii_9_reg[9]  ( .D(n4205), .CP(clk), .Q(reg_iii_9[9]) );
  dff_sg \reg_i_9_reg[8]  ( .D(n5792), .CP(clk), .Q(reg_i_9[8]) );
  dff_sg \reg_ii_9_reg[8]  ( .D(n4224), .CP(clk), .Q(reg_ii_9[8]) );
  dff_sg \reg_iii_9_reg[8]  ( .D(n4206), .CP(clk), .Q(reg_iii_9[8]) );
  dff_sg \reg_i_9_reg[7]  ( .D(n5793), .CP(clk), .Q(reg_i_9[7]) );
  dff_sg \reg_ii_9_reg[7]  ( .D(n4225), .CP(clk), .Q(reg_ii_9[7]) );
  dff_sg \reg_iii_9_reg[7]  ( .D(n4207), .CP(clk), .Q(reg_iii_9[7]) );
  dff_sg \reg_i_9_reg[6]  ( .D(n5794), .CP(clk), .Q(reg_i_9[6]) );
  dff_sg \reg_ii_9_reg[6]  ( .D(n4226), .CP(clk), .Q(reg_ii_9[6]) );
  dff_sg \reg_iii_9_reg[6]  ( .D(n4208), .CP(clk), .Q(reg_iii_9[6]) );
  dff_sg \reg_i_9_reg[5]  ( .D(n5795), .CP(clk), .Q(reg_i_9[5]) );
  dff_sg \reg_ii_9_reg[5]  ( .D(n4227), .CP(clk), .Q(reg_ii_9[5]) );
  dff_sg \reg_iii_9_reg[5]  ( .D(n4209), .CP(clk), .Q(reg_iii_9[5]) );
  dff_sg \reg_i_9_reg[4]  ( .D(n5796), .CP(clk), .Q(reg_i_9[4]) );
  dff_sg \reg_ii_9_reg[4]  ( .D(n4228), .CP(clk), .Q(reg_ii_9[4]) );
  dff_sg \reg_iii_9_reg[4]  ( .D(n4210), .CP(clk), .Q(reg_iii_9[4]) );
  dff_sg \reg_i_9_reg[3]  ( .D(n5797), .CP(clk), .Q(reg_i_9[3]) );
  dff_sg \reg_ii_9_reg[3]  ( .D(n4229), .CP(clk), .Q(reg_ii_9[3]) );
  dff_sg \reg_iii_9_reg[3]  ( .D(n4211), .CP(clk), .Q(reg_iii_9[3]) );
  dff_sg \reg_i_9_reg[2]  ( .D(n5798), .CP(clk), .Q(reg_i_9[2]) );
  dff_sg \reg_ii_9_reg[2]  ( .D(n4230), .CP(clk), .Q(reg_ii_9[2]) );
  dff_sg \reg_iii_9_reg[2]  ( .D(n4212), .CP(clk), .Q(reg_iii_9[2]) );
  dff_sg \reg_i_9_reg[1]  ( .D(n5799), .CP(clk), .Q(reg_i_9[1]) );
  dff_sg \reg_ii_9_reg[1]  ( .D(n4231), .CP(clk), .Q(reg_ii_9[1]) );
  dff_sg \reg_iii_9_reg[1]  ( .D(n4213), .CP(clk), .Q(reg_iii_9[1]) );
  dff_sg \reg_i_9_reg[0]  ( .D(n5800), .CP(clk), .Q(reg_i_9[0]) );
  dff_sg \reg_ii_9_reg[0]  ( .D(n4232), .CP(clk), .Q(reg_ii_9[0]) );
  dff_sg \reg_iii_9_reg[0]  ( .D(n4214), .CP(clk), .Q(reg_iii_9[0]) );
  dff_sg \reg_i_8_reg[19]  ( .D(n5801), .CP(clk), .Q(reg_i_8[19]) );
  dff_sg \reg_ii_8_reg[19]  ( .D(n4253), .CP(clk), .Q(reg_ii_8[19]) );
  dff_sg \reg_iii_8_reg[19]  ( .D(n4233), .CP(clk), .Q(reg_iii_8[19]) );
  dff_sg \reg_i_8_reg[18]  ( .D(n5802), .CP(clk), .Q(reg_i_8[18]) );
  dff_sg \reg_ii_8_reg[18]  ( .D(n4254), .CP(clk), .Q(reg_ii_8[18]) );
  dff_sg \reg_iii_8_reg[18]  ( .D(n4234), .CP(clk), .Q(reg_iii_8[18]) );
  dff_sg \reg_i_8_reg[17]  ( .D(n5803), .CP(clk), .Q(reg_i_8[17]) );
  dff_sg \reg_ii_8_reg[17]  ( .D(n4255), .CP(clk), .Q(reg_ii_8[17]) );
  dff_sg \reg_iii_8_reg[17]  ( .D(n4235), .CP(clk), .Q(reg_iii_8[17]) );
  dff_sg \reg_i_8_reg[16]  ( .D(n5804), .CP(clk), .Q(reg_i_8[16]) );
  dff_sg \reg_ii_8_reg[16]  ( .D(n4256), .CP(clk), .Q(reg_ii_8[16]) );
  dff_sg \reg_iii_8_reg[16]  ( .D(n4236), .CP(clk), .Q(reg_iii_8[16]) );
  dff_sg \reg_i_8_reg[15]  ( .D(n5805), .CP(clk), .Q(reg_i_8[15]) );
  dff_sg \reg_ii_8_reg[15]  ( .D(n4257), .CP(clk), .Q(reg_ii_8[15]) );
  dff_sg \reg_iii_8_reg[15]  ( .D(n4237), .CP(clk), .Q(reg_iii_8[15]) );
  dff_sg \reg_i_8_reg[14]  ( .D(n5806), .CP(clk), .Q(reg_i_8[14]) );
  dff_sg \reg_ii_8_reg[14]  ( .D(n4258), .CP(clk), .Q(reg_ii_8[14]) );
  dff_sg \reg_iii_8_reg[14]  ( .D(n4238), .CP(clk), .Q(reg_iii_8[14]) );
  dff_sg \reg_i_8_reg[13]  ( .D(n5807), .CP(clk), .Q(reg_i_8[13]) );
  dff_sg \reg_ii_8_reg[13]  ( .D(n4259), .CP(clk), .Q(reg_ii_8[13]) );
  dff_sg \reg_iii_8_reg[13]  ( .D(n4239), .CP(clk), .Q(reg_iii_8[13]) );
  dff_sg \reg_i_8_reg[12]  ( .D(n5808), .CP(clk), .Q(reg_i_8[12]) );
  dff_sg \reg_ii_8_reg[12]  ( .D(n4260), .CP(clk), .Q(reg_ii_8[12]) );
  dff_sg \reg_iii_8_reg[12]  ( .D(n4240), .CP(clk), .Q(reg_iii_8[12]) );
  dff_sg \reg_i_8_reg[11]  ( .D(n5809), .CP(clk), .Q(reg_i_8[11]) );
  dff_sg \reg_ii_8_reg[11]  ( .D(n4261), .CP(clk), .Q(reg_ii_8[11]) );
  dff_sg \reg_iii_8_reg[11]  ( .D(n4241), .CP(clk), .Q(reg_iii_8[11]) );
  dff_sg \reg_i_8_reg[10]  ( .D(n5810), .CP(clk), .Q(reg_i_8[10]) );
  dff_sg \reg_ii_8_reg[10]  ( .D(n4262), .CP(clk), .Q(reg_ii_8[10]) );
  dff_sg \reg_iii_8_reg[10]  ( .D(n4242), .CP(clk), .Q(reg_iii_8[10]) );
  dff_sg \reg_i_8_reg[9]  ( .D(n5811), .CP(clk), .Q(reg_i_8[9]) );
  dff_sg \reg_ii_8_reg[9]  ( .D(n4263), .CP(clk), .Q(reg_ii_8[9]) );
  dff_sg \reg_iii_8_reg[9]  ( .D(n4243), .CP(clk), .Q(reg_iii_8[9]) );
  dff_sg \reg_i_8_reg[8]  ( .D(n5812), .CP(clk), .Q(reg_i_8[8]) );
  dff_sg \reg_ii_8_reg[8]  ( .D(n4264), .CP(clk), .Q(reg_ii_8[8]) );
  dff_sg \reg_iii_8_reg[8]  ( .D(n4244), .CP(clk), .Q(reg_iii_8[8]) );
  dff_sg \reg_i_8_reg[7]  ( .D(n5813), .CP(clk), .Q(reg_i_8[7]) );
  dff_sg \reg_ii_8_reg[7]  ( .D(n4265), .CP(clk), .Q(reg_ii_8[7]) );
  dff_sg \reg_iii_8_reg[7]  ( .D(n4245), .CP(clk), .Q(reg_iii_8[7]) );
  dff_sg \reg_i_8_reg[6]  ( .D(n5814), .CP(clk), .Q(reg_i_8[6]) );
  dff_sg \reg_ii_8_reg[6]  ( .D(n4266), .CP(clk), .Q(reg_ii_8[6]) );
  dff_sg \reg_iii_8_reg[6]  ( .D(n4246), .CP(clk), .Q(reg_iii_8[6]) );
  dff_sg \reg_i_8_reg[5]  ( .D(n5815), .CP(clk), .Q(reg_i_8[5]) );
  dff_sg \reg_ii_8_reg[5]  ( .D(n4267), .CP(clk), .Q(reg_ii_8[5]) );
  dff_sg \reg_iii_8_reg[5]  ( .D(n4247), .CP(clk), .Q(reg_iii_8[5]) );
  dff_sg \reg_i_8_reg[4]  ( .D(n5816), .CP(clk), .Q(reg_i_8[4]) );
  dff_sg \reg_ii_8_reg[4]  ( .D(n4268), .CP(clk), .Q(reg_ii_8[4]) );
  dff_sg \reg_iii_8_reg[4]  ( .D(n4248), .CP(clk), .Q(reg_iii_8[4]) );
  dff_sg \reg_i_8_reg[3]  ( .D(n5817), .CP(clk), .Q(reg_i_8[3]) );
  dff_sg \reg_ii_8_reg[3]  ( .D(n4269), .CP(clk), .Q(reg_ii_8[3]) );
  dff_sg \reg_iii_8_reg[3]  ( .D(n4249), .CP(clk), .Q(reg_iii_8[3]) );
  dff_sg \reg_i_8_reg[2]  ( .D(n5818), .CP(clk), .Q(reg_i_8[2]) );
  dff_sg \reg_ii_8_reg[2]  ( .D(n4270), .CP(clk), .Q(reg_ii_8[2]) );
  dff_sg \reg_iii_8_reg[2]  ( .D(n4250), .CP(clk), .Q(reg_iii_8[2]) );
  dff_sg \reg_i_8_reg[1]  ( .D(n5819), .CP(clk), .Q(reg_i_8[1]) );
  dff_sg \reg_ii_8_reg[1]  ( .D(n4271), .CP(clk), .Q(reg_ii_8[1]) );
  dff_sg \reg_iii_8_reg[1]  ( .D(n4251), .CP(clk), .Q(reg_iii_8[1]) );
  dff_sg \reg_i_8_reg[0]  ( .D(n5820), .CP(clk), .Q(reg_i_8[0]) );
  dff_sg \reg_ii_8_reg[0]  ( .D(n4272), .CP(clk), .Q(reg_ii_8[0]) );
  dff_sg \reg_iii_8_reg[0]  ( .D(n4252), .CP(clk), .Q(reg_iii_8[0]) );
  dff_sg \reg_i_7_reg[19]  ( .D(n5821), .CP(clk), .Q(reg_i_7[19]) );
  dff_sg \reg_ii_7_reg[19]  ( .D(n4293), .CP(clk), .Q(reg_ii_7[19]) );
  dff_sg \reg_iii_7_reg[19]  ( .D(n4273), .CP(clk), .Q(reg_iii_7[19]) );
  dff_sg \reg_i_7_reg[18]  ( .D(n5822), .CP(clk), .Q(reg_i_7[18]) );
  dff_sg \reg_ii_7_reg[18]  ( .D(n4294), .CP(clk), .Q(reg_ii_7[18]) );
  dff_sg \reg_iii_7_reg[18]  ( .D(n4274), .CP(clk), .Q(reg_iii_7[18]) );
  dff_sg \reg_i_7_reg[17]  ( .D(n5823), .CP(clk), .Q(reg_i_7[17]) );
  dff_sg \reg_ii_7_reg[17]  ( .D(n4295), .CP(clk), .Q(reg_ii_7[17]) );
  dff_sg \reg_iii_7_reg[17]  ( .D(n4275), .CP(clk), .Q(reg_iii_7[17]) );
  dff_sg \reg_i_7_reg[16]  ( .D(n5824), .CP(clk), .Q(reg_i_7[16]) );
  dff_sg \reg_ii_7_reg[16]  ( .D(n4296), .CP(clk), .Q(reg_ii_7[16]) );
  dff_sg \reg_iii_7_reg[16]  ( .D(n4276), .CP(clk), .Q(reg_iii_7[16]) );
  dff_sg \reg_i_7_reg[15]  ( .D(n5825), .CP(clk), .Q(reg_i_7[15]) );
  dff_sg \reg_ii_7_reg[15]  ( .D(n4297), .CP(clk), .Q(reg_ii_7[15]) );
  dff_sg \reg_iii_7_reg[15]  ( .D(n4277), .CP(clk), .Q(reg_iii_7[15]) );
  dff_sg \reg_i_7_reg[14]  ( .D(n5826), .CP(clk), .Q(reg_i_7[14]) );
  dff_sg \reg_ii_7_reg[14]  ( .D(n4298), .CP(clk), .Q(reg_ii_7[14]) );
  dff_sg \reg_iii_7_reg[14]  ( .D(n4278), .CP(clk), .Q(reg_iii_7[14]) );
  dff_sg \reg_i_7_reg[13]  ( .D(n5827), .CP(clk), .Q(reg_i_7[13]) );
  dff_sg \reg_ii_7_reg[13]  ( .D(n4299), .CP(clk), .Q(reg_ii_7[13]) );
  dff_sg \reg_iii_7_reg[13]  ( .D(n4279), .CP(clk), .Q(reg_iii_7[13]) );
  dff_sg \reg_i_7_reg[12]  ( .D(n5828), .CP(clk), .Q(reg_i_7[12]) );
  dff_sg \reg_ii_7_reg[12]  ( .D(n4300), .CP(clk), .Q(reg_ii_7[12]) );
  dff_sg \reg_iii_7_reg[12]  ( .D(n4280), .CP(clk), .Q(reg_iii_7[12]) );
  dff_sg \reg_i_7_reg[11]  ( .D(n5829), .CP(clk), .Q(reg_i_7[11]) );
  dff_sg \reg_ii_7_reg[11]  ( .D(n4301), .CP(clk), .Q(reg_ii_7[11]) );
  dff_sg \reg_iii_7_reg[11]  ( .D(n4281), .CP(clk), .Q(reg_iii_7[11]) );
  dff_sg \reg_i_7_reg[10]  ( .D(n5830), .CP(clk), .Q(reg_i_7[10]) );
  dff_sg \reg_ii_7_reg[10]  ( .D(n4302), .CP(clk), .Q(reg_ii_7[10]) );
  dff_sg \reg_iii_7_reg[10]  ( .D(n4282), .CP(clk), .Q(reg_iii_7[10]) );
  dff_sg \reg_i_7_reg[9]  ( .D(n5831), .CP(clk), .Q(reg_i_7[9]) );
  dff_sg \reg_ii_7_reg[9]  ( .D(n4303), .CP(clk), .Q(reg_ii_7[9]) );
  dff_sg \reg_iii_7_reg[9]  ( .D(n4283), .CP(clk), .Q(reg_iii_7[9]) );
  dff_sg \reg_i_7_reg[8]  ( .D(n5832), .CP(clk), .Q(reg_i_7[8]) );
  dff_sg \reg_ii_7_reg[8]  ( .D(n4304), .CP(clk), .Q(reg_ii_7[8]) );
  dff_sg \reg_iii_7_reg[8]  ( .D(n4284), .CP(clk), .Q(reg_iii_7[8]) );
  dff_sg \reg_i_7_reg[7]  ( .D(n5833), .CP(clk), .Q(reg_i_7[7]) );
  dff_sg \reg_ii_7_reg[7]  ( .D(n4305), .CP(clk), .Q(reg_ii_7[7]) );
  dff_sg \reg_iii_7_reg[7]  ( .D(n4285), .CP(clk), .Q(reg_iii_7[7]) );
  dff_sg \reg_i_7_reg[6]  ( .D(n5834), .CP(clk), .Q(reg_i_7[6]) );
  dff_sg \reg_ii_7_reg[6]  ( .D(n4306), .CP(clk), .Q(reg_ii_7[6]) );
  dff_sg \reg_iii_7_reg[6]  ( .D(n4286), .CP(clk), .Q(reg_iii_7[6]) );
  dff_sg \reg_i_7_reg[5]  ( .D(n5835), .CP(clk), .Q(reg_i_7[5]) );
  dff_sg \reg_ii_7_reg[5]  ( .D(n4307), .CP(clk), .Q(reg_ii_7[5]) );
  dff_sg \reg_iii_7_reg[5]  ( .D(n4287), .CP(clk), .Q(reg_iii_7[5]) );
  dff_sg \reg_i_7_reg[4]  ( .D(n5836), .CP(clk), .Q(reg_i_7[4]) );
  dff_sg \reg_ii_7_reg[4]  ( .D(n4308), .CP(clk), .Q(reg_ii_7[4]) );
  dff_sg \reg_iii_7_reg[4]  ( .D(n4288), .CP(clk), .Q(reg_iii_7[4]) );
  dff_sg \reg_i_7_reg[3]  ( .D(n5837), .CP(clk), .Q(reg_i_7[3]) );
  dff_sg \reg_ii_7_reg[3]  ( .D(n4309), .CP(clk), .Q(reg_ii_7[3]) );
  dff_sg \reg_iii_7_reg[3]  ( .D(n4289), .CP(clk), .Q(reg_iii_7[3]) );
  dff_sg \reg_i_7_reg[2]  ( .D(n5838), .CP(clk), .Q(reg_i_7[2]) );
  dff_sg \reg_ii_7_reg[2]  ( .D(n4310), .CP(clk), .Q(reg_ii_7[2]) );
  dff_sg \reg_iii_7_reg[2]  ( .D(n4290), .CP(clk), .Q(reg_iii_7[2]) );
  dff_sg \reg_i_7_reg[1]  ( .D(n5839), .CP(clk), .Q(reg_i_7[1]) );
  dff_sg \reg_ii_7_reg[1]  ( .D(n4311), .CP(clk), .Q(reg_ii_7[1]) );
  dff_sg \reg_iii_7_reg[1]  ( .D(n4291), .CP(clk), .Q(reg_iii_7[1]) );
  dff_sg \reg_i_7_reg[0]  ( .D(n5840), .CP(clk), .Q(reg_i_7[0]) );
  dff_sg \reg_ii_7_reg[0]  ( .D(n4312), .CP(clk), .Q(reg_ii_7[0]) );
  dff_sg \reg_iii_7_reg[0]  ( .D(n4292), .CP(clk), .Q(reg_iii_7[0]) );
  dff_sg \reg_i_6_reg[19]  ( .D(n5841), .CP(clk), .Q(reg_i_6[19]) );
  dff_sg \reg_ii_6_reg[19]  ( .D(n4333), .CP(clk), .Q(reg_ii_6[19]) );
  dff_sg \reg_iii_6_reg[19]  ( .D(n4313), .CP(clk), .Q(reg_iii_6[19]) );
  dff_sg \reg_i_6_reg[18]  ( .D(n5842), .CP(clk), .Q(reg_i_6[18]) );
  dff_sg \reg_ii_6_reg[18]  ( .D(n4334), .CP(clk), .Q(reg_ii_6[18]) );
  dff_sg \reg_iii_6_reg[18]  ( .D(n4314), .CP(clk), .Q(reg_iii_6[18]) );
  dff_sg \reg_i_6_reg[17]  ( .D(n5843), .CP(clk), .Q(reg_i_6[17]) );
  dff_sg \reg_ii_6_reg[17]  ( .D(n4335), .CP(clk), .Q(reg_ii_6[17]) );
  dff_sg \reg_iii_6_reg[17]  ( .D(n4315), .CP(clk), .Q(reg_iii_6[17]) );
  dff_sg \reg_i_6_reg[16]  ( .D(n5844), .CP(clk), .Q(reg_i_6[16]) );
  dff_sg \reg_ii_6_reg[16]  ( .D(n4336), .CP(clk), .Q(reg_ii_6[16]) );
  dff_sg \reg_iii_6_reg[16]  ( .D(n4316), .CP(clk), .Q(reg_iii_6[16]) );
  dff_sg \reg_i_6_reg[15]  ( .D(n5845), .CP(clk), .Q(reg_i_6[15]) );
  dff_sg \reg_ii_6_reg[15]  ( .D(n4337), .CP(clk), .Q(reg_ii_6[15]) );
  dff_sg \reg_iii_6_reg[15]  ( .D(n4317), .CP(clk), .Q(reg_iii_6[15]) );
  dff_sg \reg_i_6_reg[14]  ( .D(n5846), .CP(clk), .Q(reg_i_6[14]) );
  dff_sg \reg_ii_6_reg[14]  ( .D(n4338), .CP(clk), .Q(reg_ii_6[14]) );
  dff_sg \reg_iii_6_reg[14]  ( .D(n4318), .CP(clk), .Q(reg_iii_6[14]) );
  dff_sg \reg_i_6_reg[13]  ( .D(n5847), .CP(clk), .Q(reg_i_6[13]) );
  dff_sg \reg_ii_6_reg[13]  ( .D(n4339), .CP(clk), .Q(reg_ii_6[13]) );
  dff_sg \reg_iii_6_reg[13]  ( .D(n4319), .CP(clk), .Q(reg_iii_6[13]) );
  dff_sg \reg_i_6_reg[12]  ( .D(n5848), .CP(clk), .Q(reg_i_6[12]) );
  dff_sg \reg_ii_6_reg[12]  ( .D(n4340), .CP(clk), .Q(reg_ii_6[12]) );
  dff_sg \reg_iii_6_reg[12]  ( .D(n4320), .CP(clk), .Q(reg_iii_6[12]) );
  dff_sg \reg_i_6_reg[11]  ( .D(n5849), .CP(clk), .Q(reg_i_6[11]) );
  dff_sg \reg_ii_6_reg[11]  ( .D(n4341), .CP(clk), .Q(reg_ii_6[11]) );
  dff_sg \reg_iii_6_reg[11]  ( .D(n4321), .CP(clk), .Q(reg_iii_6[11]) );
  dff_sg \reg_i_6_reg[10]  ( .D(n5850), .CP(clk), .Q(reg_i_6[10]) );
  dff_sg \reg_ii_6_reg[10]  ( .D(n4342), .CP(clk), .Q(reg_ii_6[10]) );
  dff_sg \reg_iii_6_reg[10]  ( .D(n4322), .CP(clk), .Q(reg_iii_6[10]) );
  dff_sg \reg_i_6_reg[9]  ( .D(n5851), .CP(clk), .Q(reg_i_6[9]) );
  dff_sg \reg_ii_6_reg[9]  ( .D(n4343), .CP(clk), .Q(reg_ii_6[9]) );
  dff_sg \reg_iii_6_reg[9]  ( .D(n4323), .CP(clk), .Q(reg_iii_6[9]) );
  dff_sg \reg_i_6_reg[8]  ( .D(n5852), .CP(clk), .Q(reg_i_6[8]) );
  dff_sg \reg_ii_6_reg[8]  ( .D(n4344), .CP(clk), .Q(reg_ii_6[8]) );
  dff_sg \reg_iii_6_reg[8]  ( .D(n4324), .CP(clk), .Q(reg_iii_6[8]) );
  dff_sg \reg_i_6_reg[7]  ( .D(n5853), .CP(clk), .Q(reg_i_6[7]) );
  dff_sg \reg_ii_6_reg[7]  ( .D(n4345), .CP(clk), .Q(reg_ii_6[7]) );
  dff_sg \reg_iii_6_reg[7]  ( .D(n4325), .CP(clk), .Q(reg_iii_6[7]) );
  dff_sg \reg_i_6_reg[6]  ( .D(n5854), .CP(clk), .Q(reg_i_6[6]) );
  dff_sg \reg_ii_6_reg[6]  ( .D(n4346), .CP(clk), .Q(reg_ii_6[6]) );
  dff_sg \reg_iii_6_reg[6]  ( .D(n4326), .CP(clk), .Q(reg_iii_6[6]) );
  dff_sg \reg_i_6_reg[5]  ( .D(n5855), .CP(clk), .Q(reg_i_6[5]) );
  dff_sg \reg_ii_6_reg[5]  ( .D(n4347), .CP(clk), .Q(reg_ii_6[5]) );
  dff_sg \reg_iii_6_reg[5]  ( .D(n4327), .CP(clk), .Q(reg_iii_6[5]) );
  dff_sg \reg_i_6_reg[4]  ( .D(n5856), .CP(clk), .Q(reg_i_6[4]) );
  dff_sg \reg_ii_6_reg[4]  ( .D(n4348), .CP(clk), .Q(reg_ii_6[4]) );
  dff_sg \reg_iii_6_reg[4]  ( .D(n4328), .CP(clk), .Q(reg_iii_6[4]) );
  dff_sg \reg_i_6_reg[3]  ( .D(n5857), .CP(clk), .Q(reg_i_6[3]) );
  dff_sg \reg_ii_6_reg[3]  ( .D(n4349), .CP(clk), .Q(reg_ii_6[3]) );
  dff_sg \reg_iii_6_reg[3]  ( .D(n4329), .CP(clk), .Q(reg_iii_6[3]) );
  dff_sg \reg_i_6_reg[2]  ( .D(n5858), .CP(clk), .Q(reg_i_6[2]) );
  dff_sg \reg_ii_6_reg[2]  ( .D(n4350), .CP(clk), .Q(reg_ii_6[2]) );
  dff_sg \reg_iii_6_reg[2]  ( .D(n4330), .CP(clk), .Q(reg_iii_6[2]) );
  dff_sg \reg_i_6_reg[1]  ( .D(n5859), .CP(clk), .Q(reg_i_6[1]) );
  dff_sg \reg_ii_6_reg[1]  ( .D(n4351), .CP(clk), .Q(reg_ii_6[1]) );
  dff_sg \reg_iii_6_reg[1]  ( .D(n4331), .CP(clk), .Q(reg_iii_6[1]) );
  dff_sg \reg_i_6_reg[0]  ( .D(n5860), .CP(clk), .Q(reg_i_6[0]) );
  dff_sg \reg_ii_6_reg[0]  ( .D(n4352), .CP(clk), .Q(reg_ii_6[0]) );
  dff_sg \reg_iii_6_reg[0]  ( .D(n4332), .CP(clk), .Q(reg_iii_6[0]) );
  dff_sg \reg_i_5_reg[19]  ( .D(n5861), .CP(clk), .Q(reg_i_5[19]) );
  dff_sg \reg_ii_5_reg[19]  ( .D(n4373), .CP(clk), .Q(reg_ii_5[19]) );
  dff_sg \reg_iii_5_reg[19]  ( .D(n4353), .CP(clk), .Q(reg_iii_5[19]) );
  dff_sg \reg_i_5_reg[18]  ( .D(n5862), .CP(clk), .Q(reg_i_5[18]) );
  dff_sg \reg_ii_5_reg[18]  ( .D(n4374), .CP(clk), .Q(reg_ii_5[18]) );
  dff_sg \reg_iii_5_reg[18]  ( .D(n4354), .CP(clk), .Q(reg_iii_5[18]) );
  dff_sg \reg_i_5_reg[17]  ( .D(n5863), .CP(clk), .Q(reg_i_5[17]) );
  dff_sg \reg_ii_5_reg[17]  ( .D(n4375), .CP(clk), .Q(reg_ii_5[17]) );
  dff_sg \reg_iii_5_reg[17]  ( .D(n4355), .CP(clk), .Q(reg_iii_5[17]) );
  dff_sg \reg_i_5_reg[16]  ( .D(n5864), .CP(clk), .Q(reg_i_5[16]) );
  dff_sg \reg_ii_5_reg[16]  ( .D(n4376), .CP(clk), .Q(reg_ii_5[16]) );
  dff_sg \reg_iii_5_reg[16]  ( .D(n4356), .CP(clk), .Q(reg_iii_5[16]) );
  dff_sg \reg_i_5_reg[15]  ( .D(n5865), .CP(clk), .Q(reg_i_5[15]) );
  dff_sg \reg_ii_5_reg[15]  ( .D(n4377), .CP(clk), .Q(reg_ii_5[15]) );
  dff_sg \reg_iii_5_reg[15]  ( .D(n4357), .CP(clk), .Q(reg_iii_5[15]) );
  dff_sg \reg_i_5_reg[14]  ( .D(n5866), .CP(clk), .Q(reg_i_5[14]) );
  dff_sg \reg_ii_5_reg[14]  ( .D(n4378), .CP(clk), .Q(reg_ii_5[14]) );
  dff_sg \reg_iii_5_reg[14]  ( .D(n4358), .CP(clk), .Q(reg_iii_5[14]) );
  dff_sg \reg_i_5_reg[13]  ( .D(n5867), .CP(clk), .Q(reg_i_5[13]) );
  dff_sg \reg_ii_5_reg[13]  ( .D(n4379), .CP(clk), .Q(reg_ii_5[13]) );
  dff_sg \reg_iii_5_reg[13]  ( .D(n4359), .CP(clk), .Q(reg_iii_5[13]) );
  dff_sg \reg_i_5_reg[12]  ( .D(n5868), .CP(clk), .Q(reg_i_5[12]) );
  dff_sg \reg_ii_5_reg[12]  ( .D(n4380), .CP(clk), .Q(reg_ii_5[12]) );
  dff_sg \reg_iii_5_reg[12]  ( .D(n4360), .CP(clk), .Q(reg_iii_5[12]) );
  dff_sg \reg_i_5_reg[11]  ( .D(n5869), .CP(clk), .Q(reg_i_5[11]) );
  dff_sg \reg_ii_5_reg[11]  ( .D(n4381), .CP(clk), .Q(reg_ii_5[11]) );
  dff_sg \reg_iii_5_reg[11]  ( .D(n4361), .CP(clk), .Q(reg_iii_5[11]) );
  dff_sg \reg_i_5_reg[10]  ( .D(n5870), .CP(clk), .Q(reg_i_5[10]) );
  dff_sg \reg_ii_5_reg[10]  ( .D(n4382), .CP(clk), .Q(reg_ii_5[10]) );
  dff_sg \reg_iii_5_reg[10]  ( .D(n4362), .CP(clk), .Q(reg_iii_5[10]) );
  dff_sg \reg_i_5_reg[9]  ( .D(n5871), .CP(clk), .Q(reg_i_5[9]) );
  dff_sg \reg_ii_5_reg[9]  ( .D(n4383), .CP(clk), .Q(reg_ii_5[9]) );
  dff_sg \reg_iii_5_reg[9]  ( .D(n4363), .CP(clk), .Q(reg_iii_5[9]) );
  dff_sg \reg_i_5_reg[8]  ( .D(n5872), .CP(clk), .Q(reg_i_5[8]) );
  dff_sg \reg_ii_5_reg[8]  ( .D(n4384), .CP(clk), .Q(reg_ii_5[8]) );
  dff_sg \reg_iii_5_reg[8]  ( .D(n4364), .CP(clk), .Q(reg_iii_5[8]) );
  dff_sg \reg_i_5_reg[7]  ( .D(n5873), .CP(clk), .Q(reg_i_5[7]) );
  dff_sg \reg_ii_5_reg[7]  ( .D(n4385), .CP(clk), .Q(reg_ii_5[7]) );
  dff_sg \reg_iii_5_reg[7]  ( .D(n4365), .CP(clk), .Q(reg_iii_5[7]) );
  dff_sg \reg_i_5_reg[6]  ( .D(n5874), .CP(clk), .Q(reg_i_5[6]) );
  dff_sg \reg_ii_5_reg[6]  ( .D(n4386), .CP(clk), .Q(reg_ii_5[6]) );
  dff_sg \reg_iii_5_reg[6]  ( .D(n4366), .CP(clk), .Q(reg_iii_5[6]) );
  dff_sg \reg_i_5_reg[5]  ( .D(n5875), .CP(clk), .Q(reg_i_5[5]) );
  dff_sg \reg_ii_5_reg[5]  ( .D(n4387), .CP(clk), .Q(reg_ii_5[5]) );
  dff_sg \reg_iii_5_reg[5]  ( .D(n4367), .CP(clk), .Q(reg_iii_5[5]) );
  dff_sg \reg_i_5_reg[4]  ( .D(n5876), .CP(clk), .Q(reg_i_5[4]) );
  dff_sg \reg_ii_5_reg[4]  ( .D(n4388), .CP(clk), .Q(reg_ii_5[4]) );
  dff_sg \reg_iii_5_reg[4]  ( .D(n4368), .CP(clk), .Q(reg_iii_5[4]) );
  dff_sg \reg_i_5_reg[3]  ( .D(n5877), .CP(clk), .Q(reg_i_5[3]) );
  dff_sg \reg_ii_5_reg[3]  ( .D(n4389), .CP(clk), .Q(reg_ii_5[3]) );
  dff_sg \reg_iii_5_reg[3]  ( .D(n4369), .CP(clk), .Q(reg_iii_5[3]) );
  dff_sg \reg_i_5_reg[2]  ( .D(n5878), .CP(clk), .Q(reg_i_5[2]) );
  dff_sg \reg_ii_5_reg[2]  ( .D(n4390), .CP(clk), .Q(reg_ii_5[2]) );
  dff_sg \reg_iii_5_reg[2]  ( .D(n4370), .CP(clk), .Q(reg_iii_5[2]) );
  dff_sg \reg_i_5_reg[1]  ( .D(n5879), .CP(clk), .Q(reg_i_5[1]) );
  dff_sg \reg_ii_5_reg[1]  ( .D(n4391), .CP(clk), .Q(reg_ii_5[1]) );
  dff_sg \reg_iii_5_reg[1]  ( .D(n4371), .CP(clk), .Q(reg_iii_5[1]) );
  dff_sg \reg_i_5_reg[0]  ( .D(n5880), .CP(clk), .Q(reg_i_5[0]) );
  dff_sg \reg_ii_5_reg[0]  ( .D(n4392), .CP(clk), .Q(reg_ii_5[0]) );
  dff_sg \reg_iii_5_reg[0]  ( .D(n4372), .CP(clk), .Q(reg_iii_5[0]) );
  dff_sg \reg_i_4_reg[19]  ( .D(n5881), .CP(clk), .Q(reg_i_4[19]) );
  dff_sg \reg_ii_4_reg[19]  ( .D(n4393), .CP(clk), .Q(reg_ii_4[19]) );
  dff_sg \reg_iii_4_reg[19]  ( .D(n3996), .CP(clk), .Q(reg_iii_4[19]) );
  dff_sg \reg_i_4_reg[18]  ( .D(n5882), .CP(clk), .Q(reg_i_4[18]) );
  dff_sg \reg_ii_4_reg[18]  ( .D(n4016), .CP(clk), .Q(reg_ii_4[18]) );
  dff_sg \reg_iii_4_reg[18]  ( .D(n3997), .CP(clk), .Q(reg_iii_4[18]) );
  dff_sg \reg_i_4_reg[17]  ( .D(n5883), .CP(clk), .Q(reg_i_4[17]) );
  dff_sg \reg_ii_4_reg[17]  ( .D(n4017), .CP(clk), .Q(reg_ii_4[17]) );
  dff_sg \reg_iii_4_reg[17]  ( .D(n3998), .CP(clk), .Q(reg_iii_4[17]) );
  dff_sg \reg_i_4_reg[16]  ( .D(n5884), .CP(clk), .Q(reg_i_4[16]) );
  dff_sg \reg_ii_4_reg[16]  ( .D(n4018), .CP(clk), .Q(reg_ii_4[16]) );
  dff_sg \reg_iii_4_reg[16]  ( .D(n3999), .CP(clk), .Q(reg_iii_4[16]) );
  dff_sg \reg_i_4_reg[15]  ( .D(n5885), .CP(clk), .Q(reg_i_4[15]) );
  dff_sg \reg_ii_4_reg[15]  ( .D(n4019), .CP(clk), .Q(reg_ii_4[15]) );
  dff_sg \reg_iii_4_reg[15]  ( .D(n4000), .CP(clk), .Q(reg_iii_4[15]) );
  dff_sg \reg_i_4_reg[14]  ( .D(n5886), .CP(clk), .Q(reg_i_4[14]) );
  dff_sg \reg_ii_4_reg[14]  ( .D(n4020), .CP(clk), .Q(reg_ii_4[14]) );
  dff_sg \reg_iii_4_reg[14]  ( .D(n4001), .CP(clk), .Q(reg_iii_4[14]) );
  dff_sg \reg_i_4_reg[13]  ( .D(n5887), .CP(clk), .Q(reg_i_4[13]) );
  dff_sg \reg_ii_4_reg[13]  ( .D(n4021), .CP(clk), .Q(reg_ii_4[13]) );
  dff_sg \reg_iii_4_reg[13]  ( .D(n4002), .CP(clk), .Q(reg_iii_4[13]) );
  dff_sg \reg_i_4_reg[12]  ( .D(n5888), .CP(clk), .Q(reg_i_4[12]) );
  dff_sg \reg_ii_4_reg[12]  ( .D(n4022), .CP(clk), .Q(reg_ii_4[12]) );
  dff_sg \reg_iii_4_reg[12]  ( .D(n4003), .CP(clk), .Q(reg_iii_4[12]) );
  dff_sg \reg_i_4_reg[11]  ( .D(n5889), .CP(clk), .Q(reg_i_4[11]) );
  dff_sg \reg_ii_4_reg[11]  ( .D(n4023), .CP(clk), .Q(reg_ii_4[11]) );
  dff_sg \reg_iii_4_reg[11]  ( .D(n4004), .CP(clk), .Q(reg_iii_4[11]) );
  dff_sg \reg_i_4_reg[10]  ( .D(n5890), .CP(clk), .Q(reg_i_4[10]) );
  dff_sg \reg_ii_4_reg[10]  ( .D(n4024), .CP(clk), .Q(reg_ii_4[10]) );
  dff_sg \reg_iii_4_reg[10]  ( .D(n4005), .CP(clk), .Q(reg_iii_4[10]) );
  dff_sg \reg_i_4_reg[9]  ( .D(n5891), .CP(clk), .Q(reg_i_4[9]) );
  dff_sg \reg_ii_4_reg[9]  ( .D(n4025), .CP(clk), .Q(reg_ii_4[9]) );
  dff_sg \reg_iii_4_reg[9]  ( .D(n4006), .CP(clk), .Q(reg_iii_4[9]) );
  dff_sg \reg_i_4_reg[8]  ( .D(n5892), .CP(clk), .Q(reg_i_4[8]) );
  dff_sg \reg_ii_4_reg[8]  ( .D(n4026), .CP(clk), .Q(reg_ii_4[8]) );
  dff_sg \reg_iii_4_reg[8]  ( .D(n4007), .CP(clk), .Q(reg_iii_4[8]) );
  dff_sg \reg_i_4_reg[7]  ( .D(n5893), .CP(clk), .Q(reg_i_4[7]) );
  dff_sg \reg_ii_4_reg[7]  ( .D(n4027), .CP(clk), .Q(reg_ii_4[7]) );
  dff_sg \reg_iii_4_reg[7]  ( .D(n4008), .CP(clk), .Q(reg_iii_4[7]) );
  dff_sg \reg_i_4_reg[6]  ( .D(n5894), .CP(clk), .Q(reg_i_4[6]) );
  dff_sg \reg_ii_4_reg[6]  ( .D(n4028), .CP(clk), .Q(reg_ii_4[6]) );
  dff_sg \reg_iii_4_reg[6]  ( .D(n4009), .CP(clk), .Q(reg_iii_4[6]) );
  dff_sg \reg_i_4_reg[5]  ( .D(n5895), .CP(clk), .Q(reg_i_4[5]) );
  dff_sg \reg_ii_4_reg[5]  ( .D(n4029), .CP(clk), .Q(reg_ii_4[5]) );
  dff_sg \reg_iii_4_reg[5]  ( .D(n4010), .CP(clk), .Q(reg_iii_4[5]) );
  dff_sg \reg_i_4_reg[4]  ( .D(n5896), .CP(clk), .Q(reg_i_4[4]) );
  dff_sg \reg_ii_4_reg[4]  ( .D(n4030), .CP(clk), .Q(reg_ii_4[4]) );
  dff_sg \reg_iii_4_reg[4]  ( .D(n4011), .CP(clk), .Q(reg_iii_4[4]) );
  dff_sg \reg_i_4_reg[3]  ( .D(n5897), .CP(clk), .Q(reg_i_4[3]) );
  dff_sg \reg_ii_4_reg[3]  ( .D(n4031), .CP(clk), .Q(reg_ii_4[3]) );
  dff_sg \reg_iii_4_reg[3]  ( .D(n4012), .CP(clk), .Q(reg_iii_4[3]) );
  dff_sg \reg_i_4_reg[2]  ( .D(n5898), .CP(clk), .Q(reg_i_4[2]) );
  dff_sg \reg_ii_4_reg[2]  ( .D(n4032), .CP(clk), .Q(reg_ii_4[2]) );
  dff_sg \reg_iii_4_reg[2]  ( .D(n4013), .CP(clk), .Q(reg_iii_4[2]) );
  dff_sg \reg_i_4_reg[1]  ( .D(n5899), .CP(clk), .Q(reg_i_4[1]) );
  dff_sg \reg_ii_4_reg[1]  ( .D(n4033), .CP(clk), .Q(reg_ii_4[1]) );
  dff_sg \reg_iii_4_reg[1]  ( .D(n4014), .CP(clk), .Q(reg_iii_4[1]) );
  dff_sg \reg_i_4_reg[0]  ( .D(n5900), .CP(clk), .Q(reg_i_4[0]) );
  dff_sg \reg_ii_4_reg[0]  ( .D(n4034), .CP(clk), .Q(reg_ii_4[0]) );
  dff_sg \reg_iii_4_reg[0]  ( .D(n4015), .CP(clk), .Q(reg_iii_4[0]) );
  dff_sg \reg_i_3_reg[19]  ( .D(n5901), .CP(clk), .Q(reg_i_3[19]) );
  dff_sg \reg_ii_3_reg[19]  ( .D(n4055), .CP(clk), .Q(reg_ii_3[19]) );
  dff_sg \reg_iii_3_reg[19]  ( .D(n4035), .CP(clk), .Q(reg_iii_3[19]) );
  dff_sg \reg_i_3_reg[18]  ( .D(n5902), .CP(clk), .Q(reg_i_3[18]) );
  dff_sg \reg_ii_3_reg[18]  ( .D(n4056), .CP(clk), .Q(reg_ii_3[18]) );
  dff_sg \reg_iii_3_reg[18]  ( .D(n4036), .CP(clk), .Q(reg_iii_3[18]) );
  dff_sg \reg_i_3_reg[17]  ( .D(n5903), .CP(clk), .Q(reg_i_3[17]) );
  dff_sg \reg_ii_3_reg[17]  ( .D(n4057), .CP(clk), .Q(reg_ii_3[17]) );
  dff_sg \reg_iii_3_reg[17]  ( .D(n4037), .CP(clk), .Q(reg_iii_3[17]) );
  dff_sg \reg_i_3_reg[16]  ( .D(n5904), .CP(clk), .Q(reg_i_3[16]) );
  dff_sg \reg_ii_3_reg[16]  ( .D(n4058), .CP(clk), .Q(reg_ii_3[16]) );
  dff_sg \reg_iii_3_reg[16]  ( .D(n4038), .CP(clk), .Q(reg_iii_3[16]) );
  dff_sg \reg_i_3_reg[15]  ( .D(n5905), .CP(clk), .Q(reg_i_3[15]) );
  dff_sg \reg_ii_3_reg[15]  ( .D(n4059), .CP(clk), .Q(reg_ii_3[15]) );
  dff_sg \reg_iii_3_reg[15]  ( .D(n4039), .CP(clk), .Q(reg_iii_3[15]) );
  dff_sg \reg_i_3_reg[14]  ( .D(n5906), .CP(clk), .Q(reg_i_3[14]) );
  dff_sg \reg_ii_3_reg[14]  ( .D(n4060), .CP(clk), .Q(reg_ii_3[14]) );
  dff_sg \reg_iii_3_reg[14]  ( .D(n4040), .CP(clk), .Q(reg_iii_3[14]) );
  dff_sg \reg_i_3_reg[13]  ( .D(n5907), .CP(clk), .Q(reg_i_3[13]) );
  dff_sg \reg_ii_3_reg[13]  ( .D(n4061), .CP(clk), .Q(reg_ii_3[13]) );
  dff_sg \reg_iii_3_reg[13]  ( .D(n4041), .CP(clk), .Q(reg_iii_3[13]) );
  dff_sg \reg_i_3_reg[12]  ( .D(n5908), .CP(clk), .Q(reg_i_3[12]) );
  dff_sg \reg_ii_3_reg[12]  ( .D(n4062), .CP(clk), .Q(reg_ii_3[12]) );
  dff_sg \reg_iii_3_reg[12]  ( .D(n4042), .CP(clk), .Q(reg_iii_3[12]) );
  dff_sg \reg_i_3_reg[11]  ( .D(n5909), .CP(clk), .Q(reg_i_3[11]) );
  dff_sg \reg_ii_3_reg[11]  ( .D(n4063), .CP(clk), .Q(reg_ii_3[11]) );
  dff_sg \reg_iii_3_reg[11]  ( .D(n4043), .CP(clk), .Q(reg_iii_3[11]) );
  dff_sg \reg_i_3_reg[10]  ( .D(n5910), .CP(clk), .Q(reg_i_3[10]) );
  dff_sg \reg_ii_3_reg[10]  ( .D(n4064), .CP(clk), .Q(reg_ii_3[10]) );
  dff_sg \reg_iii_3_reg[10]  ( .D(n4044), .CP(clk), .Q(reg_iii_3[10]) );
  dff_sg \reg_i_3_reg[9]  ( .D(n5911), .CP(clk), .Q(reg_i_3[9]) );
  dff_sg \reg_ii_3_reg[9]  ( .D(n4065), .CP(clk), .Q(reg_ii_3[9]) );
  dff_sg \reg_iii_3_reg[9]  ( .D(n4045), .CP(clk), .Q(reg_iii_3[9]) );
  dff_sg \reg_i_3_reg[8]  ( .D(n5912), .CP(clk), .Q(reg_i_3[8]) );
  dff_sg \reg_ii_3_reg[8]  ( .D(n4066), .CP(clk), .Q(reg_ii_3[8]) );
  dff_sg \reg_iii_3_reg[8]  ( .D(n4046), .CP(clk), .Q(reg_iii_3[8]) );
  dff_sg \reg_i_3_reg[7]  ( .D(n5913), .CP(clk), .Q(reg_i_3[7]) );
  dff_sg \reg_ii_3_reg[7]  ( .D(n4067), .CP(clk), .Q(reg_ii_3[7]) );
  dff_sg \reg_iii_3_reg[7]  ( .D(n4047), .CP(clk), .Q(reg_iii_3[7]) );
  dff_sg \reg_i_3_reg[6]  ( .D(n5914), .CP(clk), .Q(reg_i_3[6]) );
  dff_sg \reg_ii_3_reg[6]  ( .D(n4068), .CP(clk), .Q(reg_ii_3[6]) );
  dff_sg \reg_iii_3_reg[6]  ( .D(n4048), .CP(clk), .Q(reg_iii_3[6]) );
  dff_sg \reg_i_3_reg[5]  ( .D(n5915), .CP(clk), .Q(reg_i_3[5]) );
  dff_sg \reg_ii_3_reg[5]  ( .D(n4069), .CP(clk), .Q(reg_ii_3[5]) );
  dff_sg \reg_iii_3_reg[5]  ( .D(n4049), .CP(clk), .Q(reg_iii_3[5]) );
  dff_sg \reg_i_3_reg[4]  ( .D(n5916), .CP(clk), .Q(reg_i_3[4]) );
  dff_sg \reg_ii_3_reg[4]  ( .D(n4070), .CP(clk), .Q(reg_ii_3[4]) );
  dff_sg \reg_iii_3_reg[4]  ( .D(n4050), .CP(clk), .Q(reg_iii_3[4]) );
  dff_sg \reg_i_3_reg[3]  ( .D(n5917), .CP(clk), .Q(reg_i_3[3]) );
  dff_sg \reg_ii_3_reg[3]  ( .D(n4071), .CP(clk), .Q(reg_ii_3[3]) );
  dff_sg \reg_iii_3_reg[3]  ( .D(n4051), .CP(clk), .Q(reg_iii_3[3]) );
  dff_sg \reg_i_3_reg[2]  ( .D(n5918), .CP(clk), .Q(reg_i_3[2]) );
  dff_sg \reg_ii_3_reg[2]  ( .D(n4072), .CP(clk), .Q(reg_ii_3[2]) );
  dff_sg \reg_iii_3_reg[2]  ( .D(n4052), .CP(clk), .Q(reg_iii_3[2]) );
  dff_sg \reg_i_3_reg[1]  ( .D(n5919), .CP(clk), .Q(reg_i_3[1]) );
  dff_sg \reg_ii_3_reg[1]  ( .D(n4073), .CP(clk), .Q(reg_ii_3[1]) );
  dff_sg \reg_iii_3_reg[1]  ( .D(n4053), .CP(clk), .Q(reg_iii_3[1]) );
  dff_sg \reg_i_3_reg[0]  ( .D(n5920), .CP(clk), .Q(reg_i_3[0]) );
  dff_sg \reg_ii_3_reg[0]  ( .D(n4074), .CP(clk), .Q(reg_ii_3[0]) );
  dff_sg \reg_iii_3_reg[0]  ( .D(n4054), .CP(clk), .Q(reg_iii_3[0]) );
  dff_sg \reg_i_2_reg[19]  ( .D(n5921), .CP(clk), .Q(reg_i_2[19]) );
  dff_sg \reg_ii_2_reg[19]  ( .D(n4095), .CP(clk), .Q(reg_ii_2[19]) );
  dff_sg \reg_iii_2_reg[19]  ( .D(n4075), .CP(clk), .Q(reg_iii_2[19]) );
  dff_sg \reg_i_2_reg[18]  ( .D(n5922), .CP(clk), .Q(reg_i_2[18]) );
  dff_sg \reg_ii_2_reg[18]  ( .D(n4096), .CP(clk), .Q(reg_ii_2[18]) );
  dff_sg \reg_iii_2_reg[18]  ( .D(n4076), .CP(clk), .Q(reg_iii_2[18]) );
  dff_sg \reg_i_2_reg[17]  ( .D(n5923), .CP(clk), .Q(reg_i_2[17]) );
  dff_sg \reg_ii_2_reg[17]  ( .D(n4097), .CP(clk), .Q(reg_ii_2[17]) );
  dff_sg \reg_iii_2_reg[17]  ( .D(n4077), .CP(clk), .Q(reg_iii_2[17]) );
  dff_sg \reg_i_2_reg[16]  ( .D(n5924), .CP(clk), .Q(reg_i_2[16]) );
  dff_sg \reg_ii_2_reg[16]  ( .D(n4098), .CP(clk), .Q(reg_ii_2[16]) );
  dff_sg \reg_iii_2_reg[16]  ( .D(n4078), .CP(clk), .Q(reg_iii_2[16]) );
  dff_sg \reg_i_2_reg[15]  ( .D(n5925), .CP(clk), .Q(reg_i_2[15]) );
  dff_sg \reg_ii_2_reg[15]  ( .D(n4099), .CP(clk), .Q(reg_ii_2[15]) );
  dff_sg \reg_iii_2_reg[15]  ( .D(n4079), .CP(clk), .Q(reg_iii_2[15]) );
  dff_sg \reg_i_2_reg[14]  ( .D(n5926), .CP(clk), .Q(reg_i_2[14]) );
  dff_sg \reg_ii_2_reg[14]  ( .D(n4100), .CP(clk), .Q(reg_ii_2[14]) );
  dff_sg \reg_iii_2_reg[14]  ( .D(n4080), .CP(clk), .Q(reg_iii_2[14]) );
  dff_sg \reg_i_2_reg[13]  ( .D(n5927), .CP(clk), .Q(reg_i_2[13]) );
  dff_sg \reg_ii_2_reg[13]  ( .D(n4101), .CP(clk), .Q(reg_ii_2[13]) );
  dff_sg \reg_iii_2_reg[13]  ( .D(n4081), .CP(clk), .Q(reg_iii_2[13]) );
  dff_sg \reg_i_2_reg[12]  ( .D(n5928), .CP(clk), .Q(reg_i_2[12]) );
  dff_sg \reg_ii_2_reg[12]  ( .D(n4102), .CP(clk), .Q(reg_ii_2[12]) );
  dff_sg \reg_iii_2_reg[12]  ( .D(n4082), .CP(clk), .Q(reg_iii_2[12]) );
  dff_sg \reg_i_2_reg[11]  ( .D(n5929), .CP(clk), .Q(reg_i_2[11]) );
  dff_sg \reg_ii_2_reg[11]  ( .D(n4103), .CP(clk), .Q(reg_ii_2[11]) );
  dff_sg \reg_iii_2_reg[11]  ( .D(n4083), .CP(clk), .Q(reg_iii_2[11]) );
  dff_sg \reg_i_2_reg[10]  ( .D(n5930), .CP(clk), .Q(reg_i_2[10]) );
  dff_sg \reg_ii_2_reg[10]  ( .D(n4104), .CP(clk), .Q(reg_ii_2[10]) );
  dff_sg \reg_iii_2_reg[10]  ( .D(n4084), .CP(clk), .Q(reg_iii_2[10]) );
  dff_sg \reg_i_2_reg[9]  ( .D(n5931), .CP(clk), .Q(reg_i_2[9]) );
  dff_sg \reg_ii_2_reg[9]  ( .D(n4105), .CP(clk), .Q(reg_ii_2[9]) );
  dff_sg \reg_iii_2_reg[9]  ( .D(n4085), .CP(clk), .Q(reg_iii_2[9]) );
  dff_sg \reg_i_2_reg[8]  ( .D(n5932), .CP(clk), .Q(reg_i_2[8]) );
  dff_sg \reg_ii_2_reg[8]  ( .D(n4106), .CP(clk), .Q(reg_ii_2[8]) );
  dff_sg \reg_iii_2_reg[8]  ( .D(n4086), .CP(clk), .Q(reg_iii_2[8]) );
  dff_sg \reg_i_2_reg[7]  ( .D(n5933), .CP(clk), .Q(reg_i_2[7]) );
  dff_sg \reg_ii_2_reg[7]  ( .D(n4107), .CP(clk), .Q(reg_ii_2[7]) );
  dff_sg \reg_iii_2_reg[7]  ( .D(n4087), .CP(clk), .Q(reg_iii_2[7]) );
  dff_sg \reg_i_2_reg[6]  ( .D(n5934), .CP(clk), .Q(reg_i_2[6]) );
  dff_sg \reg_ii_2_reg[6]  ( .D(n4108), .CP(clk), .Q(reg_ii_2[6]) );
  dff_sg \reg_iii_2_reg[6]  ( .D(n4088), .CP(clk), .Q(reg_iii_2[6]) );
  dff_sg \reg_i_2_reg[5]  ( .D(n5935), .CP(clk), .Q(reg_i_2[5]) );
  dff_sg \reg_ii_2_reg[5]  ( .D(n4109), .CP(clk), .Q(reg_ii_2[5]) );
  dff_sg \reg_iii_2_reg[5]  ( .D(n4089), .CP(clk), .Q(reg_iii_2[5]) );
  dff_sg \reg_i_2_reg[4]  ( .D(n5936), .CP(clk), .Q(reg_i_2[4]) );
  dff_sg \reg_ii_2_reg[4]  ( .D(n4110), .CP(clk), .Q(reg_ii_2[4]) );
  dff_sg \reg_iii_2_reg[4]  ( .D(n4090), .CP(clk), .Q(reg_iii_2[4]) );
  dff_sg \reg_i_2_reg[3]  ( .D(n5937), .CP(clk), .Q(reg_i_2[3]) );
  dff_sg \reg_ii_2_reg[3]  ( .D(n4111), .CP(clk), .Q(reg_ii_2[3]) );
  dff_sg \reg_iii_2_reg[3]  ( .D(n4091), .CP(clk), .Q(reg_iii_2[3]) );
  dff_sg \reg_i_2_reg[2]  ( .D(n5938), .CP(clk), .Q(reg_i_2[2]) );
  dff_sg \reg_ii_2_reg[2]  ( .D(n4112), .CP(clk), .Q(reg_ii_2[2]) );
  dff_sg \reg_iii_2_reg[2]  ( .D(n4092), .CP(clk), .Q(reg_iii_2[2]) );
  dff_sg \reg_i_2_reg[1]  ( .D(n5939), .CP(clk), .Q(reg_i_2[1]) );
  dff_sg \reg_ii_2_reg[1]  ( .D(n4113), .CP(clk), .Q(reg_ii_2[1]) );
  dff_sg \reg_iii_2_reg[1]  ( .D(n4093), .CP(clk), .Q(reg_iii_2[1]) );
  dff_sg \reg_i_2_reg[0]  ( .D(n5940), .CP(clk), .Q(reg_i_2[0]) );
  dff_sg \reg_ii_2_reg[0]  ( .D(n4114), .CP(clk), .Q(reg_ii_2[0]) );
  dff_sg \reg_iii_2_reg[0]  ( .D(n4094), .CP(clk), .Q(reg_iii_2[0]) );
  dff_sg \reg_i_1_reg[19]  ( .D(n5941), .CP(clk), .Q(reg_i_1[19]) );
  dff_sg \reg_ii_1_reg[19]  ( .D(n4135), .CP(clk), .Q(reg_ii_1[19]) );
  dff_sg \reg_iii_1_reg[19]  ( .D(n4115), .CP(clk), .Q(reg_iii_1[19]) );
  dff_sg \reg_i_1_reg[18]  ( .D(n5942), .CP(clk), .Q(reg_i_1[18]) );
  dff_sg \reg_ii_1_reg[18]  ( .D(n4136), .CP(clk), .Q(reg_ii_1[18]) );
  dff_sg \reg_iii_1_reg[18]  ( .D(n4116), .CP(clk), .Q(reg_iii_1[18]) );
  dff_sg \reg_i_1_reg[17]  ( .D(n5943), .CP(clk), .Q(reg_i_1[17]) );
  dff_sg \reg_ii_1_reg[17]  ( .D(n4137), .CP(clk), .Q(reg_ii_1[17]) );
  dff_sg \reg_iii_1_reg[17]  ( .D(n4117), .CP(clk), .Q(reg_iii_1[17]) );
  dff_sg \reg_i_1_reg[16]  ( .D(n5944), .CP(clk), .Q(reg_i_1[16]) );
  dff_sg \reg_ii_1_reg[16]  ( .D(n4138), .CP(clk), .Q(reg_ii_1[16]) );
  dff_sg \reg_iii_1_reg[16]  ( .D(n4118), .CP(clk), .Q(reg_iii_1[16]) );
  dff_sg \reg_i_1_reg[15]  ( .D(n5945), .CP(clk), .Q(reg_i_1[15]) );
  dff_sg \reg_ii_1_reg[15]  ( .D(n4139), .CP(clk), .Q(reg_ii_1[15]) );
  dff_sg \reg_iii_1_reg[15]  ( .D(n4119), .CP(clk), .Q(reg_iii_1[15]) );
  dff_sg \reg_i_1_reg[14]  ( .D(n5946), .CP(clk), .Q(reg_i_1[14]) );
  dff_sg \reg_ii_1_reg[14]  ( .D(n4140), .CP(clk), .Q(reg_ii_1[14]) );
  dff_sg \reg_iii_1_reg[14]  ( .D(n4120), .CP(clk), .Q(reg_iii_1[14]) );
  dff_sg \reg_i_1_reg[13]  ( .D(n5947), .CP(clk), .Q(reg_i_1[13]) );
  dff_sg \reg_ii_1_reg[13]  ( .D(n4141), .CP(clk), .Q(reg_ii_1[13]) );
  dff_sg \reg_iii_1_reg[13]  ( .D(n4121), .CP(clk), .Q(reg_iii_1[13]) );
  dff_sg \reg_i_1_reg[12]  ( .D(n5948), .CP(clk), .Q(reg_i_1[12]) );
  dff_sg \reg_ii_1_reg[12]  ( .D(n4142), .CP(clk), .Q(reg_ii_1[12]) );
  dff_sg \reg_iii_1_reg[12]  ( .D(n4122), .CP(clk), .Q(reg_iii_1[12]) );
  dff_sg \reg_i_1_reg[11]  ( .D(n5949), .CP(clk), .Q(reg_i_1[11]) );
  dff_sg \reg_ii_1_reg[11]  ( .D(n4143), .CP(clk), .Q(reg_ii_1[11]) );
  dff_sg \reg_iii_1_reg[11]  ( .D(n4123), .CP(clk), .Q(reg_iii_1[11]) );
  dff_sg \reg_i_1_reg[10]  ( .D(n5950), .CP(clk), .Q(reg_i_1[10]) );
  dff_sg \reg_ii_1_reg[10]  ( .D(n4144), .CP(clk), .Q(reg_ii_1[10]) );
  dff_sg \reg_iii_1_reg[10]  ( .D(n4124), .CP(clk), .Q(reg_iii_1[10]) );
  dff_sg \reg_i_1_reg[9]  ( .D(n5951), .CP(clk), .Q(reg_i_1[9]) );
  dff_sg \reg_ii_1_reg[9]  ( .D(n4145), .CP(clk), .Q(reg_ii_1[9]) );
  dff_sg \reg_iii_1_reg[9]  ( .D(n4125), .CP(clk), .Q(reg_iii_1[9]) );
  dff_sg \reg_i_1_reg[8]  ( .D(n5952), .CP(clk), .Q(reg_i_1[8]) );
  dff_sg \reg_ii_1_reg[8]  ( .D(n4146), .CP(clk), .Q(reg_ii_1[8]) );
  dff_sg \reg_iii_1_reg[8]  ( .D(n4126), .CP(clk), .Q(reg_iii_1[8]) );
  dff_sg \reg_i_1_reg[7]  ( .D(n5953), .CP(clk), .Q(reg_i_1[7]) );
  dff_sg \reg_ii_1_reg[7]  ( .D(n4147), .CP(clk), .Q(reg_ii_1[7]) );
  dff_sg \reg_iii_1_reg[7]  ( .D(n4127), .CP(clk), .Q(reg_iii_1[7]) );
  dff_sg \reg_i_1_reg[6]  ( .D(n5954), .CP(clk), .Q(reg_i_1[6]) );
  dff_sg \reg_ii_1_reg[6]  ( .D(n4148), .CP(clk), .Q(reg_ii_1[6]) );
  dff_sg \reg_iii_1_reg[6]  ( .D(n4128), .CP(clk), .Q(reg_iii_1[6]) );
  dff_sg \reg_i_1_reg[5]  ( .D(n5955), .CP(clk), .Q(reg_i_1[5]) );
  dff_sg \reg_ii_1_reg[5]  ( .D(n4149), .CP(clk), .Q(reg_ii_1[5]) );
  dff_sg \reg_iii_1_reg[5]  ( .D(n4129), .CP(clk), .Q(reg_iii_1[5]) );
  dff_sg \reg_i_1_reg[4]  ( .D(n5956), .CP(clk), .Q(reg_i_1[4]) );
  dff_sg \reg_ii_1_reg[4]  ( .D(n4150), .CP(clk), .Q(reg_ii_1[4]) );
  dff_sg \reg_iii_1_reg[4]  ( .D(n4130), .CP(clk), .Q(reg_iii_1[4]) );
  dff_sg \reg_i_1_reg[3]  ( .D(n5957), .CP(clk), .Q(reg_i_1[3]) );
  dff_sg \reg_ii_1_reg[3]  ( .D(n4151), .CP(clk), .Q(reg_ii_1[3]) );
  dff_sg \reg_iii_1_reg[3]  ( .D(n4131), .CP(clk), .Q(reg_iii_1[3]) );
  dff_sg \reg_i_1_reg[2]  ( .D(n5958), .CP(clk), .Q(reg_i_1[2]) );
  dff_sg \reg_ii_1_reg[2]  ( .D(n4152), .CP(clk), .Q(reg_ii_1[2]) );
  dff_sg \reg_iii_1_reg[2]  ( .D(n4132), .CP(clk), .Q(reg_iii_1[2]) );
  dff_sg \reg_i_1_reg[1]  ( .D(n5959), .CP(clk), .Q(reg_i_1[1]) );
  dff_sg \reg_ii_1_reg[1]  ( .D(n4153), .CP(clk), .Q(reg_ii_1[1]) );
  dff_sg \reg_iii_1_reg[1]  ( .D(n4133), .CP(clk), .Q(reg_iii_1[1]) );
  dff_sg \reg_i_1_reg[0]  ( .D(n5960), .CP(clk), .Q(reg_i_1[0]) );
  dff_sg \reg_ii_1_reg[0]  ( .D(n4154), .CP(clk), .Q(reg_ii_1[0]) );
  dff_sg \reg_iii_1_reg[0]  ( .D(n4134), .CP(clk), .Q(reg_iii_1[0]) );
  dff_sg \reg_i_0_reg[19]  ( .D(n5961), .CP(clk), .Q(reg_i_0[19]) );
  dff_sg \reg_ii_0_reg[19]  ( .D(n4175), .CP(clk), .Q(reg_ii_0[19]) );
  dff_sg \reg_iii_0_reg[19]  ( .D(n4155), .CP(clk), .Q(reg_iii_0[19]) );
  dff_sg \reg_i_0_reg[18]  ( .D(n5962), .CP(clk), .Q(reg_i_0[18]) );
  dff_sg \reg_ii_0_reg[18]  ( .D(n4176), .CP(clk), .Q(reg_ii_0[18]) );
  dff_sg \reg_iii_0_reg[18]  ( .D(n4156), .CP(clk), .Q(reg_iii_0[18]) );
  dff_sg \reg_i_0_reg[17]  ( .D(n5963), .CP(clk), .Q(reg_i_0[17]) );
  dff_sg \reg_ii_0_reg[17]  ( .D(n4177), .CP(clk), .Q(reg_ii_0[17]) );
  dff_sg \reg_iii_0_reg[17]  ( .D(n4157), .CP(clk), .Q(reg_iii_0[17]) );
  dff_sg \reg_i_0_reg[16]  ( .D(n5964), .CP(clk), .Q(reg_i_0[16]) );
  dff_sg \reg_ii_0_reg[16]  ( .D(n4178), .CP(clk), .Q(reg_ii_0[16]) );
  dff_sg \reg_iii_0_reg[16]  ( .D(n4158), .CP(clk), .Q(reg_iii_0[16]) );
  dff_sg \reg_i_0_reg[15]  ( .D(n5965), .CP(clk), .Q(reg_i_0[15]) );
  dff_sg \reg_ii_0_reg[15]  ( .D(n4179), .CP(clk), .Q(reg_ii_0[15]) );
  dff_sg \reg_iii_0_reg[15]  ( .D(n4159), .CP(clk), .Q(reg_iii_0[15]) );
  dff_sg \reg_i_0_reg[14]  ( .D(n5966), .CP(clk), .Q(reg_i_0[14]) );
  dff_sg \reg_ii_0_reg[14]  ( .D(n4180), .CP(clk), .Q(reg_ii_0[14]) );
  dff_sg \reg_iii_0_reg[14]  ( .D(n4160), .CP(clk), .Q(reg_iii_0[14]) );
  dff_sg \reg_i_0_reg[13]  ( .D(n5967), .CP(clk), .Q(reg_i_0[13]) );
  dff_sg \reg_ii_0_reg[13]  ( .D(n4181), .CP(clk), .Q(reg_ii_0[13]) );
  dff_sg \reg_iii_0_reg[13]  ( .D(n4161), .CP(clk), .Q(reg_iii_0[13]) );
  dff_sg \reg_i_0_reg[12]  ( .D(n5968), .CP(clk), .Q(reg_i_0[12]) );
  dff_sg \reg_ii_0_reg[12]  ( .D(n4182), .CP(clk), .Q(reg_ii_0[12]) );
  dff_sg \reg_iii_0_reg[12]  ( .D(n4162), .CP(clk), .Q(reg_iii_0[12]) );
  dff_sg \reg_i_0_reg[11]  ( .D(n5969), .CP(clk), .Q(reg_i_0[11]) );
  dff_sg \reg_ii_0_reg[11]  ( .D(n4183), .CP(clk), .Q(reg_ii_0[11]) );
  dff_sg \reg_iii_0_reg[11]  ( .D(n4163), .CP(clk), .Q(reg_iii_0[11]) );
  dff_sg \reg_i_0_reg[10]  ( .D(n5970), .CP(clk), .Q(reg_i_0[10]) );
  dff_sg \reg_ii_0_reg[10]  ( .D(n4184), .CP(clk), .Q(reg_ii_0[10]) );
  dff_sg \reg_iii_0_reg[10]  ( .D(n4164), .CP(clk), .Q(reg_iii_0[10]) );
  dff_sg \reg_i_0_reg[9]  ( .D(n5971), .CP(clk), .Q(reg_i_0[9]) );
  dff_sg \reg_ii_0_reg[9]  ( .D(n4185), .CP(clk), .Q(reg_ii_0[9]) );
  dff_sg \reg_iii_0_reg[9]  ( .D(n4165), .CP(clk), .Q(reg_iii_0[9]) );
  dff_sg \reg_i_0_reg[8]  ( .D(n5972), .CP(clk), .Q(reg_i_0[8]) );
  dff_sg \reg_ii_0_reg[8]  ( .D(n4186), .CP(clk), .Q(reg_ii_0[8]) );
  dff_sg \reg_iii_0_reg[8]  ( .D(n4166), .CP(clk), .Q(reg_iii_0[8]) );
  dff_sg \reg_i_0_reg[7]  ( .D(n5973), .CP(clk), .Q(reg_i_0[7]) );
  dff_sg \reg_ii_0_reg[7]  ( .D(n4187), .CP(clk), .Q(reg_ii_0[7]) );
  dff_sg \reg_iii_0_reg[7]  ( .D(n4167), .CP(clk), .Q(reg_iii_0[7]) );
  dff_sg \reg_i_0_reg[6]  ( .D(n5974), .CP(clk), .Q(reg_i_0[6]) );
  dff_sg \reg_ii_0_reg[6]  ( .D(n4188), .CP(clk), .Q(reg_ii_0[6]) );
  dff_sg \reg_iii_0_reg[6]  ( .D(n4168), .CP(clk), .Q(reg_iii_0[6]) );
  dff_sg \reg_i_0_reg[5]  ( .D(n5975), .CP(clk), .Q(reg_i_0[5]) );
  dff_sg \reg_ii_0_reg[5]  ( .D(n4189), .CP(clk), .Q(reg_ii_0[5]) );
  dff_sg \reg_iii_0_reg[5]  ( .D(n4169), .CP(clk), .Q(reg_iii_0[5]) );
  dff_sg \reg_i_0_reg[4]  ( .D(n5976), .CP(clk), .Q(reg_i_0[4]) );
  dff_sg \reg_ii_0_reg[4]  ( .D(n4190), .CP(clk), .Q(reg_ii_0[4]) );
  dff_sg \reg_iii_0_reg[4]  ( .D(n4170), .CP(clk), .Q(reg_iii_0[4]) );
  dff_sg \reg_i_0_reg[3]  ( .D(n5977), .CP(clk), .Q(reg_i_0[3]) );
  dff_sg \reg_ii_0_reg[3]  ( .D(n4191), .CP(clk), .Q(reg_ii_0[3]) );
  dff_sg \reg_iii_0_reg[3]  ( .D(n4171), .CP(clk), .Q(reg_iii_0[3]) );
  dff_sg \reg_i_0_reg[2]  ( .D(n5978), .CP(clk), .Q(reg_i_0[2]) );
  dff_sg \reg_ii_0_reg[2]  ( .D(n4192), .CP(clk), .Q(reg_ii_0[2]) );
  dff_sg \reg_iii_0_reg[2]  ( .D(n4172), .CP(clk), .Q(reg_iii_0[2]) );
  dff_sg \reg_i_0_reg[1]  ( .D(n5979), .CP(clk), .Q(reg_i_0[1]) );
  dff_sg \reg_ii_0_reg[1]  ( .D(n4193), .CP(clk), .Q(reg_ii_0[1]) );
  dff_sg \reg_iii_0_reg[1]  ( .D(n4173), .CP(clk), .Q(reg_iii_0[1]) );
  dff_sg \reg_i_0_reg[0]  ( .D(n5980), .CP(clk), .Q(reg_i_0[0]) );
  dff_sg \reg_ii_0_reg[0]  ( .D(n4194), .CP(clk), .Q(reg_ii_0[0]) );
  dff_sg \reg_iii_0_reg[0]  ( .D(n4174), .CP(clk), .Q(reg_iii_0[0]) );
  dff_sg input_taken_reg ( .D(n5276), .CP(clk), .Q(input_taken) );
  dff_sg \mask_0/reg_ii_mask_reg[0]  ( .D(\mask_0/n611 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[0] ) );
  dff_sg \mask_0/reg_ii_mask_reg[1]  ( .D(\mask_0/n612 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[1] ) );
  dff_sg \mask_0/reg_ii_mask_reg[2]  ( .D(\mask_0/n613 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[2] ) );
  dff_sg \mask_0/reg_ii_mask_reg[3]  ( .D(\mask_0/n614 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[3] ) );
  dff_sg \mask_0/reg_ii_mask_reg[4]  ( .D(\mask_0/n615 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[4] ) );
  dff_sg \mask_0/reg_ii_mask_reg[5]  ( .D(\mask_0/n616 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[5] ) );
  dff_sg \mask_0/reg_ii_mask_reg[6]  ( .D(\mask_0/n617 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[6] ) );
  dff_sg \mask_0/reg_ii_mask_reg[7]  ( .D(\mask_0/n618 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[7] ) );
  dff_sg \mask_0/reg_ii_mask_reg[8]  ( .D(\mask_0/n619 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[8] ) );
  dff_sg \mask_0/reg_ii_mask_reg[9]  ( .D(\mask_0/n620 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[9] ) );
  dff_sg \mask_0/reg_ii_mask_reg[10]  ( .D(\mask_0/n621 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[10] ) );
  dff_sg \mask_0/reg_ii_mask_reg[11]  ( .D(\mask_0/n622 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[11] ) );
  dff_sg \mask_0/reg_ii_mask_reg[12]  ( .D(\mask_0/n623 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[12] ) );
  dff_sg \mask_0/reg_ii_mask_reg[13]  ( .D(\mask_0/n624 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[13] ) );
  dff_sg \mask_0/reg_ii_mask_reg[14]  ( .D(\mask_0/n625 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[14] ) );
  dff_sg \mask_0/reg_ii_mask_reg[15]  ( .D(\mask_0/n626 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[15] ) );
  dff_sg \mask_0/reg_ii_mask_reg[16]  ( .D(\mask_0/n627 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[16] ) );
  dff_sg \mask_0/reg_ii_mask_reg[17]  ( .D(\mask_0/n628 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[17] ) );
  dff_sg \mask_0/reg_ii_mask_reg[18]  ( .D(\mask_0/n629 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[18] ) );
  dff_sg \mask_0/reg_ii_mask_reg[19]  ( .D(\mask_0/n630 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[19] ) );
  dff_sg \mask_0/reg_ii_mask_reg[20]  ( .D(\mask_0/n631 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[20] ) );
  dff_sg \mask_0/reg_ii_mask_reg[21]  ( .D(\mask_0/n632 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[21] ) );
  dff_sg \mask_0/reg_ii_mask_reg[22]  ( .D(\mask_0/n633 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[22] ) );
  dff_sg \mask_0/reg_ii_mask_reg[23]  ( .D(\mask_0/n634 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[23] ) );
  dff_sg \mask_0/reg_ii_mask_reg[24]  ( .D(\mask_0/n635 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[24] ) );
  dff_sg \mask_0/reg_ii_mask_reg[25]  ( .D(\mask_0/n636 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[25] ) );
  dff_sg \mask_0/reg_ii_mask_reg[26]  ( .D(\mask_0/n637 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[26] ) );
  dff_sg \mask_0/reg_ii_mask_reg[27]  ( .D(\mask_0/n638 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[27] ) );
  dff_sg \mask_0/reg_ii_mask_reg[28]  ( .D(\mask_0/n639 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[28] ) );
  dff_sg \mask_0/reg_ii_mask_reg[29]  ( .D(\mask_0/n640 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[29] ) );
  dff_sg \mask_0/reg_ii_mask_reg[30]  ( .D(\mask_0/n641 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[30] ) );
  dff_sg \mask_0/reg_ii_mask_reg[31]  ( .D(\mask_0/n642 ), .CP(clk), .Q(
        \mask_0/reg_ii_mask[31] ) );
  dff_sg \mask_0/reg_ww_mask_reg[0]  ( .D(\mask_0/n643 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[0] ) );
  dff_sg \mask_0/reg_ww_mask_reg[1]  ( .D(\mask_0/n644 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[1] ) );
  dff_sg \mask_0/reg_ww_mask_reg[2]  ( .D(\mask_0/n645 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[2] ) );
  dff_sg \mask_0/reg_ww_mask_reg[3]  ( .D(\mask_0/n646 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[3] ) );
  dff_sg \mask_0/reg_ww_mask_reg[4]  ( .D(\mask_0/n647 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[4] ) );
  dff_sg \mask_0/reg_ww_mask_reg[5]  ( .D(\mask_0/n648 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[5] ) );
  dff_sg \mask_0/reg_ww_mask_reg[6]  ( .D(\mask_0/n649 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[6] ) );
  dff_sg \mask_0/reg_ww_mask_reg[7]  ( .D(\mask_0/n650 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[7] ) );
  dff_sg \mask_0/reg_ww_mask_reg[8]  ( .D(\mask_0/n651 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[8] ) );
  dff_sg \mask_0/reg_ww_mask_reg[9]  ( .D(\mask_0/n652 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[9] ) );
  dff_sg \mask_0/reg_ww_mask_reg[10]  ( .D(\mask_0/n653 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[10] ) );
  dff_sg \mask_0/reg_ww_mask_reg[11]  ( .D(\mask_0/n654 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[11] ) );
  dff_sg \mask_0/reg_ww_mask_reg[12]  ( .D(\mask_0/n655 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[12] ) );
  dff_sg \mask_0/reg_ww_mask_reg[13]  ( .D(\mask_0/n656 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[13] ) );
  dff_sg \mask_0/reg_ww_mask_reg[14]  ( .D(\mask_0/n657 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[14] ) );
  dff_sg \mask_0/reg_ww_mask_reg[15]  ( .D(\mask_0/n658 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[15] ) );
  dff_sg \mask_0/reg_ww_mask_reg[16]  ( .D(\mask_0/n659 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[16] ) );
  dff_sg \mask_0/reg_ww_mask_reg[17]  ( .D(\mask_0/n660 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[17] ) );
  dff_sg \mask_0/reg_ww_mask_reg[18]  ( .D(\mask_0/n661 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[18] ) );
  dff_sg \mask_0/reg_ww_mask_reg[19]  ( .D(\mask_0/n662 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[19] ) );
  dff_sg \mask_0/reg_ww_mask_reg[20]  ( .D(\mask_0/n663 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[20] ) );
  dff_sg \mask_0/reg_ww_mask_reg[21]  ( .D(\mask_0/n664 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[21] ) );
  dff_sg \mask_0/reg_ww_mask_reg[22]  ( .D(\mask_0/n665 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[22] ) );
  dff_sg \mask_0/reg_ww_mask_reg[23]  ( .D(\mask_0/n666 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[23] ) );
  dff_sg \mask_0/reg_ww_mask_reg[24]  ( .D(\mask_0/n667 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[24] ) );
  dff_sg \mask_0/reg_ww_mask_reg[25]  ( .D(\mask_0/n668 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[25] ) );
  dff_sg \mask_0/reg_ww_mask_reg[26]  ( .D(\mask_0/n669 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[26] ) );
  dff_sg \mask_0/reg_ww_mask_reg[27]  ( .D(\mask_0/n670 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[27] ) );
  dff_sg \mask_0/reg_ww_mask_reg[28]  ( .D(\mask_0/n671 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[28] ) );
  dff_sg \mask_0/reg_ww_mask_reg[29]  ( .D(\mask_0/n672 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[29] ) );
  dff_sg \mask_0/reg_ww_mask_reg[30]  ( .D(\mask_0/n673 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[30] ) );
  dff_sg \mask_0/reg_ww_mask_reg[31]  ( .D(\mask_0/n674 ), .CP(clk), .Q(
        \mask_0/reg_ww_mask[31] ) );
  dff_sg \mask_0/reg_o_mask_reg[0]  ( .D(\mask_0/n675 ), .CP(clk), .Q(
        o_mask[0]) );
  dff_sg \mask_0/reg_o_mask_reg[1]  ( .D(\mask_0/n676 ), .CP(clk), .Q(
        o_mask[1]) );
  dff_sg \mask_0/reg_o_mask_reg[2]  ( .D(\mask_0/n677 ), .CP(clk), .Q(
        o_mask[2]) );
  dff_sg \mask_0/reg_o_mask_reg[3]  ( .D(\mask_0/n678 ), .CP(clk), .Q(
        o_mask[3]) );
  dff_sg \mask_0/reg_o_mask_reg[4]  ( .D(\mask_0/n679 ), .CP(clk), .Q(
        o_mask[4]) );
  dff_sg \mask_0/reg_o_mask_reg[5]  ( .D(\mask_0/n680 ), .CP(clk), .Q(
        o_mask[5]) );
  dff_sg \mask_0/reg_o_mask_reg[6]  ( .D(\mask_0/n681 ), .CP(clk), .Q(
        o_mask[6]) );
  dff_sg \mask_0/reg_o_mask_reg[7]  ( .D(\mask_0/n682 ), .CP(clk), .Q(
        o_mask[7]) );
  dff_sg \mask_0/reg_o_mask_reg[8]  ( .D(\mask_0/n683 ), .CP(clk), .Q(
        o_mask[8]) );
  dff_sg \mask_0/reg_o_mask_reg[9]  ( .D(\mask_0/n684 ), .CP(clk), .Q(
        o_mask[9]) );
  dff_sg \mask_0/reg_o_mask_reg[10]  ( .D(\mask_0/n685 ), .CP(clk), .Q(
        o_mask[10]) );
  dff_sg \mask_0/reg_o_mask_reg[11]  ( .D(\mask_0/n686 ), .CP(clk), .Q(
        o_mask[11]) );
  dff_sg \mask_0/reg_o_mask_reg[12]  ( .D(\mask_0/n687 ), .CP(clk), .Q(
        o_mask[12]) );
  dff_sg \mask_0/reg_o_mask_reg[13]  ( .D(\mask_0/n688 ), .CP(clk), .Q(
        o_mask[13]) );
  dff_sg \mask_0/reg_o_mask_reg[14]  ( .D(\mask_0/n689 ), .CP(clk), .Q(
        o_mask[14]) );
  dff_sg \mask_0/reg_o_mask_reg[15]  ( .D(\mask_0/n690 ), .CP(clk), .Q(
        o_mask[15]) );
  dff_sg \mask_0/reg_o_mask_reg[16]  ( .D(\mask_0/n691 ), .CP(clk), .Q(
        o_mask[16]) );
  dff_sg \mask_0/reg_o_mask_reg[17]  ( .D(\mask_0/n692 ), .CP(clk), .Q(
        o_mask[17]) );
  dff_sg \mask_0/reg_o_mask_reg[18]  ( .D(\mask_0/n693 ), .CP(clk), .Q(
        o_mask[18]) );
  dff_sg \mask_0/reg_o_mask_reg[19]  ( .D(\mask_0/n694 ), .CP(clk), .Q(
        o_mask[19]) );
  dff_sg \mask_0/reg_o_mask_reg[20]  ( .D(\mask_0/n695 ), .CP(clk), .Q(
        o_mask[20]) );
  dff_sg \mask_0/reg_o_mask_reg[21]  ( .D(\mask_0/n696 ), .CP(clk), .Q(
        o_mask[21]) );
  dff_sg \mask_0/reg_o_mask_reg[22]  ( .D(\mask_0/n697 ), .CP(clk), .Q(
        o_mask[22]) );
  dff_sg \mask_0/reg_o_mask_reg[23]  ( .D(\mask_0/n698 ), .CP(clk), .Q(
        o_mask[23]) );
  dff_sg \mask_0/reg_o_mask_reg[24]  ( .D(\mask_0/n699 ), .CP(clk), .Q(
        o_mask[24]) );
  dff_sg \mask_0/reg_o_mask_reg[25]  ( .D(\mask_0/n700 ), .CP(clk), .Q(
        o_mask[25]) );
  dff_sg \mask_0/reg_o_mask_reg[26]  ( .D(\mask_0/n701 ), .CP(clk), .Q(
        o_mask[26]) );
  dff_sg \mask_0/reg_o_mask_reg[27]  ( .D(\mask_0/n702 ), .CP(clk), .Q(
        o_mask[27]) );
  dff_sg \mask_0/reg_o_mask_reg[28]  ( .D(\mask_0/n703 ), .CP(clk), .Q(
        o_mask[28]) );
  dff_sg \mask_0/reg_o_mask_reg[29]  ( .D(\mask_0/n704 ), .CP(clk), .Q(
        o_mask[29]) );
  dff_sg \mask_0/reg_o_mask_reg[30]  ( .D(\mask_0/n705 ), .CP(clk), .Q(
        o_mask[30]) );
  dff_sg \mask_0/reg_o_mask_reg[31]  ( .D(\mask_0/n706 ), .CP(clk), .Q(
        o_mask[31]) );
  dff_sg \mask_0/reg_i_mask_reg[0]  ( .D(\mask_0/n770 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[0] ) );
  dff_sg \mask_0/reg_i_mask_reg[1]  ( .D(\mask_0/n769 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[1] ) );
  dff_sg \mask_0/reg_i_mask_reg[2]  ( .D(\mask_0/n768 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[2] ) );
  dff_sg \mask_0/reg_i_mask_reg[3]  ( .D(\mask_0/n767 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[3] ) );
  dff_sg \mask_0/reg_i_mask_reg[4]  ( .D(\mask_0/n766 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[4] ) );
  dff_sg \mask_0/reg_i_mask_reg[5]  ( .D(\mask_0/n765 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[5] ) );
  dff_sg \mask_0/reg_i_mask_reg[6]  ( .D(\mask_0/n764 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[6] ) );
  dff_sg \mask_0/reg_i_mask_reg[7]  ( .D(\mask_0/n763 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[7] ) );
  dff_sg \mask_0/reg_i_mask_reg[8]  ( .D(\mask_0/n762 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[8] ) );
  dff_sg \mask_0/reg_i_mask_reg[9]  ( .D(\mask_0/n761 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[9] ) );
  dff_sg \mask_0/reg_i_mask_reg[10]  ( .D(\mask_0/n760 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[10] ) );
  dff_sg \mask_0/reg_i_mask_reg[11]  ( .D(\mask_0/n759 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[11] ) );
  dff_sg \mask_0/reg_i_mask_reg[12]  ( .D(\mask_0/n758 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[12] ) );
  dff_sg \mask_0/reg_i_mask_reg[13]  ( .D(\mask_0/n757 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[13] ) );
  dff_sg \mask_0/reg_i_mask_reg[14]  ( .D(\mask_0/n756 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[14] ) );
  dff_sg \mask_0/reg_i_mask_reg[15]  ( .D(\mask_0/n755 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[15] ) );
  dff_sg \mask_0/reg_i_mask_reg[16]  ( .D(\mask_0/n754 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[16] ) );
  dff_sg \mask_0/reg_i_mask_reg[17]  ( .D(\mask_0/n753 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[17] ) );
  dff_sg \mask_0/reg_i_mask_reg[18]  ( .D(\mask_0/n752 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[18] ) );
  dff_sg \mask_0/reg_i_mask_reg[19]  ( .D(\mask_0/n751 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[19] ) );
  dff_sg \mask_0/reg_i_mask_reg[20]  ( .D(\mask_0/n750 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[20] ) );
  dff_sg \mask_0/reg_i_mask_reg[21]  ( .D(\mask_0/n749 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[21] ) );
  dff_sg \mask_0/reg_i_mask_reg[22]  ( .D(\mask_0/n748 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[22] ) );
  dff_sg \mask_0/reg_i_mask_reg[23]  ( .D(\mask_0/n747 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[23] ) );
  dff_sg \mask_0/reg_i_mask_reg[24]  ( .D(\mask_0/n746 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[24] ) );
  dff_sg \mask_0/reg_i_mask_reg[25]  ( .D(\mask_0/n745 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[25] ) );
  dff_sg \mask_0/reg_i_mask_reg[26]  ( .D(\mask_0/n744 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[26] ) );
  dff_sg \mask_0/reg_i_mask_reg[27]  ( .D(\mask_0/n743 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[27] ) );
  dff_sg \mask_0/reg_i_mask_reg[28]  ( .D(\mask_0/n742 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[28] ) );
  dff_sg \mask_0/reg_i_mask_reg[29]  ( .D(\mask_0/n741 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[29] ) );
  dff_sg \mask_0/reg_i_mask_reg[30]  ( .D(\mask_0/n740 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[30] ) );
  dff_sg \mask_0/reg_i_mask_reg[31]  ( .D(\mask_0/n739 ), .CP(clk), .Q(
        \mask_0/reg_i_mask[31] ) );
  dff_sg \mask_0/reg_w_mask_reg[0]  ( .D(\mask_0/n738 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[0] ) );
  dff_sg \mask_0/reg_w_mask_reg[1]  ( .D(\mask_0/n737 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[1] ) );
  dff_sg \mask_0/reg_w_mask_reg[2]  ( .D(\mask_0/n736 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[2] ) );
  dff_sg \mask_0/reg_w_mask_reg[3]  ( .D(\mask_0/n735 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[3] ) );
  dff_sg \mask_0/reg_w_mask_reg[4]  ( .D(\mask_0/n734 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[4] ) );
  dff_sg \mask_0/reg_w_mask_reg[5]  ( .D(\mask_0/n733 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[5] ) );
  dff_sg \mask_0/reg_w_mask_reg[6]  ( .D(\mask_0/n732 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[6] ) );
  dff_sg \mask_0/reg_w_mask_reg[7]  ( .D(\mask_0/n731 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[7] ) );
  dff_sg \mask_0/reg_w_mask_reg[8]  ( .D(\mask_0/n730 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[8] ) );
  dff_sg \mask_0/reg_w_mask_reg[9]  ( .D(\mask_0/n729 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[9] ) );
  dff_sg \mask_0/reg_w_mask_reg[10]  ( .D(\mask_0/n728 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[10] ) );
  dff_sg \mask_0/reg_w_mask_reg[11]  ( .D(\mask_0/n727 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[11] ) );
  dff_sg \mask_0/reg_w_mask_reg[12]  ( .D(\mask_0/n726 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[12] ) );
  dff_sg \mask_0/reg_w_mask_reg[13]  ( .D(\mask_0/n725 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[13] ) );
  dff_sg \mask_0/reg_w_mask_reg[14]  ( .D(\mask_0/n724 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[14] ) );
  dff_sg \mask_0/reg_w_mask_reg[15]  ( .D(\mask_0/n723 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[15] ) );
  dff_sg \mask_0/reg_w_mask_reg[16]  ( .D(\mask_0/n722 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[16] ) );
  dff_sg \mask_0/reg_w_mask_reg[17]  ( .D(\mask_0/n721 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[17] ) );
  dff_sg \mask_0/reg_w_mask_reg[18]  ( .D(\mask_0/n720 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[18] ) );
  dff_sg \mask_0/reg_w_mask_reg[19]  ( .D(\mask_0/n719 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[19] ) );
  dff_sg \mask_0/reg_w_mask_reg[20]  ( .D(\mask_0/n718 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[20] ) );
  dff_sg \mask_0/reg_w_mask_reg[21]  ( .D(\mask_0/n717 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[21] ) );
  dff_sg \mask_0/reg_w_mask_reg[22]  ( .D(\mask_0/n716 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[22] ) );
  dff_sg \mask_0/reg_w_mask_reg[23]  ( .D(\mask_0/n715 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[23] ) );
  dff_sg \mask_0/reg_w_mask_reg[24]  ( .D(\mask_0/n714 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[24] ) );
  dff_sg \mask_0/reg_w_mask_reg[25]  ( .D(\mask_0/n713 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[25] ) );
  dff_sg \mask_0/reg_w_mask_reg[26]  ( .D(\mask_0/n712 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[26] ) );
  dff_sg \mask_0/reg_w_mask_reg[27]  ( .D(\mask_0/n711 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[27] ) );
  dff_sg \mask_0/reg_w_mask_reg[28]  ( .D(\mask_0/n710 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[28] ) );
  dff_sg \mask_0/reg_w_mask_reg[29]  ( .D(\mask_0/n709 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[29] ) );
  dff_sg \mask_0/reg_w_mask_reg[30]  ( .D(\mask_0/n708 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[30] ) );
  dff_sg \mask_0/reg_w_mask_reg[31]  ( .D(\mask_0/n707 ), .CP(clk), .Q(
        \mask_0/reg_w_mask[31] ) );
  dff_sg \mask_0/state_reg[0]  ( .D(\mask_0/n771 ), .CP(clk), .Q(
        \mask_0/state[0] ) );
  dff_sg \mask_0/state_reg[1]  ( .D(\mask_0/n772 ), .CP(clk), .Q(
        \mask_0/state[1] ) );
  dff_sg \mask_0/counter_reg[1]  ( .D(\mask_0/n773 ), .CP(clk), .Q(
        \mask_0/counter[1] ) );
  dff_sg \mask_0/counter_reg[0]  ( .D(\mask_0/n774 ), .CP(clk), .Q(
        \mask_0/counter[0] ) );
  dff_sg \filter_0/oi_8_reg[19]  ( .D(\filter_0/n8588 ), .CP(clk), .Q(
        reg_oi_8[19]) );
  dff_sg \filter_0/oi_8_reg[18]  ( .D(\filter_0/n8589 ), .CP(clk), .Q(
        reg_oi_8[18]) );
  dff_sg \filter_0/oi_8_reg[17]  ( .D(\filter_0/n8590 ), .CP(clk), .Q(
        reg_oi_8[17]) );
  dff_sg \filter_0/oi_8_reg[16]  ( .D(\filter_0/n8591 ), .CP(clk), .Q(
        reg_oi_8[16]) );
  dff_sg \filter_0/oi_8_reg[15]  ( .D(\filter_0/n8592 ), .CP(clk), .Q(
        reg_oi_8[15]) );
  dff_sg \filter_0/oi_8_reg[14]  ( .D(\filter_0/n8593 ), .CP(clk), .Q(
        reg_oi_8[14]) );
  dff_sg \filter_0/oi_8_reg[13]  ( .D(\filter_0/n8594 ), .CP(clk), .Q(
        reg_oi_8[13]) );
  dff_sg \filter_0/oi_8_reg[12]  ( .D(\filter_0/n8595 ), .CP(clk), .Q(
        reg_oi_8[12]) );
  dff_sg \filter_0/oi_8_reg[11]  ( .D(\filter_0/n8596 ), .CP(clk), .Q(
        reg_oi_8[11]) );
  dff_sg \filter_0/oi_8_reg[10]  ( .D(\filter_0/n8597 ), .CP(clk), .Q(
        reg_oi_8[10]) );
  dff_sg \filter_0/oi_8_reg[9]  ( .D(\filter_0/n8598 ), .CP(clk), .Q(
        reg_oi_8[9]) );
  dff_sg \filter_0/oi_8_reg[8]  ( .D(\filter_0/n8599 ), .CP(clk), .Q(
        reg_oi_8[8]) );
  dff_sg \filter_0/oi_8_reg[7]  ( .D(\filter_0/n8600 ), .CP(clk), .Q(
        reg_oi_8[7]) );
  dff_sg \filter_0/oi_8_reg[6]  ( .D(\filter_0/n8601 ), .CP(clk), .Q(
        reg_oi_8[6]) );
  dff_sg \filter_0/oi_8_reg[5]  ( .D(\filter_0/n8602 ), .CP(clk), .Q(
        reg_oi_8[5]) );
  dff_sg \filter_0/oi_8_reg[4]  ( .D(\filter_0/n8603 ), .CP(clk), .Q(
        reg_oi_8[4]) );
  dff_sg \filter_0/oi_8_reg[3]  ( .D(\filter_0/n8604 ), .CP(clk), .Q(
        reg_oi_8[3]) );
  dff_sg \filter_0/oi_8_reg[2]  ( .D(\filter_0/n8605 ), .CP(clk), .Q(
        reg_oi_8[2]) );
  dff_sg \filter_0/oi_8_reg[1]  ( .D(\filter_0/n8606 ), .CP(clk), .Q(
        reg_oi_8[1]) );
  dff_sg \filter_0/oi_8_reg[0]  ( .D(\filter_0/n8607 ), .CP(clk), .Q(
        reg_oi_8[0]) );
  dff_sg \filter_0/oi_9_reg[19]  ( .D(\filter_0/n8608 ), .CP(clk), .Q(
        reg_oi_9[19]) );
  dff_sg \filter_0/oi_9_reg[18]  ( .D(\filter_0/n8609 ), .CP(clk), .Q(
        reg_oi_9[18]) );
  dff_sg \filter_0/oi_9_reg[17]  ( .D(\filter_0/n8610 ), .CP(clk), .Q(
        reg_oi_9[17]) );
  dff_sg \filter_0/oi_9_reg[16]  ( .D(\filter_0/n8611 ), .CP(clk), .Q(
        reg_oi_9[16]) );
  dff_sg \filter_0/oi_9_reg[15]  ( .D(\filter_0/n8612 ), .CP(clk), .Q(
        reg_oi_9[15]) );
  dff_sg \filter_0/oi_9_reg[14]  ( .D(\filter_0/n8613 ), .CP(clk), .Q(
        reg_oi_9[14]) );
  dff_sg \filter_0/oi_9_reg[13]  ( .D(\filter_0/n8614 ), .CP(clk), .Q(
        reg_oi_9[13]) );
  dff_sg \filter_0/oi_9_reg[12]  ( .D(\filter_0/n8615 ), .CP(clk), .Q(
        reg_oi_9[12]) );
  dff_sg \filter_0/oi_9_reg[11]  ( .D(\filter_0/n8616 ), .CP(clk), .Q(
        reg_oi_9[11]) );
  dff_sg \filter_0/oi_9_reg[10]  ( .D(\filter_0/n8617 ), .CP(clk), .Q(
        reg_oi_9[10]) );
  dff_sg \filter_0/oi_9_reg[9]  ( .D(\filter_0/n8618 ), .CP(clk), .Q(
        reg_oi_9[9]) );
  dff_sg \filter_0/oi_9_reg[8]  ( .D(\filter_0/n8619 ), .CP(clk), .Q(
        reg_oi_9[8]) );
  dff_sg \filter_0/oi_9_reg[7]  ( .D(\filter_0/n8620 ), .CP(clk), .Q(
        reg_oi_9[7]) );
  dff_sg \filter_0/oi_9_reg[6]  ( .D(\filter_0/n8621 ), .CP(clk), .Q(
        reg_oi_9[6]) );
  dff_sg \filter_0/oi_9_reg[5]  ( .D(\filter_0/n8622 ), .CP(clk), .Q(
        reg_oi_9[5]) );
  dff_sg \filter_0/oi_9_reg[4]  ( .D(\filter_0/n8623 ), .CP(clk), .Q(
        reg_oi_9[4]) );
  dff_sg \filter_0/oi_9_reg[3]  ( .D(\filter_0/n8624 ), .CP(clk), .Q(
        reg_oi_9[3]) );
  dff_sg \filter_0/oi_9_reg[2]  ( .D(\filter_0/n8625 ), .CP(clk), .Q(
        reg_oi_9[2]) );
  dff_sg \filter_0/oi_9_reg[1]  ( .D(\filter_0/n8626 ), .CP(clk), .Q(
        reg_oi_9[1]) );
  dff_sg \filter_0/oi_9_reg[0]  ( .D(\filter_0/n8627 ), .CP(clk), .Q(
        reg_oi_9[0]) );
  dff_sg \filter_0/oi_10_reg[19]  ( .D(\filter_0/n8628 ), .CP(clk), .Q(
        reg_oi_10[19]) );
  dff_sg \filter_0/oi_10_reg[18]  ( .D(\filter_0/n8629 ), .CP(clk), .Q(
        reg_oi_10[18]) );
  dff_sg \filter_0/oi_10_reg[17]  ( .D(\filter_0/n8630 ), .CP(clk), .Q(
        reg_oi_10[17]) );
  dff_sg \filter_0/oi_10_reg[16]  ( .D(\filter_0/n8631 ), .CP(clk), .Q(
        reg_oi_10[16]) );
  dff_sg \filter_0/oi_10_reg[15]  ( .D(\filter_0/n8632 ), .CP(clk), .Q(
        reg_oi_10[15]) );
  dff_sg \filter_0/oi_10_reg[14]  ( .D(\filter_0/n8633 ), .CP(clk), .Q(
        reg_oi_10[14]) );
  dff_sg \filter_0/oi_10_reg[13]  ( .D(\filter_0/n8634 ), .CP(clk), .Q(
        reg_oi_10[13]) );
  dff_sg \filter_0/oi_10_reg[12]  ( .D(\filter_0/n8635 ), .CP(clk), .Q(
        reg_oi_10[12]) );
  dff_sg \filter_0/oi_10_reg[11]  ( .D(\filter_0/n8636 ), .CP(clk), .Q(
        reg_oi_10[11]) );
  dff_sg \filter_0/oi_10_reg[10]  ( .D(\filter_0/n8637 ), .CP(clk), .Q(
        reg_oi_10[10]) );
  dff_sg \filter_0/oi_10_reg[9]  ( .D(\filter_0/n8638 ), .CP(clk), .Q(
        reg_oi_10[9]) );
  dff_sg \filter_0/oi_10_reg[8]  ( .D(\filter_0/n8639 ), .CP(clk), .Q(
        reg_oi_10[8]) );
  dff_sg \filter_0/oi_10_reg[7]  ( .D(\filter_0/n8640 ), .CP(clk), .Q(
        reg_oi_10[7]) );
  dff_sg \filter_0/oi_10_reg[6]  ( .D(\filter_0/n8641 ), .CP(clk), .Q(
        reg_oi_10[6]) );
  dff_sg \filter_0/oi_10_reg[5]  ( .D(\filter_0/n8642 ), .CP(clk), .Q(
        reg_oi_10[5]) );
  dff_sg \filter_0/oi_10_reg[4]  ( .D(\filter_0/n8643 ), .CP(clk), .Q(
        reg_oi_10[4]) );
  dff_sg \filter_0/oi_10_reg[3]  ( .D(\filter_0/n8644 ), .CP(clk), .Q(
        reg_oi_10[3]) );
  dff_sg \filter_0/oi_10_reg[2]  ( .D(\filter_0/n8645 ), .CP(clk), .Q(
        reg_oi_10[2]) );
  dff_sg \filter_0/oi_10_reg[1]  ( .D(\filter_0/n8646 ), .CP(clk), .Q(
        reg_oi_10[1]) );
  dff_sg \filter_0/oi_10_reg[0]  ( .D(\filter_0/n8647 ), .CP(clk), .Q(
        reg_oi_10[0]) );
  dff_sg \filter_0/oi_11_reg[19]  ( .D(\filter_0/n8648 ), .CP(clk), .Q(
        reg_oi_11[19]) );
  dff_sg \filter_0/oi_11_reg[18]  ( .D(\filter_0/n8649 ), .CP(clk), .Q(
        reg_oi_11[18]) );
  dff_sg \filter_0/oi_11_reg[17]  ( .D(\filter_0/n8650 ), .CP(clk), .Q(
        reg_oi_11[17]) );
  dff_sg \filter_0/oi_11_reg[16]  ( .D(\filter_0/n8651 ), .CP(clk), .Q(
        reg_oi_11[16]) );
  dff_sg \filter_0/oi_11_reg[15]  ( .D(\filter_0/n8652 ), .CP(clk), .Q(
        reg_oi_11[15]) );
  dff_sg \filter_0/oi_11_reg[14]  ( .D(\filter_0/n8653 ), .CP(clk), .Q(
        reg_oi_11[14]) );
  dff_sg \filter_0/oi_11_reg[13]  ( .D(\filter_0/n8654 ), .CP(clk), .Q(
        reg_oi_11[13]) );
  dff_sg \filter_0/oi_11_reg[12]  ( .D(\filter_0/n8655 ), .CP(clk), .Q(
        reg_oi_11[12]) );
  dff_sg \filter_0/oi_11_reg[11]  ( .D(\filter_0/n8656 ), .CP(clk), .Q(
        reg_oi_11[11]) );
  dff_sg \filter_0/oi_11_reg[10]  ( .D(\filter_0/n8657 ), .CP(clk), .Q(
        reg_oi_11[10]) );
  dff_sg \filter_0/oi_11_reg[9]  ( .D(\filter_0/n8658 ), .CP(clk), .Q(
        reg_oi_11[9]) );
  dff_sg \filter_0/oi_11_reg[8]  ( .D(\filter_0/n8659 ), .CP(clk), .Q(
        reg_oi_11[8]) );
  dff_sg \filter_0/oi_11_reg[7]  ( .D(\filter_0/n8660 ), .CP(clk), .Q(
        reg_oi_11[7]) );
  dff_sg \filter_0/oi_11_reg[6]  ( .D(\filter_0/n8661 ), .CP(clk), .Q(
        reg_oi_11[6]) );
  dff_sg \filter_0/oi_11_reg[5]  ( .D(\filter_0/n8662 ), .CP(clk), .Q(
        reg_oi_11[5]) );
  dff_sg \filter_0/oi_11_reg[4]  ( .D(\filter_0/n8663 ), .CP(clk), .Q(
        reg_oi_11[4]) );
  dff_sg \filter_0/oi_11_reg[3]  ( .D(\filter_0/n8664 ), .CP(clk), .Q(
        reg_oi_11[3]) );
  dff_sg \filter_0/oi_11_reg[2]  ( .D(\filter_0/n8665 ), .CP(clk), .Q(
        reg_oi_11[2]) );
  dff_sg \filter_0/oi_11_reg[1]  ( .D(\filter_0/n8666 ), .CP(clk), .Q(
        reg_oi_11[1]) );
  dff_sg \filter_0/oi_11_reg[0]  ( .D(\filter_0/n8667 ), .CP(clk), .Q(
        reg_oi_11[0]) );
  dff_sg \filter_0/oi_15_reg[19]  ( .D(\filter_0/n8728 ), .CP(clk), .Q(
        reg_oi_15[19]) );
  dff_sg \filter_0/oi_15_reg[18]  ( .D(\filter_0/n8729 ), .CP(clk), .Q(
        reg_oi_15[18]) );
  dff_sg \filter_0/oi_15_reg[17]  ( .D(\filter_0/n8730 ), .CP(clk), .Q(
        reg_oi_15[17]) );
  dff_sg \filter_0/oi_15_reg[16]  ( .D(\filter_0/n8731 ), .CP(clk), .Q(
        reg_oi_15[16]) );
  dff_sg \filter_0/oi_15_reg[15]  ( .D(\filter_0/n8732 ), .CP(clk), .Q(
        reg_oi_15[15]) );
  dff_sg \filter_0/oi_15_reg[14]  ( .D(\filter_0/n8733 ), .CP(clk), .Q(
        reg_oi_15[14]) );
  dff_sg \filter_0/oi_15_reg[13]  ( .D(\filter_0/n8734 ), .CP(clk), .Q(
        reg_oi_15[13]) );
  dff_sg \filter_0/oi_15_reg[12]  ( .D(\filter_0/n8735 ), .CP(clk), .Q(
        reg_oi_15[12]) );
  dff_sg \filter_0/oi_15_reg[11]  ( .D(\filter_0/n8736 ), .CP(clk), .Q(
        reg_oi_15[11]) );
  dff_sg \filter_0/oi_15_reg[10]  ( .D(\filter_0/n8737 ), .CP(clk), .Q(
        reg_oi_15[10]) );
  dff_sg \filter_0/oi_15_reg[9]  ( .D(\filter_0/n8738 ), .CP(clk), .Q(
        reg_oi_15[9]) );
  dff_sg \filter_0/oi_15_reg[8]  ( .D(\filter_0/n8739 ), .CP(clk), .Q(
        reg_oi_15[8]) );
  dff_sg \filter_0/oi_15_reg[7]  ( .D(\filter_0/n8740 ), .CP(clk), .Q(
        reg_oi_15[7]) );
  dff_sg \filter_0/oi_15_reg[6]  ( .D(\filter_0/n8741 ), .CP(clk), .Q(
        reg_oi_15[6]) );
  dff_sg \filter_0/oi_15_reg[5]  ( .D(\filter_0/n8742 ), .CP(clk), .Q(
        reg_oi_15[5]) );
  dff_sg \filter_0/oi_15_reg[4]  ( .D(\filter_0/n8743 ), .CP(clk), .Q(
        reg_oi_15[4]) );
  dff_sg \filter_0/oi_15_reg[3]  ( .D(\filter_0/n8744 ), .CP(clk), .Q(
        reg_oi_15[3]) );
  dff_sg \filter_0/oi_15_reg[2]  ( .D(\filter_0/n8745 ), .CP(clk), .Q(
        reg_oi_15[2]) );
  dff_sg \filter_0/oi_15_reg[1]  ( .D(\filter_0/n8746 ), .CP(clk), .Q(
        reg_oi_15[1]) );
  dff_sg \filter_0/oi_15_reg[0]  ( .D(\filter_0/n8747 ), .CP(clk), .Q(
        reg_oi_15[0]) );
  dff_sg \filter_0/oi_12_reg[19]  ( .D(\filter_0/n8668 ), .CP(clk), .Q(
        reg_oi_12[19]) );
  dff_sg \filter_0/oi_12_reg[18]  ( .D(\filter_0/n8669 ), .CP(clk), .Q(
        reg_oi_12[18]) );
  dff_sg \filter_0/oi_12_reg[17]  ( .D(\filter_0/n8670 ), .CP(clk), .Q(
        reg_oi_12[17]) );
  dff_sg \filter_0/oi_12_reg[16]  ( .D(\filter_0/n8671 ), .CP(clk), .Q(
        reg_oi_12[16]) );
  dff_sg \filter_0/oi_12_reg[15]  ( .D(\filter_0/n8672 ), .CP(clk), .Q(
        reg_oi_12[15]) );
  dff_sg \filter_0/oi_12_reg[14]  ( .D(\filter_0/n8673 ), .CP(clk), .Q(
        reg_oi_12[14]) );
  dff_sg \filter_0/oi_12_reg[13]  ( .D(\filter_0/n8674 ), .CP(clk), .Q(
        reg_oi_12[13]) );
  dff_sg \filter_0/oi_12_reg[12]  ( .D(\filter_0/n8675 ), .CP(clk), .Q(
        reg_oi_12[12]) );
  dff_sg \filter_0/oi_12_reg[11]  ( .D(\filter_0/n8676 ), .CP(clk), .Q(
        reg_oi_12[11]) );
  dff_sg \filter_0/oi_12_reg[10]  ( .D(\filter_0/n8677 ), .CP(clk), .Q(
        reg_oi_12[10]) );
  dff_sg \filter_0/oi_12_reg[9]  ( .D(\filter_0/n8678 ), .CP(clk), .Q(
        reg_oi_12[9]) );
  dff_sg \filter_0/oi_12_reg[8]  ( .D(\filter_0/n8679 ), .CP(clk), .Q(
        reg_oi_12[8]) );
  dff_sg \filter_0/oi_12_reg[7]  ( .D(\filter_0/n8680 ), .CP(clk), .Q(
        reg_oi_12[7]) );
  dff_sg \filter_0/oi_12_reg[6]  ( .D(\filter_0/n8681 ), .CP(clk), .Q(
        reg_oi_12[6]) );
  dff_sg \filter_0/oi_12_reg[5]  ( .D(\filter_0/n8682 ), .CP(clk), .Q(
        reg_oi_12[5]) );
  dff_sg \filter_0/oi_12_reg[4]  ( .D(\filter_0/n8683 ), .CP(clk), .Q(
        reg_oi_12[4]) );
  dff_sg \filter_0/oi_12_reg[3]  ( .D(\filter_0/n8684 ), .CP(clk), .Q(
        reg_oi_12[3]) );
  dff_sg \filter_0/oi_12_reg[2]  ( .D(\filter_0/n8685 ), .CP(clk), .Q(
        reg_oi_12[2]) );
  dff_sg \filter_0/oi_12_reg[1]  ( .D(\filter_0/n8686 ), .CP(clk), .Q(
        reg_oi_12[1]) );
  dff_sg \filter_0/oi_12_reg[0]  ( .D(\filter_0/n8687 ), .CP(clk), .Q(
        reg_oi_12[0]) );
  dff_sg \filter_0/oi_13_reg[19]  ( .D(\filter_0/n8688 ), .CP(clk), .Q(
        reg_oi_13[19]) );
  dff_sg \filter_0/oi_13_reg[18]  ( .D(\filter_0/n8689 ), .CP(clk), .Q(
        reg_oi_13[18]) );
  dff_sg \filter_0/oi_13_reg[17]  ( .D(\filter_0/n8690 ), .CP(clk), .Q(
        reg_oi_13[17]) );
  dff_sg \filter_0/oi_13_reg[16]  ( .D(\filter_0/n8691 ), .CP(clk), .Q(
        reg_oi_13[16]) );
  dff_sg \filter_0/oi_13_reg[15]  ( .D(\filter_0/n8692 ), .CP(clk), .Q(
        reg_oi_13[15]) );
  dff_sg \filter_0/oi_13_reg[14]  ( .D(\filter_0/n8693 ), .CP(clk), .Q(
        reg_oi_13[14]) );
  dff_sg \filter_0/oi_13_reg[13]  ( .D(\filter_0/n8694 ), .CP(clk), .Q(
        reg_oi_13[13]) );
  dff_sg \filter_0/oi_13_reg[12]  ( .D(\filter_0/n8695 ), .CP(clk), .Q(
        reg_oi_13[12]) );
  dff_sg \filter_0/oi_13_reg[11]  ( .D(\filter_0/n8696 ), .CP(clk), .Q(
        reg_oi_13[11]) );
  dff_sg \filter_0/oi_13_reg[10]  ( .D(\filter_0/n8697 ), .CP(clk), .Q(
        reg_oi_13[10]) );
  dff_sg \filter_0/oi_13_reg[9]  ( .D(\filter_0/n8698 ), .CP(clk), .Q(
        reg_oi_13[9]) );
  dff_sg \filter_0/oi_13_reg[8]  ( .D(\filter_0/n8699 ), .CP(clk), .Q(
        reg_oi_13[8]) );
  dff_sg \filter_0/oi_13_reg[7]  ( .D(\filter_0/n8700 ), .CP(clk), .Q(
        reg_oi_13[7]) );
  dff_sg \filter_0/oi_13_reg[6]  ( .D(\filter_0/n8701 ), .CP(clk), .Q(
        reg_oi_13[6]) );
  dff_sg \filter_0/oi_13_reg[5]  ( .D(\filter_0/n8702 ), .CP(clk), .Q(
        reg_oi_13[5]) );
  dff_sg \filter_0/oi_13_reg[4]  ( .D(\filter_0/n8703 ), .CP(clk), .Q(
        reg_oi_13[4]) );
  dff_sg \filter_0/oi_13_reg[3]  ( .D(\filter_0/n8704 ), .CP(clk), .Q(
        reg_oi_13[3]) );
  dff_sg \filter_0/oi_13_reg[2]  ( .D(\filter_0/n8705 ), .CP(clk), .Q(
        reg_oi_13[2]) );
  dff_sg \filter_0/oi_13_reg[1]  ( .D(\filter_0/n8706 ), .CP(clk), .Q(
        reg_oi_13[1]) );
  dff_sg \filter_0/oi_13_reg[0]  ( .D(\filter_0/n8707 ), .CP(clk), .Q(
        reg_oi_13[0]) );
  dff_sg \filter_0/oi_14_reg[19]  ( .D(\filter_0/n8708 ), .CP(clk), .Q(
        reg_oi_14[19]) );
  dff_sg \filter_0/oi_14_reg[18]  ( .D(\filter_0/n8709 ), .CP(clk), .Q(
        reg_oi_14[18]) );
  dff_sg \filter_0/oi_14_reg[17]  ( .D(\filter_0/n8710 ), .CP(clk), .Q(
        reg_oi_14[17]) );
  dff_sg \filter_0/oi_14_reg[16]  ( .D(\filter_0/n8711 ), .CP(clk), .Q(
        reg_oi_14[16]) );
  dff_sg \filter_0/oi_14_reg[15]  ( .D(\filter_0/n8712 ), .CP(clk), .Q(
        reg_oi_14[15]) );
  dff_sg \filter_0/oi_14_reg[14]  ( .D(\filter_0/n8713 ), .CP(clk), .Q(
        reg_oi_14[14]) );
  dff_sg \filter_0/oi_14_reg[13]  ( .D(\filter_0/n8714 ), .CP(clk), .Q(
        reg_oi_14[13]) );
  dff_sg \filter_0/oi_14_reg[12]  ( .D(\filter_0/n8715 ), .CP(clk), .Q(
        reg_oi_14[12]) );
  dff_sg \filter_0/oi_14_reg[11]  ( .D(\filter_0/n8716 ), .CP(clk), .Q(
        reg_oi_14[11]) );
  dff_sg \filter_0/oi_14_reg[10]  ( .D(\filter_0/n8717 ), .CP(clk), .Q(
        reg_oi_14[10]) );
  dff_sg \filter_0/oi_14_reg[9]  ( .D(\filter_0/n8718 ), .CP(clk), .Q(
        reg_oi_14[9]) );
  dff_sg \filter_0/oi_14_reg[8]  ( .D(\filter_0/n8719 ), .CP(clk), .Q(
        reg_oi_14[8]) );
  dff_sg \filter_0/oi_14_reg[7]  ( .D(\filter_0/n8720 ), .CP(clk), .Q(
        reg_oi_14[7]) );
  dff_sg \filter_0/oi_14_reg[6]  ( .D(\filter_0/n8721 ), .CP(clk), .Q(
        reg_oi_14[6]) );
  dff_sg \filter_0/oi_14_reg[5]  ( .D(\filter_0/n8722 ), .CP(clk), .Q(
        reg_oi_14[5]) );
  dff_sg \filter_0/oi_14_reg[4]  ( .D(\filter_0/n8723 ), .CP(clk), .Q(
        reg_oi_14[4]) );
  dff_sg \filter_0/oi_14_reg[3]  ( .D(\filter_0/n8724 ), .CP(clk), .Q(
        reg_oi_14[3]) );
  dff_sg \filter_0/oi_14_reg[2]  ( .D(\filter_0/n8725 ), .CP(clk), .Q(
        reg_oi_14[2]) );
  dff_sg \filter_0/oi_14_reg[1]  ( .D(\filter_0/n8726 ), .CP(clk), .Q(
        reg_oi_14[1]) );
  dff_sg \filter_0/oi_14_reg[0]  ( .D(\filter_0/n8727 ), .CP(clk), .Q(
        reg_oi_14[0]) );
  dff_sg \filter_0/oi_4_reg[19]  ( .D(\filter_0/n8808 ), .CP(clk), .Q(
        reg_oi_4[19]) );
  dff_sg \filter_0/oi_4_reg[18]  ( .D(\filter_0/n8809 ), .CP(clk), .Q(
        reg_oi_4[18]) );
  dff_sg \filter_0/oi_4_reg[17]  ( .D(\filter_0/n8810 ), .CP(clk), .Q(
        reg_oi_4[17]) );
  dff_sg \filter_0/oi_4_reg[16]  ( .D(\filter_0/n8811 ), .CP(clk), .Q(
        reg_oi_4[16]) );
  dff_sg \filter_0/oi_4_reg[15]  ( .D(\filter_0/n8812 ), .CP(clk), .Q(
        reg_oi_4[15]) );
  dff_sg \filter_0/oi_4_reg[14]  ( .D(\filter_0/n8813 ), .CP(clk), .Q(
        reg_oi_4[14]) );
  dff_sg \filter_0/oi_4_reg[13]  ( .D(\filter_0/n8814 ), .CP(clk), .Q(
        reg_oi_4[13]) );
  dff_sg \filter_0/oi_4_reg[12]  ( .D(\filter_0/n8815 ), .CP(clk), .Q(
        reg_oi_4[12]) );
  dff_sg \filter_0/oi_4_reg[11]  ( .D(\filter_0/n8816 ), .CP(clk), .Q(
        reg_oi_4[11]) );
  dff_sg \filter_0/oi_4_reg[10]  ( .D(\filter_0/n8817 ), .CP(clk), .Q(
        reg_oi_4[10]) );
  dff_sg \filter_0/oi_4_reg[9]  ( .D(\filter_0/n8818 ), .CP(clk), .Q(
        reg_oi_4[9]) );
  dff_sg \filter_0/oi_4_reg[8]  ( .D(\filter_0/n8819 ), .CP(clk), .Q(
        reg_oi_4[8]) );
  dff_sg \filter_0/oi_4_reg[7]  ( .D(\filter_0/n8820 ), .CP(clk), .Q(
        reg_oi_4[7]) );
  dff_sg \filter_0/oi_4_reg[6]  ( .D(\filter_0/n8821 ), .CP(clk), .Q(
        reg_oi_4[6]) );
  dff_sg \filter_0/oi_4_reg[5]  ( .D(\filter_0/n8822 ), .CP(clk), .Q(
        reg_oi_4[5]) );
  dff_sg \filter_0/oi_4_reg[4]  ( .D(\filter_0/n8823 ), .CP(clk), .Q(
        reg_oi_4[4]) );
  dff_sg \filter_0/oi_4_reg[3]  ( .D(\filter_0/n8824 ), .CP(clk), .Q(
        reg_oi_4[3]) );
  dff_sg \filter_0/oi_4_reg[2]  ( .D(\filter_0/n8825 ), .CP(clk), .Q(
        reg_oi_4[2]) );
  dff_sg \filter_0/oi_4_reg[1]  ( .D(\filter_0/n8826 ), .CP(clk), .Q(
        reg_oi_4[1]) );
  dff_sg \filter_0/oi_4_reg[0]  ( .D(\filter_0/n8827 ), .CP(clk), .Q(
        reg_oi_4[0]) );
  dff_sg \filter_0/oi_5_reg[19]  ( .D(\filter_0/n8788 ), .CP(clk), .Q(
        reg_oi_5[19]) );
  dff_sg \filter_0/oi_5_reg[18]  ( .D(\filter_0/n8789 ), .CP(clk), .Q(
        reg_oi_5[18]) );
  dff_sg \filter_0/oi_5_reg[17]  ( .D(\filter_0/n8790 ), .CP(clk), .Q(
        reg_oi_5[17]) );
  dff_sg \filter_0/oi_5_reg[16]  ( .D(\filter_0/n8791 ), .CP(clk), .Q(
        reg_oi_5[16]) );
  dff_sg \filter_0/oi_5_reg[15]  ( .D(\filter_0/n8792 ), .CP(clk), .Q(
        reg_oi_5[15]) );
  dff_sg \filter_0/oi_5_reg[14]  ( .D(\filter_0/n8793 ), .CP(clk), .Q(
        reg_oi_5[14]) );
  dff_sg \filter_0/oi_5_reg[13]  ( .D(\filter_0/n8794 ), .CP(clk), .Q(
        reg_oi_5[13]) );
  dff_sg \filter_0/oi_5_reg[12]  ( .D(\filter_0/n8795 ), .CP(clk), .Q(
        reg_oi_5[12]) );
  dff_sg \filter_0/oi_5_reg[11]  ( .D(\filter_0/n8796 ), .CP(clk), .Q(
        reg_oi_5[11]) );
  dff_sg \filter_0/oi_5_reg[10]  ( .D(\filter_0/n8797 ), .CP(clk), .Q(
        reg_oi_5[10]) );
  dff_sg \filter_0/oi_5_reg[9]  ( .D(\filter_0/n8798 ), .CP(clk), .Q(
        reg_oi_5[9]) );
  dff_sg \filter_0/oi_5_reg[8]  ( .D(\filter_0/n8799 ), .CP(clk), .Q(
        reg_oi_5[8]) );
  dff_sg \filter_0/oi_5_reg[7]  ( .D(\filter_0/n8800 ), .CP(clk), .Q(
        reg_oi_5[7]) );
  dff_sg \filter_0/oi_5_reg[6]  ( .D(\filter_0/n8801 ), .CP(clk), .Q(
        reg_oi_5[6]) );
  dff_sg \filter_0/oi_5_reg[5]  ( .D(\filter_0/n8802 ), .CP(clk), .Q(
        reg_oi_5[5]) );
  dff_sg \filter_0/oi_5_reg[4]  ( .D(\filter_0/n8803 ), .CP(clk), .Q(
        reg_oi_5[4]) );
  dff_sg \filter_0/oi_5_reg[3]  ( .D(\filter_0/n8804 ), .CP(clk), .Q(
        reg_oi_5[3]) );
  dff_sg \filter_0/oi_5_reg[2]  ( .D(\filter_0/n8805 ), .CP(clk), .Q(
        reg_oi_5[2]) );
  dff_sg \filter_0/oi_5_reg[1]  ( .D(\filter_0/n8806 ), .CP(clk), .Q(
        reg_oi_5[1]) );
  dff_sg \filter_0/oi_5_reg[0]  ( .D(\filter_0/n8807 ), .CP(clk), .Q(
        reg_oi_5[0]) );
  dff_sg \filter_0/oi_6_reg[19]  ( .D(\filter_0/n8768 ), .CP(clk), .Q(
        reg_oi_6[19]) );
  dff_sg \filter_0/oi_6_reg[18]  ( .D(\filter_0/n8769 ), .CP(clk), .Q(
        reg_oi_6[18]) );
  dff_sg \filter_0/oi_6_reg[17]  ( .D(\filter_0/n8770 ), .CP(clk), .Q(
        reg_oi_6[17]) );
  dff_sg \filter_0/oi_6_reg[16]  ( .D(\filter_0/n8771 ), .CP(clk), .Q(
        reg_oi_6[16]) );
  dff_sg \filter_0/oi_6_reg[15]  ( .D(\filter_0/n8772 ), .CP(clk), .Q(
        reg_oi_6[15]) );
  dff_sg \filter_0/oi_6_reg[14]  ( .D(\filter_0/n8773 ), .CP(clk), .Q(
        reg_oi_6[14]) );
  dff_sg \filter_0/oi_6_reg[13]  ( .D(\filter_0/n8774 ), .CP(clk), .Q(
        reg_oi_6[13]) );
  dff_sg \filter_0/oi_6_reg[12]  ( .D(\filter_0/n8775 ), .CP(clk), .Q(
        reg_oi_6[12]) );
  dff_sg \filter_0/oi_6_reg[11]  ( .D(\filter_0/n8776 ), .CP(clk), .Q(
        reg_oi_6[11]) );
  dff_sg \filter_0/oi_6_reg[10]  ( .D(\filter_0/n8777 ), .CP(clk), .Q(
        reg_oi_6[10]) );
  dff_sg \filter_0/oi_6_reg[9]  ( .D(\filter_0/n8778 ), .CP(clk), .Q(
        reg_oi_6[9]) );
  dff_sg \filter_0/oi_6_reg[8]  ( .D(\filter_0/n8779 ), .CP(clk), .Q(
        reg_oi_6[8]) );
  dff_sg \filter_0/oi_6_reg[7]  ( .D(\filter_0/n8780 ), .CP(clk), .Q(
        reg_oi_6[7]) );
  dff_sg \filter_0/oi_6_reg[6]  ( .D(\filter_0/n8781 ), .CP(clk), .Q(
        reg_oi_6[6]) );
  dff_sg \filter_0/oi_6_reg[5]  ( .D(\filter_0/n8782 ), .CP(clk), .Q(
        reg_oi_6[5]) );
  dff_sg \filter_0/oi_6_reg[4]  ( .D(\filter_0/n8783 ), .CP(clk), .Q(
        reg_oi_6[4]) );
  dff_sg \filter_0/oi_6_reg[3]  ( .D(\filter_0/n8784 ), .CP(clk), .Q(
        reg_oi_6[3]) );
  dff_sg \filter_0/oi_6_reg[2]  ( .D(\filter_0/n8785 ), .CP(clk), .Q(
        reg_oi_6[2]) );
  dff_sg \filter_0/oi_6_reg[1]  ( .D(\filter_0/n8786 ), .CP(clk), .Q(
        reg_oi_6[1]) );
  dff_sg \filter_0/oi_6_reg[0]  ( .D(\filter_0/n8787 ), .CP(clk), .Q(
        reg_oi_6[0]) );
  dff_sg \filter_0/oi_7_reg[19]  ( .D(\filter_0/n8748 ), .CP(clk), .Q(
        reg_oi_7[19]) );
  dff_sg \filter_0/oi_7_reg[18]  ( .D(\filter_0/n8749 ), .CP(clk), .Q(
        reg_oi_7[18]) );
  dff_sg \filter_0/oi_7_reg[17]  ( .D(\filter_0/n8750 ), .CP(clk), .Q(
        reg_oi_7[17]) );
  dff_sg \filter_0/oi_7_reg[16]  ( .D(\filter_0/n8751 ), .CP(clk), .Q(
        reg_oi_7[16]) );
  dff_sg \filter_0/oi_7_reg[15]  ( .D(\filter_0/n8752 ), .CP(clk), .Q(
        reg_oi_7[15]) );
  dff_sg \filter_0/oi_7_reg[14]  ( .D(\filter_0/n8753 ), .CP(clk), .Q(
        reg_oi_7[14]) );
  dff_sg \filter_0/oi_7_reg[13]  ( .D(\filter_0/n8754 ), .CP(clk), .Q(
        reg_oi_7[13]) );
  dff_sg \filter_0/oi_7_reg[12]  ( .D(\filter_0/n8755 ), .CP(clk), .Q(
        reg_oi_7[12]) );
  dff_sg \filter_0/oi_7_reg[11]  ( .D(\filter_0/n8756 ), .CP(clk), .Q(
        reg_oi_7[11]) );
  dff_sg \filter_0/oi_7_reg[10]  ( .D(\filter_0/n8757 ), .CP(clk), .Q(
        reg_oi_7[10]) );
  dff_sg \filter_0/oi_7_reg[9]  ( .D(\filter_0/n8758 ), .CP(clk), .Q(
        reg_oi_7[9]) );
  dff_sg \filter_0/oi_7_reg[8]  ( .D(\filter_0/n8759 ), .CP(clk), .Q(
        reg_oi_7[8]) );
  dff_sg \filter_0/oi_7_reg[7]  ( .D(\filter_0/n8760 ), .CP(clk), .Q(
        reg_oi_7[7]) );
  dff_sg \filter_0/oi_7_reg[6]  ( .D(\filter_0/n8761 ), .CP(clk), .Q(
        reg_oi_7[6]) );
  dff_sg \filter_0/oi_7_reg[5]  ( .D(\filter_0/n8762 ), .CP(clk), .Q(
        reg_oi_7[5]) );
  dff_sg \filter_0/oi_7_reg[4]  ( .D(\filter_0/n8763 ), .CP(clk), .Q(
        reg_oi_7[4]) );
  dff_sg \filter_0/oi_7_reg[3]  ( .D(\filter_0/n8764 ), .CP(clk), .Q(
        reg_oi_7[3]) );
  dff_sg \filter_0/oi_7_reg[2]  ( .D(\filter_0/n8765 ), .CP(clk), .Q(
        reg_oi_7[2]) );
  dff_sg \filter_0/oi_7_reg[1]  ( .D(\filter_0/n8766 ), .CP(clk), .Q(
        reg_oi_7[1]) );
  dff_sg \filter_0/oi_7_reg[0]  ( .D(\filter_0/n8767 ), .CP(clk), .Q(
        reg_oi_7[0]) );
  dff_sg \filter_0/oi_0_reg[19]  ( .D(\filter_0/n8568 ), .CP(clk), .Q(
        reg_oi_0[19]) );
  dff_sg \filter_0/oi_0_reg[18]  ( .D(\filter_0/n8569 ), .CP(clk), .Q(
        reg_oi_0[18]) );
  dff_sg \filter_0/oi_0_reg[17]  ( .D(\filter_0/n8570 ), .CP(clk), .Q(
        reg_oi_0[17]) );
  dff_sg \filter_0/oi_0_reg[16]  ( .D(\filter_0/n8571 ), .CP(clk), .Q(
        reg_oi_0[16]) );
  dff_sg \filter_0/oi_0_reg[15]  ( .D(\filter_0/n8572 ), .CP(clk), .Q(
        reg_oi_0[15]) );
  dff_sg \filter_0/oi_0_reg[14]  ( .D(\filter_0/n8573 ), .CP(clk), .Q(
        reg_oi_0[14]) );
  dff_sg \filter_0/oi_0_reg[13]  ( .D(\filter_0/n8574 ), .CP(clk), .Q(
        reg_oi_0[13]) );
  dff_sg \filter_0/oi_0_reg[12]  ( .D(\filter_0/n8575 ), .CP(clk), .Q(
        reg_oi_0[12]) );
  dff_sg \filter_0/oi_0_reg[11]  ( .D(\filter_0/n8576 ), .CP(clk), .Q(
        reg_oi_0[11]) );
  dff_sg \filter_0/oi_0_reg[10]  ( .D(\filter_0/n8577 ), .CP(clk), .Q(
        reg_oi_0[10]) );
  dff_sg \filter_0/oi_0_reg[9]  ( .D(\filter_0/n8578 ), .CP(clk), .Q(
        reg_oi_0[9]) );
  dff_sg \filter_0/oi_0_reg[8]  ( .D(\filter_0/n8579 ), .CP(clk), .Q(
        reg_oi_0[8]) );
  dff_sg \filter_0/oi_0_reg[7]  ( .D(\filter_0/n8580 ), .CP(clk), .Q(
        reg_oi_0[7]) );
  dff_sg \filter_0/oi_0_reg[6]  ( .D(\filter_0/n8581 ), .CP(clk), .Q(
        reg_oi_0[6]) );
  dff_sg \filter_0/oi_0_reg[5]  ( .D(\filter_0/n8582 ), .CP(clk), .Q(
        reg_oi_0[5]) );
  dff_sg \filter_0/oi_0_reg[4]  ( .D(\filter_0/n8583 ), .CP(clk), .Q(
        reg_oi_0[4]) );
  dff_sg \filter_0/oi_0_reg[3]  ( .D(\filter_0/n8584 ), .CP(clk), .Q(
        reg_oi_0[3]) );
  dff_sg \filter_0/oi_0_reg[2]  ( .D(\filter_0/n8585 ), .CP(clk), .Q(
        reg_oi_0[2]) );
  dff_sg \filter_0/oi_0_reg[1]  ( .D(\filter_0/n8586 ), .CP(clk), .Q(
        reg_oi_0[1]) );
  dff_sg \filter_0/oi_0_reg[0]  ( .D(\filter_0/n8587 ), .CP(clk), .Q(
        reg_oi_0[0]) );
  dff_sg \filter_0/oi_1_reg[19]  ( .D(\filter_0/n8868 ), .CP(clk), .Q(
        reg_oi_1[19]) );
  dff_sg \filter_0/oi_1_reg[18]  ( .D(\filter_0/n8869 ), .CP(clk), .Q(
        reg_oi_1[18]) );
  dff_sg \filter_0/oi_1_reg[17]  ( .D(\filter_0/n8870 ), .CP(clk), .Q(
        reg_oi_1[17]) );
  dff_sg \filter_0/oi_1_reg[16]  ( .D(\filter_0/n8871 ), .CP(clk), .Q(
        reg_oi_1[16]) );
  dff_sg \filter_0/oi_1_reg[15]  ( .D(\filter_0/n8872 ), .CP(clk), .Q(
        reg_oi_1[15]) );
  dff_sg \filter_0/oi_1_reg[14]  ( .D(\filter_0/n8873 ), .CP(clk), .Q(
        reg_oi_1[14]) );
  dff_sg \filter_0/oi_1_reg[13]  ( .D(\filter_0/n8874 ), .CP(clk), .Q(
        reg_oi_1[13]) );
  dff_sg \filter_0/oi_1_reg[12]  ( .D(\filter_0/n8875 ), .CP(clk), .Q(
        reg_oi_1[12]) );
  dff_sg \filter_0/oi_1_reg[11]  ( .D(\filter_0/n8876 ), .CP(clk), .Q(
        reg_oi_1[11]) );
  dff_sg \filter_0/oi_1_reg[10]  ( .D(\filter_0/n8877 ), .CP(clk), .Q(
        reg_oi_1[10]) );
  dff_sg \filter_0/oi_1_reg[9]  ( .D(\filter_0/n8878 ), .CP(clk), .Q(
        reg_oi_1[9]) );
  dff_sg \filter_0/oi_1_reg[8]  ( .D(\filter_0/n8879 ), .CP(clk), .Q(
        reg_oi_1[8]) );
  dff_sg \filter_0/oi_1_reg[7]  ( .D(\filter_0/n8880 ), .CP(clk), .Q(
        reg_oi_1[7]) );
  dff_sg \filter_0/oi_1_reg[6]  ( .D(\filter_0/n8881 ), .CP(clk), .Q(
        reg_oi_1[6]) );
  dff_sg \filter_0/oi_1_reg[5]  ( .D(\filter_0/n8882 ), .CP(clk), .Q(
        reg_oi_1[5]) );
  dff_sg \filter_0/oi_1_reg[4]  ( .D(\filter_0/n8883 ), .CP(clk), .Q(
        reg_oi_1[4]) );
  dff_sg \filter_0/oi_1_reg[3]  ( .D(\filter_0/n8884 ), .CP(clk), .Q(
        reg_oi_1[3]) );
  dff_sg \filter_0/oi_1_reg[2]  ( .D(\filter_0/n8885 ), .CP(clk), .Q(
        reg_oi_1[2]) );
  dff_sg \filter_0/oi_1_reg[1]  ( .D(\filter_0/n8886 ), .CP(clk), .Q(
        reg_oi_1[1]) );
  dff_sg \filter_0/oi_1_reg[0]  ( .D(\filter_0/n8887 ), .CP(clk), .Q(
        reg_oi_1[0]) );
  dff_sg \filter_0/oi_2_reg[19]  ( .D(\filter_0/n8848 ), .CP(clk), .Q(
        reg_oi_2[19]) );
  dff_sg \filter_0/oi_2_reg[18]  ( .D(\filter_0/n8849 ), .CP(clk), .Q(
        reg_oi_2[18]) );
  dff_sg \filter_0/oi_2_reg[17]  ( .D(\filter_0/n8850 ), .CP(clk), .Q(
        reg_oi_2[17]) );
  dff_sg \filter_0/oi_2_reg[16]  ( .D(\filter_0/n8851 ), .CP(clk), .Q(
        reg_oi_2[16]) );
  dff_sg \filter_0/oi_2_reg[15]  ( .D(\filter_0/n8852 ), .CP(clk), .Q(
        reg_oi_2[15]) );
  dff_sg \filter_0/oi_2_reg[14]  ( .D(\filter_0/n8853 ), .CP(clk), .Q(
        reg_oi_2[14]) );
  dff_sg \filter_0/oi_2_reg[13]  ( .D(\filter_0/n8854 ), .CP(clk), .Q(
        reg_oi_2[13]) );
  dff_sg \filter_0/oi_2_reg[12]  ( .D(\filter_0/n8855 ), .CP(clk), .Q(
        reg_oi_2[12]) );
  dff_sg \filter_0/oi_2_reg[11]  ( .D(\filter_0/n8856 ), .CP(clk), .Q(
        reg_oi_2[11]) );
  dff_sg \filter_0/oi_2_reg[10]  ( .D(\filter_0/n8857 ), .CP(clk), .Q(
        reg_oi_2[10]) );
  dff_sg \filter_0/oi_2_reg[9]  ( .D(\filter_0/n8858 ), .CP(clk), .Q(
        reg_oi_2[9]) );
  dff_sg \filter_0/oi_2_reg[8]  ( .D(\filter_0/n8859 ), .CP(clk), .Q(
        reg_oi_2[8]) );
  dff_sg \filter_0/oi_2_reg[7]  ( .D(\filter_0/n8860 ), .CP(clk), .Q(
        reg_oi_2[7]) );
  dff_sg \filter_0/oi_2_reg[6]  ( .D(\filter_0/n8861 ), .CP(clk), .Q(
        reg_oi_2[6]) );
  dff_sg \filter_0/oi_2_reg[5]  ( .D(\filter_0/n8862 ), .CP(clk), .Q(
        reg_oi_2[5]) );
  dff_sg \filter_0/oi_2_reg[4]  ( .D(\filter_0/n8863 ), .CP(clk), .Q(
        reg_oi_2[4]) );
  dff_sg \filter_0/oi_2_reg[3]  ( .D(\filter_0/n8864 ), .CP(clk), .Q(
        reg_oi_2[3]) );
  dff_sg \filter_0/oi_2_reg[2]  ( .D(\filter_0/n8865 ), .CP(clk), .Q(
        reg_oi_2[2]) );
  dff_sg \filter_0/oi_2_reg[1]  ( .D(\filter_0/n8866 ), .CP(clk), .Q(
        reg_oi_2[1]) );
  dff_sg \filter_0/oi_2_reg[0]  ( .D(\filter_0/n8867 ), .CP(clk), .Q(
        reg_oi_2[0]) );
  dff_sg \filter_0/oi_3_reg[19]  ( .D(\filter_0/n8828 ), .CP(clk), .Q(
        reg_oi_3[19]) );
  dff_sg \filter_0/oi_3_reg[18]  ( .D(\filter_0/n8829 ), .CP(clk), .Q(
        reg_oi_3[18]) );
  dff_sg \filter_0/oi_3_reg[17]  ( .D(\filter_0/n8830 ), .CP(clk), .Q(
        reg_oi_3[17]) );
  dff_sg \filter_0/oi_3_reg[16]  ( .D(\filter_0/n8831 ), .CP(clk), .Q(
        reg_oi_3[16]) );
  dff_sg \filter_0/oi_3_reg[15]  ( .D(\filter_0/n8832 ), .CP(clk), .Q(
        reg_oi_3[15]) );
  dff_sg \filter_0/oi_3_reg[14]  ( .D(\filter_0/n8833 ), .CP(clk), .Q(
        reg_oi_3[14]) );
  dff_sg \filter_0/oi_3_reg[13]  ( .D(\filter_0/n8834 ), .CP(clk), .Q(
        reg_oi_3[13]) );
  dff_sg \filter_0/oi_3_reg[12]  ( .D(\filter_0/n8835 ), .CP(clk), .Q(
        reg_oi_3[12]) );
  dff_sg \filter_0/oi_3_reg[11]  ( .D(\filter_0/n8836 ), .CP(clk), .Q(
        reg_oi_3[11]) );
  dff_sg \filter_0/oi_3_reg[10]  ( .D(\filter_0/n8837 ), .CP(clk), .Q(
        reg_oi_3[10]) );
  dff_sg \filter_0/oi_3_reg[9]  ( .D(\filter_0/n8838 ), .CP(clk), .Q(
        reg_oi_3[9]) );
  dff_sg \filter_0/oi_3_reg[8]  ( .D(\filter_0/n8839 ), .CP(clk), .Q(
        reg_oi_3[8]) );
  dff_sg \filter_0/oi_3_reg[7]  ( .D(\filter_0/n8840 ), .CP(clk), .Q(
        reg_oi_3[7]) );
  dff_sg \filter_0/oi_3_reg[6]  ( .D(\filter_0/n8841 ), .CP(clk), .Q(
        reg_oi_3[6]) );
  dff_sg \filter_0/oi_3_reg[5]  ( .D(\filter_0/n8842 ), .CP(clk), .Q(
        reg_oi_3[5]) );
  dff_sg \filter_0/oi_3_reg[4]  ( .D(\filter_0/n8843 ), .CP(clk), .Q(
        reg_oi_3[4]) );
  dff_sg \filter_0/oi_3_reg[3]  ( .D(\filter_0/n8844 ), .CP(clk), .Q(
        reg_oi_3[3]) );
  dff_sg \filter_0/oi_3_reg[2]  ( .D(\filter_0/n8845 ), .CP(clk), .Q(
        reg_oi_3[2]) );
  dff_sg \filter_0/oi_3_reg[1]  ( .D(\filter_0/n8846 ), .CP(clk), .Q(
        reg_oi_3[1]) );
  dff_sg \filter_0/oi_3_reg[0]  ( .D(\filter_0/n8847 ), .CP(clk), .Q(
        reg_oi_3[0]) );
  dff_sg \filter_0/i_pointer_reg[3]  ( .D(\filter_0/n8888 ), .CP(clk), .Q(
        \filter_0/i_pointer[3] ) );
  dff_sg \filter_0/i_pointer_reg[2]  ( .D(\filter_0/n8889 ), .CP(clk), .Q(
        \filter_0/i_pointer[2] ) );
  dff_sg \filter_0/i_pointer_reg[1]  ( .D(\filter_0/n8890 ), .CP(clk), .Q(
        \filter_0/i_pointer[1] ) );
  dff_sg \filter_0/i_pointer_reg[0]  ( .D(\filter_0/n8891 ), .CP(clk), .Q(
        \filter_0/i_pointer[0] ) );
  dff_sg \filter_0/m_pointer_reg[3]  ( .D(\filter_0/n8893 ), .CP(clk), .Q(
        \filter_0/N15 ) );
  dff_sg \filter_0/m_pointer_reg[2]  ( .D(\filter_0/n8894 ), .CP(clk), .Q(
        \filter_0/N14 ) );
  dff_sg \filter_0/m_pointer_reg[1]  ( .D(\filter_0/n8895 ), .CP(clk), .Q(
        \filter_0/N13 ) );
  dff_sg \filter_0/m_pointer_reg[0]  ( .D(\filter_0/n8896 ), .CP(clk), .Q(
        \filter_0/N12 ) );
  dff_sg \filter_0/m_pointer_reg[4]  ( .D(\filter_0/n8892 ), .CP(clk), .Q(
        \filter_0/N16 ) );
  dff_sg \filter_0/ow_8_reg[19]  ( .D(\filter_0/n8264 ), .CP(clk), .Q(
        reg_ow_8[19]) );
  dff_sg \filter_0/ow_8_reg[18]  ( .D(\filter_0/n8265 ), .CP(clk), .Q(
        reg_ow_8[18]) );
  dff_sg \filter_0/ow_8_reg[17]  ( .D(\filter_0/n8266 ), .CP(clk), .Q(
        reg_ow_8[17]) );
  dff_sg \filter_0/ow_8_reg[16]  ( .D(\filter_0/n8267 ), .CP(clk), .Q(
        reg_ow_8[16]) );
  dff_sg \filter_0/ow_8_reg[15]  ( .D(\filter_0/n8268 ), .CP(clk), .Q(
        reg_ow_8[15]) );
  dff_sg \filter_0/ow_8_reg[14]  ( .D(\filter_0/n8269 ), .CP(clk), .Q(
        reg_ow_8[14]) );
  dff_sg \filter_0/ow_8_reg[13]  ( .D(\filter_0/n8270 ), .CP(clk), .Q(
        reg_ow_8[13]) );
  dff_sg \filter_0/ow_8_reg[12]  ( .D(\filter_0/n8271 ), .CP(clk), .Q(
        reg_ow_8[12]) );
  dff_sg \filter_0/ow_8_reg[11]  ( .D(\filter_0/n8272 ), .CP(clk), .Q(
        reg_ow_8[11]) );
  dff_sg \filter_0/ow_8_reg[10]  ( .D(\filter_0/n8273 ), .CP(clk), .Q(
        reg_ow_8[10]) );
  dff_sg \filter_0/ow_8_reg[9]  ( .D(\filter_0/n8274 ), .CP(clk), .Q(
        reg_ow_8[9]) );
  dff_sg \filter_0/ow_8_reg[8]  ( .D(\filter_0/n8275 ), .CP(clk), .Q(
        reg_ow_8[8]) );
  dff_sg \filter_0/ow_8_reg[7]  ( .D(\filter_0/n8276 ), .CP(clk), .Q(
        reg_ow_8[7]) );
  dff_sg \filter_0/ow_8_reg[6]  ( .D(\filter_0/n8277 ), .CP(clk), .Q(
        reg_ow_8[6]) );
  dff_sg \filter_0/ow_8_reg[5]  ( .D(\filter_0/n8278 ), .CP(clk), .Q(
        reg_ow_8[5]) );
  dff_sg \filter_0/ow_8_reg[4]  ( .D(\filter_0/n8279 ), .CP(clk), .Q(
        reg_ow_8[4]) );
  dff_sg \filter_0/ow_8_reg[3]  ( .D(\filter_0/n8280 ), .CP(clk), .Q(
        reg_ow_8[3]) );
  dff_sg \filter_0/ow_8_reg[2]  ( .D(\filter_0/n8281 ), .CP(clk), .Q(
        reg_ow_8[2]) );
  dff_sg \filter_0/ow_8_reg[1]  ( .D(\filter_0/n8282 ), .CP(clk), .Q(
        reg_ow_8[1]) );
  dff_sg \filter_0/ow_8_reg[0]  ( .D(\filter_0/n8283 ), .CP(clk), .Q(
        reg_ow_8[0]) );
  dff_sg \filter_0/ow_9_reg[19]  ( .D(\filter_0/n8284 ), .CP(clk), .Q(
        reg_ow_9[19]) );
  dff_sg \filter_0/ow_9_reg[18]  ( .D(\filter_0/n8285 ), .CP(clk), .Q(
        reg_ow_9[18]) );
  dff_sg \filter_0/ow_9_reg[17]  ( .D(\filter_0/n8286 ), .CP(clk), .Q(
        reg_ow_9[17]) );
  dff_sg \filter_0/ow_9_reg[16]  ( .D(\filter_0/n8287 ), .CP(clk), .Q(
        reg_ow_9[16]) );
  dff_sg \filter_0/ow_9_reg[15]  ( .D(\filter_0/n8288 ), .CP(clk), .Q(
        reg_ow_9[15]) );
  dff_sg \filter_0/ow_9_reg[14]  ( .D(\filter_0/n8289 ), .CP(clk), .Q(
        reg_ow_9[14]) );
  dff_sg \filter_0/ow_9_reg[13]  ( .D(\filter_0/n8290 ), .CP(clk), .Q(
        reg_ow_9[13]) );
  dff_sg \filter_0/ow_9_reg[12]  ( .D(\filter_0/n8291 ), .CP(clk), .Q(
        reg_ow_9[12]) );
  dff_sg \filter_0/ow_9_reg[11]  ( .D(\filter_0/n8292 ), .CP(clk), .Q(
        reg_ow_9[11]) );
  dff_sg \filter_0/ow_9_reg[10]  ( .D(\filter_0/n8293 ), .CP(clk), .Q(
        reg_ow_9[10]) );
  dff_sg \filter_0/ow_9_reg[9]  ( .D(\filter_0/n8294 ), .CP(clk), .Q(
        reg_ow_9[9]) );
  dff_sg \filter_0/ow_9_reg[8]  ( .D(\filter_0/n8295 ), .CP(clk), .Q(
        reg_ow_9[8]) );
  dff_sg \filter_0/ow_9_reg[7]  ( .D(\filter_0/n8296 ), .CP(clk), .Q(
        reg_ow_9[7]) );
  dff_sg \filter_0/ow_9_reg[6]  ( .D(\filter_0/n8297 ), .CP(clk), .Q(
        reg_ow_9[6]) );
  dff_sg \filter_0/ow_9_reg[5]  ( .D(\filter_0/n8298 ), .CP(clk), .Q(
        reg_ow_9[5]) );
  dff_sg \filter_0/ow_9_reg[4]  ( .D(\filter_0/n8299 ), .CP(clk), .Q(
        reg_ow_9[4]) );
  dff_sg \filter_0/ow_9_reg[3]  ( .D(\filter_0/n8300 ), .CP(clk), .Q(
        reg_ow_9[3]) );
  dff_sg \filter_0/ow_9_reg[2]  ( .D(\filter_0/n8301 ), .CP(clk), .Q(
        reg_ow_9[2]) );
  dff_sg \filter_0/ow_9_reg[1]  ( .D(\filter_0/n8302 ), .CP(clk), .Q(
        reg_ow_9[1]) );
  dff_sg \filter_0/ow_9_reg[0]  ( .D(\filter_0/n8303 ), .CP(clk), .Q(
        reg_ow_9[0]) );
  dff_sg \filter_0/ow_10_reg[19]  ( .D(\filter_0/n8304 ), .CP(clk), .Q(
        reg_ow_10[19]) );
  dff_sg \filter_0/ow_10_reg[18]  ( .D(\filter_0/n8305 ), .CP(clk), .Q(
        reg_ow_10[18]) );
  dff_sg \filter_0/ow_10_reg[17]  ( .D(\filter_0/n8306 ), .CP(clk), .Q(
        reg_ow_10[17]) );
  dff_sg \filter_0/ow_10_reg[16]  ( .D(\filter_0/n8307 ), .CP(clk), .Q(
        reg_ow_10[16]) );
  dff_sg \filter_0/ow_10_reg[15]  ( .D(\filter_0/n8308 ), .CP(clk), .Q(
        reg_ow_10[15]) );
  dff_sg \filter_0/ow_10_reg[14]  ( .D(\filter_0/n8309 ), .CP(clk), .Q(
        reg_ow_10[14]) );
  dff_sg \filter_0/ow_10_reg[13]  ( .D(\filter_0/n8310 ), .CP(clk), .Q(
        reg_ow_10[13]) );
  dff_sg \filter_0/ow_10_reg[12]  ( .D(\filter_0/n8311 ), .CP(clk), .Q(
        reg_ow_10[12]) );
  dff_sg \filter_0/ow_10_reg[11]  ( .D(\filter_0/n8312 ), .CP(clk), .Q(
        reg_ow_10[11]) );
  dff_sg \filter_0/ow_10_reg[10]  ( .D(\filter_0/n8313 ), .CP(clk), .Q(
        reg_ow_10[10]) );
  dff_sg \filter_0/ow_10_reg[9]  ( .D(\filter_0/n8314 ), .CP(clk), .Q(
        reg_ow_10[9]) );
  dff_sg \filter_0/ow_10_reg[8]  ( .D(\filter_0/n8315 ), .CP(clk), .Q(
        reg_ow_10[8]) );
  dff_sg \filter_0/ow_10_reg[7]  ( .D(\filter_0/n8316 ), .CP(clk), .Q(
        reg_ow_10[7]) );
  dff_sg \filter_0/ow_10_reg[6]  ( .D(\filter_0/n8317 ), .CP(clk), .Q(
        reg_ow_10[6]) );
  dff_sg \filter_0/ow_10_reg[5]  ( .D(\filter_0/n8318 ), .CP(clk), .Q(
        reg_ow_10[5]) );
  dff_sg \filter_0/ow_10_reg[4]  ( .D(\filter_0/n8319 ), .CP(clk), .Q(
        reg_ow_10[4]) );
  dff_sg \filter_0/ow_10_reg[3]  ( .D(\filter_0/n8320 ), .CP(clk), .Q(
        reg_ow_10[3]) );
  dff_sg \filter_0/ow_10_reg[2]  ( .D(\filter_0/n8321 ), .CP(clk), .Q(
        reg_ow_10[2]) );
  dff_sg \filter_0/ow_10_reg[1]  ( .D(\filter_0/n8322 ), .CP(clk), .Q(
        reg_ow_10[1]) );
  dff_sg \filter_0/ow_10_reg[0]  ( .D(\filter_0/n8323 ), .CP(clk), .Q(
        reg_ow_10[0]) );
  dff_sg \filter_0/ow_11_reg[19]  ( .D(\filter_0/n8324 ), .CP(clk), .Q(
        reg_ow_11[19]) );
  dff_sg \filter_0/ow_11_reg[18]  ( .D(\filter_0/n8325 ), .CP(clk), .Q(
        reg_ow_11[18]) );
  dff_sg \filter_0/ow_11_reg[17]  ( .D(\filter_0/n8326 ), .CP(clk), .Q(
        reg_ow_11[17]) );
  dff_sg \filter_0/ow_11_reg[16]  ( .D(\filter_0/n8327 ), .CP(clk), .Q(
        reg_ow_11[16]) );
  dff_sg \filter_0/ow_11_reg[15]  ( .D(\filter_0/n8328 ), .CP(clk), .Q(
        reg_ow_11[15]) );
  dff_sg \filter_0/ow_11_reg[14]  ( .D(\filter_0/n8329 ), .CP(clk), .Q(
        reg_ow_11[14]) );
  dff_sg \filter_0/ow_11_reg[13]  ( .D(\filter_0/n8330 ), .CP(clk), .Q(
        reg_ow_11[13]) );
  dff_sg \filter_0/ow_11_reg[12]  ( .D(\filter_0/n8331 ), .CP(clk), .Q(
        reg_ow_11[12]) );
  dff_sg \filter_0/ow_11_reg[11]  ( .D(\filter_0/n8332 ), .CP(clk), .Q(
        reg_ow_11[11]) );
  dff_sg \filter_0/ow_11_reg[10]  ( .D(\filter_0/n8333 ), .CP(clk), .Q(
        reg_ow_11[10]) );
  dff_sg \filter_0/ow_11_reg[9]  ( .D(\filter_0/n8334 ), .CP(clk), .Q(
        reg_ow_11[9]) );
  dff_sg \filter_0/ow_11_reg[8]  ( .D(\filter_0/n8335 ), .CP(clk), .Q(
        reg_ow_11[8]) );
  dff_sg \filter_0/ow_11_reg[7]  ( .D(\filter_0/n8336 ), .CP(clk), .Q(
        reg_ow_11[7]) );
  dff_sg \filter_0/ow_11_reg[6]  ( .D(\filter_0/n8337 ), .CP(clk), .Q(
        reg_ow_11[6]) );
  dff_sg \filter_0/ow_11_reg[5]  ( .D(\filter_0/n8338 ), .CP(clk), .Q(
        reg_ow_11[5]) );
  dff_sg \filter_0/ow_11_reg[4]  ( .D(\filter_0/n8339 ), .CP(clk), .Q(
        reg_ow_11[4]) );
  dff_sg \filter_0/ow_11_reg[3]  ( .D(\filter_0/n8340 ), .CP(clk), .Q(
        reg_ow_11[3]) );
  dff_sg \filter_0/ow_11_reg[2]  ( .D(\filter_0/n8341 ), .CP(clk), .Q(
        reg_ow_11[2]) );
  dff_sg \filter_0/ow_11_reg[1]  ( .D(\filter_0/n8342 ), .CP(clk), .Q(
        reg_ow_11[1]) );
  dff_sg \filter_0/ow_11_reg[0]  ( .D(\filter_0/n8343 ), .CP(clk), .Q(
        reg_ow_11[0]) );
  dff_sg \filter_0/ow_15_reg[19]  ( .D(\filter_0/n8404 ), .CP(clk), .Q(
        reg_ow_15[19]) );
  dff_sg \filter_0/ow_15_reg[18]  ( .D(\filter_0/n8405 ), .CP(clk), .Q(
        reg_ow_15[18]) );
  dff_sg \filter_0/ow_15_reg[17]  ( .D(\filter_0/n8406 ), .CP(clk), .Q(
        reg_ow_15[17]) );
  dff_sg \filter_0/ow_15_reg[16]  ( .D(\filter_0/n8407 ), .CP(clk), .Q(
        reg_ow_15[16]) );
  dff_sg \filter_0/ow_15_reg[15]  ( .D(\filter_0/n8408 ), .CP(clk), .Q(
        reg_ow_15[15]) );
  dff_sg \filter_0/ow_15_reg[14]  ( .D(\filter_0/n8409 ), .CP(clk), .Q(
        reg_ow_15[14]) );
  dff_sg \filter_0/ow_15_reg[13]  ( .D(\filter_0/n8410 ), .CP(clk), .Q(
        reg_ow_15[13]) );
  dff_sg \filter_0/ow_15_reg[12]  ( .D(\filter_0/n8411 ), .CP(clk), .Q(
        reg_ow_15[12]) );
  dff_sg \filter_0/ow_15_reg[11]  ( .D(\filter_0/n8412 ), .CP(clk), .Q(
        reg_ow_15[11]) );
  dff_sg \filter_0/ow_15_reg[10]  ( .D(\filter_0/n8413 ), .CP(clk), .Q(
        reg_ow_15[10]) );
  dff_sg \filter_0/ow_15_reg[9]  ( .D(\filter_0/n8414 ), .CP(clk), .Q(
        reg_ow_15[9]) );
  dff_sg \filter_0/ow_15_reg[8]  ( .D(\filter_0/n8415 ), .CP(clk), .Q(
        reg_ow_15[8]) );
  dff_sg \filter_0/ow_15_reg[7]  ( .D(\filter_0/n8416 ), .CP(clk), .Q(
        reg_ow_15[7]) );
  dff_sg \filter_0/ow_15_reg[6]  ( .D(\filter_0/n8417 ), .CP(clk), .Q(
        reg_ow_15[6]) );
  dff_sg \filter_0/ow_15_reg[5]  ( .D(\filter_0/n8418 ), .CP(clk), .Q(
        reg_ow_15[5]) );
  dff_sg \filter_0/ow_15_reg[4]  ( .D(\filter_0/n8419 ), .CP(clk), .Q(
        reg_ow_15[4]) );
  dff_sg \filter_0/ow_15_reg[3]  ( .D(\filter_0/n8420 ), .CP(clk), .Q(
        reg_ow_15[3]) );
  dff_sg \filter_0/ow_15_reg[2]  ( .D(\filter_0/n8421 ), .CP(clk), .Q(
        reg_ow_15[2]) );
  dff_sg \filter_0/ow_15_reg[1]  ( .D(\filter_0/n8422 ), .CP(clk), .Q(
        reg_ow_15[1]) );
  dff_sg \filter_0/ow_15_reg[0]  ( .D(\filter_0/n8423 ), .CP(clk), .Q(
        reg_ow_15[0]) );
  dff_sg \filter_0/ow_12_reg[19]  ( .D(\filter_0/n8344 ), .CP(clk), .Q(
        reg_ow_12[19]) );
  dff_sg \filter_0/ow_12_reg[18]  ( .D(\filter_0/n8345 ), .CP(clk), .Q(
        reg_ow_12[18]) );
  dff_sg \filter_0/ow_12_reg[17]  ( .D(\filter_0/n8346 ), .CP(clk), .Q(
        reg_ow_12[17]) );
  dff_sg \filter_0/ow_12_reg[16]  ( .D(\filter_0/n8347 ), .CP(clk), .Q(
        reg_ow_12[16]) );
  dff_sg \filter_0/ow_12_reg[15]  ( .D(\filter_0/n8348 ), .CP(clk), .Q(
        reg_ow_12[15]) );
  dff_sg \filter_0/ow_12_reg[14]  ( .D(\filter_0/n8349 ), .CP(clk), .Q(
        reg_ow_12[14]) );
  dff_sg \filter_0/ow_12_reg[13]  ( .D(\filter_0/n8350 ), .CP(clk), .Q(
        reg_ow_12[13]) );
  dff_sg \filter_0/ow_12_reg[12]  ( .D(\filter_0/n8351 ), .CP(clk), .Q(
        reg_ow_12[12]) );
  dff_sg \filter_0/ow_12_reg[11]  ( .D(\filter_0/n8352 ), .CP(clk), .Q(
        reg_ow_12[11]) );
  dff_sg \filter_0/ow_12_reg[10]  ( .D(\filter_0/n8353 ), .CP(clk), .Q(
        reg_ow_12[10]) );
  dff_sg \filter_0/ow_12_reg[9]  ( .D(\filter_0/n8354 ), .CP(clk), .Q(
        reg_ow_12[9]) );
  dff_sg \filter_0/ow_12_reg[8]  ( .D(\filter_0/n8355 ), .CP(clk), .Q(
        reg_ow_12[8]) );
  dff_sg \filter_0/ow_12_reg[7]  ( .D(\filter_0/n8356 ), .CP(clk), .Q(
        reg_ow_12[7]) );
  dff_sg \filter_0/ow_12_reg[6]  ( .D(\filter_0/n8357 ), .CP(clk), .Q(
        reg_ow_12[6]) );
  dff_sg \filter_0/ow_12_reg[5]  ( .D(\filter_0/n8358 ), .CP(clk), .Q(
        reg_ow_12[5]) );
  dff_sg \filter_0/ow_12_reg[4]  ( .D(\filter_0/n8359 ), .CP(clk), .Q(
        reg_ow_12[4]) );
  dff_sg \filter_0/ow_12_reg[3]  ( .D(\filter_0/n8360 ), .CP(clk), .Q(
        reg_ow_12[3]) );
  dff_sg \filter_0/ow_12_reg[2]  ( .D(\filter_0/n8361 ), .CP(clk), .Q(
        reg_ow_12[2]) );
  dff_sg \filter_0/ow_12_reg[1]  ( .D(\filter_0/n8362 ), .CP(clk), .Q(
        reg_ow_12[1]) );
  dff_sg \filter_0/ow_12_reg[0]  ( .D(\filter_0/n8363 ), .CP(clk), .Q(
        reg_ow_12[0]) );
  dff_sg \filter_0/ow_13_reg[19]  ( .D(\filter_0/n8364 ), .CP(clk), .Q(
        reg_ow_13[19]) );
  dff_sg \filter_0/ow_13_reg[18]  ( .D(\filter_0/n8365 ), .CP(clk), .Q(
        reg_ow_13[18]) );
  dff_sg \filter_0/ow_13_reg[17]  ( .D(\filter_0/n8366 ), .CP(clk), .Q(
        reg_ow_13[17]) );
  dff_sg \filter_0/ow_13_reg[16]  ( .D(\filter_0/n8367 ), .CP(clk), .Q(
        reg_ow_13[16]) );
  dff_sg \filter_0/ow_13_reg[15]  ( .D(\filter_0/n8368 ), .CP(clk), .Q(
        reg_ow_13[15]) );
  dff_sg \filter_0/ow_13_reg[14]  ( .D(\filter_0/n8369 ), .CP(clk), .Q(
        reg_ow_13[14]) );
  dff_sg \filter_0/ow_13_reg[13]  ( .D(\filter_0/n8370 ), .CP(clk), .Q(
        reg_ow_13[13]) );
  dff_sg \filter_0/ow_13_reg[12]  ( .D(\filter_0/n8371 ), .CP(clk), .Q(
        reg_ow_13[12]) );
  dff_sg \filter_0/ow_13_reg[11]  ( .D(\filter_0/n8372 ), .CP(clk), .Q(
        reg_ow_13[11]) );
  dff_sg \filter_0/ow_13_reg[10]  ( .D(\filter_0/n8373 ), .CP(clk), .Q(
        reg_ow_13[10]) );
  dff_sg \filter_0/ow_13_reg[9]  ( .D(\filter_0/n8374 ), .CP(clk), .Q(
        reg_ow_13[9]) );
  dff_sg \filter_0/ow_13_reg[8]  ( .D(\filter_0/n8375 ), .CP(clk), .Q(
        reg_ow_13[8]) );
  dff_sg \filter_0/ow_13_reg[7]  ( .D(\filter_0/n8376 ), .CP(clk), .Q(
        reg_ow_13[7]) );
  dff_sg \filter_0/ow_13_reg[6]  ( .D(\filter_0/n8377 ), .CP(clk), .Q(
        reg_ow_13[6]) );
  dff_sg \filter_0/ow_13_reg[5]  ( .D(\filter_0/n8378 ), .CP(clk), .Q(
        reg_ow_13[5]) );
  dff_sg \filter_0/ow_13_reg[4]  ( .D(\filter_0/n8379 ), .CP(clk), .Q(
        reg_ow_13[4]) );
  dff_sg \filter_0/ow_13_reg[3]  ( .D(\filter_0/n8380 ), .CP(clk), .Q(
        reg_ow_13[3]) );
  dff_sg \filter_0/ow_13_reg[2]  ( .D(\filter_0/n8381 ), .CP(clk), .Q(
        reg_ow_13[2]) );
  dff_sg \filter_0/ow_13_reg[1]  ( .D(\filter_0/n8382 ), .CP(clk), .Q(
        reg_ow_13[1]) );
  dff_sg \filter_0/ow_13_reg[0]  ( .D(\filter_0/n8383 ), .CP(clk), .Q(
        reg_ow_13[0]) );
  dff_sg \filter_0/ow_14_reg[19]  ( .D(\filter_0/n8384 ), .CP(clk), .Q(
        reg_ow_14[19]) );
  dff_sg \filter_0/ow_14_reg[18]  ( .D(\filter_0/n8385 ), .CP(clk), .Q(
        reg_ow_14[18]) );
  dff_sg \filter_0/ow_14_reg[17]  ( .D(\filter_0/n8386 ), .CP(clk), .Q(
        reg_ow_14[17]) );
  dff_sg \filter_0/ow_14_reg[16]  ( .D(\filter_0/n8387 ), .CP(clk), .Q(
        reg_ow_14[16]) );
  dff_sg \filter_0/ow_14_reg[15]  ( .D(\filter_0/n8388 ), .CP(clk), .Q(
        reg_ow_14[15]) );
  dff_sg \filter_0/ow_14_reg[14]  ( .D(\filter_0/n8389 ), .CP(clk), .Q(
        reg_ow_14[14]) );
  dff_sg \filter_0/ow_14_reg[13]  ( .D(\filter_0/n8390 ), .CP(clk), .Q(
        reg_ow_14[13]) );
  dff_sg \filter_0/ow_14_reg[12]  ( .D(\filter_0/n8391 ), .CP(clk), .Q(
        reg_ow_14[12]) );
  dff_sg \filter_0/ow_14_reg[11]  ( .D(\filter_0/n8392 ), .CP(clk), .Q(
        reg_ow_14[11]) );
  dff_sg \filter_0/ow_14_reg[10]  ( .D(\filter_0/n8393 ), .CP(clk), .Q(
        reg_ow_14[10]) );
  dff_sg \filter_0/ow_14_reg[9]  ( .D(\filter_0/n8394 ), .CP(clk), .Q(
        reg_ow_14[9]) );
  dff_sg \filter_0/ow_14_reg[8]  ( .D(\filter_0/n8395 ), .CP(clk), .Q(
        reg_ow_14[8]) );
  dff_sg \filter_0/ow_14_reg[7]  ( .D(\filter_0/n8396 ), .CP(clk), .Q(
        reg_ow_14[7]) );
  dff_sg \filter_0/ow_14_reg[6]  ( .D(\filter_0/n8397 ), .CP(clk), .Q(
        reg_ow_14[6]) );
  dff_sg \filter_0/ow_14_reg[5]  ( .D(\filter_0/n8398 ), .CP(clk), .Q(
        reg_ow_14[5]) );
  dff_sg \filter_0/ow_14_reg[4]  ( .D(\filter_0/n8399 ), .CP(clk), .Q(
        reg_ow_14[4]) );
  dff_sg \filter_0/ow_14_reg[3]  ( .D(\filter_0/n8400 ), .CP(clk), .Q(
        reg_ow_14[3]) );
  dff_sg \filter_0/ow_14_reg[2]  ( .D(\filter_0/n8401 ), .CP(clk), .Q(
        reg_ow_14[2]) );
  dff_sg \filter_0/ow_14_reg[1]  ( .D(\filter_0/n8402 ), .CP(clk), .Q(
        reg_ow_14[1]) );
  dff_sg \filter_0/ow_14_reg[0]  ( .D(\filter_0/n8403 ), .CP(clk), .Q(
        reg_ow_14[0]) );
  dff_sg \filter_0/ow_4_reg[19]  ( .D(\filter_0/n8484 ), .CP(clk), .Q(
        reg_ow_4[19]) );
  dff_sg \filter_0/ow_4_reg[18]  ( .D(\filter_0/n8485 ), .CP(clk), .Q(
        reg_ow_4[18]) );
  dff_sg \filter_0/ow_4_reg[17]  ( .D(\filter_0/n8486 ), .CP(clk), .Q(
        reg_ow_4[17]) );
  dff_sg \filter_0/ow_4_reg[16]  ( .D(\filter_0/n8487 ), .CP(clk), .Q(
        reg_ow_4[16]) );
  dff_sg \filter_0/ow_4_reg[15]  ( .D(\filter_0/n8488 ), .CP(clk), .Q(
        reg_ow_4[15]) );
  dff_sg \filter_0/ow_4_reg[14]  ( .D(\filter_0/n8489 ), .CP(clk), .Q(
        reg_ow_4[14]) );
  dff_sg \filter_0/ow_4_reg[13]  ( .D(\filter_0/n8490 ), .CP(clk), .Q(
        reg_ow_4[13]) );
  dff_sg \filter_0/ow_4_reg[12]  ( .D(\filter_0/n8491 ), .CP(clk), .Q(
        reg_ow_4[12]) );
  dff_sg \filter_0/ow_4_reg[11]  ( .D(\filter_0/n8492 ), .CP(clk), .Q(
        reg_ow_4[11]) );
  dff_sg \filter_0/ow_4_reg[10]  ( .D(\filter_0/n8493 ), .CP(clk), .Q(
        reg_ow_4[10]) );
  dff_sg \filter_0/ow_4_reg[9]  ( .D(\filter_0/n8494 ), .CP(clk), .Q(
        reg_ow_4[9]) );
  dff_sg \filter_0/ow_4_reg[8]  ( .D(\filter_0/n8495 ), .CP(clk), .Q(
        reg_ow_4[8]) );
  dff_sg \filter_0/ow_4_reg[7]  ( .D(\filter_0/n8496 ), .CP(clk), .Q(
        reg_ow_4[7]) );
  dff_sg \filter_0/ow_4_reg[6]  ( .D(\filter_0/n8497 ), .CP(clk), .Q(
        reg_ow_4[6]) );
  dff_sg \filter_0/ow_4_reg[5]  ( .D(\filter_0/n8498 ), .CP(clk), .Q(
        reg_ow_4[5]) );
  dff_sg \filter_0/ow_4_reg[4]  ( .D(\filter_0/n8499 ), .CP(clk), .Q(
        reg_ow_4[4]) );
  dff_sg \filter_0/ow_4_reg[3]  ( .D(\filter_0/n8500 ), .CP(clk), .Q(
        reg_ow_4[3]) );
  dff_sg \filter_0/ow_4_reg[2]  ( .D(\filter_0/n8501 ), .CP(clk), .Q(
        reg_ow_4[2]) );
  dff_sg \filter_0/ow_4_reg[1]  ( .D(\filter_0/n8502 ), .CP(clk), .Q(
        reg_ow_4[1]) );
  dff_sg \filter_0/ow_4_reg[0]  ( .D(\filter_0/n8503 ), .CP(clk), .Q(
        reg_ow_4[0]) );
  dff_sg \filter_0/ow_5_reg[19]  ( .D(\filter_0/n8464 ), .CP(clk), .Q(
        reg_ow_5[19]) );
  dff_sg \filter_0/ow_5_reg[18]  ( .D(\filter_0/n8465 ), .CP(clk), .Q(
        reg_ow_5[18]) );
  dff_sg \filter_0/ow_5_reg[17]  ( .D(\filter_0/n8466 ), .CP(clk), .Q(
        reg_ow_5[17]) );
  dff_sg \filter_0/ow_5_reg[16]  ( .D(\filter_0/n8467 ), .CP(clk), .Q(
        reg_ow_5[16]) );
  dff_sg \filter_0/ow_5_reg[15]  ( .D(\filter_0/n8468 ), .CP(clk), .Q(
        reg_ow_5[15]) );
  dff_sg \filter_0/ow_5_reg[14]  ( .D(\filter_0/n8469 ), .CP(clk), .Q(
        reg_ow_5[14]) );
  dff_sg \filter_0/ow_5_reg[13]  ( .D(\filter_0/n8470 ), .CP(clk), .Q(
        reg_ow_5[13]) );
  dff_sg \filter_0/ow_5_reg[12]  ( .D(\filter_0/n8471 ), .CP(clk), .Q(
        reg_ow_5[12]) );
  dff_sg \filter_0/ow_5_reg[11]  ( .D(\filter_0/n8472 ), .CP(clk), .Q(
        reg_ow_5[11]) );
  dff_sg \filter_0/ow_5_reg[10]  ( .D(\filter_0/n8473 ), .CP(clk), .Q(
        reg_ow_5[10]) );
  dff_sg \filter_0/ow_5_reg[9]  ( .D(\filter_0/n8474 ), .CP(clk), .Q(
        reg_ow_5[9]) );
  dff_sg \filter_0/ow_5_reg[8]  ( .D(\filter_0/n8475 ), .CP(clk), .Q(
        reg_ow_5[8]) );
  dff_sg \filter_0/ow_5_reg[7]  ( .D(\filter_0/n8476 ), .CP(clk), .Q(
        reg_ow_5[7]) );
  dff_sg \filter_0/ow_5_reg[6]  ( .D(\filter_0/n8477 ), .CP(clk), .Q(
        reg_ow_5[6]) );
  dff_sg \filter_0/ow_5_reg[5]  ( .D(\filter_0/n8478 ), .CP(clk), .Q(
        reg_ow_5[5]) );
  dff_sg \filter_0/ow_5_reg[4]  ( .D(\filter_0/n8479 ), .CP(clk), .Q(
        reg_ow_5[4]) );
  dff_sg \filter_0/ow_5_reg[3]  ( .D(\filter_0/n8480 ), .CP(clk), .Q(
        reg_ow_5[3]) );
  dff_sg \filter_0/ow_5_reg[2]  ( .D(\filter_0/n8481 ), .CP(clk), .Q(
        reg_ow_5[2]) );
  dff_sg \filter_0/ow_5_reg[1]  ( .D(\filter_0/n8482 ), .CP(clk), .Q(
        reg_ow_5[1]) );
  dff_sg \filter_0/ow_5_reg[0]  ( .D(\filter_0/n8483 ), .CP(clk), .Q(
        reg_ow_5[0]) );
  dff_sg \filter_0/ow_6_reg[19]  ( .D(\filter_0/n8444 ), .CP(clk), .Q(
        reg_ow_6[19]) );
  dff_sg \filter_0/ow_6_reg[18]  ( .D(\filter_0/n8445 ), .CP(clk), .Q(
        reg_ow_6[18]) );
  dff_sg \filter_0/ow_6_reg[17]  ( .D(\filter_0/n8446 ), .CP(clk), .Q(
        reg_ow_6[17]) );
  dff_sg \filter_0/ow_6_reg[16]  ( .D(\filter_0/n8447 ), .CP(clk), .Q(
        reg_ow_6[16]) );
  dff_sg \filter_0/ow_6_reg[15]  ( .D(\filter_0/n8448 ), .CP(clk), .Q(
        reg_ow_6[15]) );
  dff_sg \filter_0/ow_6_reg[14]  ( .D(\filter_0/n8449 ), .CP(clk), .Q(
        reg_ow_6[14]) );
  dff_sg \filter_0/ow_6_reg[13]  ( .D(\filter_0/n8450 ), .CP(clk), .Q(
        reg_ow_6[13]) );
  dff_sg \filter_0/ow_6_reg[12]  ( .D(\filter_0/n8451 ), .CP(clk), .Q(
        reg_ow_6[12]) );
  dff_sg \filter_0/ow_6_reg[11]  ( .D(\filter_0/n8452 ), .CP(clk), .Q(
        reg_ow_6[11]) );
  dff_sg \filter_0/ow_6_reg[10]  ( .D(\filter_0/n8453 ), .CP(clk), .Q(
        reg_ow_6[10]) );
  dff_sg \filter_0/ow_6_reg[9]  ( .D(\filter_0/n8454 ), .CP(clk), .Q(
        reg_ow_6[9]) );
  dff_sg \filter_0/ow_6_reg[8]  ( .D(\filter_0/n8455 ), .CP(clk), .Q(
        reg_ow_6[8]) );
  dff_sg \filter_0/ow_6_reg[7]  ( .D(\filter_0/n8456 ), .CP(clk), .Q(
        reg_ow_6[7]) );
  dff_sg \filter_0/ow_6_reg[6]  ( .D(\filter_0/n8457 ), .CP(clk), .Q(
        reg_ow_6[6]) );
  dff_sg \filter_0/ow_6_reg[5]  ( .D(\filter_0/n8458 ), .CP(clk), .Q(
        reg_ow_6[5]) );
  dff_sg \filter_0/ow_6_reg[4]  ( .D(\filter_0/n8459 ), .CP(clk), .Q(
        reg_ow_6[4]) );
  dff_sg \filter_0/ow_6_reg[3]  ( .D(\filter_0/n8460 ), .CP(clk), .Q(
        reg_ow_6[3]) );
  dff_sg \filter_0/ow_6_reg[2]  ( .D(\filter_0/n8461 ), .CP(clk), .Q(
        reg_ow_6[2]) );
  dff_sg \filter_0/ow_6_reg[1]  ( .D(\filter_0/n8462 ), .CP(clk), .Q(
        reg_ow_6[1]) );
  dff_sg \filter_0/ow_6_reg[0]  ( .D(\filter_0/n8463 ), .CP(clk), .Q(
        reg_ow_6[0]) );
  dff_sg \filter_0/ow_7_reg[19]  ( .D(\filter_0/n8424 ), .CP(clk), .Q(
        reg_ow_7[19]) );
  dff_sg \filter_0/ow_7_reg[18]  ( .D(\filter_0/n8425 ), .CP(clk), .Q(
        reg_ow_7[18]) );
  dff_sg \filter_0/ow_7_reg[17]  ( .D(\filter_0/n8426 ), .CP(clk), .Q(
        reg_ow_7[17]) );
  dff_sg \filter_0/ow_7_reg[16]  ( .D(\filter_0/n8427 ), .CP(clk), .Q(
        reg_ow_7[16]) );
  dff_sg \filter_0/ow_7_reg[15]  ( .D(\filter_0/n8428 ), .CP(clk), .Q(
        reg_ow_7[15]) );
  dff_sg \filter_0/ow_7_reg[14]  ( .D(\filter_0/n8429 ), .CP(clk), .Q(
        reg_ow_7[14]) );
  dff_sg \filter_0/ow_7_reg[13]  ( .D(\filter_0/n8430 ), .CP(clk), .Q(
        reg_ow_7[13]) );
  dff_sg \filter_0/ow_7_reg[12]  ( .D(\filter_0/n8431 ), .CP(clk), .Q(
        reg_ow_7[12]) );
  dff_sg \filter_0/ow_7_reg[11]  ( .D(\filter_0/n8432 ), .CP(clk), .Q(
        reg_ow_7[11]) );
  dff_sg \filter_0/ow_7_reg[10]  ( .D(\filter_0/n8433 ), .CP(clk), .Q(
        reg_ow_7[10]) );
  dff_sg \filter_0/ow_7_reg[9]  ( .D(\filter_0/n8434 ), .CP(clk), .Q(
        reg_ow_7[9]) );
  dff_sg \filter_0/ow_7_reg[8]  ( .D(\filter_0/n8435 ), .CP(clk), .Q(
        reg_ow_7[8]) );
  dff_sg \filter_0/ow_7_reg[7]  ( .D(\filter_0/n8436 ), .CP(clk), .Q(
        reg_ow_7[7]) );
  dff_sg \filter_0/ow_7_reg[6]  ( .D(\filter_0/n8437 ), .CP(clk), .Q(
        reg_ow_7[6]) );
  dff_sg \filter_0/ow_7_reg[5]  ( .D(\filter_0/n8438 ), .CP(clk), .Q(
        reg_ow_7[5]) );
  dff_sg \filter_0/ow_7_reg[4]  ( .D(\filter_0/n8439 ), .CP(clk), .Q(
        reg_ow_7[4]) );
  dff_sg \filter_0/ow_7_reg[3]  ( .D(\filter_0/n8440 ), .CP(clk), .Q(
        reg_ow_7[3]) );
  dff_sg \filter_0/ow_7_reg[2]  ( .D(\filter_0/n8441 ), .CP(clk), .Q(
        reg_ow_7[2]) );
  dff_sg \filter_0/ow_7_reg[1]  ( .D(\filter_0/n8442 ), .CP(clk), .Q(
        reg_ow_7[1]) );
  dff_sg \filter_0/ow_7_reg[0]  ( .D(\filter_0/n8443 ), .CP(clk), .Q(
        reg_ow_7[0]) );
  dff_sg \filter_0/ow_0_reg[19]  ( .D(\filter_0/n8244 ), .CP(clk), .Q(
        reg_ow_0[19]) );
  dff_sg \filter_0/ow_0_reg[18]  ( .D(\filter_0/n8245 ), .CP(clk), .Q(
        reg_ow_0[18]) );
  dff_sg \filter_0/ow_0_reg[17]  ( .D(\filter_0/n8246 ), .CP(clk), .Q(
        reg_ow_0[17]) );
  dff_sg \filter_0/ow_0_reg[16]  ( .D(\filter_0/n8247 ), .CP(clk), .Q(
        reg_ow_0[16]) );
  dff_sg \filter_0/ow_0_reg[15]  ( .D(\filter_0/n8248 ), .CP(clk), .Q(
        reg_ow_0[15]) );
  dff_sg \filter_0/ow_0_reg[14]  ( .D(\filter_0/n8249 ), .CP(clk), .Q(
        reg_ow_0[14]) );
  dff_sg \filter_0/ow_0_reg[13]  ( .D(\filter_0/n8250 ), .CP(clk), .Q(
        reg_ow_0[13]) );
  dff_sg \filter_0/ow_0_reg[12]  ( .D(\filter_0/n8251 ), .CP(clk), .Q(
        reg_ow_0[12]) );
  dff_sg \filter_0/ow_0_reg[11]  ( .D(\filter_0/n8252 ), .CP(clk), .Q(
        reg_ow_0[11]) );
  dff_sg \filter_0/ow_0_reg[10]  ( .D(\filter_0/n8253 ), .CP(clk), .Q(
        reg_ow_0[10]) );
  dff_sg \filter_0/ow_0_reg[9]  ( .D(\filter_0/n8254 ), .CP(clk), .Q(
        reg_ow_0[9]) );
  dff_sg \filter_0/ow_0_reg[8]  ( .D(\filter_0/n8255 ), .CP(clk), .Q(
        reg_ow_0[8]) );
  dff_sg \filter_0/ow_0_reg[7]  ( .D(\filter_0/n8256 ), .CP(clk), .Q(
        reg_ow_0[7]) );
  dff_sg \filter_0/ow_0_reg[6]  ( .D(\filter_0/n8257 ), .CP(clk), .Q(
        reg_ow_0[6]) );
  dff_sg \filter_0/ow_0_reg[5]  ( .D(\filter_0/n8258 ), .CP(clk), .Q(
        reg_ow_0[5]) );
  dff_sg \filter_0/ow_0_reg[4]  ( .D(\filter_0/n8259 ), .CP(clk), .Q(
        reg_ow_0[4]) );
  dff_sg \filter_0/ow_0_reg[3]  ( .D(\filter_0/n8260 ), .CP(clk), .Q(
        reg_ow_0[3]) );
  dff_sg \filter_0/ow_0_reg[2]  ( .D(\filter_0/n8261 ), .CP(clk), .Q(
        reg_ow_0[2]) );
  dff_sg \filter_0/ow_0_reg[1]  ( .D(\filter_0/n8262 ), .CP(clk), .Q(
        reg_ow_0[1]) );
  dff_sg \filter_0/ow_0_reg[0]  ( .D(\filter_0/n8263 ), .CP(clk), .Q(
        reg_ow_0[0]) );
  dff_sg \filter_0/ow_1_reg[19]  ( .D(\filter_0/n8544 ), .CP(clk), .Q(
        reg_ow_1[19]) );
  dff_sg \filter_0/ow_1_reg[18]  ( .D(\filter_0/n8545 ), .CP(clk), .Q(
        reg_ow_1[18]) );
  dff_sg \filter_0/ow_1_reg[17]  ( .D(\filter_0/n8546 ), .CP(clk), .Q(
        reg_ow_1[17]) );
  dff_sg \filter_0/ow_1_reg[16]  ( .D(\filter_0/n8547 ), .CP(clk), .Q(
        reg_ow_1[16]) );
  dff_sg \filter_0/ow_1_reg[15]  ( .D(\filter_0/n8548 ), .CP(clk), .Q(
        reg_ow_1[15]) );
  dff_sg \filter_0/ow_1_reg[14]  ( .D(\filter_0/n8549 ), .CP(clk), .Q(
        reg_ow_1[14]) );
  dff_sg \filter_0/ow_1_reg[13]  ( .D(\filter_0/n8550 ), .CP(clk), .Q(
        reg_ow_1[13]) );
  dff_sg \filter_0/ow_1_reg[12]  ( .D(\filter_0/n8551 ), .CP(clk), .Q(
        reg_ow_1[12]) );
  dff_sg \filter_0/ow_1_reg[11]  ( .D(\filter_0/n8552 ), .CP(clk), .Q(
        reg_ow_1[11]) );
  dff_sg \filter_0/ow_1_reg[10]  ( .D(\filter_0/n8553 ), .CP(clk), .Q(
        reg_ow_1[10]) );
  dff_sg \filter_0/ow_1_reg[9]  ( .D(\filter_0/n8554 ), .CP(clk), .Q(
        reg_ow_1[9]) );
  dff_sg \filter_0/ow_1_reg[8]  ( .D(\filter_0/n8555 ), .CP(clk), .Q(
        reg_ow_1[8]) );
  dff_sg \filter_0/ow_1_reg[7]  ( .D(\filter_0/n8556 ), .CP(clk), .Q(
        reg_ow_1[7]) );
  dff_sg \filter_0/ow_1_reg[6]  ( .D(\filter_0/n8557 ), .CP(clk), .Q(
        reg_ow_1[6]) );
  dff_sg \filter_0/ow_1_reg[5]  ( .D(\filter_0/n8558 ), .CP(clk), .Q(
        reg_ow_1[5]) );
  dff_sg \filter_0/ow_1_reg[4]  ( .D(\filter_0/n8559 ), .CP(clk), .Q(
        reg_ow_1[4]) );
  dff_sg \filter_0/ow_1_reg[3]  ( .D(\filter_0/n8560 ), .CP(clk), .Q(
        reg_ow_1[3]) );
  dff_sg \filter_0/ow_1_reg[2]  ( .D(\filter_0/n8561 ), .CP(clk), .Q(
        reg_ow_1[2]) );
  dff_sg \filter_0/ow_1_reg[1]  ( .D(\filter_0/n8562 ), .CP(clk), .Q(
        reg_ow_1[1]) );
  dff_sg \filter_0/ow_1_reg[0]  ( .D(\filter_0/n8563 ), .CP(clk), .Q(
        reg_ow_1[0]) );
  dff_sg \filter_0/ow_2_reg[19]  ( .D(\filter_0/n8524 ), .CP(clk), .Q(
        reg_ow_2[19]) );
  dff_sg \filter_0/ow_2_reg[18]  ( .D(\filter_0/n8525 ), .CP(clk), .Q(
        reg_ow_2[18]) );
  dff_sg \filter_0/ow_2_reg[17]  ( .D(\filter_0/n8526 ), .CP(clk), .Q(
        reg_ow_2[17]) );
  dff_sg \filter_0/ow_2_reg[16]  ( .D(\filter_0/n8527 ), .CP(clk), .Q(
        reg_ow_2[16]) );
  dff_sg \filter_0/ow_2_reg[15]  ( .D(\filter_0/n8528 ), .CP(clk), .Q(
        reg_ow_2[15]) );
  dff_sg \filter_0/ow_2_reg[14]  ( .D(\filter_0/n8529 ), .CP(clk), .Q(
        reg_ow_2[14]) );
  dff_sg \filter_0/ow_2_reg[13]  ( .D(\filter_0/n8530 ), .CP(clk), .Q(
        reg_ow_2[13]) );
  dff_sg \filter_0/ow_2_reg[12]  ( .D(\filter_0/n8531 ), .CP(clk), .Q(
        reg_ow_2[12]) );
  dff_sg \filter_0/ow_2_reg[11]  ( .D(\filter_0/n8532 ), .CP(clk), .Q(
        reg_ow_2[11]) );
  dff_sg \filter_0/ow_2_reg[10]  ( .D(\filter_0/n8533 ), .CP(clk), .Q(
        reg_ow_2[10]) );
  dff_sg \filter_0/ow_2_reg[9]  ( .D(\filter_0/n8534 ), .CP(clk), .Q(
        reg_ow_2[9]) );
  dff_sg \filter_0/ow_2_reg[8]  ( .D(\filter_0/n8535 ), .CP(clk), .Q(
        reg_ow_2[8]) );
  dff_sg \filter_0/ow_2_reg[7]  ( .D(\filter_0/n8536 ), .CP(clk), .Q(
        reg_ow_2[7]) );
  dff_sg \filter_0/ow_2_reg[6]  ( .D(\filter_0/n8537 ), .CP(clk), .Q(
        reg_ow_2[6]) );
  dff_sg \filter_0/ow_2_reg[5]  ( .D(\filter_0/n8538 ), .CP(clk), .Q(
        reg_ow_2[5]) );
  dff_sg \filter_0/ow_2_reg[4]  ( .D(\filter_0/n8539 ), .CP(clk), .Q(
        reg_ow_2[4]) );
  dff_sg \filter_0/ow_2_reg[3]  ( .D(\filter_0/n8540 ), .CP(clk), .Q(
        reg_ow_2[3]) );
  dff_sg \filter_0/ow_2_reg[2]  ( .D(\filter_0/n8541 ), .CP(clk), .Q(
        reg_ow_2[2]) );
  dff_sg \filter_0/ow_2_reg[1]  ( .D(\filter_0/n8542 ), .CP(clk), .Q(
        reg_ow_2[1]) );
  dff_sg \filter_0/ow_2_reg[0]  ( .D(\filter_0/n8543 ), .CP(clk), .Q(
        reg_ow_2[0]) );
  dff_sg \filter_0/ow_3_reg[19]  ( .D(\filter_0/n8504 ), .CP(clk), .Q(
        reg_ow_3[19]) );
  dff_sg \filter_0/ow_3_reg[18]  ( .D(\filter_0/n8505 ), .CP(clk), .Q(
        reg_ow_3[18]) );
  dff_sg \filter_0/ow_3_reg[17]  ( .D(\filter_0/n8506 ), .CP(clk), .Q(
        reg_ow_3[17]) );
  dff_sg \filter_0/ow_3_reg[16]  ( .D(\filter_0/n8507 ), .CP(clk), .Q(
        reg_ow_3[16]) );
  dff_sg \filter_0/ow_3_reg[15]  ( .D(\filter_0/n8508 ), .CP(clk), .Q(
        reg_ow_3[15]) );
  dff_sg \filter_0/ow_3_reg[14]  ( .D(\filter_0/n8509 ), .CP(clk), .Q(
        reg_ow_3[14]) );
  dff_sg \filter_0/ow_3_reg[13]  ( .D(\filter_0/n8510 ), .CP(clk), .Q(
        reg_ow_3[13]) );
  dff_sg \filter_0/ow_3_reg[12]  ( .D(\filter_0/n8511 ), .CP(clk), .Q(
        reg_ow_3[12]) );
  dff_sg \filter_0/ow_3_reg[11]  ( .D(\filter_0/n8512 ), .CP(clk), .Q(
        reg_ow_3[11]) );
  dff_sg \filter_0/ow_3_reg[10]  ( .D(\filter_0/n8513 ), .CP(clk), .Q(
        reg_ow_3[10]) );
  dff_sg \filter_0/ow_3_reg[9]  ( .D(\filter_0/n8514 ), .CP(clk), .Q(
        reg_ow_3[9]) );
  dff_sg \filter_0/ow_3_reg[8]  ( .D(\filter_0/n8515 ), .CP(clk), .Q(
        reg_ow_3[8]) );
  dff_sg \filter_0/ow_3_reg[7]  ( .D(\filter_0/n8516 ), .CP(clk), .Q(
        reg_ow_3[7]) );
  dff_sg \filter_0/ow_3_reg[6]  ( .D(\filter_0/n8517 ), .CP(clk), .Q(
        reg_ow_3[6]) );
  dff_sg \filter_0/ow_3_reg[5]  ( .D(\filter_0/n8518 ), .CP(clk), .Q(
        reg_ow_3[5]) );
  dff_sg \filter_0/ow_3_reg[4]  ( .D(\filter_0/n8519 ), .CP(clk), .Q(
        reg_ow_3[4]) );
  dff_sg \filter_0/ow_3_reg[3]  ( .D(\filter_0/n8520 ), .CP(clk), .Q(
        reg_ow_3[3]) );
  dff_sg \filter_0/ow_3_reg[2]  ( .D(\filter_0/n8521 ), .CP(clk), .Q(
        reg_ow_3[2]) );
  dff_sg \filter_0/ow_3_reg[1]  ( .D(\filter_0/n8522 ), .CP(clk), .Q(
        reg_ow_3[1]) );
  dff_sg \filter_0/ow_3_reg[0]  ( .D(\filter_0/n8523 ), .CP(clk), .Q(
        reg_ow_3[0]) );
  dff_sg \filter_0/w_pointer_reg[3]  ( .D(\filter_0/n8564 ), .CP(clk), .Q(
        \filter_0/w_pointer[3] ) );
  dff_sg \filter_0/w_pointer_reg[2]  ( .D(\filter_0/n8565 ), .CP(clk), .Q(
        \filter_0/w_pointer[2] ) );
  dff_sg \filter_0/w_pointer_reg[1]  ( .D(\filter_0/n8566 ), .CP(clk), .Q(
        \filter_0/w_pointer[1] ) );
  dff_sg \filter_0/w_pointer_reg[0]  ( .D(\filter_0/n8567 ), .CP(clk), .Q(
        \filter_0/w_pointer[0] ) );
  dff_sg \filter_0/input_taken_reg  ( .D(\filter_0/n9633 ), .CP(clk), .Q(
        mask_output_filter_input_taken) );
  dff_sg \filter_0/reg_i_0_reg[0]  ( .D(\filter_0/n9632 ), .CP(clk), .Q(
        \filter_0/reg_i_0[0] ) );
  dff_sg \filter_0/reg_i_0_reg[1]  ( .D(\filter_0/n9631 ), .CP(clk), .Q(
        \filter_0/reg_i_0[1] ) );
  dff_sg \filter_0/reg_i_0_reg[2]  ( .D(\filter_0/n9630 ), .CP(clk), .Q(
        \filter_0/reg_i_0[2] ) );
  dff_sg \filter_0/reg_i_0_reg[3]  ( .D(\filter_0/n9629 ), .CP(clk), .Q(
        \filter_0/reg_i_0[3] ) );
  dff_sg \filter_0/reg_i_0_reg[4]  ( .D(\filter_0/n9628 ), .CP(clk), .Q(
        \filter_0/reg_i_0[4] ) );
  dff_sg \filter_0/reg_i_0_reg[5]  ( .D(\filter_0/n9627 ), .CP(clk), .Q(
        \filter_0/reg_i_0[5] ) );
  dff_sg \filter_0/reg_i_0_reg[6]  ( .D(\filter_0/n9626 ), .CP(clk), .Q(
        \filter_0/reg_i_0[6] ) );
  dff_sg \filter_0/reg_i_0_reg[7]  ( .D(\filter_0/n9625 ), .CP(clk), .Q(
        \filter_0/reg_i_0[7] ) );
  dff_sg \filter_0/reg_i_0_reg[8]  ( .D(\filter_0/n9624 ), .CP(clk), .Q(
        \filter_0/reg_i_0[8] ) );
  dff_sg \filter_0/reg_i_0_reg[9]  ( .D(\filter_0/n9623 ), .CP(clk), .Q(
        \filter_0/reg_i_0[9] ) );
  dff_sg \filter_0/reg_i_0_reg[10]  ( .D(\filter_0/n9622 ), .CP(clk), .Q(
        \filter_0/reg_i_0[10] ) );
  dff_sg \filter_0/reg_i_0_reg[11]  ( .D(\filter_0/n9621 ), .CP(clk), .Q(
        \filter_0/reg_i_0[11] ) );
  dff_sg \filter_0/reg_i_0_reg[12]  ( .D(\filter_0/n9620 ), .CP(clk), .Q(
        \filter_0/reg_i_0[12] ) );
  dff_sg \filter_0/reg_i_0_reg[13]  ( .D(\filter_0/n9619 ), .CP(clk), .Q(
        \filter_0/reg_i_0[13] ) );
  dff_sg \filter_0/reg_i_0_reg[14]  ( .D(\filter_0/n9618 ), .CP(clk), .Q(
        \filter_0/reg_i_0[14] ) );
  dff_sg \filter_0/reg_i_0_reg[15]  ( .D(\filter_0/n9617 ), .CP(clk), .Q(
        \filter_0/reg_i_0[15] ) );
  dff_sg \filter_0/reg_i_0_reg[16]  ( .D(\filter_0/n9616 ), .CP(clk), .Q(
        \filter_0/reg_i_0[16] ) );
  dff_sg \filter_0/reg_i_0_reg[17]  ( .D(\filter_0/n9615 ), .CP(clk), .Q(
        \filter_0/reg_i_0[17] ) );
  dff_sg \filter_0/reg_i_0_reg[18]  ( .D(\filter_0/n9614 ), .CP(clk), .Q(
        \filter_0/reg_i_0[18] ) );
  dff_sg \filter_0/reg_i_0_reg[19]  ( .D(\filter_0/n9613 ), .CP(clk), .Q(
        \filter_0/reg_i_0[19] ) );
  dff_sg \filter_0/reg_i_1_reg[0]  ( .D(\filter_0/n9612 ), .CP(clk), .Q(
        \filter_0/reg_i_1[0] ) );
  dff_sg \filter_0/reg_i_1_reg[1]  ( .D(\filter_0/n9611 ), .CP(clk), .Q(
        \filter_0/reg_i_1[1] ) );
  dff_sg \filter_0/reg_i_1_reg[2]  ( .D(\filter_0/n9610 ), .CP(clk), .Q(
        \filter_0/reg_i_1[2] ) );
  dff_sg \filter_0/reg_i_1_reg[3]  ( .D(\filter_0/n9609 ), .CP(clk), .Q(
        \filter_0/reg_i_1[3] ) );
  dff_sg \filter_0/reg_i_1_reg[4]  ( .D(\filter_0/n9608 ), .CP(clk), .Q(
        \filter_0/reg_i_1[4] ) );
  dff_sg \filter_0/reg_i_1_reg[5]  ( .D(\filter_0/n9607 ), .CP(clk), .Q(
        \filter_0/reg_i_1[5] ) );
  dff_sg \filter_0/reg_i_1_reg[6]  ( .D(\filter_0/n9606 ), .CP(clk), .Q(
        \filter_0/reg_i_1[6] ) );
  dff_sg \filter_0/reg_i_1_reg[7]  ( .D(\filter_0/n9605 ), .CP(clk), .Q(
        \filter_0/reg_i_1[7] ) );
  dff_sg \filter_0/reg_i_1_reg[8]  ( .D(\filter_0/n9604 ), .CP(clk), .Q(
        \filter_0/reg_i_1[8] ) );
  dff_sg \filter_0/reg_i_1_reg[9]  ( .D(\filter_0/n9603 ), .CP(clk), .Q(
        \filter_0/reg_i_1[9] ) );
  dff_sg \filter_0/reg_i_1_reg[10]  ( .D(\filter_0/n9602 ), .CP(clk), .Q(
        \filter_0/reg_i_1[10] ) );
  dff_sg \filter_0/reg_i_1_reg[11]  ( .D(\filter_0/n9601 ), .CP(clk), .Q(
        \filter_0/reg_i_1[11] ) );
  dff_sg \filter_0/reg_i_1_reg[12]  ( .D(\filter_0/n9600 ), .CP(clk), .Q(
        \filter_0/reg_i_1[12] ) );
  dff_sg \filter_0/reg_i_1_reg[13]  ( .D(\filter_0/n9599 ), .CP(clk), .Q(
        \filter_0/reg_i_1[13] ) );
  dff_sg \filter_0/reg_i_1_reg[14]  ( .D(\filter_0/n9598 ), .CP(clk), .Q(
        \filter_0/reg_i_1[14] ) );
  dff_sg \filter_0/reg_i_1_reg[15]  ( .D(\filter_0/n9597 ), .CP(clk), .Q(
        \filter_0/reg_i_1[15] ) );
  dff_sg \filter_0/reg_i_1_reg[16]  ( .D(\filter_0/n9596 ), .CP(clk), .Q(
        \filter_0/reg_i_1[16] ) );
  dff_sg \filter_0/reg_i_1_reg[17]  ( .D(\filter_0/n9595 ), .CP(clk), .Q(
        \filter_0/reg_i_1[17] ) );
  dff_sg \filter_0/reg_i_1_reg[18]  ( .D(\filter_0/n9594 ), .CP(clk), .Q(
        \filter_0/reg_i_1[18] ) );
  dff_sg \filter_0/reg_i_1_reg[19]  ( .D(\filter_0/n9593 ), .CP(clk), .Q(
        \filter_0/reg_i_1[19] ) );
  dff_sg \filter_0/reg_i_2_reg[0]  ( .D(\filter_0/n9592 ), .CP(clk), .Q(
        \filter_0/reg_i_2[0] ) );
  dff_sg \filter_0/reg_i_2_reg[1]  ( .D(\filter_0/n9591 ), .CP(clk), .Q(
        \filter_0/reg_i_2[1] ) );
  dff_sg \filter_0/reg_i_2_reg[2]  ( .D(\filter_0/n9590 ), .CP(clk), .Q(
        \filter_0/reg_i_2[2] ) );
  dff_sg \filter_0/reg_i_2_reg[3]  ( .D(\filter_0/n9589 ), .CP(clk), .Q(
        \filter_0/reg_i_2[3] ) );
  dff_sg \filter_0/reg_i_2_reg[4]  ( .D(\filter_0/n9588 ), .CP(clk), .Q(
        \filter_0/reg_i_2[4] ) );
  dff_sg \filter_0/reg_i_2_reg[5]  ( .D(\filter_0/n9587 ), .CP(clk), .Q(
        \filter_0/reg_i_2[5] ) );
  dff_sg \filter_0/reg_i_2_reg[6]  ( .D(\filter_0/n9586 ), .CP(clk), .Q(
        \filter_0/reg_i_2[6] ) );
  dff_sg \filter_0/reg_i_2_reg[7]  ( .D(\filter_0/n9585 ), .CP(clk), .Q(
        \filter_0/reg_i_2[7] ) );
  dff_sg \filter_0/reg_i_2_reg[8]  ( .D(\filter_0/n9584 ), .CP(clk), .Q(
        \filter_0/reg_i_2[8] ) );
  dff_sg \filter_0/reg_i_2_reg[9]  ( .D(\filter_0/n9583 ), .CP(clk), .Q(
        \filter_0/reg_i_2[9] ) );
  dff_sg \filter_0/reg_i_2_reg[10]  ( .D(\filter_0/n9582 ), .CP(clk), .Q(
        \filter_0/reg_i_2[10] ) );
  dff_sg \filter_0/reg_i_2_reg[11]  ( .D(\filter_0/n9581 ), .CP(clk), .Q(
        \filter_0/reg_i_2[11] ) );
  dff_sg \filter_0/reg_i_2_reg[12]  ( .D(\filter_0/n9580 ), .CP(clk), .Q(
        \filter_0/reg_i_2[12] ) );
  dff_sg \filter_0/reg_i_2_reg[13]  ( .D(\filter_0/n9579 ), .CP(clk), .Q(
        \filter_0/reg_i_2[13] ) );
  dff_sg \filter_0/reg_i_2_reg[14]  ( .D(\filter_0/n9578 ), .CP(clk), .Q(
        \filter_0/reg_i_2[14] ) );
  dff_sg \filter_0/reg_i_2_reg[15]  ( .D(\filter_0/n9577 ), .CP(clk), .Q(
        \filter_0/reg_i_2[15] ) );
  dff_sg \filter_0/reg_i_2_reg[16]  ( .D(\filter_0/n9576 ), .CP(clk), .Q(
        \filter_0/reg_i_2[16] ) );
  dff_sg \filter_0/reg_i_2_reg[17]  ( .D(\filter_0/n9575 ), .CP(clk), .Q(
        \filter_0/reg_i_2[17] ) );
  dff_sg \filter_0/reg_i_2_reg[18]  ( .D(\filter_0/n9574 ), .CP(clk), .Q(
        \filter_0/reg_i_2[18] ) );
  dff_sg \filter_0/reg_i_2_reg[19]  ( .D(\filter_0/n9573 ), .CP(clk), .Q(
        \filter_0/reg_i_2[19] ) );
  dff_sg \filter_0/reg_i_3_reg[0]  ( .D(\filter_0/n9572 ), .CP(clk), .Q(
        \filter_0/reg_i_3[0] ) );
  dff_sg \filter_0/reg_i_3_reg[1]  ( .D(\filter_0/n9571 ), .CP(clk), .Q(
        \filter_0/reg_i_3[1] ) );
  dff_sg \filter_0/reg_i_3_reg[2]  ( .D(\filter_0/n9570 ), .CP(clk), .Q(
        \filter_0/reg_i_3[2] ) );
  dff_sg \filter_0/reg_i_3_reg[3]  ( .D(\filter_0/n9569 ), .CP(clk), .Q(
        \filter_0/reg_i_3[3] ) );
  dff_sg \filter_0/reg_i_3_reg[4]  ( .D(\filter_0/n9568 ), .CP(clk), .Q(
        \filter_0/reg_i_3[4] ) );
  dff_sg \filter_0/reg_i_3_reg[5]  ( .D(\filter_0/n9567 ), .CP(clk), .Q(
        \filter_0/reg_i_3[5] ) );
  dff_sg \filter_0/reg_i_3_reg[6]  ( .D(\filter_0/n9566 ), .CP(clk), .Q(
        \filter_0/reg_i_3[6] ) );
  dff_sg \filter_0/reg_i_3_reg[7]  ( .D(\filter_0/n9565 ), .CP(clk), .Q(
        \filter_0/reg_i_3[7] ) );
  dff_sg \filter_0/reg_i_3_reg[8]  ( .D(\filter_0/n9564 ), .CP(clk), .Q(
        \filter_0/reg_i_3[8] ) );
  dff_sg \filter_0/reg_i_3_reg[9]  ( .D(\filter_0/n9563 ), .CP(clk), .Q(
        \filter_0/reg_i_3[9] ) );
  dff_sg \filter_0/reg_i_3_reg[10]  ( .D(\filter_0/n9562 ), .CP(clk), .Q(
        \filter_0/reg_i_3[10] ) );
  dff_sg \filter_0/reg_i_3_reg[11]  ( .D(\filter_0/n9561 ), .CP(clk), .Q(
        \filter_0/reg_i_3[11] ) );
  dff_sg \filter_0/reg_i_3_reg[12]  ( .D(\filter_0/n9560 ), .CP(clk), .Q(
        \filter_0/reg_i_3[12] ) );
  dff_sg \filter_0/reg_i_3_reg[13]  ( .D(\filter_0/n9559 ), .CP(clk), .Q(
        \filter_0/reg_i_3[13] ) );
  dff_sg \filter_0/reg_i_3_reg[14]  ( .D(\filter_0/n9558 ), .CP(clk), .Q(
        \filter_0/reg_i_3[14] ) );
  dff_sg \filter_0/reg_i_3_reg[15]  ( .D(\filter_0/n9557 ), .CP(clk), .Q(
        \filter_0/reg_i_3[15] ) );
  dff_sg \filter_0/reg_i_3_reg[16]  ( .D(\filter_0/n9556 ), .CP(clk), .Q(
        \filter_0/reg_i_3[16] ) );
  dff_sg \filter_0/reg_i_3_reg[17]  ( .D(\filter_0/n9555 ), .CP(clk), .Q(
        \filter_0/reg_i_3[17] ) );
  dff_sg \filter_0/reg_i_3_reg[18]  ( .D(\filter_0/n9554 ), .CP(clk), .Q(
        \filter_0/reg_i_3[18] ) );
  dff_sg \filter_0/reg_i_3_reg[19]  ( .D(\filter_0/n9553 ), .CP(clk), .Q(
        \filter_0/reg_i_3[19] ) );
  dff_sg \filter_0/reg_i_4_reg[0]  ( .D(\filter_0/n9552 ), .CP(clk), .Q(
        \filter_0/reg_i_4[0] ) );
  dff_sg \filter_0/reg_i_4_reg[1]  ( .D(\filter_0/n9551 ), .CP(clk), .Q(
        \filter_0/reg_i_4[1] ) );
  dff_sg \filter_0/reg_i_4_reg[2]  ( .D(\filter_0/n9550 ), .CP(clk), .Q(
        \filter_0/reg_i_4[2] ) );
  dff_sg \filter_0/reg_i_4_reg[3]  ( .D(\filter_0/n9549 ), .CP(clk), .Q(
        \filter_0/reg_i_4[3] ) );
  dff_sg \filter_0/reg_i_4_reg[4]  ( .D(\filter_0/n9548 ), .CP(clk), .Q(
        \filter_0/reg_i_4[4] ) );
  dff_sg \filter_0/reg_i_4_reg[5]  ( .D(\filter_0/n9547 ), .CP(clk), .Q(
        \filter_0/reg_i_4[5] ) );
  dff_sg \filter_0/reg_i_4_reg[6]  ( .D(\filter_0/n9546 ), .CP(clk), .Q(
        \filter_0/reg_i_4[6] ) );
  dff_sg \filter_0/reg_i_4_reg[7]  ( .D(\filter_0/n9545 ), .CP(clk), .Q(
        \filter_0/reg_i_4[7] ) );
  dff_sg \filter_0/reg_i_4_reg[8]  ( .D(\filter_0/n9544 ), .CP(clk), .Q(
        \filter_0/reg_i_4[8] ) );
  dff_sg \filter_0/reg_i_4_reg[9]  ( .D(\filter_0/n9543 ), .CP(clk), .Q(
        \filter_0/reg_i_4[9] ) );
  dff_sg \filter_0/reg_i_4_reg[10]  ( .D(\filter_0/n9542 ), .CP(clk), .Q(
        \filter_0/reg_i_4[10] ) );
  dff_sg \filter_0/reg_i_4_reg[11]  ( .D(\filter_0/n9541 ), .CP(clk), .Q(
        \filter_0/reg_i_4[11] ) );
  dff_sg \filter_0/reg_i_4_reg[12]  ( .D(\filter_0/n9540 ), .CP(clk), .Q(
        \filter_0/reg_i_4[12] ) );
  dff_sg \filter_0/reg_i_4_reg[13]  ( .D(\filter_0/n9539 ), .CP(clk), .Q(
        \filter_0/reg_i_4[13] ) );
  dff_sg \filter_0/reg_i_4_reg[14]  ( .D(\filter_0/n9538 ), .CP(clk), .Q(
        \filter_0/reg_i_4[14] ) );
  dff_sg \filter_0/reg_i_4_reg[15]  ( .D(\filter_0/n9537 ), .CP(clk), .Q(
        \filter_0/reg_i_4[15] ) );
  dff_sg \filter_0/reg_i_4_reg[16]  ( .D(\filter_0/n9536 ), .CP(clk), .Q(
        \filter_0/reg_i_4[16] ) );
  dff_sg \filter_0/reg_i_4_reg[17]  ( .D(\filter_0/n9535 ), .CP(clk), .Q(
        \filter_0/reg_i_4[17] ) );
  dff_sg \filter_0/reg_i_4_reg[18]  ( .D(\filter_0/n9534 ), .CP(clk), .Q(
        \filter_0/reg_i_4[18] ) );
  dff_sg \filter_0/reg_i_4_reg[19]  ( .D(\filter_0/n9533 ), .CP(clk), .Q(
        \filter_0/reg_i_4[19] ) );
  dff_sg \filter_0/reg_i_5_reg[0]  ( .D(\filter_0/n9532 ), .CP(clk), .Q(
        \filter_0/reg_i_5[0] ) );
  dff_sg \filter_0/reg_i_5_reg[1]  ( .D(\filter_0/n9531 ), .CP(clk), .Q(
        \filter_0/reg_i_5[1] ) );
  dff_sg \filter_0/reg_i_5_reg[2]  ( .D(\filter_0/n9530 ), .CP(clk), .Q(
        \filter_0/reg_i_5[2] ) );
  dff_sg \filter_0/reg_i_5_reg[3]  ( .D(\filter_0/n9529 ), .CP(clk), .Q(
        \filter_0/reg_i_5[3] ) );
  dff_sg \filter_0/reg_i_5_reg[4]  ( .D(\filter_0/n9528 ), .CP(clk), .Q(
        \filter_0/reg_i_5[4] ) );
  dff_sg \filter_0/reg_i_5_reg[5]  ( .D(\filter_0/n9527 ), .CP(clk), .Q(
        \filter_0/reg_i_5[5] ) );
  dff_sg \filter_0/reg_i_5_reg[6]  ( .D(\filter_0/n9526 ), .CP(clk), .Q(
        \filter_0/reg_i_5[6] ) );
  dff_sg \filter_0/reg_i_5_reg[7]  ( .D(\filter_0/n9525 ), .CP(clk), .Q(
        \filter_0/reg_i_5[7] ) );
  dff_sg \filter_0/reg_i_5_reg[8]  ( .D(\filter_0/n9524 ), .CP(clk), .Q(
        \filter_0/reg_i_5[8] ) );
  dff_sg \filter_0/reg_i_5_reg[9]  ( .D(\filter_0/n9523 ), .CP(clk), .Q(
        \filter_0/reg_i_5[9] ) );
  dff_sg \filter_0/reg_i_5_reg[10]  ( .D(\filter_0/n9522 ), .CP(clk), .Q(
        \filter_0/reg_i_5[10] ) );
  dff_sg \filter_0/reg_i_5_reg[11]  ( .D(\filter_0/n9521 ), .CP(clk), .Q(
        \filter_0/reg_i_5[11] ) );
  dff_sg \filter_0/reg_i_5_reg[12]  ( .D(\filter_0/n9520 ), .CP(clk), .Q(
        \filter_0/reg_i_5[12] ) );
  dff_sg \filter_0/reg_i_5_reg[13]  ( .D(\filter_0/n9519 ), .CP(clk), .Q(
        \filter_0/reg_i_5[13] ) );
  dff_sg \filter_0/reg_i_5_reg[14]  ( .D(\filter_0/n9518 ), .CP(clk), .Q(
        \filter_0/reg_i_5[14] ) );
  dff_sg \filter_0/reg_i_5_reg[15]  ( .D(\filter_0/n9517 ), .CP(clk), .Q(
        \filter_0/reg_i_5[15] ) );
  dff_sg \filter_0/reg_i_5_reg[16]  ( .D(\filter_0/n9516 ), .CP(clk), .Q(
        \filter_0/reg_i_5[16] ) );
  dff_sg \filter_0/reg_i_5_reg[17]  ( .D(\filter_0/n9515 ), .CP(clk), .Q(
        \filter_0/reg_i_5[17] ) );
  dff_sg \filter_0/reg_i_5_reg[18]  ( .D(\filter_0/n9514 ), .CP(clk), .Q(
        \filter_0/reg_i_5[18] ) );
  dff_sg \filter_0/reg_i_5_reg[19]  ( .D(\filter_0/n9513 ), .CP(clk), .Q(
        \filter_0/reg_i_5[19] ) );
  dff_sg \filter_0/reg_i_6_reg[0]  ( .D(\filter_0/n9512 ), .CP(clk), .Q(
        \filter_0/reg_i_6[0] ) );
  dff_sg \filter_0/reg_i_6_reg[1]  ( .D(\filter_0/n9511 ), .CP(clk), .Q(
        \filter_0/reg_i_6[1] ) );
  dff_sg \filter_0/reg_i_6_reg[2]  ( .D(\filter_0/n9510 ), .CP(clk), .Q(
        \filter_0/reg_i_6[2] ) );
  dff_sg \filter_0/reg_i_6_reg[3]  ( .D(\filter_0/n9509 ), .CP(clk), .Q(
        \filter_0/reg_i_6[3] ) );
  dff_sg \filter_0/reg_i_6_reg[4]  ( .D(\filter_0/n9508 ), .CP(clk), .Q(
        \filter_0/reg_i_6[4] ) );
  dff_sg \filter_0/reg_i_6_reg[5]  ( .D(\filter_0/n9507 ), .CP(clk), .Q(
        \filter_0/reg_i_6[5] ) );
  dff_sg \filter_0/reg_i_6_reg[6]  ( .D(\filter_0/n9506 ), .CP(clk), .Q(
        \filter_0/reg_i_6[6] ) );
  dff_sg \filter_0/reg_i_6_reg[7]  ( .D(\filter_0/n9505 ), .CP(clk), .Q(
        \filter_0/reg_i_6[7] ) );
  dff_sg \filter_0/reg_i_6_reg[8]  ( .D(\filter_0/n9504 ), .CP(clk), .Q(
        \filter_0/reg_i_6[8] ) );
  dff_sg \filter_0/reg_i_6_reg[9]  ( .D(\filter_0/n9503 ), .CP(clk), .Q(
        \filter_0/reg_i_6[9] ) );
  dff_sg \filter_0/reg_i_6_reg[10]  ( .D(\filter_0/n9502 ), .CP(clk), .Q(
        \filter_0/reg_i_6[10] ) );
  dff_sg \filter_0/reg_i_6_reg[11]  ( .D(\filter_0/n9501 ), .CP(clk), .Q(
        \filter_0/reg_i_6[11] ) );
  dff_sg \filter_0/reg_i_6_reg[12]  ( .D(\filter_0/n9500 ), .CP(clk), .Q(
        \filter_0/reg_i_6[12] ) );
  dff_sg \filter_0/reg_i_6_reg[13]  ( .D(\filter_0/n9499 ), .CP(clk), .Q(
        \filter_0/reg_i_6[13] ) );
  dff_sg \filter_0/reg_i_6_reg[14]  ( .D(\filter_0/n9498 ), .CP(clk), .Q(
        \filter_0/reg_i_6[14] ) );
  dff_sg \filter_0/reg_i_6_reg[15]  ( .D(\filter_0/n9497 ), .CP(clk), .Q(
        \filter_0/reg_i_6[15] ) );
  dff_sg \filter_0/reg_i_6_reg[16]  ( .D(\filter_0/n9496 ), .CP(clk), .Q(
        \filter_0/reg_i_6[16] ) );
  dff_sg \filter_0/reg_i_6_reg[17]  ( .D(\filter_0/n9495 ), .CP(clk), .Q(
        \filter_0/reg_i_6[17] ) );
  dff_sg \filter_0/reg_i_6_reg[18]  ( .D(\filter_0/n9494 ), .CP(clk), .Q(
        \filter_0/reg_i_6[18] ) );
  dff_sg \filter_0/reg_i_6_reg[19]  ( .D(\filter_0/n9493 ), .CP(clk), .Q(
        \filter_0/reg_i_6[19] ) );
  dff_sg \filter_0/reg_i_7_reg[0]  ( .D(\filter_0/n9492 ), .CP(clk), .Q(
        \filter_0/reg_i_7[0] ) );
  dff_sg \filter_0/reg_i_7_reg[1]  ( .D(\filter_0/n9491 ), .CP(clk), .Q(
        \filter_0/reg_i_7[1] ) );
  dff_sg \filter_0/reg_i_7_reg[2]  ( .D(\filter_0/n9490 ), .CP(clk), .Q(
        \filter_0/reg_i_7[2] ) );
  dff_sg \filter_0/reg_i_7_reg[3]  ( .D(\filter_0/n9489 ), .CP(clk), .Q(
        \filter_0/reg_i_7[3] ) );
  dff_sg \filter_0/reg_i_7_reg[4]  ( .D(\filter_0/n9488 ), .CP(clk), .Q(
        \filter_0/reg_i_7[4] ) );
  dff_sg \filter_0/reg_i_7_reg[5]  ( .D(\filter_0/n9487 ), .CP(clk), .Q(
        \filter_0/reg_i_7[5] ) );
  dff_sg \filter_0/reg_i_7_reg[6]  ( .D(\filter_0/n9486 ), .CP(clk), .Q(
        \filter_0/reg_i_7[6] ) );
  dff_sg \filter_0/reg_i_7_reg[7]  ( .D(\filter_0/n9485 ), .CP(clk), .Q(
        \filter_0/reg_i_7[7] ) );
  dff_sg \filter_0/reg_i_7_reg[8]  ( .D(\filter_0/n9484 ), .CP(clk), .Q(
        \filter_0/reg_i_7[8] ) );
  dff_sg \filter_0/reg_i_7_reg[9]  ( .D(\filter_0/n9483 ), .CP(clk), .Q(
        \filter_0/reg_i_7[9] ) );
  dff_sg \filter_0/reg_i_7_reg[10]  ( .D(\filter_0/n9482 ), .CP(clk), .Q(
        \filter_0/reg_i_7[10] ) );
  dff_sg \filter_0/reg_i_7_reg[11]  ( .D(\filter_0/n9481 ), .CP(clk), .Q(
        \filter_0/reg_i_7[11] ) );
  dff_sg \filter_0/reg_i_7_reg[12]  ( .D(\filter_0/n9480 ), .CP(clk), .Q(
        \filter_0/reg_i_7[12] ) );
  dff_sg \filter_0/reg_i_7_reg[13]  ( .D(\filter_0/n9479 ), .CP(clk), .Q(
        \filter_0/reg_i_7[13] ) );
  dff_sg \filter_0/reg_i_7_reg[14]  ( .D(\filter_0/n9478 ), .CP(clk), .Q(
        \filter_0/reg_i_7[14] ) );
  dff_sg \filter_0/reg_i_7_reg[15]  ( .D(\filter_0/n9477 ), .CP(clk), .Q(
        \filter_0/reg_i_7[15] ) );
  dff_sg \filter_0/reg_i_7_reg[16]  ( .D(\filter_0/n9476 ), .CP(clk), .Q(
        \filter_0/reg_i_7[16] ) );
  dff_sg \filter_0/reg_i_7_reg[17]  ( .D(\filter_0/n9475 ), .CP(clk), .Q(
        \filter_0/reg_i_7[17] ) );
  dff_sg \filter_0/reg_i_7_reg[18]  ( .D(\filter_0/n9474 ), .CP(clk), .Q(
        \filter_0/reg_i_7[18] ) );
  dff_sg \filter_0/reg_i_7_reg[19]  ( .D(\filter_0/n9473 ), .CP(clk), .Q(
        \filter_0/reg_i_7[19] ) );
  dff_sg \filter_0/reg_i_8_reg[0]  ( .D(\filter_0/n9472 ), .CP(clk), .Q(
        \filter_0/reg_i_8[0] ) );
  dff_sg \filter_0/reg_i_8_reg[1]  ( .D(\filter_0/n9471 ), .CP(clk), .Q(
        \filter_0/reg_i_8[1] ) );
  dff_sg \filter_0/reg_i_8_reg[2]  ( .D(\filter_0/n9470 ), .CP(clk), .Q(
        \filter_0/reg_i_8[2] ) );
  dff_sg \filter_0/reg_i_8_reg[3]  ( .D(\filter_0/n9469 ), .CP(clk), .Q(
        \filter_0/reg_i_8[3] ) );
  dff_sg \filter_0/reg_i_8_reg[4]  ( .D(\filter_0/n9468 ), .CP(clk), .Q(
        \filter_0/reg_i_8[4] ) );
  dff_sg \filter_0/reg_i_8_reg[5]  ( .D(\filter_0/n9467 ), .CP(clk), .Q(
        \filter_0/reg_i_8[5] ) );
  dff_sg \filter_0/reg_i_8_reg[6]  ( .D(\filter_0/n9466 ), .CP(clk), .Q(
        \filter_0/reg_i_8[6] ) );
  dff_sg \filter_0/reg_i_8_reg[7]  ( .D(\filter_0/n9465 ), .CP(clk), .Q(
        \filter_0/reg_i_8[7] ) );
  dff_sg \filter_0/reg_i_8_reg[8]  ( .D(\filter_0/n9464 ), .CP(clk), .Q(
        \filter_0/reg_i_8[8] ) );
  dff_sg \filter_0/reg_i_8_reg[9]  ( .D(\filter_0/n9463 ), .CP(clk), .Q(
        \filter_0/reg_i_8[9] ) );
  dff_sg \filter_0/reg_i_8_reg[10]  ( .D(\filter_0/n9462 ), .CP(clk), .Q(
        \filter_0/reg_i_8[10] ) );
  dff_sg \filter_0/reg_i_8_reg[11]  ( .D(\filter_0/n9461 ), .CP(clk), .Q(
        \filter_0/reg_i_8[11] ) );
  dff_sg \filter_0/reg_i_8_reg[12]  ( .D(\filter_0/n9460 ), .CP(clk), .Q(
        \filter_0/reg_i_8[12] ) );
  dff_sg \filter_0/reg_i_8_reg[13]  ( .D(\filter_0/n9459 ), .CP(clk), .Q(
        \filter_0/reg_i_8[13] ) );
  dff_sg \filter_0/reg_i_8_reg[14]  ( .D(\filter_0/n9458 ), .CP(clk), .Q(
        \filter_0/reg_i_8[14] ) );
  dff_sg \filter_0/reg_i_8_reg[15]  ( .D(\filter_0/n9457 ), .CP(clk), .Q(
        \filter_0/reg_i_8[15] ) );
  dff_sg \filter_0/reg_i_8_reg[16]  ( .D(\filter_0/n9456 ), .CP(clk), .Q(
        \filter_0/reg_i_8[16] ) );
  dff_sg \filter_0/reg_i_8_reg[17]  ( .D(\filter_0/n9455 ), .CP(clk), .Q(
        \filter_0/reg_i_8[17] ) );
  dff_sg \filter_0/reg_i_8_reg[18]  ( .D(\filter_0/n9454 ), .CP(clk), .Q(
        \filter_0/reg_i_8[18] ) );
  dff_sg \filter_0/reg_i_8_reg[19]  ( .D(\filter_0/n9453 ), .CP(clk), .Q(
        \filter_0/reg_i_8[19] ) );
  dff_sg \filter_0/reg_i_9_reg[0]  ( .D(\filter_0/n9452 ), .CP(clk), .Q(
        \filter_0/reg_i_9[0] ) );
  dff_sg \filter_0/reg_i_9_reg[1]  ( .D(\filter_0/n9451 ), .CP(clk), .Q(
        \filter_0/reg_i_9[1] ) );
  dff_sg \filter_0/reg_i_9_reg[2]  ( .D(\filter_0/n9450 ), .CP(clk), .Q(
        \filter_0/reg_i_9[2] ) );
  dff_sg \filter_0/reg_i_9_reg[3]  ( .D(\filter_0/n9449 ), .CP(clk), .Q(
        \filter_0/reg_i_9[3] ) );
  dff_sg \filter_0/reg_i_9_reg[4]  ( .D(\filter_0/n9448 ), .CP(clk), .Q(
        \filter_0/reg_i_9[4] ) );
  dff_sg \filter_0/reg_i_9_reg[5]  ( .D(\filter_0/n9447 ), .CP(clk), .Q(
        \filter_0/reg_i_9[5] ) );
  dff_sg \filter_0/reg_i_9_reg[6]  ( .D(\filter_0/n9446 ), .CP(clk), .Q(
        \filter_0/reg_i_9[6] ) );
  dff_sg \filter_0/reg_i_9_reg[7]  ( .D(\filter_0/n9445 ), .CP(clk), .Q(
        \filter_0/reg_i_9[7] ) );
  dff_sg \filter_0/reg_i_9_reg[8]  ( .D(\filter_0/n9444 ), .CP(clk), .Q(
        \filter_0/reg_i_9[8] ) );
  dff_sg \filter_0/reg_i_9_reg[9]  ( .D(\filter_0/n9443 ), .CP(clk), .Q(
        \filter_0/reg_i_9[9] ) );
  dff_sg \filter_0/reg_i_9_reg[10]  ( .D(\filter_0/n9442 ), .CP(clk), .Q(
        \filter_0/reg_i_9[10] ) );
  dff_sg \filter_0/reg_i_9_reg[11]  ( .D(\filter_0/n9441 ), .CP(clk), .Q(
        \filter_0/reg_i_9[11] ) );
  dff_sg \filter_0/reg_i_9_reg[12]  ( .D(\filter_0/n9440 ), .CP(clk), .Q(
        \filter_0/reg_i_9[12] ) );
  dff_sg \filter_0/reg_i_9_reg[13]  ( .D(\filter_0/n9439 ), .CP(clk), .Q(
        \filter_0/reg_i_9[13] ) );
  dff_sg \filter_0/reg_i_9_reg[14]  ( .D(\filter_0/n9438 ), .CP(clk), .Q(
        \filter_0/reg_i_9[14] ) );
  dff_sg \filter_0/reg_i_9_reg[15]  ( .D(\filter_0/n9437 ), .CP(clk), .Q(
        \filter_0/reg_i_9[15] ) );
  dff_sg \filter_0/reg_i_9_reg[16]  ( .D(\filter_0/n9436 ), .CP(clk), .Q(
        \filter_0/reg_i_9[16] ) );
  dff_sg \filter_0/reg_i_9_reg[17]  ( .D(\filter_0/n9435 ), .CP(clk), .Q(
        \filter_0/reg_i_9[17] ) );
  dff_sg \filter_0/reg_i_9_reg[18]  ( .D(\filter_0/n9434 ), .CP(clk), .Q(
        \filter_0/reg_i_9[18] ) );
  dff_sg \filter_0/reg_i_9_reg[19]  ( .D(\filter_0/n9433 ), .CP(clk), .Q(
        \filter_0/reg_i_9[19] ) );
  dff_sg \filter_0/reg_i_10_reg[0]  ( .D(\filter_0/n9432 ), .CP(clk), .Q(
        \filter_0/reg_i_10[0] ) );
  dff_sg \filter_0/reg_i_10_reg[1]  ( .D(\filter_0/n9431 ), .CP(clk), .Q(
        \filter_0/reg_i_10[1] ) );
  dff_sg \filter_0/reg_i_10_reg[2]  ( .D(\filter_0/n9430 ), .CP(clk), .Q(
        \filter_0/reg_i_10[2] ) );
  dff_sg \filter_0/reg_i_10_reg[3]  ( .D(\filter_0/n9429 ), .CP(clk), .Q(
        \filter_0/reg_i_10[3] ) );
  dff_sg \filter_0/reg_i_10_reg[4]  ( .D(\filter_0/n9428 ), .CP(clk), .Q(
        \filter_0/reg_i_10[4] ) );
  dff_sg \filter_0/reg_i_10_reg[5]  ( .D(\filter_0/n9427 ), .CP(clk), .Q(
        \filter_0/reg_i_10[5] ) );
  dff_sg \filter_0/reg_i_10_reg[6]  ( .D(\filter_0/n9426 ), .CP(clk), .Q(
        \filter_0/reg_i_10[6] ) );
  dff_sg \filter_0/reg_i_10_reg[7]  ( .D(\filter_0/n9425 ), .CP(clk), .Q(
        \filter_0/reg_i_10[7] ) );
  dff_sg \filter_0/reg_i_10_reg[8]  ( .D(\filter_0/n9424 ), .CP(clk), .Q(
        \filter_0/reg_i_10[8] ) );
  dff_sg \filter_0/reg_i_10_reg[9]  ( .D(\filter_0/n9423 ), .CP(clk), .Q(
        \filter_0/reg_i_10[9] ) );
  dff_sg \filter_0/reg_i_10_reg[10]  ( .D(\filter_0/n9422 ), .CP(clk), .Q(
        \filter_0/reg_i_10[10] ) );
  dff_sg \filter_0/reg_i_10_reg[11]  ( .D(\filter_0/n9421 ), .CP(clk), .Q(
        \filter_0/reg_i_10[11] ) );
  dff_sg \filter_0/reg_i_10_reg[12]  ( .D(\filter_0/n9420 ), .CP(clk), .Q(
        \filter_0/reg_i_10[12] ) );
  dff_sg \filter_0/reg_i_10_reg[13]  ( .D(\filter_0/n9419 ), .CP(clk), .Q(
        \filter_0/reg_i_10[13] ) );
  dff_sg \filter_0/reg_i_10_reg[14]  ( .D(\filter_0/n9418 ), .CP(clk), .Q(
        \filter_0/reg_i_10[14] ) );
  dff_sg \filter_0/reg_i_10_reg[15]  ( .D(\filter_0/n9417 ), .CP(clk), .Q(
        \filter_0/reg_i_10[15] ) );
  dff_sg \filter_0/reg_i_10_reg[16]  ( .D(\filter_0/n9416 ), .CP(clk), .Q(
        \filter_0/reg_i_10[16] ) );
  dff_sg \filter_0/reg_i_10_reg[17]  ( .D(\filter_0/n9415 ), .CP(clk), .Q(
        \filter_0/reg_i_10[17] ) );
  dff_sg \filter_0/reg_i_10_reg[18]  ( .D(\filter_0/n9414 ), .CP(clk), .Q(
        \filter_0/reg_i_10[18] ) );
  dff_sg \filter_0/reg_i_10_reg[19]  ( .D(\filter_0/n9413 ), .CP(clk), .Q(
        \filter_0/reg_i_10[19] ) );
  dff_sg \filter_0/reg_i_11_reg[0]  ( .D(\filter_0/n9412 ), .CP(clk), .Q(
        \filter_0/reg_i_11[0] ) );
  dff_sg \filter_0/reg_i_11_reg[1]  ( .D(\filter_0/n9411 ), .CP(clk), .Q(
        \filter_0/reg_i_11[1] ) );
  dff_sg \filter_0/reg_i_11_reg[2]  ( .D(\filter_0/n9410 ), .CP(clk), .Q(
        \filter_0/reg_i_11[2] ) );
  dff_sg \filter_0/reg_i_11_reg[3]  ( .D(\filter_0/n9409 ), .CP(clk), .Q(
        \filter_0/reg_i_11[3] ) );
  dff_sg \filter_0/reg_i_11_reg[4]  ( .D(\filter_0/n9408 ), .CP(clk), .Q(
        \filter_0/reg_i_11[4] ) );
  dff_sg \filter_0/reg_i_11_reg[5]  ( .D(\filter_0/n9407 ), .CP(clk), .Q(
        \filter_0/reg_i_11[5] ) );
  dff_sg \filter_0/reg_i_11_reg[6]  ( .D(\filter_0/n9406 ), .CP(clk), .Q(
        \filter_0/reg_i_11[6] ) );
  dff_sg \filter_0/reg_i_11_reg[7]  ( .D(\filter_0/n9405 ), .CP(clk), .Q(
        \filter_0/reg_i_11[7] ) );
  dff_sg \filter_0/reg_i_11_reg[8]  ( .D(\filter_0/n9404 ), .CP(clk), .Q(
        \filter_0/reg_i_11[8] ) );
  dff_sg \filter_0/reg_i_11_reg[9]  ( .D(\filter_0/n9403 ), .CP(clk), .Q(
        \filter_0/reg_i_11[9] ) );
  dff_sg \filter_0/reg_i_11_reg[10]  ( .D(\filter_0/n9402 ), .CP(clk), .Q(
        \filter_0/reg_i_11[10] ) );
  dff_sg \filter_0/reg_i_11_reg[11]  ( .D(\filter_0/n9401 ), .CP(clk), .Q(
        \filter_0/reg_i_11[11] ) );
  dff_sg \filter_0/reg_i_11_reg[12]  ( .D(\filter_0/n9400 ), .CP(clk), .Q(
        \filter_0/reg_i_11[12] ) );
  dff_sg \filter_0/reg_i_11_reg[13]  ( .D(\filter_0/n9399 ), .CP(clk), .Q(
        \filter_0/reg_i_11[13] ) );
  dff_sg \filter_0/reg_i_11_reg[14]  ( .D(\filter_0/n9398 ), .CP(clk), .Q(
        \filter_0/reg_i_11[14] ) );
  dff_sg \filter_0/reg_i_11_reg[15]  ( .D(\filter_0/n9397 ), .CP(clk), .Q(
        \filter_0/reg_i_11[15] ) );
  dff_sg \filter_0/reg_i_11_reg[16]  ( .D(\filter_0/n9396 ), .CP(clk), .Q(
        \filter_0/reg_i_11[16] ) );
  dff_sg \filter_0/reg_i_11_reg[17]  ( .D(\filter_0/n9395 ), .CP(clk), .Q(
        \filter_0/reg_i_11[17] ) );
  dff_sg \filter_0/reg_i_11_reg[18]  ( .D(\filter_0/n9394 ), .CP(clk), .Q(
        \filter_0/reg_i_11[18] ) );
  dff_sg \filter_0/reg_i_11_reg[19]  ( .D(\filter_0/n9393 ), .CP(clk), .Q(
        \filter_0/reg_i_11[19] ) );
  dff_sg \filter_0/reg_i_12_reg[0]  ( .D(\filter_0/n9392 ), .CP(clk), .Q(
        \filter_0/reg_i_12[0] ) );
  dff_sg \filter_0/reg_i_12_reg[1]  ( .D(\filter_0/n9391 ), .CP(clk), .Q(
        \filter_0/reg_i_12[1] ) );
  dff_sg \filter_0/reg_i_12_reg[2]  ( .D(\filter_0/n9390 ), .CP(clk), .Q(
        \filter_0/reg_i_12[2] ) );
  dff_sg \filter_0/reg_i_12_reg[3]  ( .D(\filter_0/n9389 ), .CP(clk), .Q(
        \filter_0/reg_i_12[3] ) );
  dff_sg \filter_0/reg_i_12_reg[4]  ( .D(\filter_0/n9388 ), .CP(clk), .Q(
        \filter_0/reg_i_12[4] ) );
  dff_sg \filter_0/reg_i_12_reg[5]  ( .D(\filter_0/n9387 ), .CP(clk), .Q(
        \filter_0/reg_i_12[5] ) );
  dff_sg \filter_0/reg_i_12_reg[6]  ( .D(\filter_0/n9386 ), .CP(clk), .Q(
        \filter_0/reg_i_12[6] ) );
  dff_sg \filter_0/reg_i_12_reg[7]  ( .D(\filter_0/n9385 ), .CP(clk), .Q(
        \filter_0/reg_i_12[7] ) );
  dff_sg \filter_0/reg_i_12_reg[8]  ( .D(\filter_0/n9384 ), .CP(clk), .Q(
        \filter_0/reg_i_12[8] ) );
  dff_sg \filter_0/reg_i_12_reg[9]  ( .D(\filter_0/n9383 ), .CP(clk), .Q(
        \filter_0/reg_i_12[9] ) );
  dff_sg \filter_0/reg_i_12_reg[10]  ( .D(\filter_0/n9382 ), .CP(clk), .Q(
        \filter_0/reg_i_12[10] ) );
  dff_sg \filter_0/reg_i_12_reg[11]  ( .D(\filter_0/n9381 ), .CP(clk), .Q(
        \filter_0/reg_i_12[11] ) );
  dff_sg \filter_0/reg_i_12_reg[12]  ( .D(\filter_0/n9380 ), .CP(clk), .Q(
        \filter_0/reg_i_12[12] ) );
  dff_sg \filter_0/reg_i_12_reg[13]  ( .D(\filter_0/n9379 ), .CP(clk), .Q(
        \filter_0/reg_i_12[13] ) );
  dff_sg \filter_0/reg_i_12_reg[14]  ( .D(\filter_0/n9378 ), .CP(clk), .Q(
        \filter_0/reg_i_12[14] ) );
  dff_sg \filter_0/reg_i_12_reg[15]  ( .D(\filter_0/n9377 ), .CP(clk), .Q(
        \filter_0/reg_i_12[15] ) );
  dff_sg \filter_0/reg_i_12_reg[16]  ( .D(\filter_0/n9376 ), .CP(clk), .Q(
        \filter_0/reg_i_12[16] ) );
  dff_sg \filter_0/reg_i_12_reg[17]  ( .D(\filter_0/n9375 ), .CP(clk), .Q(
        \filter_0/reg_i_12[17] ) );
  dff_sg \filter_0/reg_i_12_reg[18]  ( .D(\filter_0/n9374 ), .CP(clk), .Q(
        \filter_0/reg_i_12[18] ) );
  dff_sg \filter_0/reg_i_12_reg[19]  ( .D(\filter_0/n9373 ), .CP(clk), .Q(
        \filter_0/reg_i_12[19] ) );
  dff_sg \filter_0/reg_i_13_reg[0]  ( .D(\filter_0/n9372 ), .CP(clk), .Q(
        \filter_0/reg_i_13[0] ) );
  dff_sg \filter_0/reg_i_13_reg[1]  ( .D(\filter_0/n9371 ), .CP(clk), .Q(
        \filter_0/reg_i_13[1] ) );
  dff_sg \filter_0/reg_i_13_reg[2]  ( .D(\filter_0/n9370 ), .CP(clk), .Q(
        \filter_0/reg_i_13[2] ) );
  dff_sg \filter_0/reg_i_13_reg[3]  ( .D(\filter_0/n9369 ), .CP(clk), .Q(
        \filter_0/reg_i_13[3] ) );
  dff_sg \filter_0/reg_i_13_reg[4]  ( .D(\filter_0/n9368 ), .CP(clk), .Q(
        \filter_0/reg_i_13[4] ) );
  dff_sg \filter_0/reg_i_13_reg[5]  ( .D(\filter_0/n9367 ), .CP(clk), .Q(
        \filter_0/reg_i_13[5] ) );
  dff_sg \filter_0/reg_i_13_reg[6]  ( .D(\filter_0/n9366 ), .CP(clk), .Q(
        \filter_0/reg_i_13[6] ) );
  dff_sg \filter_0/reg_i_13_reg[7]  ( .D(\filter_0/n9365 ), .CP(clk), .Q(
        \filter_0/reg_i_13[7] ) );
  dff_sg \filter_0/reg_i_13_reg[8]  ( .D(\filter_0/n9364 ), .CP(clk), .Q(
        \filter_0/reg_i_13[8] ) );
  dff_sg \filter_0/reg_i_13_reg[9]  ( .D(\filter_0/n9363 ), .CP(clk), .Q(
        \filter_0/reg_i_13[9] ) );
  dff_sg \filter_0/reg_i_13_reg[10]  ( .D(\filter_0/n9362 ), .CP(clk), .Q(
        \filter_0/reg_i_13[10] ) );
  dff_sg \filter_0/reg_i_13_reg[11]  ( .D(\filter_0/n9361 ), .CP(clk), .Q(
        \filter_0/reg_i_13[11] ) );
  dff_sg \filter_0/reg_i_13_reg[12]  ( .D(\filter_0/n9360 ), .CP(clk), .Q(
        \filter_0/reg_i_13[12] ) );
  dff_sg \filter_0/reg_i_13_reg[13]  ( .D(\filter_0/n9359 ), .CP(clk), .Q(
        \filter_0/reg_i_13[13] ) );
  dff_sg \filter_0/reg_i_13_reg[14]  ( .D(\filter_0/n9358 ), .CP(clk), .Q(
        \filter_0/reg_i_13[14] ) );
  dff_sg \filter_0/reg_i_13_reg[15]  ( .D(\filter_0/n9357 ), .CP(clk), .Q(
        \filter_0/reg_i_13[15] ) );
  dff_sg \filter_0/reg_i_13_reg[16]  ( .D(\filter_0/n9356 ), .CP(clk), .Q(
        \filter_0/reg_i_13[16] ) );
  dff_sg \filter_0/reg_i_13_reg[17]  ( .D(\filter_0/n9355 ), .CP(clk), .Q(
        \filter_0/reg_i_13[17] ) );
  dff_sg \filter_0/reg_i_13_reg[18]  ( .D(\filter_0/n9354 ), .CP(clk), .Q(
        \filter_0/reg_i_13[18] ) );
  dff_sg \filter_0/reg_i_13_reg[19]  ( .D(\filter_0/n9353 ), .CP(clk), .Q(
        \filter_0/reg_i_13[19] ) );
  dff_sg \filter_0/reg_i_14_reg[0]  ( .D(\filter_0/n9352 ), .CP(clk), .Q(
        \filter_0/reg_i_14[0] ) );
  dff_sg \filter_0/reg_i_14_reg[1]  ( .D(\filter_0/n9351 ), .CP(clk), .Q(
        \filter_0/reg_i_14[1] ) );
  dff_sg \filter_0/reg_i_14_reg[2]  ( .D(\filter_0/n9350 ), .CP(clk), .Q(
        \filter_0/reg_i_14[2] ) );
  dff_sg \filter_0/reg_i_14_reg[3]  ( .D(\filter_0/n9349 ), .CP(clk), .Q(
        \filter_0/reg_i_14[3] ) );
  dff_sg \filter_0/reg_i_14_reg[4]  ( .D(\filter_0/n9348 ), .CP(clk), .Q(
        \filter_0/reg_i_14[4] ) );
  dff_sg \filter_0/reg_i_14_reg[5]  ( .D(\filter_0/n9347 ), .CP(clk), .Q(
        \filter_0/reg_i_14[5] ) );
  dff_sg \filter_0/reg_i_14_reg[6]  ( .D(\filter_0/n9346 ), .CP(clk), .Q(
        \filter_0/reg_i_14[6] ) );
  dff_sg \filter_0/reg_i_14_reg[7]  ( .D(\filter_0/n9345 ), .CP(clk), .Q(
        \filter_0/reg_i_14[7] ) );
  dff_sg \filter_0/reg_i_14_reg[8]  ( .D(\filter_0/n9344 ), .CP(clk), .Q(
        \filter_0/reg_i_14[8] ) );
  dff_sg \filter_0/reg_i_14_reg[9]  ( .D(\filter_0/n9343 ), .CP(clk), .Q(
        \filter_0/reg_i_14[9] ) );
  dff_sg \filter_0/reg_i_14_reg[10]  ( .D(\filter_0/n9342 ), .CP(clk), .Q(
        \filter_0/reg_i_14[10] ) );
  dff_sg \filter_0/reg_i_14_reg[11]  ( .D(\filter_0/n9341 ), .CP(clk), .Q(
        \filter_0/reg_i_14[11] ) );
  dff_sg \filter_0/reg_i_14_reg[12]  ( .D(\filter_0/n9340 ), .CP(clk), .Q(
        \filter_0/reg_i_14[12] ) );
  dff_sg \filter_0/reg_i_14_reg[13]  ( .D(\filter_0/n9339 ), .CP(clk), .Q(
        \filter_0/reg_i_14[13] ) );
  dff_sg \filter_0/reg_i_14_reg[14]  ( .D(\filter_0/n9338 ), .CP(clk), .Q(
        \filter_0/reg_i_14[14] ) );
  dff_sg \filter_0/reg_i_14_reg[15]  ( .D(\filter_0/n9337 ), .CP(clk), .Q(
        \filter_0/reg_i_14[15] ) );
  dff_sg \filter_0/reg_i_14_reg[16]  ( .D(\filter_0/n9336 ), .CP(clk), .Q(
        \filter_0/reg_i_14[16] ) );
  dff_sg \filter_0/reg_i_14_reg[17]  ( .D(\filter_0/n9335 ), .CP(clk), .Q(
        \filter_0/reg_i_14[17] ) );
  dff_sg \filter_0/reg_i_14_reg[18]  ( .D(\filter_0/n9334 ), .CP(clk), .Q(
        \filter_0/reg_i_14[18] ) );
  dff_sg \filter_0/reg_i_14_reg[19]  ( .D(\filter_0/n9333 ), .CP(clk), .Q(
        \filter_0/reg_i_14[19] ) );
  dff_sg \filter_0/reg_i_15_reg[0]  ( .D(\filter_0/n9332 ), .CP(clk), .Q(
        \filter_0/reg_i_15[0] ) );
  dff_sg \filter_0/reg_i_15_reg[1]  ( .D(\filter_0/n9331 ), .CP(clk), .Q(
        \filter_0/reg_i_15[1] ) );
  dff_sg \filter_0/reg_i_15_reg[2]  ( .D(\filter_0/n9330 ), .CP(clk), .Q(
        \filter_0/reg_i_15[2] ) );
  dff_sg \filter_0/reg_i_15_reg[3]  ( .D(\filter_0/n9329 ), .CP(clk), .Q(
        \filter_0/reg_i_15[3] ) );
  dff_sg \filter_0/reg_i_15_reg[4]  ( .D(\filter_0/n9328 ), .CP(clk), .Q(
        \filter_0/reg_i_15[4] ) );
  dff_sg \filter_0/reg_i_15_reg[5]  ( .D(\filter_0/n9327 ), .CP(clk), .Q(
        \filter_0/reg_i_15[5] ) );
  dff_sg \filter_0/reg_i_15_reg[6]  ( .D(\filter_0/n9326 ), .CP(clk), .Q(
        \filter_0/reg_i_15[6] ) );
  dff_sg \filter_0/reg_i_15_reg[7]  ( .D(\filter_0/n9325 ), .CP(clk), .Q(
        \filter_0/reg_i_15[7] ) );
  dff_sg \filter_0/reg_i_15_reg[8]  ( .D(\filter_0/n9324 ), .CP(clk), .Q(
        \filter_0/reg_i_15[8] ) );
  dff_sg \filter_0/reg_i_15_reg[9]  ( .D(\filter_0/n9323 ), .CP(clk), .Q(
        \filter_0/reg_i_15[9] ) );
  dff_sg \filter_0/reg_i_15_reg[10]  ( .D(\filter_0/n9322 ), .CP(clk), .Q(
        \filter_0/reg_i_15[10] ) );
  dff_sg \filter_0/reg_i_15_reg[11]  ( .D(\filter_0/n9321 ), .CP(clk), .Q(
        \filter_0/reg_i_15[11] ) );
  dff_sg \filter_0/reg_i_15_reg[12]  ( .D(\filter_0/n9320 ), .CP(clk), .Q(
        \filter_0/reg_i_15[12] ) );
  dff_sg \filter_0/reg_i_15_reg[13]  ( .D(\filter_0/n9319 ), .CP(clk), .Q(
        \filter_0/reg_i_15[13] ) );
  dff_sg \filter_0/reg_i_15_reg[14]  ( .D(\filter_0/n9318 ), .CP(clk), .Q(
        \filter_0/reg_i_15[14] ) );
  dff_sg \filter_0/reg_i_15_reg[15]  ( .D(\filter_0/n9317 ), .CP(clk), .Q(
        \filter_0/reg_i_15[15] ) );
  dff_sg \filter_0/reg_i_15_reg[16]  ( .D(\filter_0/n9316 ), .CP(clk), .Q(
        \filter_0/reg_i_15[16] ) );
  dff_sg \filter_0/reg_i_15_reg[17]  ( .D(\filter_0/n9315 ), .CP(clk), .Q(
        \filter_0/reg_i_15[17] ) );
  dff_sg \filter_0/reg_i_15_reg[18]  ( .D(\filter_0/n9314 ), .CP(clk), .Q(
        \filter_0/reg_i_15[18] ) );
  dff_sg \filter_0/reg_i_15_reg[19]  ( .D(\filter_0/n9313 ), .CP(clk), .Q(
        \filter_0/reg_i_15[19] ) );
  dff_sg \filter_0/reg_w_0_reg[0]  ( .D(\filter_0/n9312 ), .CP(clk), .Q(
        \filter_0/reg_w_0[0] ) );
  dff_sg \filter_0/reg_w_0_reg[1]  ( .D(\filter_0/n9311 ), .CP(clk), .Q(
        \filter_0/reg_w_0[1] ) );
  dff_sg \filter_0/reg_w_0_reg[2]  ( .D(\filter_0/n9310 ), .CP(clk), .Q(
        \filter_0/reg_w_0[2] ) );
  dff_sg \filter_0/reg_w_0_reg[3]  ( .D(\filter_0/n9309 ), .CP(clk), .Q(
        \filter_0/reg_w_0[3] ) );
  dff_sg \filter_0/reg_w_0_reg[4]  ( .D(\filter_0/n9308 ), .CP(clk), .Q(
        \filter_0/reg_w_0[4] ) );
  dff_sg \filter_0/reg_w_0_reg[5]  ( .D(\filter_0/n9307 ), .CP(clk), .Q(
        \filter_0/reg_w_0[5] ) );
  dff_sg \filter_0/reg_w_0_reg[6]  ( .D(\filter_0/n9306 ), .CP(clk), .Q(
        \filter_0/reg_w_0[6] ) );
  dff_sg \filter_0/reg_w_0_reg[7]  ( .D(\filter_0/n9305 ), .CP(clk), .Q(
        \filter_0/reg_w_0[7] ) );
  dff_sg \filter_0/reg_w_0_reg[8]  ( .D(\filter_0/n9304 ), .CP(clk), .Q(
        \filter_0/reg_w_0[8] ) );
  dff_sg \filter_0/reg_w_0_reg[9]  ( .D(\filter_0/n9303 ), .CP(clk), .Q(
        \filter_0/reg_w_0[9] ) );
  dff_sg \filter_0/reg_w_0_reg[10]  ( .D(\filter_0/n9302 ), .CP(clk), .Q(
        \filter_0/reg_w_0[10] ) );
  dff_sg \filter_0/reg_w_0_reg[11]  ( .D(\filter_0/n9301 ), .CP(clk), .Q(
        \filter_0/reg_w_0[11] ) );
  dff_sg \filter_0/reg_w_0_reg[12]  ( .D(\filter_0/n9300 ), .CP(clk), .Q(
        \filter_0/reg_w_0[12] ) );
  dff_sg \filter_0/reg_w_0_reg[13]  ( .D(\filter_0/n9299 ), .CP(clk), .Q(
        \filter_0/reg_w_0[13] ) );
  dff_sg \filter_0/reg_w_0_reg[14]  ( .D(\filter_0/n9298 ), .CP(clk), .Q(
        \filter_0/reg_w_0[14] ) );
  dff_sg \filter_0/reg_w_0_reg[15]  ( .D(\filter_0/n9297 ), .CP(clk), .Q(
        \filter_0/reg_w_0[15] ) );
  dff_sg \filter_0/reg_w_0_reg[16]  ( .D(\filter_0/n9296 ), .CP(clk), .Q(
        \filter_0/reg_w_0[16] ) );
  dff_sg \filter_0/reg_w_0_reg[17]  ( .D(\filter_0/n9295 ), .CP(clk), .Q(
        \filter_0/reg_w_0[17] ) );
  dff_sg \filter_0/reg_w_0_reg[18]  ( .D(\filter_0/n9294 ), .CP(clk), .Q(
        \filter_0/reg_w_0[18] ) );
  dff_sg \filter_0/reg_w_0_reg[19]  ( .D(\filter_0/n9293 ), .CP(clk), .Q(
        \filter_0/reg_w_0[19] ) );
  dff_sg \filter_0/reg_w_1_reg[0]  ( .D(\filter_0/n9292 ), .CP(clk), .Q(
        \filter_0/reg_w_1[0] ) );
  dff_sg \filter_0/reg_w_1_reg[1]  ( .D(\filter_0/n9291 ), .CP(clk), .Q(
        \filter_0/reg_w_1[1] ) );
  dff_sg \filter_0/reg_w_1_reg[2]  ( .D(\filter_0/n9290 ), .CP(clk), .Q(
        \filter_0/reg_w_1[2] ) );
  dff_sg \filter_0/reg_w_1_reg[3]  ( .D(\filter_0/n9289 ), .CP(clk), .Q(
        \filter_0/reg_w_1[3] ) );
  dff_sg \filter_0/reg_w_1_reg[4]  ( .D(\filter_0/n9288 ), .CP(clk), .Q(
        \filter_0/reg_w_1[4] ) );
  dff_sg \filter_0/reg_w_1_reg[5]  ( .D(\filter_0/n9287 ), .CP(clk), .Q(
        \filter_0/reg_w_1[5] ) );
  dff_sg \filter_0/reg_w_1_reg[6]  ( .D(\filter_0/n9286 ), .CP(clk), .Q(
        \filter_0/reg_w_1[6] ) );
  dff_sg \filter_0/reg_w_1_reg[7]  ( .D(\filter_0/n9285 ), .CP(clk), .Q(
        \filter_0/reg_w_1[7] ) );
  dff_sg \filter_0/reg_w_1_reg[8]  ( .D(\filter_0/n9284 ), .CP(clk), .Q(
        \filter_0/reg_w_1[8] ) );
  dff_sg \filter_0/reg_w_1_reg[9]  ( .D(\filter_0/n9283 ), .CP(clk), .Q(
        \filter_0/reg_w_1[9] ) );
  dff_sg \filter_0/reg_w_1_reg[10]  ( .D(\filter_0/n9282 ), .CP(clk), .Q(
        \filter_0/reg_w_1[10] ) );
  dff_sg \filter_0/reg_w_1_reg[11]  ( .D(\filter_0/n9281 ), .CP(clk), .Q(
        \filter_0/reg_w_1[11] ) );
  dff_sg \filter_0/reg_w_1_reg[12]  ( .D(\filter_0/n9280 ), .CP(clk), .Q(
        \filter_0/reg_w_1[12] ) );
  dff_sg \filter_0/reg_w_1_reg[13]  ( .D(\filter_0/n9279 ), .CP(clk), .Q(
        \filter_0/reg_w_1[13] ) );
  dff_sg \filter_0/reg_w_1_reg[14]  ( .D(\filter_0/n9278 ), .CP(clk), .Q(
        \filter_0/reg_w_1[14] ) );
  dff_sg \filter_0/reg_w_1_reg[15]  ( .D(\filter_0/n9277 ), .CP(clk), .Q(
        \filter_0/reg_w_1[15] ) );
  dff_sg \filter_0/reg_w_1_reg[16]  ( .D(\filter_0/n9276 ), .CP(clk), .Q(
        \filter_0/reg_w_1[16] ) );
  dff_sg \filter_0/reg_w_1_reg[17]  ( .D(\filter_0/n9275 ), .CP(clk), .Q(
        \filter_0/reg_w_1[17] ) );
  dff_sg \filter_0/reg_w_1_reg[18]  ( .D(\filter_0/n9274 ), .CP(clk), .Q(
        \filter_0/reg_w_1[18] ) );
  dff_sg \filter_0/reg_w_1_reg[19]  ( .D(\filter_0/n9273 ), .CP(clk), .Q(
        \filter_0/reg_w_1[19] ) );
  dff_sg \filter_0/reg_w_2_reg[0]  ( .D(\filter_0/n9272 ), .CP(clk), .Q(
        \filter_0/reg_w_2[0] ) );
  dff_sg \filter_0/reg_w_2_reg[1]  ( .D(\filter_0/n9271 ), .CP(clk), .Q(
        \filter_0/reg_w_2[1] ) );
  dff_sg \filter_0/reg_w_2_reg[2]  ( .D(\filter_0/n9270 ), .CP(clk), .Q(
        \filter_0/reg_w_2[2] ) );
  dff_sg \filter_0/reg_w_2_reg[3]  ( .D(\filter_0/n9269 ), .CP(clk), .Q(
        \filter_0/reg_w_2[3] ) );
  dff_sg \filter_0/reg_w_2_reg[4]  ( .D(\filter_0/n9268 ), .CP(clk), .Q(
        \filter_0/reg_w_2[4] ) );
  dff_sg \filter_0/reg_w_2_reg[5]  ( .D(\filter_0/n9267 ), .CP(clk), .Q(
        \filter_0/reg_w_2[5] ) );
  dff_sg \filter_0/reg_w_2_reg[6]  ( .D(\filter_0/n9266 ), .CP(clk), .Q(
        \filter_0/reg_w_2[6] ) );
  dff_sg \filter_0/reg_w_2_reg[7]  ( .D(\filter_0/n9265 ), .CP(clk), .Q(
        \filter_0/reg_w_2[7] ) );
  dff_sg \filter_0/reg_w_2_reg[8]  ( .D(\filter_0/n9264 ), .CP(clk), .Q(
        \filter_0/reg_w_2[8] ) );
  dff_sg \filter_0/reg_w_2_reg[9]  ( .D(\filter_0/n9263 ), .CP(clk), .Q(
        \filter_0/reg_w_2[9] ) );
  dff_sg \filter_0/reg_w_2_reg[10]  ( .D(\filter_0/n9262 ), .CP(clk), .Q(
        \filter_0/reg_w_2[10] ) );
  dff_sg \filter_0/reg_w_2_reg[11]  ( .D(\filter_0/n9261 ), .CP(clk), .Q(
        \filter_0/reg_w_2[11] ) );
  dff_sg \filter_0/reg_w_2_reg[12]  ( .D(\filter_0/n9260 ), .CP(clk), .Q(
        \filter_0/reg_w_2[12] ) );
  dff_sg \filter_0/reg_w_2_reg[13]  ( .D(\filter_0/n9259 ), .CP(clk), .Q(
        \filter_0/reg_w_2[13] ) );
  dff_sg \filter_0/reg_w_2_reg[14]  ( .D(\filter_0/n9258 ), .CP(clk), .Q(
        \filter_0/reg_w_2[14] ) );
  dff_sg \filter_0/reg_w_2_reg[15]  ( .D(\filter_0/n9257 ), .CP(clk), .Q(
        \filter_0/reg_w_2[15] ) );
  dff_sg \filter_0/reg_w_2_reg[16]  ( .D(\filter_0/n9256 ), .CP(clk), .Q(
        \filter_0/reg_w_2[16] ) );
  dff_sg \filter_0/reg_w_2_reg[17]  ( .D(\filter_0/n9255 ), .CP(clk), .Q(
        \filter_0/reg_w_2[17] ) );
  dff_sg \filter_0/reg_w_2_reg[18]  ( .D(\filter_0/n9254 ), .CP(clk), .Q(
        \filter_0/reg_w_2[18] ) );
  dff_sg \filter_0/reg_w_2_reg[19]  ( .D(\filter_0/n9253 ), .CP(clk), .Q(
        \filter_0/reg_w_2[19] ) );
  dff_sg \filter_0/reg_w_3_reg[0]  ( .D(\filter_0/n9252 ), .CP(clk), .Q(
        \filter_0/reg_w_3[0] ) );
  dff_sg \filter_0/reg_w_3_reg[1]  ( .D(\filter_0/n9251 ), .CP(clk), .Q(
        \filter_0/reg_w_3[1] ) );
  dff_sg \filter_0/reg_w_3_reg[2]  ( .D(\filter_0/n9250 ), .CP(clk), .Q(
        \filter_0/reg_w_3[2] ) );
  dff_sg \filter_0/reg_w_3_reg[3]  ( .D(\filter_0/n9249 ), .CP(clk), .Q(
        \filter_0/reg_w_3[3] ) );
  dff_sg \filter_0/reg_w_3_reg[4]  ( .D(\filter_0/n9248 ), .CP(clk), .Q(
        \filter_0/reg_w_3[4] ) );
  dff_sg \filter_0/reg_w_3_reg[5]  ( .D(\filter_0/n9247 ), .CP(clk), .Q(
        \filter_0/reg_w_3[5] ) );
  dff_sg \filter_0/reg_w_3_reg[6]  ( .D(\filter_0/n9246 ), .CP(clk), .Q(
        \filter_0/reg_w_3[6] ) );
  dff_sg \filter_0/reg_w_3_reg[7]  ( .D(\filter_0/n9245 ), .CP(clk), .Q(
        \filter_0/reg_w_3[7] ) );
  dff_sg \filter_0/reg_w_3_reg[8]  ( .D(\filter_0/n9244 ), .CP(clk), .Q(
        \filter_0/reg_w_3[8] ) );
  dff_sg \filter_0/reg_w_3_reg[9]  ( .D(\filter_0/n9243 ), .CP(clk), .Q(
        \filter_0/reg_w_3[9] ) );
  dff_sg \filter_0/reg_w_3_reg[10]  ( .D(\filter_0/n9242 ), .CP(clk), .Q(
        \filter_0/reg_w_3[10] ) );
  dff_sg \filter_0/reg_w_3_reg[11]  ( .D(\filter_0/n9241 ), .CP(clk), .Q(
        \filter_0/reg_w_3[11] ) );
  dff_sg \filter_0/reg_w_3_reg[12]  ( .D(\filter_0/n9240 ), .CP(clk), .Q(
        \filter_0/reg_w_3[12] ) );
  dff_sg \filter_0/reg_w_3_reg[13]  ( .D(\filter_0/n9239 ), .CP(clk), .Q(
        \filter_0/reg_w_3[13] ) );
  dff_sg \filter_0/reg_w_3_reg[14]  ( .D(\filter_0/n9238 ), .CP(clk), .Q(
        \filter_0/reg_w_3[14] ) );
  dff_sg \filter_0/reg_w_3_reg[15]  ( .D(\filter_0/n9237 ), .CP(clk), .Q(
        \filter_0/reg_w_3[15] ) );
  dff_sg \filter_0/reg_w_3_reg[16]  ( .D(\filter_0/n9236 ), .CP(clk), .Q(
        \filter_0/reg_w_3[16] ) );
  dff_sg \filter_0/reg_w_3_reg[17]  ( .D(\filter_0/n9235 ), .CP(clk), .Q(
        \filter_0/reg_w_3[17] ) );
  dff_sg \filter_0/reg_w_3_reg[18]  ( .D(\filter_0/n9234 ), .CP(clk), .Q(
        \filter_0/reg_w_3[18] ) );
  dff_sg \filter_0/reg_w_3_reg[19]  ( .D(\filter_0/n9233 ), .CP(clk), .Q(
        \filter_0/reg_w_3[19] ) );
  dff_sg \filter_0/reg_w_4_reg[0]  ( .D(\filter_0/n9232 ), .CP(clk), .Q(
        \filter_0/reg_w_4[0] ) );
  dff_sg \filter_0/reg_w_4_reg[1]  ( .D(\filter_0/n9231 ), .CP(clk), .Q(
        \filter_0/reg_w_4[1] ) );
  dff_sg \filter_0/reg_w_4_reg[2]  ( .D(\filter_0/n9230 ), .CP(clk), .Q(
        \filter_0/reg_w_4[2] ) );
  dff_sg \filter_0/reg_w_4_reg[3]  ( .D(\filter_0/n9229 ), .CP(clk), .Q(
        \filter_0/reg_w_4[3] ) );
  dff_sg \filter_0/reg_w_4_reg[4]  ( .D(\filter_0/n9228 ), .CP(clk), .Q(
        \filter_0/reg_w_4[4] ) );
  dff_sg \filter_0/reg_w_4_reg[5]  ( .D(\filter_0/n9227 ), .CP(clk), .Q(
        \filter_0/reg_w_4[5] ) );
  dff_sg \filter_0/reg_w_4_reg[6]  ( .D(\filter_0/n9226 ), .CP(clk), .Q(
        \filter_0/reg_w_4[6] ) );
  dff_sg \filter_0/reg_w_4_reg[7]  ( .D(\filter_0/n9225 ), .CP(clk), .Q(
        \filter_0/reg_w_4[7] ) );
  dff_sg \filter_0/reg_w_4_reg[8]  ( .D(\filter_0/n9224 ), .CP(clk), .Q(
        \filter_0/reg_w_4[8] ) );
  dff_sg \filter_0/reg_w_4_reg[9]  ( .D(\filter_0/n9223 ), .CP(clk), .Q(
        \filter_0/reg_w_4[9] ) );
  dff_sg \filter_0/reg_w_4_reg[10]  ( .D(\filter_0/n9222 ), .CP(clk), .Q(
        \filter_0/reg_w_4[10] ) );
  dff_sg \filter_0/reg_w_4_reg[11]  ( .D(\filter_0/n9221 ), .CP(clk), .Q(
        \filter_0/reg_w_4[11] ) );
  dff_sg \filter_0/reg_w_4_reg[12]  ( .D(\filter_0/n9220 ), .CP(clk), .Q(
        \filter_0/reg_w_4[12] ) );
  dff_sg \filter_0/reg_w_4_reg[13]  ( .D(\filter_0/n9219 ), .CP(clk), .Q(
        \filter_0/reg_w_4[13] ) );
  dff_sg \filter_0/reg_w_4_reg[14]  ( .D(\filter_0/n9218 ), .CP(clk), .Q(
        \filter_0/reg_w_4[14] ) );
  dff_sg \filter_0/reg_w_4_reg[15]  ( .D(\filter_0/n9217 ), .CP(clk), .Q(
        \filter_0/reg_w_4[15] ) );
  dff_sg \filter_0/reg_w_4_reg[16]  ( .D(\filter_0/n9216 ), .CP(clk), .Q(
        \filter_0/reg_w_4[16] ) );
  dff_sg \filter_0/reg_w_4_reg[17]  ( .D(\filter_0/n9215 ), .CP(clk), .Q(
        \filter_0/reg_w_4[17] ) );
  dff_sg \filter_0/reg_w_4_reg[18]  ( .D(\filter_0/n9214 ), .CP(clk), .Q(
        \filter_0/reg_w_4[18] ) );
  dff_sg \filter_0/reg_w_4_reg[19]  ( .D(\filter_0/n9213 ), .CP(clk), .Q(
        \filter_0/reg_w_4[19] ) );
  dff_sg \filter_0/reg_w_5_reg[0]  ( .D(\filter_0/n9212 ), .CP(clk), .Q(
        \filter_0/reg_w_5[0] ) );
  dff_sg \filter_0/reg_w_5_reg[1]  ( .D(\filter_0/n9211 ), .CP(clk), .Q(
        \filter_0/reg_w_5[1] ) );
  dff_sg \filter_0/reg_w_5_reg[2]  ( .D(\filter_0/n9210 ), .CP(clk), .Q(
        \filter_0/reg_w_5[2] ) );
  dff_sg \filter_0/reg_w_5_reg[3]  ( .D(\filter_0/n9209 ), .CP(clk), .Q(
        \filter_0/reg_w_5[3] ) );
  dff_sg \filter_0/reg_w_5_reg[4]  ( .D(\filter_0/n9208 ), .CP(clk), .Q(
        \filter_0/reg_w_5[4] ) );
  dff_sg \filter_0/reg_w_5_reg[5]  ( .D(\filter_0/n9207 ), .CP(clk), .Q(
        \filter_0/reg_w_5[5] ) );
  dff_sg \filter_0/reg_w_5_reg[6]  ( .D(\filter_0/n9206 ), .CP(clk), .Q(
        \filter_0/reg_w_5[6] ) );
  dff_sg \filter_0/reg_w_5_reg[7]  ( .D(\filter_0/n9205 ), .CP(clk), .Q(
        \filter_0/reg_w_5[7] ) );
  dff_sg \filter_0/reg_w_5_reg[8]  ( .D(\filter_0/n9204 ), .CP(clk), .Q(
        \filter_0/reg_w_5[8] ) );
  dff_sg \filter_0/reg_w_5_reg[9]  ( .D(\filter_0/n9203 ), .CP(clk), .Q(
        \filter_0/reg_w_5[9] ) );
  dff_sg \filter_0/reg_w_5_reg[10]  ( .D(\filter_0/n9202 ), .CP(clk), .Q(
        \filter_0/reg_w_5[10] ) );
  dff_sg \filter_0/reg_w_5_reg[11]  ( .D(\filter_0/n9201 ), .CP(clk), .Q(
        \filter_0/reg_w_5[11] ) );
  dff_sg \filter_0/reg_w_5_reg[12]  ( .D(\filter_0/n9200 ), .CP(clk), .Q(
        \filter_0/reg_w_5[12] ) );
  dff_sg \filter_0/reg_w_5_reg[13]  ( .D(\filter_0/n9199 ), .CP(clk), .Q(
        \filter_0/reg_w_5[13] ) );
  dff_sg \filter_0/reg_w_5_reg[14]  ( .D(\filter_0/n9198 ), .CP(clk), .Q(
        \filter_0/reg_w_5[14] ) );
  dff_sg \filter_0/reg_w_5_reg[15]  ( .D(\filter_0/n9197 ), .CP(clk), .Q(
        \filter_0/reg_w_5[15] ) );
  dff_sg \filter_0/reg_w_5_reg[16]  ( .D(\filter_0/n9196 ), .CP(clk), .Q(
        \filter_0/reg_w_5[16] ) );
  dff_sg \filter_0/reg_w_5_reg[17]  ( .D(\filter_0/n9195 ), .CP(clk), .Q(
        \filter_0/reg_w_5[17] ) );
  dff_sg \filter_0/reg_w_5_reg[18]  ( .D(\filter_0/n9194 ), .CP(clk), .Q(
        \filter_0/reg_w_5[18] ) );
  dff_sg \filter_0/reg_w_5_reg[19]  ( .D(\filter_0/n9193 ), .CP(clk), .Q(
        \filter_0/reg_w_5[19] ) );
  dff_sg \filter_0/reg_w_6_reg[0]  ( .D(\filter_0/n9192 ), .CP(clk), .Q(
        \filter_0/reg_w_6[0] ) );
  dff_sg \filter_0/reg_w_6_reg[1]  ( .D(\filter_0/n9191 ), .CP(clk), .Q(
        \filter_0/reg_w_6[1] ) );
  dff_sg \filter_0/reg_w_6_reg[2]  ( .D(\filter_0/n9190 ), .CP(clk), .Q(
        \filter_0/reg_w_6[2] ) );
  dff_sg \filter_0/reg_w_6_reg[3]  ( .D(\filter_0/n9189 ), .CP(clk), .Q(
        \filter_0/reg_w_6[3] ) );
  dff_sg \filter_0/reg_w_6_reg[4]  ( .D(\filter_0/n9188 ), .CP(clk), .Q(
        \filter_0/reg_w_6[4] ) );
  dff_sg \filter_0/reg_w_6_reg[5]  ( .D(\filter_0/n9187 ), .CP(clk), .Q(
        \filter_0/reg_w_6[5] ) );
  dff_sg \filter_0/reg_w_6_reg[6]  ( .D(\filter_0/n9186 ), .CP(clk), .Q(
        \filter_0/reg_w_6[6] ) );
  dff_sg \filter_0/reg_w_6_reg[7]  ( .D(\filter_0/n9185 ), .CP(clk), .Q(
        \filter_0/reg_w_6[7] ) );
  dff_sg \filter_0/reg_w_6_reg[8]  ( .D(\filter_0/n9184 ), .CP(clk), .Q(
        \filter_0/reg_w_6[8] ) );
  dff_sg \filter_0/reg_w_6_reg[9]  ( .D(\filter_0/n9183 ), .CP(clk), .Q(
        \filter_0/reg_w_6[9] ) );
  dff_sg \filter_0/reg_w_6_reg[10]  ( .D(\filter_0/n9182 ), .CP(clk), .Q(
        \filter_0/reg_w_6[10] ) );
  dff_sg \filter_0/reg_w_6_reg[11]  ( .D(\filter_0/n9181 ), .CP(clk), .Q(
        \filter_0/reg_w_6[11] ) );
  dff_sg \filter_0/reg_w_6_reg[12]  ( .D(\filter_0/n9180 ), .CP(clk), .Q(
        \filter_0/reg_w_6[12] ) );
  dff_sg \filter_0/reg_w_6_reg[13]  ( .D(\filter_0/n9179 ), .CP(clk), .Q(
        \filter_0/reg_w_6[13] ) );
  dff_sg \filter_0/reg_w_6_reg[14]  ( .D(\filter_0/n9178 ), .CP(clk), .Q(
        \filter_0/reg_w_6[14] ) );
  dff_sg \filter_0/reg_w_6_reg[15]  ( .D(\filter_0/n9177 ), .CP(clk), .Q(
        \filter_0/reg_w_6[15] ) );
  dff_sg \filter_0/reg_w_6_reg[16]  ( .D(\filter_0/n9176 ), .CP(clk), .Q(
        \filter_0/reg_w_6[16] ) );
  dff_sg \filter_0/reg_w_6_reg[17]  ( .D(\filter_0/n9175 ), .CP(clk), .Q(
        \filter_0/reg_w_6[17] ) );
  dff_sg \filter_0/reg_w_6_reg[18]  ( .D(\filter_0/n9174 ), .CP(clk), .Q(
        \filter_0/reg_w_6[18] ) );
  dff_sg \filter_0/reg_w_6_reg[19]  ( .D(\filter_0/n9173 ), .CP(clk), .Q(
        \filter_0/reg_w_6[19] ) );
  dff_sg \filter_0/reg_w_7_reg[0]  ( .D(\filter_0/n9172 ), .CP(clk), .Q(
        \filter_0/reg_w_7[0] ) );
  dff_sg \filter_0/reg_w_7_reg[1]  ( .D(\filter_0/n9171 ), .CP(clk), .Q(
        \filter_0/reg_w_7[1] ) );
  dff_sg \filter_0/reg_w_7_reg[2]  ( .D(\filter_0/n9170 ), .CP(clk), .Q(
        \filter_0/reg_w_7[2] ) );
  dff_sg \filter_0/reg_w_7_reg[3]  ( .D(\filter_0/n9169 ), .CP(clk), .Q(
        \filter_0/reg_w_7[3] ) );
  dff_sg \filter_0/reg_w_7_reg[4]  ( .D(\filter_0/n9168 ), .CP(clk), .Q(
        \filter_0/reg_w_7[4] ) );
  dff_sg \filter_0/reg_w_7_reg[5]  ( .D(\filter_0/n9167 ), .CP(clk), .Q(
        \filter_0/reg_w_7[5] ) );
  dff_sg \filter_0/reg_w_7_reg[6]  ( .D(\filter_0/n9166 ), .CP(clk), .Q(
        \filter_0/reg_w_7[6] ) );
  dff_sg \filter_0/reg_w_7_reg[7]  ( .D(\filter_0/n9165 ), .CP(clk), .Q(
        \filter_0/reg_w_7[7] ) );
  dff_sg \filter_0/reg_w_7_reg[8]  ( .D(\filter_0/n9164 ), .CP(clk), .Q(
        \filter_0/reg_w_7[8] ) );
  dff_sg \filter_0/reg_w_7_reg[9]  ( .D(\filter_0/n9163 ), .CP(clk), .Q(
        \filter_0/reg_w_7[9] ) );
  dff_sg \filter_0/reg_w_7_reg[10]  ( .D(\filter_0/n9162 ), .CP(clk), .Q(
        \filter_0/reg_w_7[10] ) );
  dff_sg \filter_0/reg_w_7_reg[11]  ( .D(\filter_0/n9161 ), .CP(clk), .Q(
        \filter_0/reg_w_7[11] ) );
  dff_sg \filter_0/reg_w_7_reg[12]  ( .D(\filter_0/n9160 ), .CP(clk), .Q(
        \filter_0/reg_w_7[12] ) );
  dff_sg \filter_0/reg_w_7_reg[13]  ( .D(\filter_0/n9159 ), .CP(clk), .Q(
        \filter_0/reg_w_7[13] ) );
  dff_sg \filter_0/reg_w_7_reg[14]  ( .D(\filter_0/n9158 ), .CP(clk), .Q(
        \filter_0/reg_w_7[14] ) );
  dff_sg \filter_0/reg_w_7_reg[15]  ( .D(\filter_0/n9157 ), .CP(clk), .Q(
        \filter_0/reg_w_7[15] ) );
  dff_sg \filter_0/reg_w_7_reg[16]  ( .D(\filter_0/n9156 ), .CP(clk), .Q(
        \filter_0/reg_w_7[16] ) );
  dff_sg \filter_0/reg_w_7_reg[17]  ( .D(\filter_0/n9155 ), .CP(clk), .Q(
        \filter_0/reg_w_7[17] ) );
  dff_sg \filter_0/reg_w_7_reg[18]  ( .D(\filter_0/n9154 ), .CP(clk), .Q(
        \filter_0/reg_w_7[18] ) );
  dff_sg \filter_0/reg_w_7_reg[19]  ( .D(\filter_0/n9153 ), .CP(clk), .Q(
        \filter_0/reg_w_7[19] ) );
  dff_sg \filter_0/reg_w_8_reg[0]  ( .D(\filter_0/n9152 ), .CP(clk), .Q(
        \filter_0/reg_w_8[0] ) );
  dff_sg \filter_0/reg_w_8_reg[1]  ( .D(\filter_0/n9151 ), .CP(clk), .Q(
        \filter_0/reg_w_8[1] ) );
  dff_sg \filter_0/reg_w_8_reg[2]  ( .D(\filter_0/n9150 ), .CP(clk), .Q(
        \filter_0/reg_w_8[2] ) );
  dff_sg \filter_0/reg_w_8_reg[3]  ( .D(\filter_0/n9149 ), .CP(clk), .Q(
        \filter_0/reg_w_8[3] ) );
  dff_sg \filter_0/reg_w_8_reg[4]  ( .D(\filter_0/n9148 ), .CP(clk), .Q(
        \filter_0/reg_w_8[4] ) );
  dff_sg \filter_0/reg_w_8_reg[5]  ( .D(\filter_0/n9147 ), .CP(clk), .Q(
        \filter_0/reg_w_8[5] ) );
  dff_sg \filter_0/reg_w_8_reg[6]  ( .D(\filter_0/n9146 ), .CP(clk), .Q(
        \filter_0/reg_w_8[6] ) );
  dff_sg \filter_0/reg_w_8_reg[7]  ( .D(\filter_0/n9145 ), .CP(clk), .Q(
        \filter_0/reg_w_8[7] ) );
  dff_sg \filter_0/reg_w_8_reg[8]  ( .D(\filter_0/n9144 ), .CP(clk), .Q(
        \filter_0/reg_w_8[8] ) );
  dff_sg \filter_0/reg_w_8_reg[9]  ( .D(\filter_0/n9143 ), .CP(clk), .Q(
        \filter_0/reg_w_8[9] ) );
  dff_sg \filter_0/reg_w_8_reg[10]  ( .D(\filter_0/n9142 ), .CP(clk), .Q(
        \filter_0/reg_w_8[10] ) );
  dff_sg \filter_0/reg_w_8_reg[11]  ( .D(\filter_0/n9141 ), .CP(clk), .Q(
        \filter_0/reg_w_8[11] ) );
  dff_sg \filter_0/reg_w_8_reg[12]  ( .D(\filter_0/n9140 ), .CP(clk), .Q(
        \filter_0/reg_w_8[12] ) );
  dff_sg \filter_0/reg_w_8_reg[13]  ( .D(\filter_0/n9139 ), .CP(clk), .Q(
        \filter_0/reg_w_8[13] ) );
  dff_sg \filter_0/reg_w_8_reg[14]  ( .D(\filter_0/n9138 ), .CP(clk), .Q(
        \filter_0/reg_w_8[14] ) );
  dff_sg \filter_0/reg_w_8_reg[15]  ( .D(\filter_0/n9137 ), .CP(clk), .Q(
        \filter_0/reg_w_8[15] ) );
  dff_sg \filter_0/reg_w_8_reg[16]  ( .D(\filter_0/n9136 ), .CP(clk), .Q(
        \filter_0/reg_w_8[16] ) );
  dff_sg \filter_0/reg_w_8_reg[17]  ( .D(\filter_0/n9135 ), .CP(clk), .Q(
        \filter_0/reg_w_8[17] ) );
  dff_sg \filter_0/reg_w_8_reg[18]  ( .D(\filter_0/n9134 ), .CP(clk), .Q(
        \filter_0/reg_w_8[18] ) );
  dff_sg \filter_0/reg_w_8_reg[19]  ( .D(\filter_0/n9133 ), .CP(clk), .Q(
        \filter_0/reg_w_8[19] ) );
  dff_sg \filter_0/reg_w_9_reg[0]  ( .D(\filter_0/n9132 ), .CP(clk), .Q(
        \filter_0/reg_w_9[0] ) );
  dff_sg \filter_0/reg_w_9_reg[1]  ( .D(\filter_0/n9131 ), .CP(clk), .Q(
        \filter_0/reg_w_9[1] ) );
  dff_sg \filter_0/reg_w_9_reg[2]  ( .D(\filter_0/n9130 ), .CP(clk), .Q(
        \filter_0/reg_w_9[2] ) );
  dff_sg \filter_0/reg_w_9_reg[3]  ( .D(\filter_0/n9129 ), .CP(clk), .Q(
        \filter_0/reg_w_9[3] ) );
  dff_sg \filter_0/reg_w_9_reg[4]  ( .D(\filter_0/n9128 ), .CP(clk), .Q(
        \filter_0/reg_w_9[4] ) );
  dff_sg \filter_0/reg_w_9_reg[5]  ( .D(\filter_0/n9127 ), .CP(clk), .Q(
        \filter_0/reg_w_9[5] ) );
  dff_sg \filter_0/reg_w_9_reg[6]  ( .D(\filter_0/n9126 ), .CP(clk), .Q(
        \filter_0/reg_w_9[6] ) );
  dff_sg \filter_0/reg_w_9_reg[7]  ( .D(\filter_0/n9125 ), .CP(clk), .Q(
        \filter_0/reg_w_9[7] ) );
  dff_sg \filter_0/reg_w_9_reg[8]  ( .D(\filter_0/n9124 ), .CP(clk), .Q(
        \filter_0/reg_w_9[8] ) );
  dff_sg \filter_0/reg_w_9_reg[9]  ( .D(\filter_0/n9123 ), .CP(clk), .Q(
        \filter_0/reg_w_9[9] ) );
  dff_sg \filter_0/reg_w_9_reg[10]  ( .D(\filter_0/n9122 ), .CP(clk), .Q(
        \filter_0/reg_w_9[10] ) );
  dff_sg \filter_0/reg_w_9_reg[11]  ( .D(\filter_0/n9121 ), .CP(clk), .Q(
        \filter_0/reg_w_9[11] ) );
  dff_sg \filter_0/reg_w_9_reg[12]  ( .D(\filter_0/n9120 ), .CP(clk), .Q(
        \filter_0/reg_w_9[12] ) );
  dff_sg \filter_0/reg_w_9_reg[13]  ( .D(\filter_0/n9119 ), .CP(clk), .Q(
        \filter_0/reg_w_9[13] ) );
  dff_sg \filter_0/reg_w_9_reg[14]  ( .D(\filter_0/n9118 ), .CP(clk), .Q(
        \filter_0/reg_w_9[14] ) );
  dff_sg \filter_0/reg_w_9_reg[15]  ( .D(\filter_0/n9117 ), .CP(clk), .Q(
        \filter_0/reg_w_9[15] ) );
  dff_sg \filter_0/reg_w_9_reg[16]  ( .D(\filter_0/n9116 ), .CP(clk), .Q(
        \filter_0/reg_w_9[16] ) );
  dff_sg \filter_0/reg_w_9_reg[17]  ( .D(\filter_0/n9115 ), .CP(clk), .Q(
        \filter_0/reg_w_9[17] ) );
  dff_sg \filter_0/reg_w_9_reg[18]  ( .D(\filter_0/n9114 ), .CP(clk), .Q(
        \filter_0/reg_w_9[18] ) );
  dff_sg \filter_0/reg_w_9_reg[19]  ( .D(\filter_0/n9113 ), .CP(clk), .Q(
        \filter_0/reg_w_9[19] ) );
  dff_sg \filter_0/reg_w_10_reg[0]  ( .D(\filter_0/n9112 ), .CP(clk), .Q(
        \filter_0/reg_w_10[0] ) );
  dff_sg \filter_0/reg_w_10_reg[1]  ( .D(\filter_0/n9111 ), .CP(clk), .Q(
        \filter_0/reg_w_10[1] ) );
  dff_sg \filter_0/reg_w_10_reg[2]  ( .D(\filter_0/n9110 ), .CP(clk), .Q(
        \filter_0/reg_w_10[2] ) );
  dff_sg \filter_0/reg_w_10_reg[3]  ( .D(\filter_0/n9109 ), .CP(clk), .Q(
        \filter_0/reg_w_10[3] ) );
  dff_sg \filter_0/reg_w_10_reg[4]  ( .D(\filter_0/n9108 ), .CP(clk), .Q(
        \filter_0/reg_w_10[4] ) );
  dff_sg \filter_0/reg_w_10_reg[5]  ( .D(\filter_0/n9107 ), .CP(clk), .Q(
        \filter_0/reg_w_10[5] ) );
  dff_sg \filter_0/reg_w_10_reg[6]  ( .D(\filter_0/n9106 ), .CP(clk), .Q(
        \filter_0/reg_w_10[6] ) );
  dff_sg \filter_0/reg_w_10_reg[7]  ( .D(\filter_0/n9105 ), .CP(clk), .Q(
        \filter_0/reg_w_10[7] ) );
  dff_sg \filter_0/reg_w_10_reg[8]  ( .D(\filter_0/n9104 ), .CP(clk), .Q(
        \filter_0/reg_w_10[8] ) );
  dff_sg \filter_0/reg_w_10_reg[9]  ( .D(\filter_0/n9103 ), .CP(clk), .Q(
        \filter_0/reg_w_10[9] ) );
  dff_sg \filter_0/reg_w_10_reg[10]  ( .D(\filter_0/n9102 ), .CP(clk), .Q(
        \filter_0/reg_w_10[10] ) );
  dff_sg \filter_0/reg_w_10_reg[11]  ( .D(\filter_0/n9101 ), .CP(clk), .Q(
        \filter_0/reg_w_10[11] ) );
  dff_sg \filter_0/reg_w_10_reg[12]  ( .D(\filter_0/n9100 ), .CP(clk), .Q(
        \filter_0/reg_w_10[12] ) );
  dff_sg \filter_0/reg_w_10_reg[13]  ( .D(\filter_0/n9099 ), .CP(clk), .Q(
        \filter_0/reg_w_10[13] ) );
  dff_sg \filter_0/reg_w_10_reg[14]  ( .D(\filter_0/n9098 ), .CP(clk), .Q(
        \filter_0/reg_w_10[14] ) );
  dff_sg \filter_0/reg_w_10_reg[15]  ( .D(\filter_0/n9097 ), .CP(clk), .Q(
        \filter_0/reg_w_10[15] ) );
  dff_sg \filter_0/reg_w_10_reg[16]  ( .D(\filter_0/n9096 ), .CP(clk), .Q(
        \filter_0/reg_w_10[16] ) );
  dff_sg \filter_0/reg_w_10_reg[17]  ( .D(\filter_0/n9095 ), .CP(clk), .Q(
        \filter_0/reg_w_10[17] ) );
  dff_sg \filter_0/reg_w_10_reg[18]  ( .D(\filter_0/n9094 ), .CP(clk), .Q(
        \filter_0/reg_w_10[18] ) );
  dff_sg \filter_0/reg_w_10_reg[19]  ( .D(\filter_0/n9093 ), .CP(clk), .Q(
        \filter_0/reg_w_10[19] ) );
  dff_sg \filter_0/reg_w_11_reg[0]  ( .D(\filter_0/n9092 ), .CP(clk), .Q(
        \filter_0/reg_w_11[0] ) );
  dff_sg \filter_0/reg_w_11_reg[1]  ( .D(\filter_0/n9091 ), .CP(clk), .Q(
        \filter_0/reg_w_11[1] ) );
  dff_sg \filter_0/reg_w_11_reg[2]  ( .D(\filter_0/n9090 ), .CP(clk), .Q(
        \filter_0/reg_w_11[2] ) );
  dff_sg \filter_0/reg_w_11_reg[3]  ( .D(\filter_0/n9089 ), .CP(clk), .Q(
        \filter_0/reg_w_11[3] ) );
  dff_sg \filter_0/reg_w_11_reg[4]  ( .D(\filter_0/n9088 ), .CP(clk), .Q(
        \filter_0/reg_w_11[4] ) );
  dff_sg \filter_0/reg_w_11_reg[5]  ( .D(\filter_0/n9087 ), .CP(clk), .Q(
        \filter_0/reg_w_11[5] ) );
  dff_sg \filter_0/reg_w_11_reg[6]  ( .D(\filter_0/n9086 ), .CP(clk), .Q(
        \filter_0/reg_w_11[6] ) );
  dff_sg \filter_0/reg_w_11_reg[7]  ( .D(\filter_0/n9085 ), .CP(clk), .Q(
        \filter_0/reg_w_11[7] ) );
  dff_sg \filter_0/reg_w_11_reg[8]  ( .D(\filter_0/n9084 ), .CP(clk), .Q(
        \filter_0/reg_w_11[8] ) );
  dff_sg \filter_0/reg_w_11_reg[9]  ( .D(\filter_0/n9083 ), .CP(clk), .Q(
        \filter_0/reg_w_11[9] ) );
  dff_sg \filter_0/reg_w_11_reg[10]  ( .D(\filter_0/n9082 ), .CP(clk), .Q(
        \filter_0/reg_w_11[10] ) );
  dff_sg \filter_0/reg_w_11_reg[11]  ( .D(\filter_0/n9081 ), .CP(clk), .Q(
        \filter_0/reg_w_11[11] ) );
  dff_sg \filter_0/reg_w_11_reg[12]  ( .D(\filter_0/n9080 ), .CP(clk), .Q(
        \filter_0/reg_w_11[12] ) );
  dff_sg \filter_0/reg_w_11_reg[13]  ( .D(\filter_0/n9079 ), .CP(clk), .Q(
        \filter_0/reg_w_11[13] ) );
  dff_sg \filter_0/reg_w_11_reg[14]  ( .D(\filter_0/n9078 ), .CP(clk), .Q(
        \filter_0/reg_w_11[14] ) );
  dff_sg \filter_0/reg_w_11_reg[15]  ( .D(\filter_0/n9077 ), .CP(clk), .Q(
        \filter_0/reg_w_11[15] ) );
  dff_sg \filter_0/reg_w_11_reg[16]  ( .D(\filter_0/n9076 ), .CP(clk), .Q(
        \filter_0/reg_w_11[16] ) );
  dff_sg \filter_0/reg_w_11_reg[17]  ( .D(\filter_0/n9075 ), .CP(clk), .Q(
        \filter_0/reg_w_11[17] ) );
  dff_sg \filter_0/reg_w_11_reg[18]  ( .D(\filter_0/n9074 ), .CP(clk), .Q(
        \filter_0/reg_w_11[18] ) );
  dff_sg \filter_0/reg_w_11_reg[19]  ( .D(\filter_0/n9073 ), .CP(clk), .Q(
        \filter_0/reg_w_11[19] ) );
  dff_sg \filter_0/reg_w_12_reg[0]  ( .D(\filter_0/n9072 ), .CP(clk), .Q(
        \filter_0/reg_w_12[0] ) );
  dff_sg \filter_0/reg_w_12_reg[1]  ( .D(\filter_0/n9071 ), .CP(clk), .Q(
        \filter_0/reg_w_12[1] ) );
  dff_sg \filter_0/reg_w_12_reg[2]  ( .D(\filter_0/n9070 ), .CP(clk), .Q(
        \filter_0/reg_w_12[2] ) );
  dff_sg \filter_0/reg_w_12_reg[3]  ( .D(\filter_0/n9069 ), .CP(clk), .Q(
        \filter_0/reg_w_12[3] ) );
  dff_sg \filter_0/reg_w_12_reg[4]  ( .D(\filter_0/n9068 ), .CP(clk), .Q(
        \filter_0/reg_w_12[4] ) );
  dff_sg \filter_0/reg_w_12_reg[5]  ( .D(\filter_0/n9067 ), .CP(clk), .Q(
        \filter_0/reg_w_12[5] ) );
  dff_sg \filter_0/reg_w_12_reg[6]  ( .D(\filter_0/n9066 ), .CP(clk), .Q(
        \filter_0/reg_w_12[6] ) );
  dff_sg \filter_0/reg_w_12_reg[7]  ( .D(\filter_0/n9065 ), .CP(clk), .Q(
        \filter_0/reg_w_12[7] ) );
  dff_sg \filter_0/reg_w_12_reg[8]  ( .D(\filter_0/n9064 ), .CP(clk), .Q(
        \filter_0/reg_w_12[8] ) );
  dff_sg \filter_0/reg_w_12_reg[9]  ( .D(\filter_0/n9063 ), .CP(clk), .Q(
        \filter_0/reg_w_12[9] ) );
  dff_sg \filter_0/reg_w_12_reg[10]  ( .D(\filter_0/n9062 ), .CP(clk), .Q(
        \filter_0/reg_w_12[10] ) );
  dff_sg \filter_0/reg_w_12_reg[11]  ( .D(\filter_0/n9061 ), .CP(clk), .Q(
        \filter_0/reg_w_12[11] ) );
  dff_sg \filter_0/reg_w_12_reg[12]  ( .D(\filter_0/n9060 ), .CP(clk), .Q(
        \filter_0/reg_w_12[12] ) );
  dff_sg \filter_0/reg_w_12_reg[13]  ( .D(\filter_0/n9059 ), .CP(clk), .Q(
        \filter_0/reg_w_12[13] ) );
  dff_sg \filter_0/reg_w_12_reg[14]  ( .D(\filter_0/n9058 ), .CP(clk), .Q(
        \filter_0/reg_w_12[14] ) );
  dff_sg \filter_0/reg_w_12_reg[15]  ( .D(\filter_0/n9057 ), .CP(clk), .Q(
        \filter_0/reg_w_12[15] ) );
  dff_sg \filter_0/reg_w_12_reg[16]  ( .D(\filter_0/n9056 ), .CP(clk), .Q(
        \filter_0/reg_w_12[16] ) );
  dff_sg \filter_0/reg_w_12_reg[17]  ( .D(\filter_0/n9055 ), .CP(clk), .Q(
        \filter_0/reg_w_12[17] ) );
  dff_sg \filter_0/reg_w_12_reg[18]  ( .D(\filter_0/n9054 ), .CP(clk), .Q(
        \filter_0/reg_w_12[18] ) );
  dff_sg \filter_0/reg_w_12_reg[19]  ( .D(\filter_0/n9053 ), .CP(clk), .Q(
        \filter_0/reg_w_12[19] ) );
  dff_sg \filter_0/reg_w_13_reg[0]  ( .D(\filter_0/n9052 ), .CP(clk), .Q(
        \filter_0/reg_w_13[0] ) );
  dff_sg \filter_0/reg_w_13_reg[1]  ( .D(\filter_0/n9051 ), .CP(clk), .Q(
        \filter_0/reg_w_13[1] ) );
  dff_sg \filter_0/reg_w_13_reg[2]  ( .D(\filter_0/n9050 ), .CP(clk), .Q(
        \filter_0/reg_w_13[2] ) );
  dff_sg \filter_0/reg_w_13_reg[3]  ( .D(\filter_0/n9049 ), .CP(clk), .Q(
        \filter_0/reg_w_13[3] ) );
  dff_sg \filter_0/reg_w_13_reg[4]  ( .D(\filter_0/n9048 ), .CP(clk), .Q(
        \filter_0/reg_w_13[4] ) );
  dff_sg \filter_0/reg_w_13_reg[5]  ( .D(\filter_0/n9047 ), .CP(clk), .Q(
        \filter_0/reg_w_13[5] ) );
  dff_sg \filter_0/reg_w_13_reg[6]  ( .D(\filter_0/n9046 ), .CP(clk), .Q(
        \filter_0/reg_w_13[6] ) );
  dff_sg \filter_0/reg_w_13_reg[7]  ( .D(\filter_0/n9045 ), .CP(clk), .Q(
        \filter_0/reg_w_13[7] ) );
  dff_sg \filter_0/reg_w_13_reg[8]  ( .D(\filter_0/n9044 ), .CP(clk), .Q(
        \filter_0/reg_w_13[8] ) );
  dff_sg \filter_0/reg_w_13_reg[9]  ( .D(\filter_0/n9043 ), .CP(clk), .Q(
        \filter_0/reg_w_13[9] ) );
  dff_sg \filter_0/reg_w_13_reg[10]  ( .D(\filter_0/n9042 ), .CP(clk), .Q(
        \filter_0/reg_w_13[10] ) );
  dff_sg \filter_0/reg_w_13_reg[11]  ( .D(\filter_0/n9041 ), .CP(clk), .Q(
        \filter_0/reg_w_13[11] ) );
  dff_sg \filter_0/reg_w_13_reg[12]  ( .D(\filter_0/n9040 ), .CP(clk), .Q(
        \filter_0/reg_w_13[12] ) );
  dff_sg \filter_0/reg_w_13_reg[13]  ( .D(\filter_0/n9039 ), .CP(clk), .Q(
        \filter_0/reg_w_13[13] ) );
  dff_sg \filter_0/reg_w_13_reg[14]  ( .D(\filter_0/n9038 ), .CP(clk), .Q(
        \filter_0/reg_w_13[14] ) );
  dff_sg \filter_0/reg_w_13_reg[15]  ( .D(\filter_0/n9037 ), .CP(clk), .Q(
        \filter_0/reg_w_13[15] ) );
  dff_sg \filter_0/reg_w_13_reg[16]  ( .D(\filter_0/n9036 ), .CP(clk), .Q(
        \filter_0/reg_w_13[16] ) );
  dff_sg \filter_0/reg_w_13_reg[17]  ( .D(\filter_0/n9035 ), .CP(clk), .Q(
        \filter_0/reg_w_13[17] ) );
  dff_sg \filter_0/reg_w_13_reg[18]  ( .D(\filter_0/n9034 ), .CP(clk), .Q(
        \filter_0/reg_w_13[18] ) );
  dff_sg \filter_0/reg_w_13_reg[19]  ( .D(\filter_0/n9033 ), .CP(clk), .Q(
        \filter_0/reg_w_13[19] ) );
  dff_sg \filter_0/reg_w_14_reg[0]  ( .D(\filter_0/n9032 ), .CP(clk), .Q(
        \filter_0/reg_w_14[0] ) );
  dff_sg \filter_0/reg_w_14_reg[1]  ( .D(\filter_0/n9031 ), .CP(clk), .Q(
        \filter_0/reg_w_14[1] ) );
  dff_sg \filter_0/reg_w_14_reg[2]  ( .D(\filter_0/n9030 ), .CP(clk), .Q(
        \filter_0/reg_w_14[2] ) );
  dff_sg \filter_0/reg_w_14_reg[3]  ( .D(\filter_0/n9029 ), .CP(clk), .Q(
        \filter_0/reg_w_14[3] ) );
  dff_sg \filter_0/reg_w_14_reg[4]  ( .D(\filter_0/n9028 ), .CP(clk), .Q(
        \filter_0/reg_w_14[4] ) );
  dff_sg \filter_0/reg_w_14_reg[5]  ( .D(\filter_0/n9027 ), .CP(clk), .Q(
        \filter_0/reg_w_14[5] ) );
  dff_sg \filter_0/reg_w_14_reg[6]  ( .D(\filter_0/n9026 ), .CP(clk), .Q(
        \filter_0/reg_w_14[6] ) );
  dff_sg \filter_0/reg_w_14_reg[7]  ( .D(\filter_0/n9025 ), .CP(clk), .Q(
        \filter_0/reg_w_14[7] ) );
  dff_sg \filter_0/reg_w_14_reg[8]  ( .D(\filter_0/n9024 ), .CP(clk), .Q(
        \filter_0/reg_w_14[8] ) );
  dff_sg \filter_0/reg_w_14_reg[9]  ( .D(\filter_0/n9023 ), .CP(clk), .Q(
        \filter_0/reg_w_14[9] ) );
  dff_sg \filter_0/reg_w_14_reg[10]  ( .D(\filter_0/n9022 ), .CP(clk), .Q(
        \filter_0/reg_w_14[10] ) );
  dff_sg \filter_0/reg_w_14_reg[11]  ( .D(\filter_0/n9021 ), .CP(clk), .Q(
        \filter_0/reg_w_14[11] ) );
  dff_sg \filter_0/reg_w_14_reg[12]  ( .D(\filter_0/n9020 ), .CP(clk), .Q(
        \filter_0/reg_w_14[12] ) );
  dff_sg \filter_0/reg_w_14_reg[13]  ( .D(\filter_0/n9019 ), .CP(clk), .Q(
        \filter_0/reg_w_14[13] ) );
  dff_sg \filter_0/reg_w_14_reg[14]  ( .D(\filter_0/n9018 ), .CP(clk), .Q(
        \filter_0/reg_w_14[14] ) );
  dff_sg \filter_0/reg_w_14_reg[15]  ( .D(\filter_0/n9017 ), .CP(clk), .Q(
        \filter_0/reg_w_14[15] ) );
  dff_sg \filter_0/reg_w_14_reg[16]  ( .D(\filter_0/n9016 ), .CP(clk), .Q(
        \filter_0/reg_w_14[16] ) );
  dff_sg \filter_0/reg_w_14_reg[17]  ( .D(\filter_0/n9015 ), .CP(clk), .Q(
        \filter_0/reg_w_14[17] ) );
  dff_sg \filter_0/reg_w_14_reg[18]  ( .D(\filter_0/n9014 ), .CP(clk), .Q(
        \filter_0/reg_w_14[18] ) );
  dff_sg \filter_0/reg_w_14_reg[19]  ( .D(\filter_0/n9013 ), .CP(clk), .Q(
        \filter_0/reg_w_14[19] ) );
  dff_sg \filter_0/reg_w_15_reg[0]  ( .D(\filter_0/n9012 ), .CP(clk), .Q(
        \filter_0/reg_w_15[0] ) );
  dff_sg \filter_0/reg_w_15_reg[1]  ( .D(\filter_0/n9011 ), .CP(clk), .Q(
        \filter_0/reg_w_15[1] ) );
  dff_sg \filter_0/reg_w_15_reg[2]  ( .D(\filter_0/n9010 ), .CP(clk), .Q(
        \filter_0/reg_w_15[2] ) );
  dff_sg \filter_0/reg_w_15_reg[3]  ( .D(\filter_0/n9009 ), .CP(clk), .Q(
        \filter_0/reg_w_15[3] ) );
  dff_sg \filter_0/reg_w_15_reg[4]  ( .D(\filter_0/n9008 ), .CP(clk), .Q(
        \filter_0/reg_w_15[4] ) );
  dff_sg \filter_0/reg_w_15_reg[5]  ( .D(\filter_0/n9007 ), .CP(clk), .Q(
        \filter_0/reg_w_15[5] ) );
  dff_sg \filter_0/reg_w_15_reg[6]  ( .D(\filter_0/n9006 ), .CP(clk), .Q(
        \filter_0/reg_w_15[6] ) );
  dff_sg \filter_0/reg_w_15_reg[7]  ( .D(\filter_0/n9005 ), .CP(clk), .Q(
        \filter_0/reg_w_15[7] ) );
  dff_sg \filter_0/reg_w_15_reg[8]  ( .D(\filter_0/n9004 ), .CP(clk), .Q(
        \filter_0/reg_w_15[8] ) );
  dff_sg \filter_0/reg_w_15_reg[9]  ( .D(\filter_0/n9003 ), .CP(clk), .Q(
        \filter_0/reg_w_15[9] ) );
  dff_sg \filter_0/reg_w_15_reg[10]  ( .D(\filter_0/n9002 ), .CP(clk), .Q(
        \filter_0/reg_w_15[10] ) );
  dff_sg \filter_0/reg_w_15_reg[11]  ( .D(\filter_0/n9001 ), .CP(clk), .Q(
        \filter_0/reg_w_15[11] ) );
  dff_sg \filter_0/reg_w_15_reg[12]  ( .D(\filter_0/n9000 ), .CP(clk), .Q(
        \filter_0/reg_w_15[12] ) );
  dff_sg \filter_0/reg_w_15_reg[13]  ( .D(\filter_0/n8999 ), .CP(clk), .Q(
        \filter_0/reg_w_15[13] ) );
  dff_sg \filter_0/reg_w_15_reg[14]  ( .D(\filter_0/n8998 ), .CP(clk), .Q(
        \filter_0/reg_w_15[14] ) );
  dff_sg \filter_0/reg_w_15_reg[15]  ( .D(\filter_0/n8997 ), .CP(clk), .Q(
        \filter_0/reg_w_15[15] ) );
  dff_sg \filter_0/reg_w_15_reg[16]  ( .D(\filter_0/n8996 ), .CP(clk), .Q(
        \filter_0/reg_w_15[16] ) );
  dff_sg \filter_0/reg_w_15_reg[17]  ( .D(\filter_0/n8995 ), .CP(clk), .Q(
        \filter_0/reg_w_15[17] ) );
  dff_sg \filter_0/reg_w_15_reg[18]  ( .D(\filter_0/n8994 ), .CP(clk), .Q(
        \filter_0/reg_w_15[18] ) );
  dff_sg \filter_0/reg_w_15_reg[19]  ( .D(\filter_0/n8993 ), .CP(clk), .Q(
        \filter_0/reg_w_15[19] ) );
  dff_sg \filter_0/reg_o_mask_reg[0]  ( .D(\filter_0/n8992 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[0] ) );
  dff_sg \filter_0/reg_o_mask_reg[1]  ( .D(\filter_0/n8991 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[1] ) );
  dff_sg \filter_0/reg_o_mask_reg[2]  ( .D(\filter_0/n8990 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[2] ) );
  dff_sg \filter_0/reg_o_mask_reg[3]  ( .D(\filter_0/n8989 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[3] ) );
  dff_sg \filter_0/reg_o_mask_reg[4]  ( .D(\filter_0/n8988 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[4] ) );
  dff_sg \filter_0/reg_o_mask_reg[5]  ( .D(\filter_0/n8987 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[5] ) );
  dff_sg \filter_0/reg_o_mask_reg[6]  ( .D(\filter_0/n8986 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[6] ) );
  dff_sg \filter_0/reg_o_mask_reg[7]  ( .D(\filter_0/n8985 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[7] ) );
  dff_sg \filter_0/reg_o_mask_reg[8]  ( .D(\filter_0/n8984 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[8] ) );
  dff_sg \filter_0/reg_o_mask_reg[9]  ( .D(\filter_0/n8983 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[9] ) );
  dff_sg \filter_0/reg_o_mask_reg[10]  ( .D(\filter_0/n8982 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[10] ) );
  dff_sg \filter_0/reg_o_mask_reg[11]  ( .D(\filter_0/n8981 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[11] ) );
  dff_sg \filter_0/reg_o_mask_reg[12]  ( .D(\filter_0/n8980 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[12] ) );
  dff_sg \filter_0/reg_o_mask_reg[13]  ( .D(\filter_0/n8979 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[13] ) );
  dff_sg \filter_0/reg_o_mask_reg[14]  ( .D(\filter_0/n8978 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[14] ) );
  dff_sg \filter_0/reg_o_mask_reg[15]  ( .D(\filter_0/n8977 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[15] ) );
  dff_sg \filter_0/reg_o_mask_reg[16]  ( .D(\filter_0/n8976 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[16] ) );
  dff_sg \filter_0/reg_o_mask_reg[17]  ( .D(\filter_0/n8975 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[17] ) );
  dff_sg \filter_0/reg_o_mask_reg[18]  ( .D(\filter_0/n8974 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[18] ) );
  dff_sg \filter_0/reg_o_mask_reg[19]  ( .D(\filter_0/n8973 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[19] ) );
  dff_sg \filter_0/reg_o_mask_reg[20]  ( .D(\filter_0/n8972 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[20] ) );
  dff_sg \filter_0/reg_o_mask_reg[21]  ( .D(\filter_0/n8971 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[21] ) );
  dff_sg \filter_0/reg_o_mask_reg[22]  ( .D(\filter_0/n8970 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[22] ) );
  dff_sg \filter_0/reg_o_mask_reg[23]  ( .D(\filter_0/n8969 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[23] ) );
  dff_sg \filter_0/reg_o_mask_reg[24]  ( .D(\filter_0/n8968 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[24] ) );
  dff_sg \filter_0/reg_o_mask_reg[25]  ( .D(\filter_0/n8967 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[25] ) );
  dff_sg \filter_0/reg_o_mask_reg[26]  ( .D(\filter_0/n8966 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[26] ) );
  dff_sg \filter_0/reg_o_mask_reg[27]  ( .D(\filter_0/n8965 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[27] ) );
  dff_sg \filter_0/reg_o_mask_reg[28]  ( .D(\filter_0/n8964 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[28] ) );
  dff_sg \filter_0/reg_o_mask_reg[29]  ( .D(\filter_0/n8963 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[29] ) );
  dff_sg \filter_0/reg_o_mask_reg[30]  ( .D(\filter_0/n8962 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[30] ) );
  dff_sg \filter_0/reg_o_mask_reg[31]  ( .D(\filter_0/n8961 ), .CP(clk), .Q(
        \filter_0/reg_o_mask[31] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[0]  ( .D(\filter_0/n8960 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[0] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[1]  ( .D(\filter_0/n8959 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[1] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[2]  ( .D(\filter_0/n8958 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[2] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[3]  ( .D(\filter_0/n8957 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[3] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[4]  ( .D(\filter_0/n8956 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[4] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[5]  ( .D(\filter_0/n8955 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[5] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[6]  ( .D(\filter_0/n8954 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[6] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[7]  ( .D(\filter_0/n8953 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[7] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[8]  ( .D(\filter_0/n8952 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[8] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[9]  ( .D(\filter_0/n8951 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[9] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[10]  ( .D(\filter_0/n8950 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[10] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[11]  ( .D(\filter_0/n8949 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[11] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[12]  ( .D(\filter_0/n8948 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[12] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[13]  ( .D(\filter_0/n8947 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[13] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[14]  ( .D(\filter_0/n8946 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[14] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[15]  ( .D(\filter_0/n8945 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[15] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[16]  ( .D(\filter_0/n8944 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[16] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[17]  ( .D(\filter_0/n8943 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[17] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[18]  ( .D(\filter_0/n8942 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[18] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[19]  ( .D(\filter_0/n8941 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[19] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[20]  ( .D(\filter_0/n8940 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[20] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[21]  ( .D(\filter_0/n8939 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[21] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[22]  ( .D(\filter_0/n8938 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[22] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[23]  ( .D(\filter_0/n8937 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[23] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[24]  ( .D(\filter_0/n8936 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[24] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[25]  ( .D(\filter_0/n8935 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[25] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[26]  ( .D(\filter_0/n8934 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[26] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[27]  ( .D(\filter_0/n8933 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[27] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[28]  ( .D(\filter_0/n8932 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[28] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[29]  ( .D(\filter_0/n8931 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[29] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[30]  ( .D(\filter_0/n8930 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[30] ) );
  dff_sg \filter_0/reg_xor_i_mask_reg[31]  ( .D(\filter_0/n8929 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask[31] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[0]  ( .D(\filter_0/n8928 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[0] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[1]  ( .D(\filter_0/n8927 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[1] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[2]  ( .D(\filter_0/n8926 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[2] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[3]  ( .D(\filter_0/n8925 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[3] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[4]  ( .D(\filter_0/n8924 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[4] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[5]  ( .D(\filter_0/n8923 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[5] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[6]  ( .D(\filter_0/n8922 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[6] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[7]  ( .D(\filter_0/n8921 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[7] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[8]  ( .D(\filter_0/n8920 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[8] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[9]  ( .D(\filter_0/n8919 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[9] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[10]  ( .D(\filter_0/n8918 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[10] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[11]  ( .D(\filter_0/n8917 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[11] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[12]  ( .D(\filter_0/n8916 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[12] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[13]  ( .D(\filter_0/n8915 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[13] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[14]  ( .D(\filter_0/n8914 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[14] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[15]  ( .D(\filter_0/n8913 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[15] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[16]  ( .D(\filter_0/n8912 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[16] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[17]  ( .D(\filter_0/n8911 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[17] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[18]  ( .D(\filter_0/n8910 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[18] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[19]  ( .D(\filter_0/n8909 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[19] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[20]  ( .D(\filter_0/n8908 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[20] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[21]  ( .D(\filter_0/n8907 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[21] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[22]  ( .D(\filter_0/n8906 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[22] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[23]  ( .D(\filter_0/n8905 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[23] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[24]  ( .D(\filter_0/n8904 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[24] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[25]  ( .D(\filter_0/n8903 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[25] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[26]  ( .D(\filter_0/n8902 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[26] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[27]  ( .D(\filter_0/n8901 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[27] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[28]  ( .D(\filter_0/n8900 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[28] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[29]  ( .D(\filter_0/n8899 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[29] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[30]  ( .D(\filter_0/n8898 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[30] ) );
  dff_sg \filter_0/reg_xor_w_mask_reg[31]  ( .D(\filter_0/n8897 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask[31] ) );
  dff_sg \filter_0/state_reg[0]  ( .D(\filter_0/n9634 ), .CP(clk), .Q(
        filter_state[0]) );
  dff_sg \filter_0/state_reg[1]  ( .D(\filter_0/n9635 ), .CP(clk), .Q(
        filter_state[1]) );
  dff_sg \filter_0/done_reg  ( .D(\filter_0/N1845 ), .CP(clk), .Q(
        \filter_0/done ) );
  dff_sg \shifter_0/ow_14_reg[0]  ( .D(\shifter_0/n9592 ), .CP(clk), .Q(
        ow_14[0]) );
  dff_sg \shifter_0/ow_14_reg[1]  ( .D(\shifter_0/n9593 ), .CP(clk), .Q(
        ow_14[1]) );
  dff_sg \shifter_0/ow_14_reg[2]  ( .D(\shifter_0/n9594 ), .CP(clk), .Q(
        ow_14[2]) );
  dff_sg \shifter_0/ow_14_reg[3]  ( .D(\shifter_0/n9595 ), .CP(clk), .Q(
        ow_14[3]) );
  dff_sg \shifter_0/ow_14_reg[4]  ( .D(\shifter_0/n9596 ), .CP(clk), .Q(
        ow_14[4]) );
  dff_sg \shifter_0/ow_14_reg[5]  ( .D(\shifter_0/n9597 ), .CP(clk), .Q(
        ow_14[5]) );
  dff_sg \shifter_0/ow_14_reg[6]  ( .D(\shifter_0/n9598 ), .CP(clk), .Q(
        ow_14[6]) );
  dff_sg \shifter_0/ow_14_reg[7]  ( .D(\shifter_0/n9599 ), .CP(clk), .Q(
        ow_14[7]) );
  dff_sg \shifter_0/ow_14_reg[8]  ( .D(\shifter_0/n9600 ), .CP(clk), .Q(
        ow_14[8]) );
  dff_sg \shifter_0/ow_14_reg[9]  ( .D(\shifter_0/n9601 ), .CP(clk), .Q(
        ow_14[9]) );
  dff_sg \shifter_0/ow_14_reg[10]  ( .D(\shifter_0/n9602 ), .CP(clk), .Q(
        ow_14[10]) );
  dff_sg \shifter_0/ow_14_reg[11]  ( .D(\shifter_0/n9603 ), .CP(clk), .Q(
        ow_14[11]) );
  dff_sg \shifter_0/ow_14_reg[12]  ( .D(\shifter_0/n9604 ), .CP(clk), .Q(
        ow_14[12]) );
  dff_sg \shifter_0/ow_14_reg[13]  ( .D(\shifter_0/n9605 ), .CP(clk), .Q(
        ow_14[13]) );
  dff_sg \shifter_0/ow_14_reg[14]  ( .D(\shifter_0/n9606 ), .CP(clk), .Q(
        ow_14[14]) );
  dff_sg \shifter_0/ow_14_reg[15]  ( .D(\shifter_0/n9607 ), .CP(clk), .Q(
        ow_14[15]) );
  dff_sg \shifter_0/ow_14_reg[16]  ( .D(\shifter_0/n9608 ), .CP(clk), .Q(
        ow_14[16]) );
  dff_sg \shifter_0/ow_14_reg[17]  ( .D(\shifter_0/n9609 ), .CP(clk), .Q(
        ow_14[17]) );
  dff_sg \shifter_0/ow_14_reg[18]  ( .D(\shifter_0/n9610 ), .CP(clk), .Q(
        ow_14[18]) );
  dff_sg \shifter_0/ow_14_reg[19]  ( .D(\shifter_0/n9611 ), .CP(clk), .Q(
        ow_14[19]) );
  dff_sg \shifter_0/ow_13_reg[0]  ( .D(\shifter_0/n9612 ), .CP(clk), .Q(
        ow_13[0]) );
  dff_sg \shifter_0/ow_13_reg[1]  ( .D(\shifter_0/n9613 ), .CP(clk), .Q(
        ow_13[1]) );
  dff_sg \shifter_0/ow_13_reg[2]  ( .D(\shifter_0/n9614 ), .CP(clk), .Q(
        ow_13[2]) );
  dff_sg \shifter_0/ow_13_reg[3]  ( .D(\shifter_0/n9615 ), .CP(clk), .Q(
        ow_13[3]) );
  dff_sg \shifter_0/ow_13_reg[4]  ( .D(\shifter_0/n9616 ), .CP(clk), .Q(
        ow_13[4]) );
  dff_sg \shifter_0/ow_13_reg[5]  ( .D(\shifter_0/n9617 ), .CP(clk), .Q(
        ow_13[5]) );
  dff_sg \shifter_0/ow_13_reg[6]  ( .D(\shifter_0/n9618 ), .CP(clk), .Q(
        ow_13[6]) );
  dff_sg \shifter_0/ow_13_reg[7]  ( .D(\shifter_0/n9619 ), .CP(clk), .Q(
        ow_13[7]) );
  dff_sg \shifter_0/ow_13_reg[8]  ( .D(\shifter_0/n9620 ), .CP(clk), .Q(
        ow_13[8]) );
  dff_sg \shifter_0/ow_13_reg[9]  ( .D(\shifter_0/n9621 ), .CP(clk), .Q(
        ow_13[9]) );
  dff_sg \shifter_0/ow_13_reg[10]  ( .D(\shifter_0/n9622 ), .CP(clk), .Q(
        ow_13[10]) );
  dff_sg \shifter_0/ow_13_reg[11]  ( .D(\shifter_0/n9623 ), .CP(clk), .Q(
        ow_13[11]) );
  dff_sg \shifter_0/ow_13_reg[12]  ( .D(\shifter_0/n9624 ), .CP(clk), .Q(
        ow_13[12]) );
  dff_sg \shifter_0/ow_13_reg[13]  ( .D(\shifter_0/n9625 ), .CP(clk), .Q(
        ow_13[13]) );
  dff_sg \shifter_0/ow_13_reg[14]  ( .D(\shifter_0/n9626 ), .CP(clk), .Q(
        ow_13[14]) );
  dff_sg \shifter_0/ow_13_reg[15]  ( .D(\shifter_0/n9627 ), .CP(clk), .Q(
        ow_13[15]) );
  dff_sg \shifter_0/ow_13_reg[16]  ( .D(\shifter_0/n9628 ), .CP(clk), .Q(
        ow_13[16]) );
  dff_sg \shifter_0/ow_13_reg[17]  ( .D(\shifter_0/n9629 ), .CP(clk), .Q(
        ow_13[17]) );
  dff_sg \shifter_0/ow_13_reg[18]  ( .D(\shifter_0/n9630 ), .CP(clk), .Q(
        ow_13[18]) );
  dff_sg \shifter_0/ow_13_reg[19]  ( .D(\shifter_0/n9631 ), .CP(clk), .Q(
        ow_13[19]) );
  dff_sg \shifter_0/ow_12_reg[0]  ( .D(\shifter_0/n9632 ), .CP(clk), .Q(
        ow_12[0]) );
  dff_sg \shifter_0/ow_12_reg[1]  ( .D(\shifter_0/n9633 ), .CP(clk), .Q(
        ow_12[1]) );
  dff_sg \shifter_0/ow_12_reg[2]  ( .D(\shifter_0/n9634 ), .CP(clk), .Q(
        ow_12[2]) );
  dff_sg \shifter_0/ow_12_reg[3]  ( .D(\shifter_0/n9635 ), .CP(clk), .Q(
        ow_12[3]) );
  dff_sg \shifter_0/ow_12_reg[4]  ( .D(\shifter_0/n9636 ), .CP(clk), .Q(
        ow_12[4]) );
  dff_sg \shifter_0/ow_12_reg[5]  ( .D(\shifter_0/n9637 ), .CP(clk), .Q(
        ow_12[5]) );
  dff_sg \shifter_0/ow_12_reg[6]  ( .D(\shifter_0/n9638 ), .CP(clk), .Q(
        ow_12[6]) );
  dff_sg \shifter_0/ow_12_reg[7]  ( .D(\shifter_0/n9639 ), .CP(clk), .Q(
        ow_12[7]) );
  dff_sg \shifter_0/ow_12_reg[8]  ( .D(\shifter_0/n9640 ), .CP(clk), .Q(
        ow_12[8]) );
  dff_sg \shifter_0/ow_12_reg[9]  ( .D(\shifter_0/n9641 ), .CP(clk), .Q(
        ow_12[9]) );
  dff_sg \shifter_0/ow_12_reg[10]  ( .D(\shifter_0/n9642 ), .CP(clk), .Q(
        ow_12[10]) );
  dff_sg \shifter_0/ow_12_reg[11]  ( .D(\shifter_0/n9643 ), .CP(clk), .Q(
        ow_12[11]) );
  dff_sg \shifter_0/ow_12_reg[12]  ( .D(\shifter_0/n9644 ), .CP(clk), .Q(
        ow_12[12]) );
  dff_sg \shifter_0/ow_12_reg[13]  ( .D(\shifter_0/n9645 ), .CP(clk), .Q(
        ow_12[13]) );
  dff_sg \shifter_0/ow_12_reg[14]  ( .D(\shifter_0/n9646 ), .CP(clk), .Q(
        ow_12[14]) );
  dff_sg \shifter_0/ow_12_reg[15]  ( .D(\shifter_0/n9647 ), .CP(clk), .Q(
        ow_12[15]) );
  dff_sg \shifter_0/ow_12_reg[16]  ( .D(\shifter_0/n9648 ), .CP(clk), .Q(
        ow_12[16]) );
  dff_sg \shifter_0/ow_12_reg[17]  ( .D(\shifter_0/n9649 ), .CP(clk), .Q(
        ow_12[17]) );
  dff_sg \shifter_0/ow_12_reg[18]  ( .D(\shifter_0/n9650 ), .CP(clk), .Q(
        ow_12[18]) );
  dff_sg \shifter_0/ow_12_reg[19]  ( .D(\shifter_0/n9651 ), .CP(clk), .Q(
        ow_12[19]) );
  dff_sg \shifter_0/ow_11_reg[0]  ( .D(\shifter_0/n9652 ), .CP(clk), .Q(
        ow_11[0]) );
  dff_sg \shifter_0/ow_11_reg[1]  ( .D(\shifter_0/n9653 ), .CP(clk), .Q(
        ow_11[1]) );
  dff_sg \shifter_0/ow_11_reg[2]  ( .D(\shifter_0/n9654 ), .CP(clk), .Q(
        ow_11[2]) );
  dff_sg \shifter_0/ow_11_reg[3]  ( .D(\shifter_0/n9655 ), .CP(clk), .Q(
        ow_11[3]) );
  dff_sg \shifter_0/ow_11_reg[4]  ( .D(\shifter_0/n9656 ), .CP(clk), .Q(
        ow_11[4]) );
  dff_sg \shifter_0/ow_11_reg[5]  ( .D(\shifter_0/n9657 ), .CP(clk), .Q(
        ow_11[5]) );
  dff_sg \shifter_0/ow_11_reg[6]  ( .D(\shifter_0/n9658 ), .CP(clk), .Q(
        ow_11[6]) );
  dff_sg \shifter_0/ow_11_reg[7]  ( .D(\shifter_0/n9659 ), .CP(clk), .Q(
        ow_11[7]) );
  dff_sg \shifter_0/ow_11_reg[8]  ( .D(\shifter_0/n9660 ), .CP(clk), .Q(
        ow_11[8]) );
  dff_sg \shifter_0/ow_11_reg[9]  ( .D(\shifter_0/n9661 ), .CP(clk), .Q(
        ow_11[9]) );
  dff_sg \shifter_0/ow_11_reg[10]  ( .D(\shifter_0/n9662 ), .CP(clk), .Q(
        ow_11[10]) );
  dff_sg \shifter_0/ow_11_reg[11]  ( .D(\shifter_0/n9663 ), .CP(clk), .Q(
        ow_11[11]) );
  dff_sg \shifter_0/ow_11_reg[12]  ( .D(\shifter_0/n9664 ), .CP(clk), .Q(
        ow_11[12]) );
  dff_sg \shifter_0/ow_11_reg[13]  ( .D(\shifter_0/n9665 ), .CP(clk), .Q(
        ow_11[13]) );
  dff_sg \shifter_0/ow_11_reg[14]  ( .D(\shifter_0/n9666 ), .CP(clk), .Q(
        ow_11[14]) );
  dff_sg \shifter_0/ow_11_reg[15]  ( .D(\shifter_0/n9667 ), .CP(clk), .Q(
        ow_11[15]) );
  dff_sg \shifter_0/ow_11_reg[16]  ( .D(\shifter_0/n9668 ), .CP(clk), .Q(
        ow_11[16]) );
  dff_sg \shifter_0/ow_11_reg[17]  ( .D(\shifter_0/n9669 ), .CP(clk), .Q(
        ow_11[17]) );
  dff_sg \shifter_0/ow_11_reg[18]  ( .D(\shifter_0/n9670 ), .CP(clk), .Q(
        ow_11[18]) );
  dff_sg \shifter_0/ow_11_reg[19]  ( .D(\shifter_0/n9671 ), .CP(clk), .Q(
        ow_11[19]) );
  dff_sg \shifter_0/ow_10_reg[0]  ( .D(\shifter_0/n9672 ), .CP(clk), .Q(
        ow_10[0]) );
  dff_sg \shifter_0/ow_10_reg[1]  ( .D(\shifter_0/n9673 ), .CP(clk), .Q(
        ow_10[1]) );
  dff_sg \shifter_0/ow_10_reg[2]  ( .D(\shifter_0/n9674 ), .CP(clk), .Q(
        ow_10[2]) );
  dff_sg \shifter_0/ow_10_reg[3]  ( .D(\shifter_0/n9675 ), .CP(clk), .Q(
        ow_10[3]) );
  dff_sg \shifter_0/ow_10_reg[4]  ( .D(\shifter_0/n9676 ), .CP(clk), .Q(
        ow_10[4]) );
  dff_sg \shifter_0/ow_10_reg[5]  ( .D(\shifter_0/n9677 ), .CP(clk), .Q(
        ow_10[5]) );
  dff_sg \shifter_0/ow_10_reg[6]  ( .D(\shifter_0/n9678 ), .CP(clk), .Q(
        ow_10[6]) );
  dff_sg \shifter_0/ow_10_reg[7]  ( .D(\shifter_0/n9679 ), .CP(clk), .Q(
        ow_10[7]) );
  dff_sg \shifter_0/ow_10_reg[8]  ( .D(\shifter_0/n9680 ), .CP(clk), .Q(
        ow_10[8]) );
  dff_sg \shifter_0/ow_10_reg[9]  ( .D(\shifter_0/n9681 ), .CP(clk), .Q(
        ow_10[9]) );
  dff_sg \shifter_0/ow_10_reg[10]  ( .D(\shifter_0/n9682 ), .CP(clk), .Q(
        ow_10[10]) );
  dff_sg \shifter_0/ow_10_reg[11]  ( .D(\shifter_0/n9683 ), .CP(clk), .Q(
        ow_10[11]) );
  dff_sg \shifter_0/ow_10_reg[12]  ( .D(\shifter_0/n9684 ), .CP(clk), .Q(
        ow_10[12]) );
  dff_sg \shifter_0/ow_10_reg[13]  ( .D(\shifter_0/n9685 ), .CP(clk), .Q(
        ow_10[13]) );
  dff_sg \shifter_0/ow_10_reg[14]  ( .D(\shifter_0/n9686 ), .CP(clk), .Q(
        ow_10[14]) );
  dff_sg \shifter_0/ow_10_reg[15]  ( .D(\shifter_0/n9687 ), .CP(clk), .Q(
        ow_10[15]) );
  dff_sg \shifter_0/ow_10_reg[16]  ( .D(\shifter_0/n9688 ), .CP(clk), .Q(
        ow_10[16]) );
  dff_sg \shifter_0/ow_10_reg[17]  ( .D(\shifter_0/n9689 ), .CP(clk), .Q(
        ow_10[17]) );
  dff_sg \shifter_0/ow_10_reg[18]  ( .D(\shifter_0/n9690 ), .CP(clk), .Q(
        ow_10[18]) );
  dff_sg \shifter_0/ow_10_reg[19]  ( .D(\shifter_0/n9691 ), .CP(clk), .Q(
        ow_10[19]) );
  dff_sg \shifter_0/ow_9_reg[0]  ( .D(\shifter_0/n9692 ), .CP(clk), .Q(ow_9[0]) );
  dff_sg \shifter_0/ow_9_reg[1]  ( .D(\shifter_0/n9693 ), .CP(clk), .Q(ow_9[1]) );
  dff_sg \shifter_0/ow_9_reg[2]  ( .D(\shifter_0/n9694 ), .CP(clk), .Q(ow_9[2]) );
  dff_sg \shifter_0/ow_9_reg[3]  ( .D(\shifter_0/n9695 ), .CP(clk), .Q(ow_9[3]) );
  dff_sg \shifter_0/ow_9_reg[4]  ( .D(\shifter_0/n9696 ), .CP(clk), .Q(ow_9[4]) );
  dff_sg \shifter_0/ow_9_reg[5]  ( .D(\shifter_0/n9697 ), .CP(clk), .Q(ow_9[5]) );
  dff_sg \shifter_0/ow_9_reg[6]  ( .D(\shifter_0/n9698 ), .CP(clk), .Q(ow_9[6]) );
  dff_sg \shifter_0/ow_9_reg[7]  ( .D(\shifter_0/n9699 ), .CP(clk), .Q(ow_9[7]) );
  dff_sg \shifter_0/ow_9_reg[8]  ( .D(\shifter_0/n9700 ), .CP(clk), .Q(ow_9[8]) );
  dff_sg \shifter_0/ow_9_reg[9]  ( .D(\shifter_0/n9701 ), .CP(clk), .Q(ow_9[9]) );
  dff_sg \shifter_0/ow_9_reg[10]  ( .D(\shifter_0/n9702 ), .CP(clk), .Q(
        ow_9[10]) );
  dff_sg \shifter_0/ow_9_reg[11]  ( .D(\shifter_0/n9703 ), .CP(clk), .Q(
        ow_9[11]) );
  dff_sg \shifter_0/ow_9_reg[12]  ( .D(\shifter_0/n9704 ), .CP(clk), .Q(
        ow_9[12]) );
  dff_sg \shifter_0/ow_9_reg[13]  ( .D(\shifter_0/n9705 ), .CP(clk), .Q(
        ow_9[13]) );
  dff_sg \shifter_0/ow_9_reg[14]  ( .D(\shifter_0/n9706 ), .CP(clk), .Q(
        ow_9[14]) );
  dff_sg \shifter_0/ow_9_reg[15]  ( .D(\shifter_0/n9707 ), .CP(clk), .Q(
        ow_9[15]) );
  dff_sg \shifter_0/ow_9_reg[16]  ( .D(\shifter_0/n9708 ), .CP(clk), .Q(
        ow_9[16]) );
  dff_sg \shifter_0/ow_9_reg[17]  ( .D(\shifter_0/n9709 ), .CP(clk), .Q(
        ow_9[17]) );
  dff_sg \shifter_0/ow_9_reg[18]  ( .D(\shifter_0/n9710 ), .CP(clk), .Q(
        ow_9[18]) );
  dff_sg \shifter_0/ow_9_reg[19]  ( .D(\shifter_0/n9711 ), .CP(clk), .Q(
        ow_9[19]) );
  dff_sg \shifter_0/ow_8_reg[0]  ( .D(\shifter_0/n9712 ), .CP(clk), .Q(ow_8[0]) );
  dff_sg \shifter_0/ow_8_reg[1]  ( .D(\shifter_0/n9713 ), .CP(clk), .Q(ow_8[1]) );
  dff_sg \shifter_0/ow_8_reg[2]  ( .D(\shifter_0/n9714 ), .CP(clk), .Q(ow_8[2]) );
  dff_sg \shifter_0/ow_8_reg[3]  ( .D(\shifter_0/n9715 ), .CP(clk), .Q(ow_8[3]) );
  dff_sg \shifter_0/ow_8_reg[4]  ( .D(\shifter_0/n9716 ), .CP(clk), .Q(ow_8[4]) );
  dff_sg \shifter_0/ow_8_reg[5]  ( .D(\shifter_0/n9717 ), .CP(clk), .Q(ow_8[5]) );
  dff_sg \shifter_0/ow_8_reg[6]  ( .D(\shifter_0/n9718 ), .CP(clk), .Q(ow_8[6]) );
  dff_sg \shifter_0/ow_8_reg[7]  ( .D(\shifter_0/n9719 ), .CP(clk), .Q(ow_8[7]) );
  dff_sg \shifter_0/ow_8_reg[8]  ( .D(\shifter_0/n9720 ), .CP(clk), .Q(ow_8[8]) );
  dff_sg \shifter_0/ow_8_reg[9]  ( .D(\shifter_0/n9721 ), .CP(clk), .Q(ow_8[9]) );
  dff_sg \shifter_0/ow_8_reg[10]  ( .D(\shifter_0/n9722 ), .CP(clk), .Q(
        ow_8[10]) );
  dff_sg \shifter_0/ow_8_reg[11]  ( .D(\shifter_0/n9723 ), .CP(clk), .Q(
        ow_8[11]) );
  dff_sg \shifter_0/ow_8_reg[12]  ( .D(\shifter_0/n9724 ), .CP(clk), .Q(
        ow_8[12]) );
  dff_sg \shifter_0/ow_8_reg[13]  ( .D(\shifter_0/n9725 ), .CP(clk), .Q(
        ow_8[13]) );
  dff_sg \shifter_0/ow_8_reg[14]  ( .D(\shifter_0/n9726 ), .CP(clk), .Q(
        ow_8[14]) );
  dff_sg \shifter_0/ow_8_reg[15]  ( .D(\shifter_0/n9727 ), .CP(clk), .Q(
        ow_8[15]) );
  dff_sg \shifter_0/ow_8_reg[16]  ( .D(\shifter_0/n9728 ), .CP(clk), .Q(
        ow_8[16]) );
  dff_sg \shifter_0/ow_8_reg[17]  ( .D(\shifter_0/n9729 ), .CP(clk), .Q(
        ow_8[17]) );
  dff_sg \shifter_0/ow_8_reg[18]  ( .D(\shifter_0/n9730 ), .CP(clk), .Q(
        ow_8[18]) );
  dff_sg \shifter_0/ow_8_reg[19]  ( .D(\shifter_0/n9731 ), .CP(clk), .Q(
        ow_8[19]) );
  dff_sg \shifter_0/ow_7_reg[0]  ( .D(\shifter_0/n9732 ), .CP(clk), .Q(ow_7[0]) );
  dff_sg \shifter_0/ow_7_reg[1]  ( .D(\shifter_0/n9733 ), .CP(clk), .Q(ow_7[1]) );
  dff_sg \shifter_0/ow_7_reg[2]  ( .D(\shifter_0/n9734 ), .CP(clk), .Q(ow_7[2]) );
  dff_sg \shifter_0/ow_7_reg[3]  ( .D(\shifter_0/n9735 ), .CP(clk), .Q(ow_7[3]) );
  dff_sg \shifter_0/ow_7_reg[4]  ( .D(\shifter_0/n9736 ), .CP(clk), .Q(ow_7[4]) );
  dff_sg \shifter_0/ow_7_reg[5]  ( .D(\shifter_0/n9737 ), .CP(clk), .Q(ow_7[5]) );
  dff_sg \shifter_0/ow_7_reg[6]  ( .D(\shifter_0/n9738 ), .CP(clk), .Q(ow_7[6]) );
  dff_sg \shifter_0/ow_7_reg[7]  ( .D(\shifter_0/n9739 ), .CP(clk), .Q(ow_7[7]) );
  dff_sg \shifter_0/ow_7_reg[8]  ( .D(\shifter_0/n9740 ), .CP(clk), .Q(ow_7[8]) );
  dff_sg \shifter_0/ow_7_reg[9]  ( .D(\shifter_0/n9741 ), .CP(clk), .Q(ow_7[9]) );
  dff_sg \shifter_0/ow_7_reg[10]  ( .D(\shifter_0/n9742 ), .CP(clk), .Q(
        ow_7[10]) );
  dff_sg \shifter_0/ow_7_reg[11]  ( .D(\shifter_0/n9743 ), .CP(clk), .Q(
        ow_7[11]) );
  dff_sg \shifter_0/ow_7_reg[12]  ( .D(\shifter_0/n9744 ), .CP(clk), .Q(
        ow_7[12]) );
  dff_sg \shifter_0/ow_7_reg[13]  ( .D(\shifter_0/n9745 ), .CP(clk), .Q(
        ow_7[13]) );
  dff_sg \shifter_0/ow_7_reg[14]  ( .D(\shifter_0/n9746 ), .CP(clk), .Q(
        ow_7[14]) );
  dff_sg \shifter_0/ow_7_reg[15]  ( .D(\shifter_0/n9747 ), .CP(clk), .Q(
        ow_7[15]) );
  dff_sg \shifter_0/ow_7_reg[16]  ( .D(\shifter_0/n9748 ), .CP(clk), .Q(
        ow_7[16]) );
  dff_sg \shifter_0/ow_7_reg[17]  ( .D(\shifter_0/n9749 ), .CP(clk), .Q(
        ow_7[17]) );
  dff_sg \shifter_0/ow_7_reg[18]  ( .D(\shifter_0/n9750 ), .CP(clk), .Q(
        ow_7[18]) );
  dff_sg \shifter_0/ow_7_reg[19]  ( .D(\shifter_0/n9751 ), .CP(clk), .Q(
        ow_7[19]) );
  dff_sg \shifter_0/ow_6_reg[0]  ( .D(\shifter_0/n9752 ), .CP(clk), .Q(ow_6[0]) );
  dff_sg \shifter_0/ow_6_reg[1]  ( .D(\shifter_0/n9753 ), .CP(clk), .Q(ow_6[1]) );
  dff_sg \shifter_0/ow_6_reg[2]  ( .D(\shifter_0/n9754 ), .CP(clk), .Q(ow_6[2]) );
  dff_sg \shifter_0/ow_6_reg[3]  ( .D(\shifter_0/n9755 ), .CP(clk), .Q(ow_6[3]) );
  dff_sg \shifter_0/ow_6_reg[4]  ( .D(\shifter_0/n9756 ), .CP(clk), .Q(ow_6[4]) );
  dff_sg \shifter_0/ow_6_reg[5]  ( .D(\shifter_0/n9757 ), .CP(clk), .Q(ow_6[5]) );
  dff_sg \shifter_0/ow_6_reg[6]  ( .D(\shifter_0/n9758 ), .CP(clk), .Q(ow_6[6]) );
  dff_sg \shifter_0/ow_6_reg[7]  ( .D(\shifter_0/n9759 ), .CP(clk), .Q(ow_6[7]) );
  dff_sg \shifter_0/ow_6_reg[8]  ( .D(\shifter_0/n9760 ), .CP(clk), .Q(ow_6[8]) );
  dff_sg \shifter_0/ow_6_reg[9]  ( .D(\shifter_0/n9761 ), .CP(clk), .Q(ow_6[9]) );
  dff_sg \shifter_0/ow_6_reg[10]  ( .D(\shifter_0/n9762 ), .CP(clk), .Q(
        ow_6[10]) );
  dff_sg \shifter_0/ow_6_reg[11]  ( .D(\shifter_0/n9763 ), .CP(clk), .Q(
        ow_6[11]) );
  dff_sg \shifter_0/ow_6_reg[12]  ( .D(\shifter_0/n9764 ), .CP(clk), .Q(
        ow_6[12]) );
  dff_sg \shifter_0/ow_6_reg[13]  ( .D(\shifter_0/n9765 ), .CP(clk), .Q(
        ow_6[13]) );
  dff_sg \shifter_0/ow_6_reg[14]  ( .D(\shifter_0/n9766 ), .CP(clk), .Q(
        ow_6[14]) );
  dff_sg \shifter_0/ow_6_reg[15]  ( .D(\shifter_0/n9767 ), .CP(clk), .Q(
        ow_6[15]) );
  dff_sg \shifter_0/ow_6_reg[16]  ( .D(\shifter_0/n9768 ), .CP(clk), .Q(
        ow_6[16]) );
  dff_sg \shifter_0/ow_6_reg[17]  ( .D(\shifter_0/n9769 ), .CP(clk), .Q(
        ow_6[17]) );
  dff_sg \shifter_0/ow_6_reg[18]  ( .D(\shifter_0/n9770 ), .CP(clk), .Q(
        ow_6[18]) );
  dff_sg \shifter_0/ow_6_reg[19]  ( .D(\shifter_0/n9771 ), .CP(clk), .Q(
        ow_6[19]) );
  dff_sg \shifter_0/ow_5_reg[0]  ( .D(\shifter_0/n9772 ), .CP(clk), .Q(ow_5[0]) );
  dff_sg \shifter_0/ow_5_reg[1]  ( .D(\shifter_0/n9773 ), .CP(clk), .Q(ow_5[1]) );
  dff_sg \shifter_0/ow_5_reg[2]  ( .D(\shifter_0/n9774 ), .CP(clk), .Q(ow_5[2]) );
  dff_sg \shifter_0/ow_5_reg[3]  ( .D(\shifter_0/n9775 ), .CP(clk), .Q(ow_5[3]) );
  dff_sg \shifter_0/ow_5_reg[4]  ( .D(\shifter_0/n9776 ), .CP(clk), .Q(ow_5[4]) );
  dff_sg \shifter_0/ow_5_reg[5]  ( .D(\shifter_0/n9777 ), .CP(clk), .Q(ow_5[5]) );
  dff_sg \shifter_0/ow_5_reg[6]  ( .D(\shifter_0/n9778 ), .CP(clk), .Q(ow_5[6]) );
  dff_sg \shifter_0/ow_5_reg[7]  ( .D(\shifter_0/n9779 ), .CP(clk), .Q(ow_5[7]) );
  dff_sg \shifter_0/ow_5_reg[8]  ( .D(\shifter_0/n9780 ), .CP(clk), .Q(ow_5[8]) );
  dff_sg \shifter_0/ow_5_reg[9]  ( .D(\shifter_0/n9781 ), .CP(clk), .Q(ow_5[9]) );
  dff_sg \shifter_0/ow_5_reg[10]  ( .D(\shifter_0/n9782 ), .CP(clk), .Q(
        ow_5[10]) );
  dff_sg \shifter_0/ow_5_reg[11]  ( .D(\shifter_0/n9783 ), .CP(clk), .Q(
        ow_5[11]) );
  dff_sg \shifter_0/ow_5_reg[12]  ( .D(\shifter_0/n9784 ), .CP(clk), .Q(
        ow_5[12]) );
  dff_sg \shifter_0/ow_5_reg[13]  ( .D(\shifter_0/n9785 ), .CP(clk), .Q(
        ow_5[13]) );
  dff_sg \shifter_0/ow_5_reg[14]  ( .D(\shifter_0/n9786 ), .CP(clk), .Q(
        ow_5[14]) );
  dff_sg \shifter_0/ow_5_reg[15]  ( .D(\shifter_0/n9787 ), .CP(clk), .Q(
        ow_5[15]) );
  dff_sg \shifter_0/ow_5_reg[16]  ( .D(\shifter_0/n9788 ), .CP(clk), .Q(
        ow_5[16]) );
  dff_sg \shifter_0/ow_5_reg[17]  ( .D(\shifter_0/n9789 ), .CP(clk), .Q(
        ow_5[17]) );
  dff_sg \shifter_0/ow_5_reg[18]  ( .D(\shifter_0/n9790 ), .CP(clk), .Q(
        ow_5[18]) );
  dff_sg \shifter_0/ow_5_reg[19]  ( .D(\shifter_0/n9791 ), .CP(clk), .Q(
        ow_5[19]) );
  dff_sg \shifter_0/ow_4_reg[0]  ( .D(\shifter_0/n9792 ), .CP(clk), .Q(ow_4[0]) );
  dff_sg \shifter_0/ow_4_reg[1]  ( .D(\shifter_0/n9793 ), .CP(clk), .Q(ow_4[1]) );
  dff_sg \shifter_0/ow_4_reg[2]  ( .D(\shifter_0/n9794 ), .CP(clk), .Q(ow_4[2]) );
  dff_sg \shifter_0/ow_4_reg[3]  ( .D(\shifter_0/n9795 ), .CP(clk), .Q(ow_4[3]) );
  dff_sg \shifter_0/ow_4_reg[4]  ( .D(\shifter_0/n9796 ), .CP(clk), .Q(ow_4[4]) );
  dff_sg \shifter_0/ow_4_reg[5]  ( .D(\shifter_0/n9797 ), .CP(clk), .Q(ow_4[5]) );
  dff_sg \shifter_0/ow_4_reg[6]  ( .D(\shifter_0/n9798 ), .CP(clk), .Q(ow_4[6]) );
  dff_sg \shifter_0/ow_4_reg[7]  ( .D(\shifter_0/n9799 ), .CP(clk), .Q(ow_4[7]) );
  dff_sg \shifter_0/ow_4_reg[8]  ( .D(\shifter_0/n9800 ), .CP(clk), .Q(ow_4[8]) );
  dff_sg \shifter_0/ow_4_reg[9]  ( .D(\shifter_0/n9801 ), .CP(clk), .Q(ow_4[9]) );
  dff_sg \shifter_0/ow_4_reg[10]  ( .D(\shifter_0/n9802 ), .CP(clk), .Q(
        ow_4[10]) );
  dff_sg \shifter_0/ow_4_reg[11]  ( .D(\shifter_0/n9803 ), .CP(clk), .Q(
        ow_4[11]) );
  dff_sg \shifter_0/ow_4_reg[12]  ( .D(\shifter_0/n9804 ), .CP(clk), .Q(
        ow_4[12]) );
  dff_sg \shifter_0/ow_4_reg[13]  ( .D(\shifter_0/n9805 ), .CP(clk), .Q(
        ow_4[13]) );
  dff_sg \shifter_0/ow_4_reg[14]  ( .D(\shifter_0/n9806 ), .CP(clk), .Q(
        ow_4[14]) );
  dff_sg \shifter_0/ow_4_reg[15]  ( .D(\shifter_0/n9807 ), .CP(clk), .Q(
        ow_4[15]) );
  dff_sg \shifter_0/ow_4_reg[16]  ( .D(\shifter_0/n9808 ), .CP(clk), .Q(
        ow_4[16]) );
  dff_sg \shifter_0/ow_4_reg[17]  ( .D(\shifter_0/n9809 ), .CP(clk), .Q(
        ow_4[17]) );
  dff_sg \shifter_0/ow_4_reg[18]  ( .D(\shifter_0/n9810 ), .CP(clk), .Q(
        ow_4[18]) );
  dff_sg \shifter_0/ow_4_reg[19]  ( .D(\shifter_0/n9811 ), .CP(clk), .Q(
        ow_4[19]) );
  dff_sg \shifter_0/ow_3_reg[0]  ( .D(\shifter_0/n9812 ), .CP(clk), .Q(ow_3[0]) );
  dff_sg \shifter_0/ow_3_reg[1]  ( .D(\shifter_0/n9813 ), .CP(clk), .Q(ow_3[1]) );
  dff_sg \shifter_0/ow_3_reg[2]  ( .D(\shifter_0/n9814 ), .CP(clk), .Q(ow_3[2]) );
  dff_sg \shifter_0/ow_3_reg[3]  ( .D(\shifter_0/n9815 ), .CP(clk), .Q(ow_3[3]) );
  dff_sg \shifter_0/ow_3_reg[4]  ( .D(\shifter_0/n9816 ), .CP(clk), .Q(ow_3[4]) );
  dff_sg \shifter_0/ow_3_reg[5]  ( .D(\shifter_0/n9817 ), .CP(clk), .Q(ow_3[5]) );
  dff_sg \shifter_0/ow_3_reg[6]  ( .D(\shifter_0/n9818 ), .CP(clk), .Q(ow_3[6]) );
  dff_sg \shifter_0/ow_3_reg[7]  ( .D(\shifter_0/n9819 ), .CP(clk), .Q(ow_3[7]) );
  dff_sg \shifter_0/ow_3_reg[8]  ( .D(\shifter_0/n9820 ), .CP(clk), .Q(ow_3[8]) );
  dff_sg \shifter_0/ow_3_reg[9]  ( .D(\shifter_0/n9821 ), .CP(clk), .Q(ow_3[9]) );
  dff_sg \shifter_0/ow_3_reg[10]  ( .D(\shifter_0/n9822 ), .CP(clk), .Q(
        ow_3[10]) );
  dff_sg \shifter_0/ow_3_reg[11]  ( .D(\shifter_0/n9823 ), .CP(clk), .Q(
        ow_3[11]) );
  dff_sg \shifter_0/ow_3_reg[12]  ( .D(\shifter_0/n9824 ), .CP(clk), .Q(
        ow_3[12]) );
  dff_sg \shifter_0/ow_3_reg[13]  ( .D(\shifter_0/n9825 ), .CP(clk), .Q(
        ow_3[13]) );
  dff_sg \shifter_0/ow_3_reg[14]  ( .D(\shifter_0/n9826 ), .CP(clk), .Q(
        ow_3[14]) );
  dff_sg \shifter_0/ow_3_reg[15]  ( .D(\shifter_0/n9827 ), .CP(clk), .Q(
        ow_3[15]) );
  dff_sg \shifter_0/ow_3_reg[16]  ( .D(\shifter_0/n9828 ), .CP(clk), .Q(
        ow_3[16]) );
  dff_sg \shifter_0/ow_3_reg[17]  ( .D(\shifter_0/n9829 ), .CP(clk), .Q(
        ow_3[17]) );
  dff_sg \shifter_0/ow_3_reg[18]  ( .D(\shifter_0/n9830 ), .CP(clk), .Q(
        ow_3[18]) );
  dff_sg \shifter_0/ow_3_reg[19]  ( .D(\shifter_0/n9831 ), .CP(clk), .Q(
        ow_3[19]) );
  dff_sg \shifter_0/ow_2_reg[0]  ( .D(\shifter_0/n9832 ), .CP(clk), .Q(ow_2[0]) );
  dff_sg \shifter_0/ow_2_reg[1]  ( .D(\shifter_0/n9833 ), .CP(clk), .Q(ow_2[1]) );
  dff_sg \shifter_0/ow_2_reg[2]  ( .D(\shifter_0/n9834 ), .CP(clk), .Q(ow_2[2]) );
  dff_sg \shifter_0/ow_2_reg[3]  ( .D(\shifter_0/n9835 ), .CP(clk), .Q(ow_2[3]) );
  dff_sg \shifter_0/ow_2_reg[4]  ( .D(\shifter_0/n9836 ), .CP(clk), .Q(ow_2[4]) );
  dff_sg \shifter_0/ow_2_reg[5]  ( .D(\shifter_0/n9837 ), .CP(clk), .Q(ow_2[5]) );
  dff_sg \shifter_0/ow_2_reg[6]  ( .D(\shifter_0/n9838 ), .CP(clk), .Q(ow_2[6]) );
  dff_sg \shifter_0/ow_2_reg[7]  ( .D(\shifter_0/n9839 ), .CP(clk), .Q(ow_2[7]) );
  dff_sg \shifter_0/ow_2_reg[8]  ( .D(\shifter_0/n9840 ), .CP(clk), .Q(ow_2[8]) );
  dff_sg \shifter_0/ow_2_reg[9]  ( .D(\shifter_0/n9841 ), .CP(clk), .Q(ow_2[9]) );
  dff_sg \shifter_0/ow_2_reg[10]  ( .D(\shifter_0/n9842 ), .CP(clk), .Q(
        ow_2[10]) );
  dff_sg \shifter_0/ow_2_reg[11]  ( .D(\shifter_0/n9843 ), .CP(clk), .Q(
        ow_2[11]) );
  dff_sg \shifter_0/ow_2_reg[12]  ( .D(\shifter_0/n9844 ), .CP(clk), .Q(
        ow_2[12]) );
  dff_sg \shifter_0/ow_2_reg[13]  ( .D(\shifter_0/n9845 ), .CP(clk), .Q(
        ow_2[13]) );
  dff_sg \shifter_0/ow_2_reg[14]  ( .D(\shifter_0/n9846 ), .CP(clk), .Q(
        ow_2[14]) );
  dff_sg \shifter_0/ow_2_reg[15]  ( .D(\shifter_0/n9847 ), .CP(clk), .Q(
        ow_2[15]) );
  dff_sg \shifter_0/ow_2_reg[16]  ( .D(\shifter_0/n9848 ), .CP(clk), .Q(
        ow_2[16]) );
  dff_sg \shifter_0/ow_2_reg[17]  ( .D(\shifter_0/n9849 ), .CP(clk), .Q(
        ow_2[17]) );
  dff_sg \shifter_0/ow_2_reg[18]  ( .D(\shifter_0/n9850 ), .CP(clk), .Q(
        ow_2[18]) );
  dff_sg \shifter_0/ow_2_reg[19]  ( .D(\shifter_0/n9851 ), .CP(clk), .Q(
        ow_2[19]) );
  dff_sg \shifter_0/ow_1_reg[0]  ( .D(\shifter_0/n9852 ), .CP(clk), .Q(ow_1[0]) );
  dff_sg \shifter_0/ow_1_reg[1]  ( .D(\shifter_0/n9853 ), .CP(clk), .Q(ow_1[1]) );
  dff_sg \shifter_0/ow_1_reg[2]  ( .D(\shifter_0/n9854 ), .CP(clk), .Q(ow_1[2]) );
  dff_sg \shifter_0/ow_1_reg[3]  ( .D(\shifter_0/n9855 ), .CP(clk), .Q(ow_1[3]) );
  dff_sg \shifter_0/ow_1_reg[4]  ( .D(\shifter_0/n9856 ), .CP(clk), .Q(ow_1[4]) );
  dff_sg \shifter_0/ow_1_reg[5]  ( .D(\shifter_0/n9857 ), .CP(clk), .Q(ow_1[5]) );
  dff_sg \shifter_0/ow_1_reg[6]  ( .D(\shifter_0/n9858 ), .CP(clk), .Q(ow_1[6]) );
  dff_sg \shifter_0/ow_1_reg[7]  ( .D(\shifter_0/n9859 ), .CP(clk), .Q(ow_1[7]) );
  dff_sg \shifter_0/ow_1_reg[8]  ( .D(\shifter_0/n9860 ), .CP(clk), .Q(ow_1[8]) );
  dff_sg \shifter_0/ow_1_reg[9]  ( .D(\shifter_0/n9861 ), .CP(clk), .Q(ow_1[9]) );
  dff_sg \shifter_0/ow_1_reg[10]  ( .D(\shifter_0/n9862 ), .CP(clk), .Q(
        ow_1[10]) );
  dff_sg \shifter_0/ow_1_reg[11]  ( .D(\shifter_0/n9863 ), .CP(clk), .Q(
        ow_1[11]) );
  dff_sg \shifter_0/ow_1_reg[12]  ( .D(\shifter_0/n9864 ), .CP(clk), .Q(
        ow_1[12]) );
  dff_sg \shifter_0/ow_1_reg[13]  ( .D(\shifter_0/n9865 ), .CP(clk), .Q(
        ow_1[13]) );
  dff_sg \shifter_0/ow_1_reg[14]  ( .D(\shifter_0/n9866 ), .CP(clk), .Q(
        ow_1[14]) );
  dff_sg \shifter_0/ow_1_reg[15]  ( .D(\shifter_0/n9867 ), .CP(clk), .Q(
        ow_1[15]) );
  dff_sg \shifter_0/ow_1_reg[16]  ( .D(\shifter_0/n9868 ), .CP(clk), .Q(
        ow_1[16]) );
  dff_sg \shifter_0/ow_1_reg[17]  ( .D(\shifter_0/n9869 ), .CP(clk), .Q(
        ow_1[17]) );
  dff_sg \shifter_0/ow_1_reg[18]  ( .D(\shifter_0/n9870 ), .CP(clk), .Q(
        ow_1[18]) );
  dff_sg \shifter_0/ow_1_reg[19]  ( .D(\shifter_0/n9871 ), .CP(clk), .Q(
        ow_1[19]) );
  dff_sg \shifter_0/ow_0_reg[0]  ( .D(\shifter_0/n9872 ), .CP(clk), .Q(ow_0[0]) );
  dff_sg \shifter_0/ow_0_reg[1]  ( .D(\shifter_0/n9873 ), .CP(clk), .Q(ow_0[1]) );
  dff_sg \shifter_0/ow_0_reg[2]  ( .D(\shifter_0/n9874 ), .CP(clk), .Q(ow_0[2]) );
  dff_sg \shifter_0/ow_0_reg[3]  ( .D(\shifter_0/n9875 ), .CP(clk), .Q(ow_0[3]) );
  dff_sg \shifter_0/ow_0_reg[4]  ( .D(\shifter_0/n9876 ), .CP(clk), .Q(ow_0[4]) );
  dff_sg \shifter_0/ow_0_reg[5]  ( .D(\shifter_0/n9877 ), .CP(clk), .Q(ow_0[5]) );
  dff_sg \shifter_0/ow_0_reg[6]  ( .D(\shifter_0/n9878 ), .CP(clk), .Q(ow_0[6]) );
  dff_sg \shifter_0/ow_0_reg[7]  ( .D(\shifter_0/n9879 ), .CP(clk), .Q(ow_0[7]) );
  dff_sg \shifter_0/ow_0_reg[8]  ( .D(\shifter_0/n9880 ), .CP(clk), .Q(ow_0[8]) );
  dff_sg \shifter_0/ow_0_reg[9]  ( .D(\shifter_0/n9881 ), .CP(clk), .Q(ow_0[9]) );
  dff_sg \shifter_0/ow_0_reg[10]  ( .D(\shifter_0/n9882 ), .CP(clk), .Q(
        ow_0[10]) );
  dff_sg \shifter_0/ow_0_reg[11]  ( .D(\shifter_0/n9883 ), .CP(clk), .Q(
        ow_0[11]) );
  dff_sg \shifter_0/ow_0_reg[12]  ( .D(\shifter_0/n9884 ), .CP(clk), .Q(
        ow_0[12]) );
  dff_sg \shifter_0/ow_0_reg[13]  ( .D(\shifter_0/n9885 ), .CP(clk), .Q(
        ow_0[13]) );
  dff_sg \shifter_0/ow_0_reg[14]  ( .D(\shifter_0/n9886 ), .CP(clk), .Q(
        ow_0[14]) );
  dff_sg \shifter_0/ow_0_reg[15]  ( .D(\shifter_0/n9887 ), .CP(clk), .Q(
        ow_0[15]) );
  dff_sg \shifter_0/ow_0_reg[16]  ( .D(\shifter_0/n9888 ), .CP(clk), .Q(
        ow_0[16]) );
  dff_sg \shifter_0/ow_0_reg[17]  ( .D(\shifter_0/n9889 ), .CP(clk), .Q(
        ow_0[17]) );
  dff_sg \shifter_0/ow_0_reg[18]  ( .D(\shifter_0/n9890 ), .CP(clk), .Q(
        ow_0[18]) );
  dff_sg \shifter_0/ow_0_reg[19]  ( .D(\shifter_0/n9891 ), .CP(clk), .Q(
        ow_0[19]) );
  dff_sg \shifter_0/oi_15_reg[0]  ( .D(\shifter_0/n9892 ), .CP(clk), .Q(
        oi_15[0]) );
  dff_sg \shifter_0/oi_15_reg[1]  ( .D(\shifter_0/n9893 ), .CP(clk), .Q(
        oi_15[1]) );
  dff_sg \shifter_0/oi_15_reg[2]  ( .D(\shifter_0/n9894 ), .CP(clk), .Q(
        oi_15[2]) );
  dff_sg \shifter_0/oi_15_reg[3]  ( .D(\shifter_0/n9895 ), .CP(clk), .Q(
        oi_15[3]) );
  dff_sg \shifter_0/oi_15_reg[4]  ( .D(\shifter_0/n9896 ), .CP(clk), .Q(
        oi_15[4]) );
  dff_sg \shifter_0/oi_15_reg[5]  ( .D(\shifter_0/n9897 ), .CP(clk), .Q(
        oi_15[5]) );
  dff_sg \shifter_0/oi_15_reg[6]  ( .D(\shifter_0/n9898 ), .CP(clk), .Q(
        oi_15[6]) );
  dff_sg \shifter_0/oi_15_reg[7]  ( .D(\shifter_0/n9899 ), .CP(clk), .Q(
        oi_15[7]) );
  dff_sg \shifter_0/oi_15_reg[8]  ( .D(\shifter_0/n9900 ), .CP(clk), .Q(
        oi_15[8]) );
  dff_sg \shifter_0/oi_15_reg[9]  ( .D(\shifter_0/n9901 ), .CP(clk), .Q(
        oi_15[9]) );
  dff_sg \shifter_0/oi_15_reg[10]  ( .D(\shifter_0/n9902 ), .CP(clk), .Q(
        oi_15[10]) );
  dff_sg \shifter_0/oi_15_reg[11]  ( .D(\shifter_0/n9903 ), .CP(clk), .Q(
        oi_15[11]) );
  dff_sg \shifter_0/oi_15_reg[12]  ( .D(\shifter_0/n9904 ), .CP(clk), .Q(
        oi_15[12]) );
  dff_sg \shifter_0/oi_15_reg[13]  ( .D(\shifter_0/n9905 ), .CP(clk), .Q(
        oi_15[13]) );
  dff_sg \shifter_0/oi_15_reg[14]  ( .D(\shifter_0/n9906 ), .CP(clk), .Q(
        oi_15[14]) );
  dff_sg \shifter_0/oi_15_reg[15]  ( .D(\shifter_0/n9907 ), .CP(clk), .Q(
        oi_15[15]) );
  dff_sg \shifter_0/oi_15_reg[16]  ( .D(\shifter_0/n9908 ), .CP(clk), .Q(
        oi_15[16]) );
  dff_sg \shifter_0/oi_15_reg[17]  ( .D(\shifter_0/n9909 ), .CP(clk), .Q(
        oi_15[17]) );
  dff_sg \shifter_0/oi_15_reg[18]  ( .D(\shifter_0/n9910 ), .CP(clk), .Q(
        oi_15[18]) );
  dff_sg \shifter_0/oi_15_reg[19]  ( .D(\shifter_0/n9911 ), .CP(clk), .Q(
        oi_15[19]) );
  dff_sg \shifter_0/oi_14_reg[0]  ( .D(\shifter_0/n9912 ), .CP(clk), .Q(
        oi_14[0]) );
  dff_sg \shifter_0/oi_14_reg[1]  ( .D(\shifter_0/n9913 ), .CP(clk), .Q(
        oi_14[1]) );
  dff_sg \shifter_0/oi_14_reg[2]  ( .D(\shifter_0/n9914 ), .CP(clk), .Q(
        oi_14[2]) );
  dff_sg \shifter_0/oi_14_reg[3]  ( .D(\shifter_0/n9915 ), .CP(clk), .Q(
        oi_14[3]) );
  dff_sg \shifter_0/oi_14_reg[4]  ( .D(\shifter_0/n9916 ), .CP(clk), .Q(
        oi_14[4]) );
  dff_sg \shifter_0/oi_14_reg[5]  ( .D(\shifter_0/n9917 ), .CP(clk), .Q(
        oi_14[5]) );
  dff_sg \shifter_0/oi_14_reg[6]  ( .D(\shifter_0/n9918 ), .CP(clk), .Q(
        oi_14[6]) );
  dff_sg \shifter_0/oi_14_reg[7]  ( .D(\shifter_0/n9919 ), .CP(clk), .Q(
        oi_14[7]) );
  dff_sg \shifter_0/oi_14_reg[8]  ( .D(\shifter_0/n9920 ), .CP(clk), .Q(
        oi_14[8]) );
  dff_sg \shifter_0/oi_14_reg[9]  ( .D(\shifter_0/n9921 ), .CP(clk), .Q(
        oi_14[9]) );
  dff_sg \shifter_0/oi_14_reg[10]  ( .D(\shifter_0/n9922 ), .CP(clk), .Q(
        oi_14[10]) );
  dff_sg \shifter_0/oi_14_reg[11]  ( .D(\shifter_0/n9923 ), .CP(clk), .Q(
        oi_14[11]) );
  dff_sg \shifter_0/oi_14_reg[12]  ( .D(\shifter_0/n9924 ), .CP(clk), .Q(
        oi_14[12]) );
  dff_sg \shifter_0/oi_14_reg[13]  ( .D(\shifter_0/n9925 ), .CP(clk), .Q(
        oi_14[13]) );
  dff_sg \shifter_0/oi_14_reg[14]  ( .D(\shifter_0/n9926 ), .CP(clk), .Q(
        oi_14[14]) );
  dff_sg \shifter_0/oi_14_reg[15]  ( .D(\shifter_0/n9927 ), .CP(clk), .Q(
        oi_14[15]) );
  dff_sg \shifter_0/oi_14_reg[16]  ( .D(\shifter_0/n9928 ), .CP(clk), .Q(
        oi_14[16]) );
  dff_sg \shifter_0/oi_14_reg[17]  ( .D(\shifter_0/n9929 ), .CP(clk), .Q(
        oi_14[17]) );
  dff_sg \shifter_0/oi_14_reg[18]  ( .D(\shifter_0/n9930 ), .CP(clk), .Q(
        oi_14[18]) );
  dff_sg \shifter_0/oi_14_reg[19]  ( .D(\shifter_0/n9931 ), .CP(clk), .Q(
        oi_14[19]) );
  dff_sg \shifter_0/oi_13_reg[0]  ( .D(\shifter_0/n9932 ), .CP(clk), .Q(
        oi_13[0]) );
  dff_sg \shifter_0/oi_13_reg[1]  ( .D(\shifter_0/n9933 ), .CP(clk), .Q(
        oi_13[1]) );
  dff_sg \shifter_0/oi_13_reg[2]  ( .D(\shifter_0/n9934 ), .CP(clk), .Q(
        oi_13[2]) );
  dff_sg \shifter_0/oi_13_reg[3]  ( .D(\shifter_0/n9935 ), .CP(clk), .Q(
        oi_13[3]) );
  dff_sg \shifter_0/oi_13_reg[4]  ( .D(\shifter_0/n9936 ), .CP(clk), .Q(
        oi_13[4]) );
  dff_sg \shifter_0/oi_13_reg[5]  ( .D(\shifter_0/n9937 ), .CP(clk), .Q(
        oi_13[5]) );
  dff_sg \shifter_0/oi_13_reg[6]  ( .D(\shifter_0/n9938 ), .CP(clk), .Q(
        oi_13[6]) );
  dff_sg \shifter_0/oi_13_reg[7]  ( .D(\shifter_0/n9939 ), .CP(clk), .Q(
        oi_13[7]) );
  dff_sg \shifter_0/oi_13_reg[8]  ( .D(\shifter_0/n9940 ), .CP(clk), .Q(
        oi_13[8]) );
  dff_sg \shifter_0/oi_13_reg[9]  ( .D(\shifter_0/n9941 ), .CP(clk), .Q(
        oi_13[9]) );
  dff_sg \shifter_0/oi_13_reg[10]  ( .D(\shifter_0/n9942 ), .CP(clk), .Q(
        oi_13[10]) );
  dff_sg \shifter_0/oi_13_reg[11]  ( .D(\shifter_0/n9943 ), .CP(clk), .Q(
        oi_13[11]) );
  dff_sg \shifter_0/oi_13_reg[12]  ( .D(\shifter_0/n9944 ), .CP(clk), .Q(
        oi_13[12]) );
  dff_sg \shifter_0/oi_13_reg[13]  ( .D(\shifter_0/n9945 ), .CP(clk), .Q(
        oi_13[13]) );
  dff_sg \shifter_0/oi_13_reg[14]  ( .D(\shifter_0/n9946 ), .CP(clk), .Q(
        oi_13[14]) );
  dff_sg \shifter_0/oi_13_reg[15]  ( .D(\shifter_0/n9947 ), .CP(clk), .Q(
        oi_13[15]) );
  dff_sg \shifter_0/oi_13_reg[16]  ( .D(\shifter_0/n9948 ), .CP(clk), .Q(
        oi_13[16]) );
  dff_sg \shifter_0/oi_13_reg[17]  ( .D(\shifter_0/n9949 ), .CP(clk), .Q(
        oi_13[17]) );
  dff_sg \shifter_0/oi_13_reg[18]  ( .D(\shifter_0/n9950 ), .CP(clk), .Q(
        oi_13[18]) );
  dff_sg \shifter_0/oi_13_reg[19]  ( .D(\shifter_0/n9951 ), .CP(clk), .Q(
        oi_13[19]) );
  dff_sg \shifter_0/oi_12_reg[0]  ( .D(\shifter_0/n9952 ), .CP(clk), .Q(
        oi_12[0]) );
  dff_sg \shifter_0/oi_12_reg[1]  ( .D(\shifter_0/n9953 ), .CP(clk), .Q(
        oi_12[1]) );
  dff_sg \shifter_0/oi_12_reg[2]  ( .D(\shifter_0/n9954 ), .CP(clk), .Q(
        oi_12[2]) );
  dff_sg \shifter_0/oi_12_reg[3]  ( .D(\shifter_0/n9955 ), .CP(clk), .Q(
        oi_12[3]) );
  dff_sg \shifter_0/oi_12_reg[4]  ( .D(\shifter_0/n9956 ), .CP(clk), .Q(
        oi_12[4]) );
  dff_sg \shifter_0/oi_12_reg[5]  ( .D(\shifter_0/n9957 ), .CP(clk), .Q(
        oi_12[5]) );
  dff_sg \shifter_0/oi_12_reg[6]  ( .D(\shifter_0/n9958 ), .CP(clk), .Q(
        oi_12[6]) );
  dff_sg \shifter_0/oi_12_reg[7]  ( .D(\shifter_0/n9959 ), .CP(clk), .Q(
        oi_12[7]) );
  dff_sg \shifter_0/oi_12_reg[8]  ( .D(\shifter_0/n9960 ), .CP(clk), .Q(
        oi_12[8]) );
  dff_sg \shifter_0/oi_12_reg[9]  ( .D(\shifter_0/n9961 ), .CP(clk), .Q(
        oi_12[9]) );
  dff_sg \shifter_0/oi_12_reg[10]  ( .D(\shifter_0/n9962 ), .CP(clk), .Q(
        oi_12[10]) );
  dff_sg \shifter_0/oi_12_reg[11]  ( .D(\shifter_0/n9963 ), .CP(clk), .Q(
        oi_12[11]) );
  dff_sg \shifter_0/oi_12_reg[12]  ( .D(\shifter_0/n9964 ), .CP(clk), .Q(
        oi_12[12]) );
  dff_sg \shifter_0/oi_12_reg[13]  ( .D(\shifter_0/n9965 ), .CP(clk), .Q(
        oi_12[13]) );
  dff_sg \shifter_0/oi_12_reg[14]  ( .D(\shifter_0/n9966 ), .CP(clk), .Q(
        oi_12[14]) );
  dff_sg \shifter_0/oi_12_reg[15]  ( .D(\shifter_0/n9967 ), .CP(clk), .Q(
        oi_12[15]) );
  dff_sg \shifter_0/oi_12_reg[16]  ( .D(\shifter_0/n9968 ), .CP(clk), .Q(
        oi_12[16]) );
  dff_sg \shifter_0/oi_12_reg[17]  ( .D(\shifter_0/n9969 ), .CP(clk), .Q(
        oi_12[17]) );
  dff_sg \shifter_0/oi_12_reg[18]  ( .D(\shifter_0/n9970 ), .CP(clk), .Q(
        oi_12[18]) );
  dff_sg \shifter_0/oi_12_reg[19]  ( .D(\shifter_0/n9971 ), .CP(clk), .Q(
        oi_12[19]) );
  dff_sg \shifter_0/oi_11_reg[0]  ( .D(\shifter_0/n9972 ), .CP(clk), .Q(
        oi_11[0]) );
  dff_sg \shifter_0/oi_11_reg[1]  ( .D(\shifter_0/n9973 ), .CP(clk), .Q(
        oi_11[1]) );
  dff_sg \shifter_0/oi_11_reg[2]  ( .D(\shifter_0/n9974 ), .CP(clk), .Q(
        oi_11[2]) );
  dff_sg \shifter_0/oi_11_reg[3]  ( .D(\shifter_0/n9975 ), .CP(clk), .Q(
        oi_11[3]) );
  dff_sg \shifter_0/oi_11_reg[4]  ( .D(\shifter_0/n9976 ), .CP(clk), .Q(
        oi_11[4]) );
  dff_sg \shifter_0/oi_11_reg[5]  ( .D(\shifter_0/n9977 ), .CP(clk), .Q(
        oi_11[5]) );
  dff_sg \shifter_0/oi_11_reg[6]  ( .D(\shifter_0/n9978 ), .CP(clk), .Q(
        oi_11[6]) );
  dff_sg \shifter_0/oi_11_reg[7]  ( .D(\shifter_0/n9979 ), .CP(clk), .Q(
        oi_11[7]) );
  dff_sg \shifter_0/oi_11_reg[8]  ( .D(\shifter_0/n9980 ), .CP(clk), .Q(
        oi_11[8]) );
  dff_sg \shifter_0/oi_11_reg[9]  ( .D(\shifter_0/n9981 ), .CP(clk), .Q(
        oi_11[9]) );
  dff_sg \shifter_0/oi_11_reg[10]  ( .D(\shifter_0/n9982 ), .CP(clk), .Q(
        oi_11[10]) );
  dff_sg \shifter_0/oi_11_reg[11]  ( .D(\shifter_0/n9983 ), .CP(clk), .Q(
        oi_11[11]) );
  dff_sg \shifter_0/oi_11_reg[12]  ( .D(\shifter_0/n9984 ), .CP(clk), .Q(
        oi_11[12]) );
  dff_sg \shifter_0/oi_11_reg[13]  ( .D(\shifter_0/n9985 ), .CP(clk), .Q(
        oi_11[13]) );
  dff_sg \shifter_0/oi_11_reg[14]  ( .D(\shifter_0/n9986 ), .CP(clk), .Q(
        oi_11[14]) );
  dff_sg \shifter_0/oi_11_reg[15]  ( .D(\shifter_0/n9987 ), .CP(clk), .Q(
        oi_11[15]) );
  dff_sg \shifter_0/oi_11_reg[16]  ( .D(\shifter_0/n9988 ), .CP(clk), .Q(
        oi_11[16]) );
  dff_sg \shifter_0/oi_11_reg[17]  ( .D(\shifter_0/n9989 ), .CP(clk), .Q(
        oi_11[17]) );
  dff_sg \shifter_0/oi_11_reg[18]  ( .D(\shifter_0/n9990 ), .CP(clk), .Q(
        oi_11[18]) );
  dff_sg \shifter_0/oi_11_reg[19]  ( .D(\shifter_0/n9991 ), .CP(clk), .Q(
        oi_11[19]) );
  dff_sg \shifter_0/oi_10_reg[0]  ( .D(\shifter_0/n9992 ), .CP(clk), .Q(
        oi_10[0]) );
  dff_sg \shifter_0/oi_10_reg[1]  ( .D(\shifter_0/n9993 ), .CP(clk), .Q(
        oi_10[1]) );
  dff_sg \shifter_0/oi_10_reg[2]  ( .D(\shifter_0/n9994 ), .CP(clk), .Q(
        oi_10[2]) );
  dff_sg \shifter_0/oi_10_reg[3]  ( .D(\shifter_0/n9995 ), .CP(clk), .Q(
        oi_10[3]) );
  dff_sg \shifter_0/oi_10_reg[4]  ( .D(\shifter_0/n9996 ), .CP(clk), .Q(
        oi_10[4]) );
  dff_sg \shifter_0/oi_10_reg[5]  ( .D(\shifter_0/n9997 ), .CP(clk), .Q(
        oi_10[5]) );
  dff_sg \shifter_0/oi_10_reg[6]  ( .D(\shifter_0/n9998 ), .CP(clk), .Q(
        oi_10[6]) );
  dff_sg \shifter_0/oi_10_reg[7]  ( .D(\shifter_0/n9999 ), .CP(clk), .Q(
        oi_10[7]) );
  dff_sg \shifter_0/oi_10_reg[8]  ( .D(\shifter_0/n10000 ), .CP(clk), .Q(
        oi_10[8]) );
  dff_sg \shifter_0/oi_10_reg[9]  ( .D(\shifter_0/n10001 ), .CP(clk), .Q(
        oi_10[9]) );
  dff_sg \shifter_0/oi_10_reg[10]  ( .D(\shifter_0/n10002 ), .CP(clk), .Q(
        oi_10[10]) );
  dff_sg \shifter_0/oi_10_reg[11]  ( .D(\shifter_0/n10003 ), .CP(clk), .Q(
        oi_10[11]) );
  dff_sg \shifter_0/oi_10_reg[12]  ( .D(\shifter_0/n10004 ), .CP(clk), .Q(
        oi_10[12]) );
  dff_sg \shifter_0/oi_10_reg[13]  ( .D(\shifter_0/n10005 ), .CP(clk), .Q(
        oi_10[13]) );
  dff_sg \shifter_0/oi_10_reg[14]  ( .D(\shifter_0/n10006 ), .CP(clk), .Q(
        oi_10[14]) );
  dff_sg \shifter_0/oi_10_reg[15]  ( .D(\shifter_0/n10007 ), .CP(clk), .Q(
        oi_10[15]) );
  dff_sg \shifter_0/oi_10_reg[16]  ( .D(\shifter_0/n10008 ), .CP(clk), .Q(
        oi_10[16]) );
  dff_sg \shifter_0/oi_10_reg[17]  ( .D(\shifter_0/n10009 ), .CP(clk), .Q(
        oi_10[17]) );
  dff_sg \shifter_0/oi_10_reg[18]  ( .D(\shifter_0/n10010 ), .CP(clk), .Q(
        oi_10[18]) );
  dff_sg \shifter_0/oi_10_reg[19]  ( .D(\shifter_0/n10011 ), .CP(clk), .Q(
        oi_10[19]) );
  dff_sg \shifter_0/oi_9_reg[0]  ( .D(\shifter_0/n10012 ), .CP(clk), .Q(
        oi_9[0]) );
  dff_sg \shifter_0/oi_9_reg[1]  ( .D(\shifter_0/n10013 ), .CP(clk), .Q(
        oi_9[1]) );
  dff_sg \shifter_0/oi_9_reg[2]  ( .D(\shifter_0/n10014 ), .CP(clk), .Q(
        oi_9[2]) );
  dff_sg \shifter_0/oi_9_reg[3]  ( .D(\shifter_0/n10015 ), .CP(clk), .Q(
        oi_9[3]) );
  dff_sg \shifter_0/oi_9_reg[4]  ( .D(\shifter_0/n10016 ), .CP(clk), .Q(
        oi_9[4]) );
  dff_sg \shifter_0/oi_9_reg[5]  ( .D(\shifter_0/n10017 ), .CP(clk), .Q(
        oi_9[5]) );
  dff_sg \shifter_0/oi_9_reg[6]  ( .D(\shifter_0/n10018 ), .CP(clk), .Q(
        oi_9[6]) );
  dff_sg \shifter_0/oi_9_reg[7]  ( .D(\shifter_0/n10019 ), .CP(clk), .Q(
        oi_9[7]) );
  dff_sg \shifter_0/oi_9_reg[8]  ( .D(\shifter_0/n10020 ), .CP(clk), .Q(
        oi_9[8]) );
  dff_sg \shifter_0/oi_9_reg[9]  ( .D(\shifter_0/n10021 ), .CP(clk), .Q(
        oi_9[9]) );
  dff_sg \shifter_0/oi_9_reg[10]  ( .D(\shifter_0/n10022 ), .CP(clk), .Q(
        oi_9[10]) );
  dff_sg \shifter_0/oi_9_reg[11]  ( .D(\shifter_0/n10023 ), .CP(clk), .Q(
        oi_9[11]) );
  dff_sg \shifter_0/oi_9_reg[12]  ( .D(\shifter_0/n10024 ), .CP(clk), .Q(
        oi_9[12]) );
  dff_sg \shifter_0/oi_9_reg[13]  ( .D(\shifter_0/n10025 ), .CP(clk), .Q(
        oi_9[13]) );
  dff_sg \shifter_0/oi_9_reg[14]  ( .D(\shifter_0/n10026 ), .CP(clk), .Q(
        oi_9[14]) );
  dff_sg \shifter_0/oi_9_reg[15]  ( .D(\shifter_0/n10027 ), .CP(clk), .Q(
        oi_9[15]) );
  dff_sg \shifter_0/oi_9_reg[16]  ( .D(\shifter_0/n10028 ), .CP(clk), .Q(
        oi_9[16]) );
  dff_sg \shifter_0/oi_9_reg[17]  ( .D(\shifter_0/n10029 ), .CP(clk), .Q(
        oi_9[17]) );
  dff_sg \shifter_0/oi_9_reg[18]  ( .D(\shifter_0/n10030 ), .CP(clk), .Q(
        oi_9[18]) );
  dff_sg \shifter_0/oi_9_reg[19]  ( .D(\shifter_0/n10031 ), .CP(clk), .Q(
        oi_9[19]) );
  dff_sg \shifter_0/oi_8_reg[0]  ( .D(\shifter_0/n10032 ), .CP(clk), .Q(
        oi_8[0]) );
  dff_sg \shifter_0/oi_8_reg[1]  ( .D(\shifter_0/n10033 ), .CP(clk), .Q(
        oi_8[1]) );
  dff_sg \shifter_0/oi_8_reg[2]  ( .D(\shifter_0/n10034 ), .CP(clk), .Q(
        oi_8[2]) );
  dff_sg \shifter_0/oi_8_reg[3]  ( .D(\shifter_0/n10035 ), .CP(clk), .Q(
        oi_8[3]) );
  dff_sg \shifter_0/oi_8_reg[4]  ( .D(\shifter_0/n10036 ), .CP(clk), .Q(
        oi_8[4]) );
  dff_sg \shifter_0/oi_8_reg[5]  ( .D(\shifter_0/n10037 ), .CP(clk), .Q(
        oi_8[5]) );
  dff_sg \shifter_0/oi_8_reg[6]  ( .D(\shifter_0/n10038 ), .CP(clk), .Q(
        oi_8[6]) );
  dff_sg \shifter_0/oi_8_reg[7]  ( .D(\shifter_0/n10039 ), .CP(clk), .Q(
        oi_8[7]) );
  dff_sg \shifter_0/oi_8_reg[8]  ( .D(\shifter_0/n10040 ), .CP(clk), .Q(
        oi_8[8]) );
  dff_sg \shifter_0/oi_8_reg[9]  ( .D(\shifter_0/n10041 ), .CP(clk), .Q(
        oi_8[9]) );
  dff_sg \shifter_0/oi_8_reg[10]  ( .D(\shifter_0/n10042 ), .CP(clk), .Q(
        oi_8[10]) );
  dff_sg \shifter_0/oi_8_reg[11]  ( .D(\shifter_0/n10043 ), .CP(clk), .Q(
        oi_8[11]) );
  dff_sg \shifter_0/oi_8_reg[12]  ( .D(\shifter_0/n10044 ), .CP(clk), .Q(
        oi_8[12]) );
  dff_sg \shifter_0/oi_8_reg[13]  ( .D(\shifter_0/n10045 ), .CP(clk), .Q(
        oi_8[13]) );
  dff_sg \shifter_0/oi_8_reg[14]  ( .D(\shifter_0/n10046 ), .CP(clk), .Q(
        oi_8[14]) );
  dff_sg \shifter_0/oi_8_reg[15]  ( .D(\shifter_0/n10047 ), .CP(clk), .Q(
        oi_8[15]) );
  dff_sg \shifter_0/oi_8_reg[16]  ( .D(\shifter_0/n10048 ), .CP(clk), .Q(
        oi_8[16]) );
  dff_sg \shifter_0/oi_8_reg[17]  ( .D(\shifter_0/n10049 ), .CP(clk), .Q(
        oi_8[17]) );
  dff_sg \shifter_0/oi_8_reg[18]  ( .D(\shifter_0/n10050 ), .CP(clk), .Q(
        oi_8[18]) );
  dff_sg \shifter_0/oi_8_reg[19]  ( .D(\shifter_0/n10051 ), .CP(clk), .Q(
        oi_8[19]) );
  dff_sg \shifter_0/oi_7_reg[0]  ( .D(\shifter_0/n10052 ), .CP(clk), .Q(
        oi_7[0]) );
  dff_sg \shifter_0/oi_7_reg[1]  ( .D(\shifter_0/n10053 ), .CP(clk), .Q(
        oi_7[1]) );
  dff_sg \shifter_0/oi_7_reg[2]  ( .D(\shifter_0/n10054 ), .CP(clk), .Q(
        oi_7[2]) );
  dff_sg \shifter_0/oi_7_reg[3]  ( .D(\shifter_0/n10055 ), .CP(clk), .Q(
        oi_7[3]) );
  dff_sg \shifter_0/oi_7_reg[4]  ( .D(\shifter_0/n10056 ), .CP(clk), .Q(
        oi_7[4]) );
  dff_sg \shifter_0/oi_7_reg[5]  ( .D(\shifter_0/n10057 ), .CP(clk), .Q(
        oi_7[5]) );
  dff_sg \shifter_0/oi_7_reg[6]  ( .D(\shifter_0/n10058 ), .CP(clk), .Q(
        oi_7[6]) );
  dff_sg \shifter_0/oi_7_reg[7]  ( .D(\shifter_0/n10059 ), .CP(clk), .Q(
        oi_7[7]) );
  dff_sg \shifter_0/oi_7_reg[8]  ( .D(\shifter_0/n10060 ), .CP(clk), .Q(
        oi_7[8]) );
  dff_sg \shifter_0/oi_7_reg[9]  ( .D(\shifter_0/n10061 ), .CP(clk), .Q(
        oi_7[9]) );
  dff_sg \shifter_0/oi_7_reg[10]  ( .D(\shifter_0/n10062 ), .CP(clk), .Q(
        oi_7[10]) );
  dff_sg \shifter_0/oi_7_reg[11]  ( .D(\shifter_0/n10063 ), .CP(clk), .Q(
        oi_7[11]) );
  dff_sg \shifter_0/oi_7_reg[12]  ( .D(\shifter_0/n10064 ), .CP(clk), .Q(
        oi_7[12]) );
  dff_sg \shifter_0/oi_7_reg[13]  ( .D(\shifter_0/n10065 ), .CP(clk), .Q(
        oi_7[13]) );
  dff_sg \shifter_0/oi_7_reg[14]  ( .D(\shifter_0/n10066 ), .CP(clk), .Q(
        oi_7[14]) );
  dff_sg \shifter_0/oi_7_reg[15]  ( .D(\shifter_0/n10067 ), .CP(clk), .Q(
        oi_7[15]) );
  dff_sg \shifter_0/oi_7_reg[16]  ( .D(\shifter_0/n10068 ), .CP(clk), .Q(
        oi_7[16]) );
  dff_sg \shifter_0/oi_7_reg[17]  ( .D(\shifter_0/n10069 ), .CP(clk), .Q(
        oi_7[17]) );
  dff_sg \shifter_0/oi_7_reg[18]  ( .D(\shifter_0/n10070 ), .CP(clk), .Q(
        oi_7[18]) );
  dff_sg \shifter_0/oi_7_reg[19]  ( .D(\shifter_0/n10071 ), .CP(clk), .Q(
        oi_7[19]) );
  dff_sg \shifter_0/oi_6_reg[0]  ( .D(\shifter_0/n10072 ), .CP(clk), .Q(
        oi_6[0]) );
  dff_sg \shifter_0/oi_6_reg[1]  ( .D(\shifter_0/n10073 ), .CP(clk), .Q(
        oi_6[1]) );
  dff_sg \shifter_0/oi_6_reg[2]  ( .D(\shifter_0/n10074 ), .CP(clk), .Q(
        oi_6[2]) );
  dff_sg \shifter_0/oi_6_reg[3]  ( .D(\shifter_0/n10075 ), .CP(clk), .Q(
        oi_6[3]) );
  dff_sg \shifter_0/oi_6_reg[4]  ( .D(\shifter_0/n10076 ), .CP(clk), .Q(
        oi_6[4]) );
  dff_sg \shifter_0/oi_6_reg[5]  ( .D(\shifter_0/n10077 ), .CP(clk), .Q(
        oi_6[5]) );
  dff_sg \shifter_0/oi_6_reg[6]  ( .D(\shifter_0/n10078 ), .CP(clk), .Q(
        oi_6[6]) );
  dff_sg \shifter_0/oi_6_reg[7]  ( .D(\shifter_0/n10079 ), .CP(clk), .Q(
        oi_6[7]) );
  dff_sg \shifter_0/oi_6_reg[8]  ( .D(\shifter_0/n10080 ), .CP(clk), .Q(
        oi_6[8]) );
  dff_sg \shifter_0/oi_6_reg[9]  ( .D(\shifter_0/n10081 ), .CP(clk), .Q(
        oi_6[9]) );
  dff_sg \shifter_0/oi_6_reg[10]  ( .D(\shifter_0/n10082 ), .CP(clk), .Q(
        oi_6[10]) );
  dff_sg \shifter_0/oi_6_reg[11]  ( .D(\shifter_0/n10083 ), .CP(clk), .Q(
        oi_6[11]) );
  dff_sg \shifter_0/oi_6_reg[12]  ( .D(\shifter_0/n10084 ), .CP(clk), .Q(
        oi_6[12]) );
  dff_sg \shifter_0/oi_6_reg[13]  ( .D(\shifter_0/n10085 ), .CP(clk), .Q(
        oi_6[13]) );
  dff_sg \shifter_0/oi_6_reg[14]  ( .D(\shifter_0/n10086 ), .CP(clk), .Q(
        oi_6[14]) );
  dff_sg \shifter_0/oi_6_reg[15]  ( .D(\shifter_0/n10087 ), .CP(clk), .Q(
        oi_6[15]) );
  dff_sg \shifter_0/oi_6_reg[16]  ( .D(\shifter_0/n10088 ), .CP(clk), .Q(
        oi_6[16]) );
  dff_sg \shifter_0/oi_6_reg[17]  ( .D(\shifter_0/n10089 ), .CP(clk), .Q(
        oi_6[17]) );
  dff_sg \shifter_0/oi_6_reg[18]  ( .D(\shifter_0/n10090 ), .CP(clk), .Q(
        oi_6[18]) );
  dff_sg \shifter_0/oi_6_reg[19]  ( .D(\shifter_0/n10091 ), .CP(clk), .Q(
        oi_6[19]) );
  dff_sg \shifter_0/oi_5_reg[0]  ( .D(\shifter_0/n10092 ), .CP(clk), .Q(
        oi_5[0]) );
  dff_sg \shifter_0/oi_5_reg[1]  ( .D(\shifter_0/n10093 ), .CP(clk), .Q(
        oi_5[1]) );
  dff_sg \shifter_0/oi_5_reg[2]  ( .D(\shifter_0/n10094 ), .CP(clk), .Q(
        oi_5[2]) );
  dff_sg \shifter_0/oi_5_reg[3]  ( .D(\shifter_0/n10095 ), .CP(clk), .Q(
        oi_5[3]) );
  dff_sg \shifter_0/oi_5_reg[4]  ( .D(\shifter_0/n10096 ), .CP(clk), .Q(
        oi_5[4]) );
  dff_sg \shifter_0/oi_5_reg[5]  ( .D(\shifter_0/n10097 ), .CP(clk), .Q(
        oi_5[5]) );
  dff_sg \shifter_0/oi_5_reg[6]  ( .D(\shifter_0/n10098 ), .CP(clk), .Q(
        oi_5[6]) );
  dff_sg \shifter_0/oi_5_reg[7]  ( .D(\shifter_0/n10099 ), .CP(clk), .Q(
        oi_5[7]) );
  dff_sg \shifter_0/oi_5_reg[8]  ( .D(\shifter_0/n10100 ), .CP(clk), .Q(
        oi_5[8]) );
  dff_sg \shifter_0/oi_5_reg[9]  ( .D(\shifter_0/n10101 ), .CP(clk), .Q(
        oi_5[9]) );
  dff_sg \shifter_0/oi_5_reg[10]  ( .D(\shifter_0/n10102 ), .CP(clk), .Q(
        oi_5[10]) );
  dff_sg \shifter_0/oi_5_reg[11]  ( .D(\shifter_0/n10103 ), .CP(clk), .Q(
        oi_5[11]) );
  dff_sg \shifter_0/oi_5_reg[12]  ( .D(\shifter_0/n10104 ), .CP(clk), .Q(
        oi_5[12]) );
  dff_sg \shifter_0/oi_5_reg[13]  ( .D(\shifter_0/n10105 ), .CP(clk), .Q(
        oi_5[13]) );
  dff_sg \shifter_0/oi_5_reg[14]  ( .D(\shifter_0/n10106 ), .CP(clk), .Q(
        oi_5[14]) );
  dff_sg \shifter_0/oi_5_reg[15]  ( .D(\shifter_0/n10107 ), .CP(clk), .Q(
        oi_5[15]) );
  dff_sg \shifter_0/oi_5_reg[16]  ( .D(\shifter_0/n10108 ), .CP(clk), .Q(
        oi_5[16]) );
  dff_sg \shifter_0/oi_5_reg[17]  ( .D(\shifter_0/n10109 ), .CP(clk), .Q(
        oi_5[17]) );
  dff_sg \shifter_0/oi_5_reg[18]  ( .D(\shifter_0/n10110 ), .CP(clk), .Q(
        oi_5[18]) );
  dff_sg \shifter_0/oi_5_reg[19]  ( .D(\shifter_0/n10111 ), .CP(clk), .Q(
        oi_5[19]) );
  dff_sg \shifter_0/oi_4_reg[0]  ( .D(\shifter_0/n10112 ), .CP(clk), .Q(
        oi_4[0]) );
  dff_sg \shifter_0/oi_4_reg[1]  ( .D(\shifter_0/n10113 ), .CP(clk), .Q(
        oi_4[1]) );
  dff_sg \shifter_0/oi_4_reg[2]  ( .D(\shifter_0/n10114 ), .CP(clk), .Q(
        oi_4[2]) );
  dff_sg \shifter_0/oi_4_reg[3]  ( .D(\shifter_0/n10115 ), .CP(clk), .Q(
        oi_4[3]) );
  dff_sg \shifter_0/oi_4_reg[4]  ( .D(\shifter_0/n10116 ), .CP(clk), .Q(
        oi_4[4]) );
  dff_sg \shifter_0/oi_4_reg[5]  ( .D(\shifter_0/n10117 ), .CP(clk), .Q(
        oi_4[5]) );
  dff_sg \shifter_0/oi_4_reg[6]  ( .D(\shifter_0/n10118 ), .CP(clk), .Q(
        oi_4[6]) );
  dff_sg \shifter_0/oi_4_reg[7]  ( .D(\shifter_0/n10119 ), .CP(clk), .Q(
        oi_4[7]) );
  dff_sg \shifter_0/oi_4_reg[8]  ( .D(\shifter_0/n10120 ), .CP(clk), .Q(
        oi_4[8]) );
  dff_sg \shifter_0/oi_4_reg[9]  ( .D(\shifter_0/n10121 ), .CP(clk), .Q(
        oi_4[9]) );
  dff_sg \shifter_0/oi_4_reg[10]  ( .D(\shifter_0/n10122 ), .CP(clk), .Q(
        oi_4[10]) );
  dff_sg \shifter_0/oi_4_reg[11]  ( .D(\shifter_0/n10123 ), .CP(clk), .Q(
        oi_4[11]) );
  dff_sg \shifter_0/oi_4_reg[12]  ( .D(\shifter_0/n10124 ), .CP(clk), .Q(
        oi_4[12]) );
  dff_sg \shifter_0/oi_4_reg[13]  ( .D(\shifter_0/n10125 ), .CP(clk), .Q(
        oi_4[13]) );
  dff_sg \shifter_0/oi_4_reg[14]  ( .D(\shifter_0/n10126 ), .CP(clk), .Q(
        oi_4[14]) );
  dff_sg \shifter_0/oi_4_reg[15]  ( .D(\shifter_0/n10127 ), .CP(clk), .Q(
        oi_4[15]) );
  dff_sg \shifter_0/oi_4_reg[16]  ( .D(\shifter_0/n10128 ), .CP(clk), .Q(
        oi_4[16]) );
  dff_sg \shifter_0/oi_4_reg[17]  ( .D(\shifter_0/n10129 ), .CP(clk), .Q(
        oi_4[17]) );
  dff_sg \shifter_0/oi_4_reg[18]  ( .D(\shifter_0/n10130 ), .CP(clk), .Q(
        oi_4[18]) );
  dff_sg \shifter_0/oi_4_reg[19]  ( .D(\shifter_0/n10131 ), .CP(clk), .Q(
        oi_4[19]) );
  dff_sg \shifter_0/oi_3_reg[0]  ( .D(\shifter_0/n10132 ), .CP(clk), .Q(
        oi_3[0]) );
  dff_sg \shifter_0/oi_3_reg[1]  ( .D(\shifter_0/n10133 ), .CP(clk), .Q(
        oi_3[1]) );
  dff_sg \shifter_0/oi_3_reg[2]  ( .D(\shifter_0/n10134 ), .CP(clk), .Q(
        oi_3[2]) );
  dff_sg \shifter_0/oi_3_reg[3]  ( .D(\shifter_0/n10135 ), .CP(clk), .Q(
        oi_3[3]) );
  dff_sg \shifter_0/oi_3_reg[4]  ( .D(\shifter_0/n10136 ), .CP(clk), .Q(
        oi_3[4]) );
  dff_sg \shifter_0/oi_3_reg[5]  ( .D(\shifter_0/n10137 ), .CP(clk), .Q(
        oi_3[5]) );
  dff_sg \shifter_0/oi_3_reg[6]  ( .D(\shifter_0/n10138 ), .CP(clk), .Q(
        oi_3[6]) );
  dff_sg \shifter_0/oi_3_reg[7]  ( .D(\shifter_0/n10139 ), .CP(clk), .Q(
        oi_3[7]) );
  dff_sg \shifter_0/oi_3_reg[8]  ( .D(\shifter_0/n10140 ), .CP(clk), .Q(
        oi_3[8]) );
  dff_sg \shifter_0/oi_3_reg[9]  ( .D(\shifter_0/n10141 ), .CP(clk), .Q(
        oi_3[9]) );
  dff_sg \shifter_0/oi_3_reg[10]  ( .D(\shifter_0/n10142 ), .CP(clk), .Q(
        oi_3[10]) );
  dff_sg \shifter_0/oi_3_reg[11]  ( .D(\shifter_0/n10143 ), .CP(clk), .Q(
        oi_3[11]) );
  dff_sg \shifter_0/oi_3_reg[12]  ( .D(\shifter_0/n10144 ), .CP(clk), .Q(
        oi_3[12]) );
  dff_sg \shifter_0/oi_3_reg[13]  ( .D(\shifter_0/n10145 ), .CP(clk), .Q(
        oi_3[13]) );
  dff_sg \shifter_0/oi_3_reg[14]  ( .D(\shifter_0/n10146 ), .CP(clk), .Q(
        oi_3[14]) );
  dff_sg \shifter_0/oi_3_reg[15]  ( .D(\shifter_0/n10147 ), .CP(clk), .Q(
        oi_3[15]) );
  dff_sg \shifter_0/oi_3_reg[16]  ( .D(\shifter_0/n10148 ), .CP(clk), .Q(
        oi_3[16]) );
  dff_sg \shifter_0/oi_3_reg[17]  ( .D(\shifter_0/n10149 ), .CP(clk), .Q(
        oi_3[17]) );
  dff_sg \shifter_0/oi_3_reg[18]  ( .D(\shifter_0/n10150 ), .CP(clk), .Q(
        oi_3[18]) );
  dff_sg \shifter_0/oi_3_reg[19]  ( .D(\shifter_0/n10151 ), .CP(clk), .Q(
        oi_3[19]) );
  dff_sg \shifter_0/oi_2_reg[0]  ( .D(\shifter_0/n10152 ), .CP(clk), .Q(
        oi_2[0]) );
  dff_sg \shifter_0/oi_2_reg[1]  ( .D(\shifter_0/n10153 ), .CP(clk), .Q(
        oi_2[1]) );
  dff_sg \shifter_0/oi_2_reg[2]  ( .D(\shifter_0/n10154 ), .CP(clk), .Q(
        oi_2[2]) );
  dff_sg \shifter_0/oi_2_reg[3]  ( .D(\shifter_0/n10155 ), .CP(clk), .Q(
        oi_2[3]) );
  dff_sg \shifter_0/oi_2_reg[4]  ( .D(\shifter_0/n10156 ), .CP(clk), .Q(
        oi_2[4]) );
  dff_sg \shifter_0/oi_2_reg[5]  ( .D(\shifter_0/n10157 ), .CP(clk), .Q(
        oi_2[5]) );
  dff_sg \shifter_0/oi_2_reg[6]  ( .D(\shifter_0/n10158 ), .CP(clk), .Q(
        oi_2[6]) );
  dff_sg \shifter_0/oi_2_reg[7]  ( .D(\shifter_0/n10159 ), .CP(clk), .Q(
        oi_2[7]) );
  dff_sg \shifter_0/oi_2_reg[8]  ( .D(\shifter_0/n10160 ), .CP(clk), .Q(
        oi_2[8]) );
  dff_sg \shifter_0/oi_2_reg[9]  ( .D(\shifter_0/n10161 ), .CP(clk), .Q(
        oi_2[9]) );
  dff_sg \shifter_0/oi_2_reg[10]  ( .D(\shifter_0/n10162 ), .CP(clk), .Q(
        oi_2[10]) );
  dff_sg \shifter_0/oi_2_reg[11]  ( .D(\shifter_0/n10163 ), .CP(clk), .Q(
        oi_2[11]) );
  dff_sg \shifter_0/oi_2_reg[12]  ( .D(\shifter_0/n10164 ), .CP(clk), .Q(
        oi_2[12]) );
  dff_sg \shifter_0/oi_2_reg[13]  ( .D(\shifter_0/n10165 ), .CP(clk), .Q(
        oi_2[13]) );
  dff_sg \shifter_0/oi_2_reg[14]  ( .D(\shifter_0/n10166 ), .CP(clk), .Q(
        oi_2[14]) );
  dff_sg \shifter_0/oi_2_reg[15]  ( .D(\shifter_0/n10167 ), .CP(clk), .Q(
        oi_2[15]) );
  dff_sg \shifter_0/oi_2_reg[16]  ( .D(\shifter_0/n10168 ), .CP(clk), .Q(
        oi_2[16]) );
  dff_sg \shifter_0/oi_2_reg[17]  ( .D(\shifter_0/n10169 ), .CP(clk), .Q(
        oi_2[17]) );
  dff_sg \shifter_0/oi_2_reg[18]  ( .D(\shifter_0/n10170 ), .CP(clk), .Q(
        oi_2[18]) );
  dff_sg \shifter_0/oi_2_reg[19]  ( .D(\shifter_0/n10171 ), .CP(clk), .Q(
        oi_2[19]) );
  dff_sg \shifter_0/oi_1_reg[0]  ( .D(\shifter_0/n10172 ), .CP(clk), .Q(
        oi_1[0]) );
  dff_sg \shifter_0/oi_1_reg[1]  ( .D(\shifter_0/n10173 ), .CP(clk), .Q(
        oi_1[1]) );
  dff_sg \shifter_0/oi_1_reg[2]  ( .D(\shifter_0/n10174 ), .CP(clk), .Q(
        oi_1[2]) );
  dff_sg \shifter_0/oi_1_reg[3]  ( .D(\shifter_0/n10175 ), .CP(clk), .Q(
        oi_1[3]) );
  dff_sg \shifter_0/oi_1_reg[4]  ( .D(\shifter_0/n10176 ), .CP(clk), .Q(
        oi_1[4]) );
  dff_sg \shifter_0/oi_1_reg[5]  ( .D(\shifter_0/n10177 ), .CP(clk), .Q(
        oi_1[5]) );
  dff_sg \shifter_0/oi_1_reg[6]  ( .D(\shifter_0/n10178 ), .CP(clk), .Q(
        oi_1[6]) );
  dff_sg \shifter_0/oi_1_reg[7]  ( .D(\shifter_0/n10179 ), .CP(clk), .Q(
        oi_1[7]) );
  dff_sg \shifter_0/oi_1_reg[8]  ( .D(\shifter_0/n10180 ), .CP(clk), .Q(
        oi_1[8]) );
  dff_sg \shifter_0/oi_1_reg[9]  ( .D(\shifter_0/n10181 ), .CP(clk), .Q(
        oi_1[9]) );
  dff_sg \shifter_0/oi_1_reg[10]  ( .D(\shifter_0/n10182 ), .CP(clk), .Q(
        oi_1[10]) );
  dff_sg \shifter_0/oi_1_reg[11]  ( .D(\shifter_0/n10183 ), .CP(clk), .Q(
        oi_1[11]) );
  dff_sg \shifter_0/oi_1_reg[12]  ( .D(\shifter_0/n10184 ), .CP(clk), .Q(
        oi_1[12]) );
  dff_sg \shifter_0/oi_1_reg[13]  ( .D(\shifter_0/n10185 ), .CP(clk), .Q(
        oi_1[13]) );
  dff_sg \shifter_0/oi_1_reg[14]  ( .D(\shifter_0/n10186 ), .CP(clk), .Q(
        oi_1[14]) );
  dff_sg \shifter_0/oi_1_reg[15]  ( .D(\shifter_0/n10187 ), .CP(clk), .Q(
        oi_1[15]) );
  dff_sg \shifter_0/oi_1_reg[16]  ( .D(\shifter_0/n10188 ), .CP(clk), .Q(
        oi_1[16]) );
  dff_sg \shifter_0/oi_1_reg[17]  ( .D(\shifter_0/n10189 ), .CP(clk), .Q(
        oi_1[17]) );
  dff_sg \shifter_0/oi_1_reg[18]  ( .D(\shifter_0/n10190 ), .CP(clk), .Q(
        oi_1[18]) );
  dff_sg \shifter_0/oi_1_reg[19]  ( .D(\shifter_0/n10191 ), .CP(clk), .Q(
        oi_1[19]) );
  dff_sg \shifter_0/oi_0_reg[0]  ( .D(\shifter_0/n10192 ), .CP(clk), .Q(
        oi_0[0]) );
  dff_sg \shifter_0/oi_0_reg[1]  ( .D(\shifter_0/n10193 ), .CP(clk), .Q(
        oi_0[1]) );
  dff_sg \shifter_0/oi_0_reg[2]  ( .D(\shifter_0/n10194 ), .CP(clk), .Q(
        oi_0[2]) );
  dff_sg \shifter_0/oi_0_reg[3]  ( .D(\shifter_0/n10195 ), .CP(clk), .Q(
        oi_0[3]) );
  dff_sg \shifter_0/oi_0_reg[4]  ( .D(\shifter_0/n10196 ), .CP(clk), .Q(
        oi_0[4]) );
  dff_sg \shifter_0/oi_0_reg[5]  ( .D(\shifter_0/n10197 ), .CP(clk), .Q(
        oi_0[5]) );
  dff_sg \shifter_0/oi_0_reg[6]  ( .D(\shifter_0/n10198 ), .CP(clk), .Q(
        oi_0[6]) );
  dff_sg \shifter_0/oi_0_reg[7]  ( .D(\shifter_0/n10199 ), .CP(clk), .Q(
        oi_0[7]) );
  dff_sg \shifter_0/oi_0_reg[8]  ( .D(\shifter_0/n10200 ), .CP(clk), .Q(
        oi_0[8]) );
  dff_sg \shifter_0/oi_0_reg[9]  ( .D(\shifter_0/n10201 ), .CP(clk), .Q(
        oi_0[9]) );
  dff_sg \shifter_0/oi_0_reg[10]  ( .D(\shifter_0/n10202 ), .CP(clk), .Q(
        oi_0[10]) );
  dff_sg \shifter_0/oi_0_reg[11]  ( .D(\shifter_0/n10203 ), .CP(clk), .Q(
        oi_0[11]) );
  dff_sg \shifter_0/oi_0_reg[12]  ( .D(\shifter_0/n10204 ), .CP(clk), .Q(
        oi_0[12]) );
  dff_sg \shifter_0/oi_0_reg[13]  ( .D(\shifter_0/n10205 ), .CP(clk), .Q(
        oi_0[13]) );
  dff_sg \shifter_0/oi_0_reg[14]  ( .D(\shifter_0/n10206 ), .CP(clk), .Q(
        oi_0[14]) );
  dff_sg \shifter_0/oi_0_reg[15]  ( .D(\shifter_0/n10207 ), .CP(clk), .Q(
        oi_0[15]) );
  dff_sg \shifter_0/oi_0_reg[16]  ( .D(\shifter_0/n10208 ), .CP(clk), .Q(
        oi_0[16]) );
  dff_sg \shifter_0/oi_0_reg[17]  ( .D(\shifter_0/n10209 ), .CP(clk), .Q(
        oi_0[17]) );
  dff_sg \shifter_0/oi_0_reg[18]  ( .D(\shifter_0/n10210 ), .CP(clk), .Q(
        oi_0[18]) );
  dff_sg \shifter_0/oi_0_reg[19]  ( .D(\shifter_0/n10211 ), .CP(clk), .Q(
        oi_0[19]) );
  dff_sg \shifter_0/ow_15_reg[0]  ( .D(\shifter_0/n10212 ), .CP(clk), .Q(
        ow_15[0]) );
  dff_sg \shifter_0/ow_15_reg[1]  ( .D(\shifter_0/n10213 ), .CP(clk), .Q(
        ow_15[1]) );
  dff_sg \shifter_0/ow_15_reg[2]  ( .D(\shifter_0/n10214 ), .CP(clk), .Q(
        ow_15[2]) );
  dff_sg \shifter_0/ow_15_reg[3]  ( .D(\shifter_0/n10215 ), .CP(clk), .Q(
        ow_15[3]) );
  dff_sg \shifter_0/ow_15_reg[4]  ( .D(\shifter_0/n10216 ), .CP(clk), .Q(
        ow_15[4]) );
  dff_sg \shifter_0/ow_15_reg[5]  ( .D(\shifter_0/n10217 ), .CP(clk), .Q(
        ow_15[5]) );
  dff_sg \shifter_0/ow_15_reg[6]  ( .D(\shifter_0/n10218 ), .CP(clk), .Q(
        ow_15[6]) );
  dff_sg \shifter_0/ow_15_reg[7]  ( .D(\shifter_0/n10219 ), .CP(clk), .Q(
        ow_15[7]) );
  dff_sg \shifter_0/ow_15_reg[8]  ( .D(\shifter_0/n10220 ), .CP(clk), .Q(
        ow_15[8]) );
  dff_sg \shifter_0/ow_15_reg[9]  ( .D(\shifter_0/n10221 ), .CP(clk), .Q(
        ow_15[9]) );
  dff_sg \shifter_0/ow_15_reg[10]  ( .D(\shifter_0/n10222 ), .CP(clk), .Q(
        ow_15[10]) );
  dff_sg \shifter_0/ow_15_reg[11]  ( .D(\shifter_0/n10223 ), .CP(clk), .Q(
        ow_15[11]) );
  dff_sg \shifter_0/ow_15_reg[12]  ( .D(\shifter_0/n10224 ), .CP(clk), .Q(
        ow_15[12]) );
  dff_sg \shifter_0/ow_15_reg[13]  ( .D(\shifter_0/n10225 ), .CP(clk), .Q(
        ow_15[13]) );
  dff_sg \shifter_0/ow_15_reg[14]  ( .D(\shifter_0/n10226 ), .CP(clk), .Q(
        ow_15[14]) );
  dff_sg \shifter_0/ow_15_reg[15]  ( .D(\shifter_0/n10227 ), .CP(clk), .Q(
        ow_15[15]) );
  dff_sg \shifter_0/ow_15_reg[16]  ( .D(\shifter_0/n10228 ), .CP(clk), .Q(
        ow_15[16]) );
  dff_sg \shifter_0/ow_15_reg[17]  ( .D(\shifter_0/n10229 ), .CP(clk), .Q(
        ow_15[17]) );
  dff_sg \shifter_0/ow_15_reg[18]  ( .D(\shifter_0/n10230 ), .CP(clk), .Q(
        ow_15[18]) );
  dff_sg \shifter_0/ow_15_reg[19]  ( .D(\shifter_0/n10231 ), .CP(clk), .Q(
        ow_15[19]) );
  dff_sg \shifter_0/i_pointer_reg[0]  ( .D(\shifter_0/n10232 ), .CP(clk), .Q(
        \shifter_0/i_pointer[0] ) );
  dff_sg \shifter_0/i_pointer_reg[1]  ( .D(\shifter_0/n10233 ), .CP(clk), .Q(
        \shifter_0/i_pointer[1] ) );
  dff_sg \shifter_0/i_pointer_reg[2]  ( .D(\shifter_0/n10234 ), .CP(clk), .Q(
        \shifter_0/i_pointer[2] ) );
  dff_sg \shifter_0/i_pointer_reg[3]  ( .D(\shifter_0/n10235 ), .CP(clk), .Q(
        \shifter_0/i_pointer[3] ) );
  dff_sg \shifter_0/pointer_reg[3]  ( .D(\shifter_0/n10885 ), .CP(clk), .Q(
        \shifter_0/pointer[3] ) );
  dff_sg \shifter_0/pointer_reg[2]  ( .D(\shifter_0/n10240 ), .CP(clk), .Q(
        \shifter_0/pointer[2] ) );
  dff_sg \shifter_0/pointer_reg[1]  ( .D(\shifter_0/n10241 ), .CP(clk), .Q(
        \shifter_0/pointer[1] ) );
  dff_sg \shifter_0/w_pointer_reg[0]  ( .D(\shifter_0/n10239 ), .CP(clk), .Q(
        \shifter_0/w_pointer[0] ) );
  dff_sg \shifter_0/w_pointer_reg[1]  ( .D(\shifter_0/n10238 ), .CP(clk), .Q(
        \shifter_0/w_pointer[1] ) );
  dff_sg \shifter_0/w_pointer_reg[2]  ( .D(\shifter_0/n10237 ), .CP(clk), .Q(
        \shifter_0/w_pointer[2] ) );
  dff_sg \shifter_0/w_pointer_reg[3]  ( .D(\shifter_0/n10236 ), .CP(clk), .Q(
        \shifter_0/w_pointer[3] ) );
  dff_sg \shifter_0/input_taken_reg  ( .D(\shifter_0/n10882 ), .CP(clk), .Q(
        filter_output_shifter_input_taken) );
  dff_sg \shifter_0/reg_i_0_reg[0]  ( .D(\shifter_0/n10881 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[0] ) );
  dff_sg \shifter_0/reg_i_0_reg[1]  ( .D(\shifter_0/n10880 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[1] ) );
  dff_sg \shifter_0/reg_i_0_reg[2]  ( .D(\shifter_0/n10879 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[2] ) );
  dff_sg \shifter_0/reg_i_0_reg[3]  ( .D(\shifter_0/n10878 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[3] ) );
  dff_sg \shifter_0/reg_i_0_reg[4]  ( .D(\shifter_0/n10877 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[4] ) );
  dff_sg \shifter_0/reg_i_0_reg[5]  ( .D(\shifter_0/n10876 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[5] ) );
  dff_sg \shifter_0/reg_i_0_reg[6]  ( .D(\shifter_0/n10875 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[6] ) );
  dff_sg \shifter_0/reg_i_0_reg[7]  ( .D(\shifter_0/n10874 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[7] ) );
  dff_sg \shifter_0/reg_i_0_reg[8]  ( .D(\shifter_0/n10873 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[8] ) );
  dff_sg \shifter_0/reg_i_0_reg[9]  ( .D(\shifter_0/n10872 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[9] ) );
  dff_sg \shifter_0/reg_i_0_reg[10]  ( .D(\shifter_0/n10871 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[10] ) );
  dff_sg \shifter_0/reg_i_0_reg[11]  ( .D(\shifter_0/n10870 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[11] ) );
  dff_sg \shifter_0/reg_i_0_reg[12]  ( .D(\shifter_0/n10869 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[12] ) );
  dff_sg \shifter_0/reg_i_0_reg[13]  ( .D(\shifter_0/n10868 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[13] ) );
  dff_sg \shifter_0/reg_i_0_reg[14]  ( .D(\shifter_0/n10867 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[14] ) );
  dff_sg \shifter_0/reg_i_0_reg[15]  ( .D(\shifter_0/n10866 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[15] ) );
  dff_sg \shifter_0/reg_i_0_reg[16]  ( .D(\shifter_0/n10865 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[16] ) );
  dff_sg \shifter_0/reg_i_0_reg[17]  ( .D(\shifter_0/n10864 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[17] ) );
  dff_sg \shifter_0/reg_i_0_reg[18]  ( .D(\shifter_0/n10863 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[18] ) );
  dff_sg \shifter_0/reg_i_0_reg[19]  ( .D(\shifter_0/n10862 ), .CP(clk), .Q(
        \shifter_0/reg_i_0[19] ) );
  dff_sg \shifter_0/reg_i_1_reg[0]  ( .D(\shifter_0/n10861 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[0] ) );
  dff_sg \shifter_0/reg_i_1_reg[1]  ( .D(\shifter_0/n10860 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[1] ) );
  dff_sg \shifter_0/reg_i_1_reg[2]  ( .D(\shifter_0/n10859 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[2] ) );
  dff_sg \shifter_0/reg_i_1_reg[3]  ( .D(\shifter_0/n10858 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[3] ) );
  dff_sg \shifter_0/reg_i_1_reg[4]  ( .D(\shifter_0/n10857 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[4] ) );
  dff_sg \shifter_0/reg_i_1_reg[5]  ( .D(\shifter_0/n10856 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[5] ) );
  dff_sg \shifter_0/reg_i_1_reg[6]  ( .D(\shifter_0/n10855 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[6] ) );
  dff_sg \shifter_0/reg_i_1_reg[7]  ( .D(\shifter_0/n10854 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[7] ) );
  dff_sg \shifter_0/reg_i_1_reg[8]  ( .D(\shifter_0/n10853 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[8] ) );
  dff_sg \shifter_0/reg_i_1_reg[9]  ( .D(\shifter_0/n10852 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[9] ) );
  dff_sg \shifter_0/reg_i_1_reg[10]  ( .D(\shifter_0/n10851 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[10] ) );
  dff_sg \shifter_0/reg_i_1_reg[11]  ( .D(\shifter_0/n10850 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[11] ) );
  dff_sg \shifter_0/reg_i_1_reg[12]  ( .D(\shifter_0/n10849 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[12] ) );
  dff_sg \shifter_0/reg_i_1_reg[13]  ( .D(\shifter_0/n10848 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[13] ) );
  dff_sg \shifter_0/reg_i_1_reg[14]  ( .D(\shifter_0/n10847 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[14] ) );
  dff_sg \shifter_0/reg_i_1_reg[15]  ( .D(\shifter_0/n10846 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[15] ) );
  dff_sg \shifter_0/reg_i_1_reg[16]  ( .D(\shifter_0/n10845 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[16] ) );
  dff_sg \shifter_0/reg_i_1_reg[17]  ( .D(\shifter_0/n10844 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[17] ) );
  dff_sg \shifter_0/reg_i_1_reg[18]  ( .D(\shifter_0/n10843 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[18] ) );
  dff_sg \shifter_0/reg_i_1_reg[19]  ( .D(\shifter_0/n10842 ), .CP(clk), .Q(
        \shifter_0/reg_i_1[19] ) );
  dff_sg \shifter_0/reg_i_2_reg[0]  ( .D(\shifter_0/n10841 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[0] ) );
  dff_sg \shifter_0/reg_i_2_reg[1]  ( .D(\shifter_0/n10840 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[1] ) );
  dff_sg \shifter_0/reg_i_2_reg[2]  ( .D(\shifter_0/n10839 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[2] ) );
  dff_sg \shifter_0/reg_i_2_reg[3]  ( .D(\shifter_0/n10838 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[3] ) );
  dff_sg \shifter_0/reg_i_2_reg[4]  ( .D(\shifter_0/n10837 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[4] ) );
  dff_sg \shifter_0/reg_i_2_reg[5]  ( .D(\shifter_0/n10836 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[5] ) );
  dff_sg \shifter_0/reg_i_2_reg[6]  ( .D(\shifter_0/n10835 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[6] ) );
  dff_sg \shifter_0/reg_i_2_reg[7]  ( .D(\shifter_0/n10834 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[7] ) );
  dff_sg \shifter_0/reg_i_2_reg[8]  ( .D(\shifter_0/n10833 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[8] ) );
  dff_sg \shifter_0/reg_i_2_reg[9]  ( .D(\shifter_0/n10832 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[9] ) );
  dff_sg \shifter_0/reg_i_2_reg[10]  ( .D(\shifter_0/n10831 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[10] ) );
  dff_sg \shifter_0/reg_i_2_reg[11]  ( .D(\shifter_0/n10830 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[11] ) );
  dff_sg \shifter_0/reg_i_2_reg[12]  ( .D(\shifter_0/n10829 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[12] ) );
  dff_sg \shifter_0/reg_i_2_reg[13]  ( .D(\shifter_0/n10828 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[13] ) );
  dff_sg \shifter_0/reg_i_2_reg[14]  ( .D(\shifter_0/n10827 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[14] ) );
  dff_sg \shifter_0/reg_i_2_reg[15]  ( .D(\shifter_0/n10826 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[15] ) );
  dff_sg \shifter_0/reg_i_2_reg[16]  ( .D(\shifter_0/n10825 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[16] ) );
  dff_sg \shifter_0/reg_i_2_reg[17]  ( .D(\shifter_0/n10824 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[17] ) );
  dff_sg \shifter_0/reg_i_2_reg[18]  ( .D(\shifter_0/n10823 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[18] ) );
  dff_sg \shifter_0/reg_i_2_reg[19]  ( .D(\shifter_0/n10822 ), .CP(clk), .Q(
        \shifter_0/reg_i_2[19] ) );
  dff_sg \shifter_0/reg_i_3_reg[0]  ( .D(\shifter_0/n10821 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[0] ) );
  dff_sg \shifter_0/reg_i_3_reg[1]  ( .D(\shifter_0/n10820 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[1] ) );
  dff_sg \shifter_0/reg_i_3_reg[2]  ( .D(\shifter_0/n10819 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[2] ) );
  dff_sg \shifter_0/reg_i_3_reg[3]  ( .D(\shifter_0/n10818 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[3] ) );
  dff_sg \shifter_0/reg_i_3_reg[4]  ( .D(\shifter_0/n10817 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[4] ) );
  dff_sg \shifter_0/reg_i_3_reg[5]  ( .D(\shifter_0/n10816 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[5] ) );
  dff_sg \shifter_0/reg_i_3_reg[6]  ( .D(\shifter_0/n10815 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[6] ) );
  dff_sg \shifter_0/reg_i_3_reg[7]  ( .D(\shifter_0/n10814 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[7] ) );
  dff_sg \shifter_0/reg_i_3_reg[8]  ( .D(\shifter_0/n10813 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[8] ) );
  dff_sg \shifter_0/reg_i_3_reg[9]  ( .D(\shifter_0/n10812 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[9] ) );
  dff_sg \shifter_0/reg_i_3_reg[10]  ( .D(\shifter_0/n10811 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[10] ) );
  dff_sg \shifter_0/reg_i_3_reg[11]  ( .D(\shifter_0/n10810 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[11] ) );
  dff_sg \shifter_0/reg_i_3_reg[12]  ( .D(\shifter_0/n10809 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[12] ) );
  dff_sg \shifter_0/reg_i_3_reg[13]  ( .D(\shifter_0/n10808 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[13] ) );
  dff_sg \shifter_0/reg_i_3_reg[14]  ( .D(\shifter_0/n10807 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[14] ) );
  dff_sg \shifter_0/reg_i_3_reg[15]  ( .D(\shifter_0/n10806 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[15] ) );
  dff_sg \shifter_0/reg_i_3_reg[16]  ( .D(\shifter_0/n10805 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[16] ) );
  dff_sg \shifter_0/reg_i_3_reg[17]  ( .D(\shifter_0/n10804 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[17] ) );
  dff_sg \shifter_0/reg_i_3_reg[18]  ( .D(\shifter_0/n10803 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[18] ) );
  dff_sg \shifter_0/reg_i_3_reg[19]  ( .D(\shifter_0/n10802 ), .CP(clk), .Q(
        \shifter_0/reg_i_3[19] ) );
  dff_sg \shifter_0/reg_i_4_reg[0]  ( .D(\shifter_0/n10801 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[0] ) );
  dff_sg \shifter_0/reg_i_4_reg[1]  ( .D(\shifter_0/n10800 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[1] ) );
  dff_sg \shifter_0/reg_i_4_reg[2]  ( .D(\shifter_0/n10799 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[2] ) );
  dff_sg \shifter_0/reg_i_4_reg[3]  ( .D(\shifter_0/n10798 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[3] ) );
  dff_sg \shifter_0/reg_i_4_reg[4]  ( .D(\shifter_0/n10797 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[4] ) );
  dff_sg \shifter_0/reg_i_4_reg[5]  ( .D(\shifter_0/n10796 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[5] ) );
  dff_sg \shifter_0/reg_i_4_reg[6]  ( .D(\shifter_0/n10795 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[6] ) );
  dff_sg \shifter_0/reg_i_4_reg[7]  ( .D(\shifter_0/n10794 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[7] ) );
  dff_sg \shifter_0/reg_i_4_reg[8]  ( .D(\shifter_0/n10793 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[8] ) );
  dff_sg \shifter_0/reg_i_4_reg[9]  ( .D(\shifter_0/n10792 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[9] ) );
  dff_sg \shifter_0/reg_i_4_reg[10]  ( .D(\shifter_0/n10791 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[10] ) );
  dff_sg \shifter_0/reg_i_4_reg[11]  ( .D(\shifter_0/n10790 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[11] ) );
  dff_sg \shifter_0/reg_i_4_reg[12]  ( .D(\shifter_0/n10789 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[12] ) );
  dff_sg \shifter_0/reg_i_4_reg[13]  ( .D(\shifter_0/n10788 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[13] ) );
  dff_sg \shifter_0/reg_i_4_reg[14]  ( .D(\shifter_0/n10787 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[14] ) );
  dff_sg \shifter_0/reg_i_4_reg[15]  ( .D(\shifter_0/n10786 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[15] ) );
  dff_sg \shifter_0/reg_i_4_reg[16]  ( .D(\shifter_0/n10785 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[16] ) );
  dff_sg \shifter_0/reg_i_4_reg[17]  ( .D(\shifter_0/n10784 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[17] ) );
  dff_sg \shifter_0/reg_i_4_reg[18]  ( .D(\shifter_0/n10783 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[18] ) );
  dff_sg \shifter_0/reg_i_4_reg[19]  ( .D(\shifter_0/n10782 ), .CP(clk), .Q(
        \shifter_0/reg_i_4[19] ) );
  dff_sg \shifter_0/reg_i_5_reg[0]  ( .D(\shifter_0/n10781 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[0] ) );
  dff_sg \shifter_0/reg_i_5_reg[1]  ( .D(\shifter_0/n10780 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[1] ) );
  dff_sg \shifter_0/reg_i_5_reg[2]  ( .D(\shifter_0/n10779 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[2] ) );
  dff_sg \shifter_0/reg_i_5_reg[3]  ( .D(\shifter_0/n10778 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[3] ) );
  dff_sg \shifter_0/reg_i_5_reg[4]  ( .D(\shifter_0/n10777 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[4] ) );
  dff_sg \shifter_0/reg_i_5_reg[5]  ( .D(\shifter_0/n10776 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[5] ) );
  dff_sg \shifter_0/reg_i_5_reg[6]  ( .D(\shifter_0/n10775 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[6] ) );
  dff_sg \shifter_0/reg_i_5_reg[7]  ( .D(\shifter_0/n10774 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[7] ) );
  dff_sg \shifter_0/reg_i_5_reg[8]  ( .D(\shifter_0/n10773 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[8] ) );
  dff_sg \shifter_0/reg_i_5_reg[9]  ( .D(\shifter_0/n10772 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[9] ) );
  dff_sg \shifter_0/reg_i_5_reg[10]  ( .D(\shifter_0/n10771 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[10] ) );
  dff_sg \shifter_0/reg_i_5_reg[11]  ( .D(\shifter_0/n10770 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[11] ) );
  dff_sg \shifter_0/reg_i_5_reg[12]  ( .D(\shifter_0/n10769 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[12] ) );
  dff_sg \shifter_0/reg_i_5_reg[13]  ( .D(\shifter_0/n10768 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[13] ) );
  dff_sg \shifter_0/reg_i_5_reg[14]  ( .D(\shifter_0/n10767 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[14] ) );
  dff_sg \shifter_0/reg_i_5_reg[15]  ( .D(\shifter_0/n10766 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[15] ) );
  dff_sg \shifter_0/reg_i_5_reg[16]  ( .D(\shifter_0/n10765 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[16] ) );
  dff_sg \shifter_0/reg_i_5_reg[17]  ( .D(\shifter_0/n10764 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[17] ) );
  dff_sg \shifter_0/reg_i_5_reg[18]  ( .D(\shifter_0/n10763 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[18] ) );
  dff_sg \shifter_0/reg_i_5_reg[19]  ( .D(\shifter_0/n10762 ), .CP(clk), .Q(
        \shifter_0/reg_i_5[19] ) );
  dff_sg \shifter_0/reg_i_6_reg[0]  ( .D(\shifter_0/n10761 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[0] ) );
  dff_sg \shifter_0/reg_i_6_reg[1]  ( .D(\shifter_0/n10760 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[1] ) );
  dff_sg \shifter_0/reg_i_6_reg[2]  ( .D(\shifter_0/n10759 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[2] ) );
  dff_sg \shifter_0/reg_i_6_reg[3]  ( .D(\shifter_0/n10758 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[3] ) );
  dff_sg \shifter_0/reg_i_6_reg[4]  ( .D(\shifter_0/n10757 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[4] ) );
  dff_sg \shifter_0/reg_i_6_reg[5]  ( .D(\shifter_0/n10756 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[5] ) );
  dff_sg \shifter_0/reg_i_6_reg[6]  ( .D(\shifter_0/n10755 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[6] ) );
  dff_sg \shifter_0/reg_i_6_reg[7]  ( .D(\shifter_0/n10754 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[7] ) );
  dff_sg \shifter_0/reg_i_6_reg[8]  ( .D(\shifter_0/n10753 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[8] ) );
  dff_sg \shifter_0/reg_i_6_reg[9]  ( .D(\shifter_0/n10752 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[9] ) );
  dff_sg \shifter_0/reg_i_6_reg[10]  ( .D(\shifter_0/n10751 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[10] ) );
  dff_sg \shifter_0/reg_i_6_reg[11]  ( .D(\shifter_0/n10750 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[11] ) );
  dff_sg \shifter_0/reg_i_6_reg[12]  ( .D(\shifter_0/n10749 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[12] ) );
  dff_sg \shifter_0/reg_i_6_reg[13]  ( .D(\shifter_0/n10748 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[13] ) );
  dff_sg \shifter_0/reg_i_6_reg[14]  ( .D(\shifter_0/n10747 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[14] ) );
  dff_sg \shifter_0/reg_i_6_reg[15]  ( .D(\shifter_0/n10746 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[15] ) );
  dff_sg \shifter_0/reg_i_6_reg[16]  ( .D(\shifter_0/n10745 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[16] ) );
  dff_sg \shifter_0/reg_i_6_reg[17]  ( .D(\shifter_0/n10744 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[17] ) );
  dff_sg \shifter_0/reg_i_6_reg[18]  ( .D(\shifter_0/n10743 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[18] ) );
  dff_sg \shifter_0/reg_i_6_reg[19]  ( .D(\shifter_0/n10742 ), .CP(clk), .Q(
        \shifter_0/reg_i_6[19] ) );
  dff_sg \shifter_0/reg_i_7_reg[0]  ( .D(\shifter_0/n10741 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[0] ) );
  dff_sg \shifter_0/reg_i_7_reg[1]  ( .D(\shifter_0/n10740 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[1] ) );
  dff_sg \shifter_0/reg_i_7_reg[2]  ( .D(\shifter_0/n10739 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[2] ) );
  dff_sg \shifter_0/reg_i_7_reg[3]  ( .D(\shifter_0/n10738 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[3] ) );
  dff_sg \shifter_0/reg_i_7_reg[4]  ( .D(\shifter_0/n10737 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[4] ) );
  dff_sg \shifter_0/reg_i_7_reg[5]  ( .D(\shifter_0/n10736 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[5] ) );
  dff_sg \shifter_0/reg_i_7_reg[6]  ( .D(\shifter_0/n10735 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[6] ) );
  dff_sg \shifter_0/reg_i_7_reg[7]  ( .D(\shifter_0/n10734 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[7] ) );
  dff_sg \shifter_0/reg_i_7_reg[8]  ( .D(\shifter_0/n10733 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[8] ) );
  dff_sg \shifter_0/reg_i_7_reg[9]  ( .D(\shifter_0/n10732 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[9] ) );
  dff_sg \shifter_0/reg_i_7_reg[10]  ( .D(\shifter_0/n10731 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[10] ) );
  dff_sg \shifter_0/reg_i_7_reg[11]  ( .D(\shifter_0/n10730 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[11] ) );
  dff_sg \shifter_0/reg_i_7_reg[12]  ( .D(\shifter_0/n10729 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[12] ) );
  dff_sg \shifter_0/reg_i_7_reg[13]  ( .D(\shifter_0/n10728 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[13] ) );
  dff_sg \shifter_0/reg_i_7_reg[14]  ( .D(\shifter_0/n10727 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[14] ) );
  dff_sg \shifter_0/reg_i_7_reg[15]  ( .D(\shifter_0/n10726 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[15] ) );
  dff_sg \shifter_0/reg_i_7_reg[16]  ( .D(\shifter_0/n10725 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[16] ) );
  dff_sg \shifter_0/reg_i_7_reg[17]  ( .D(\shifter_0/n10724 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[17] ) );
  dff_sg \shifter_0/reg_i_7_reg[18]  ( .D(\shifter_0/n10723 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[18] ) );
  dff_sg \shifter_0/reg_i_7_reg[19]  ( .D(\shifter_0/n10722 ), .CP(clk), .Q(
        \shifter_0/reg_i_7[19] ) );
  dff_sg \shifter_0/reg_i_8_reg[0]  ( .D(\shifter_0/n10721 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[0] ) );
  dff_sg \shifter_0/reg_i_8_reg[1]  ( .D(\shifter_0/n10720 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[1] ) );
  dff_sg \shifter_0/reg_i_8_reg[2]  ( .D(\shifter_0/n10719 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[2] ) );
  dff_sg \shifter_0/reg_i_8_reg[3]  ( .D(\shifter_0/n10718 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[3] ) );
  dff_sg \shifter_0/reg_i_8_reg[4]  ( .D(\shifter_0/n10717 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[4] ) );
  dff_sg \shifter_0/reg_i_8_reg[5]  ( .D(\shifter_0/n10716 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[5] ) );
  dff_sg \shifter_0/reg_i_8_reg[6]  ( .D(\shifter_0/n10715 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[6] ) );
  dff_sg \shifter_0/reg_i_8_reg[7]  ( .D(\shifter_0/n10714 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[7] ) );
  dff_sg \shifter_0/reg_i_8_reg[8]  ( .D(\shifter_0/n10713 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[8] ) );
  dff_sg \shifter_0/reg_i_8_reg[9]  ( .D(\shifter_0/n10712 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[9] ) );
  dff_sg \shifter_0/reg_i_8_reg[10]  ( .D(\shifter_0/n10711 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[10] ) );
  dff_sg \shifter_0/reg_i_8_reg[11]  ( .D(\shifter_0/n10710 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[11] ) );
  dff_sg \shifter_0/reg_i_8_reg[12]  ( .D(\shifter_0/n10709 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[12] ) );
  dff_sg \shifter_0/reg_i_8_reg[13]  ( .D(\shifter_0/n10708 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[13] ) );
  dff_sg \shifter_0/reg_i_8_reg[14]  ( .D(\shifter_0/n10707 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[14] ) );
  dff_sg \shifter_0/reg_i_8_reg[15]  ( .D(\shifter_0/n10706 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[15] ) );
  dff_sg \shifter_0/reg_i_8_reg[16]  ( .D(\shifter_0/n10705 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[16] ) );
  dff_sg \shifter_0/reg_i_8_reg[17]  ( .D(\shifter_0/n10704 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[17] ) );
  dff_sg \shifter_0/reg_i_8_reg[18]  ( .D(\shifter_0/n10703 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[18] ) );
  dff_sg \shifter_0/reg_i_8_reg[19]  ( .D(\shifter_0/n10702 ), .CP(clk), .Q(
        \shifter_0/reg_i_8[19] ) );
  dff_sg \shifter_0/reg_i_9_reg[0]  ( .D(\shifter_0/n10701 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[0] ) );
  dff_sg \shifter_0/reg_i_9_reg[1]  ( .D(\shifter_0/n10700 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[1] ) );
  dff_sg \shifter_0/reg_i_9_reg[2]  ( .D(\shifter_0/n10699 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[2] ) );
  dff_sg \shifter_0/reg_i_9_reg[3]  ( .D(\shifter_0/n10698 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[3] ) );
  dff_sg \shifter_0/reg_i_9_reg[4]  ( .D(\shifter_0/n10697 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[4] ) );
  dff_sg \shifter_0/reg_i_9_reg[5]  ( .D(\shifter_0/n10696 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[5] ) );
  dff_sg \shifter_0/reg_i_9_reg[6]  ( .D(\shifter_0/n10695 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[6] ) );
  dff_sg \shifter_0/reg_i_9_reg[7]  ( .D(\shifter_0/n10694 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[7] ) );
  dff_sg \shifter_0/reg_i_9_reg[8]  ( .D(\shifter_0/n10693 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[8] ) );
  dff_sg \shifter_0/reg_i_9_reg[9]  ( .D(\shifter_0/n10692 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[9] ) );
  dff_sg \shifter_0/reg_i_9_reg[10]  ( .D(\shifter_0/n10691 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[10] ) );
  dff_sg \shifter_0/reg_i_9_reg[11]  ( .D(\shifter_0/n10690 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[11] ) );
  dff_sg \shifter_0/reg_i_9_reg[12]  ( .D(\shifter_0/n10689 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[12] ) );
  dff_sg \shifter_0/reg_i_9_reg[13]  ( .D(\shifter_0/n10688 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[13] ) );
  dff_sg \shifter_0/reg_i_9_reg[14]  ( .D(\shifter_0/n10687 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[14] ) );
  dff_sg \shifter_0/reg_i_9_reg[15]  ( .D(\shifter_0/n10686 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[15] ) );
  dff_sg \shifter_0/reg_i_9_reg[16]  ( .D(\shifter_0/n10685 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[16] ) );
  dff_sg \shifter_0/reg_i_9_reg[17]  ( .D(\shifter_0/n10684 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[17] ) );
  dff_sg \shifter_0/reg_i_9_reg[18]  ( .D(\shifter_0/n10683 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[18] ) );
  dff_sg \shifter_0/reg_i_9_reg[19]  ( .D(\shifter_0/n10682 ), .CP(clk), .Q(
        \shifter_0/reg_i_9[19] ) );
  dff_sg \shifter_0/reg_i_10_reg[0]  ( .D(\shifter_0/n10681 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[0] ) );
  dff_sg \shifter_0/reg_i_10_reg[1]  ( .D(\shifter_0/n10680 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[1] ) );
  dff_sg \shifter_0/reg_i_10_reg[2]  ( .D(\shifter_0/n10679 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[2] ) );
  dff_sg \shifter_0/reg_i_10_reg[3]  ( .D(\shifter_0/n10678 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[3] ) );
  dff_sg \shifter_0/reg_i_10_reg[4]  ( .D(\shifter_0/n10677 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[4] ) );
  dff_sg \shifter_0/reg_i_10_reg[5]  ( .D(\shifter_0/n10676 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[5] ) );
  dff_sg \shifter_0/reg_i_10_reg[6]  ( .D(\shifter_0/n10675 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[6] ) );
  dff_sg \shifter_0/reg_i_10_reg[7]  ( .D(\shifter_0/n10674 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[7] ) );
  dff_sg \shifter_0/reg_i_10_reg[8]  ( .D(\shifter_0/n10673 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[8] ) );
  dff_sg \shifter_0/reg_i_10_reg[9]  ( .D(\shifter_0/n10672 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[9] ) );
  dff_sg \shifter_0/reg_i_10_reg[10]  ( .D(\shifter_0/n10671 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[10] ) );
  dff_sg \shifter_0/reg_i_10_reg[11]  ( .D(\shifter_0/n10670 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[11] ) );
  dff_sg \shifter_0/reg_i_10_reg[12]  ( .D(\shifter_0/n10669 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[12] ) );
  dff_sg \shifter_0/reg_i_10_reg[13]  ( .D(\shifter_0/n10668 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[13] ) );
  dff_sg \shifter_0/reg_i_10_reg[14]  ( .D(\shifter_0/n10667 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[14] ) );
  dff_sg \shifter_0/reg_i_10_reg[15]  ( .D(\shifter_0/n10666 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[15] ) );
  dff_sg \shifter_0/reg_i_10_reg[16]  ( .D(\shifter_0/n10665 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[16] ) );
  dff_sg \shifter_0/reg_i_10_reg[17]  ( .D(\shifter_0/n10664 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[17] ) );
  dff_sg \shifter_0/reg_i_10_reg[18]  ( .D(\shifter_0/n10663 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[18] ) );
  dff_sg \shifter_0/reg_i_10_reg[19]  ( .D(\shifter_0/n10662 ), .CP(clk), .Q(
        \shifter_0/reg_i_10[19] ) );
  dff_sg \shifter_0/reg_i_11_reg[0]  ( .D(\shifter_0/n10661 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[0] ) );
  dff_sg \shifter_0/reg_i_11_reg[1]  ( .D(\shifter_0/n10660 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[1] ) );
  dff_sg \shifter_0/reg_i_11_reg[2]  ( .D(\shifter_0/n10659 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[2] ) );
  dff_sg \shifter_0/reg_i_11_reg[3]  ( .D(\shifter_0/n10658 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[3] ) );
  dff_sg \shifter_0/reg_i_11_reg[4]  ( .D(\shifter_0/n10657 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[4] ) );
  dff_sg \shifter_0/reg_i_11_reg[5]  ( .D(\shifter_0/n10656 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[5] ) );
  dff_sg \shifter_0/reg_i_11_reg[6]  ( .D(\shifter_0/n10655 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[6] ) );
  dff_sg \shifter_0/reg_i_11_reg[7]  ( .D(\shifter_0/n10654 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[7] ) );
  dff_sg \shifter_0/reg_i_11_reg[8]  ( .D(\shifter_0/n10653 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[8] ) );
  dff_sg \shifter_0/reg_i_11_reg[9]  ( .D(\shifter_0/n10652 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[9] ) );
  dff_sg \shifter_0/reg_i_11_reg[10]  ( .D(\shifter_0/n10651 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[10] ) );
  dff_sg \shifter_0/reg_i_11_reg[11]  ( .D(\shifter_0/n10650 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[11] ) );
  dff_sg \shifter_0/reg_i_11_reg[12]  ( .D(\shifter_0/n10649 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[12] ) );
  dff_sg \shifter_0/reg_i_11_reg[13]  ( .D(\shifter_0/n10648 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[13] ) );
  dff_sg \shifter_0/reg_i_11_reg[14]  ( .D(\shifter_0/n10647 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[14] ) );
  dff_sg \shifter_0/reg_i_11_reg[15]  ( .D(\shifter_0/n10646 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[15] ) );
  dff_sg \shifter_0/reg_i_11_reg[16]  ( .D(\shifter_0/n10645 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[16] ) );
  dff_sg \shifter_0/reg_i_11_reg[17]  ( .D(\shifter_0/n10644 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[17] ) );
  dff_sg \shifter_0/reg_i_11_reg[18]  ( .D(\shifter_0/n10643 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[18] ) );
  dff_sg \shifter_0/reg_i_11_reg[19]  ( .D(\shifter_0/n10642 ), .CP(clk), .Q(
        \shifter_0/reg_i_11[19] ) );
  dff_sg \shifter_0/reg_i_12_reg[0]  ( .D(\shifter_0/n10641 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[0] ) );
  dff_sg \shifter_0/reg_i_12_reg[1]  ( .D(\shifter_0/n10640 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[1] ) );
  dff_sg \shifter_0/reg_i_12_reg[2]  ( .D(\shifter_0/n10639 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[2] ) );
  dff_sg \shifter_0/reg_i_12_reg[3]  ( .D(\shifter_0/n10638 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[3] ) );
  dff_sg \shifter_0/reg_i_12_reg[4]  ( .D(\shifter_0/n10637 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[4] ) );
  dff_sg \shifter_0/reg_i_12_reg[5]  ( .D(\shifter_0/n10636 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[5] ) );
  dff_sg \shifter_0/reg_i_12_reg[6]  ( .D(\shifter_0/n10635 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[6] ) );
  dff_sg \shifter_0/reg_i_12_reg[7]  ( .D(\shifter_0/n10634 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[7] ) );
  dff_sg \shifter_0/reg_i_12_reg[8]  ( .D(\shifter_0/n10633 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[8] ) );
  dff_sg \shifter_0/reg_i_12_reg[9]  ( .D(\shifter_0/n10632 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[9] ) );
  dff_sg \shifter_0/reg_i_12_reg[10]  ( .D(\shifter_0/n10631 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[10] ) );
  dff_sg \shifter_0/reg_i_12_reg[11]  ( .D(\shifter_0/n10630 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[11] ) );
  dff_sg \shifter_0/reg_i_12_reg[12]  ( .D(\shifter_0/n10629 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[12] ) );
  dff_sg \shifter_0/reg_i_12_reg[13]  ( .D(\shifter_0/n10628 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[13] ) );
  dff_sg \shifter_0/reg_i_12_reg[14]  ( .D(\shifter_0/n10627 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[14] ) );
  dff_sg \shifter_0/reg_i_12_reg[15]  ( .D(\shifter_0/n10626 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[15] ) );
  dff_sg \shifter_0/reg_i_12_reg[16]  ( .D(\shifter_0/n10625 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[16] ) );
  dff_sg \shifter_0/reg_i_12_reg[17]  ( .D(\shifter_0/n10624 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[17] ) );
  dff_sg \shifter_0/reg_i_12_reg[18]  ( .D(\shifter_0/n10623 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[18] ) );
  dff_sg \shifter_0/reg_i_12_reg[19]  ( .D(\shifter_0/n10622 ), .CP(clk), .Q(
        \shifter_0/reg_i_12[19] ) );
  dff_sg \shifter_0/reg_i_13_reg[0]  ( .D(\shifter_0/n10621 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[0] ) );
  dff_sg \shifter_0/reg_i_13_reg[1]  ( .D(\shifter_0/n10620 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[1] ) );
  dff_sg \shifter_0/reg_i_13_reg[2]  ( .D(\shifter_0/n10619 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[2] ) );
  dff_sg \shifter_0/reg_i_13_reg[3]  ( .D(\shifter_0/n10618 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[3] ) );
  dff_sg \shifter_0/reg_i_13_reg[4]  ( .D(\shifter_0/n10617 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[4] ) );
  dff_sg \shifter_0/reg_i_13_reg[5]  ( .D(\shifter_0/n10616 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[5] ) );
  dff_sg \shifter_0/reg_i_13_reg[6]  ( .D(\shifter_0/n10615 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[6] ) );
  dff_sg \shifter_0/reg_i_13_reg[7]  ( .D(\shifter_0/n10614 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[7] ) );
  dff_sg \shifter_0/reg_i_13_reg[8]  ( .D(\shifter_0/n10613 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[8] ) );
  dff_sg \shifter_0/reg_i_13_reg[9]  ( .D(\shifter_0/n10612 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[9] ) );
  dff_sg \shifter_0/reg_i_13_reg[10]  ( .D(\shifter_0/n10611 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[10] ) );
  dff_sg \shifter_0/reg_i_13_reg[11]  ( .D(\shifter_0/n10610 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[11] ) );
  dff_sg \shifter_0/reg_i_13_reg[12]  ( .D(\shifter_0/n10609 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[12] ) );
  dff_sg \shifter_0/reg_i_13_reg[13]  ( .D(\shifter_0/n10608 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[13] ) );
  dff_sg \shifter_0/reg_i_13_reg[14]  ( .D(\shifter_0/n10607 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[14] ) );
  dff_sg \shifter_0/reg_i_13_reg[15]  ( .D(\shifter_0/n10606 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[15] ) );
  dff_sg \shifter_0/reg_i_13_reg[16]  ( .D(\shifter_0/n10605 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[16] ) );
  dff_sg \shifter_0/reg_i_13_reg[17]  ( .D(\shifter_0/n10604 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[17] ) );
  dff_sg \shifter_0/reg_i_13_reg[18]  ( .D(\shifter_0/n10603 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[18] ) );
  dff_sg \shifter_0/reg_i_13_reg[19]  ( .D(\shifter_0/n10602 ), .CP(clk), .Q(
        \shifter_0/reg_i_13[19] ) );
  dff_sg \shifter_0/reg_i_14_reg[0]  ( .D(\shifter_0/n10601 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[0] ) );
  dff_sg \shifter_0/reg_i_14_reg[1]  ( .D(\shifter_0/n10600 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[1] ) );
  dff_sg \shifter_0/reg_i_14_reg[2]  ( .D(\shifter_0/n10599 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[2] ) );
  dff_sg \shifter_0/reg_i_14_reg[3]  ( .D(\shifter_0/n10598 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[3] ) );
  dff_sg \shifter_0/reg_i_14_reg[4]  ( .D(\shifter_0/n10597 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[4] ) );
  dff_sg \shifter_0/reg_i_14_reg[5]  ( .D(\shifter_0/n10596 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[5] ) );
  dff_sg \shifter_0/reg_i_14_reg[6]  ( .D(\shifter_0/n10595 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[6] ) );
  dff_sg \shifter_0/reg_i_14_reg[7]  ( .D(\shifter_0/n10594 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[7] ) );
  dff_sg \shifter_0/reg_i_14_reg[8]  ( .D(\shifter_0/n10593 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[8] ) );
  dff_sg \shifter_0/reg_i_14_reg[9]  ( .D(\shifter_0/n10592 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[9] ) );
  dff_sg \shifter_0/reg_i_14_reg[10]  ( .D(\shifter_0/n10591 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[10] ) );
  dff_sg \shifter_0/reg_i_14_reg[11]  ( .D(\shifter_0/n10590 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[11] ) );
  dff_sg \shifter_0/reg_i_14_reg[12]  ( .D(\shifter_0/n10589 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[12] ) );
  dff_sg \shifter_0/reg_i_14_reg[13]  ( .D(\shifter_0/n10588 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[13] ) );
  dff_sg \shifter_0/reg_i_14_reg[14]  ( .D(\shifter_0/n10587 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[14] ) );
  dff_sg \shifter_0/reg_i_14_reg[15]  ( .D(\shifter_0/n10586 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[15] ) );
  dff_sg \shifter_0/reg_i_14_reg[16]  ( .D(\shifter_0/n10585 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[16] ) );
  dff_sg \shifter_0/reg_i_14_reg[17]  ( .D(\shifter_0/n10584 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[17] ) );
  dff_sg \shifter_0/reg_i_14_reg[18]  ( .D(\shifter_0/n10583 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[18] ) );
  dff_sg \shifter_0/reg_i_14_reg[19]  ( .D(\shifter_0/n10582 ), .CP(clk), .Q(
        \shifter_0/reg_i_14[19] ) );
  dff_sg \shifter_0/reg_i_15_reg[0]  ( .D(\shifter_0/n10581 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[0] ) );
  dff_sg \shifter_0/reg_i_15_reg[1]  ( .D(\shifter_0/n10580 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[1] ) );
  dff_sg \shifter_0/reg_i_15_reg[2]  ( .D(\shifter_0/n10579 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[2] ) );
  dff_sg \shifter_0/reg_i_15_reg[3]  ( .D(\shifter_0/n10578 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[3] ) );
  dff_sg \shifter_0/reg_i_15_reg[4]  ( .D(\shifter_0/n10577 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[4] ) );
  dff_sg \shifter_0/reg_i_15_reg[5]  ( .D(\shifter_0/n10576 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[5] ) );
  dff_sg \shifter_0/reg_i_15_reg[6]  ( .D(\shifter_0/n10575 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[6] ) );
  dff_sg \shifter_0/reg_i_15_reg[7]  ( .D(\shifter_0/n10574 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[7] ) );
  dff_sg \shifter_0/reg_i_15_reg[8]  ( .D(\shifter_0/n10573 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[8] ) );
  dff_sg \shifter_0/reg_i_15_reg[9]  ( .D(\shifter_0/n10572 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[9] ) );
  dff_sg \shifter_0/reg_i_15_reg[10]  ( .D(\shifter_0/n10571 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[10] ) );
  dff_sg \shifter_0/reg_i_15_reg[11]  ( .D(\shifter_0/n10570 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[11] ) );
  dff_sg \shifter_0/reg_i_15_reg[12]  ( .D(\shifter_0/n10569 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[12] ) );
  dff_sg \shifter_0/reg_i_15_reg[13]  ( .D(\shifter_0/n10568 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[13] ) );
  dff_sg \shifter_0/reg_i_15_reg[14]  ( .D(\shifter_0/n10567 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[14] ) );
  dff_sg \shifter_0/reg_i_15_reg[15]  ( .D(\shifter_0/n10566 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[15] ) );
  dff_sg \shifter_0/reg_i_15_reg[16]  ( .D(\shifter_0/n10565 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[16] ) );
  dff_sg \shifter_0/reg_i_15_reg[17]  ( .D(\shifter_0/n10564 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[17] ) );
  dff_sg \shifter_0/reg_i_15_reg[18]  ( .D(\shifter_0/n10563 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[18] ) );
  dff_sg \shifter_0/reg_i_15_reg[19]  ( .D(\shifter_0/n10562 ), .CP(clk), .Q(
        \shifter_0/reg_i_15[19] ) );
  dff_sg \shifter_0/reg_w_0_reg[0]  ( .D(\shifter_0/n10561 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[0] ) );
  dff_sg \shifter_0/reg_w_0_reg[1]  ( .D(\shifter_0/n10560 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[1] ) );
  dff_sg \shifter_0/reg_w_0_reg[2]  ( .D(\shifter_0/n10559 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[2] ) );
  dff_sg \shifter_0/reg_w_0_reg[3]  ( .D(\shifter_0/n10558 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[3] ) );
  dff_sg \shifter_0/reg_w_0_reg[4]  ( .D(\shifter_0/n10557 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[4] ) );
  dff_sg \shifter_0/reg_w_0_reg[5]  ( .D(\shifter_0/n10556 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[5] ) );
  dff_sg \shifter_0/reg_w_0_reg[6]  ( .D(\shifter_0/n10555 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[6] ) );
  dff_sg \shifter_0/reg_w_0_reg[7]  ( .D(\shifter_0/n10554 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[7] ) );
  dff_sg \shifter_0/reg_w_0_reg[8]  ( .D(\shifter_0/n10553 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[8] ) );
  dff_sg \shifter_0/reg_w_0_reg[9]  ( .D(\shifter_0/n10552 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[9] ) );
  dff_sg \shifter_0/reg_w_0_reg[10]  ( .D(\shifter_0/n10551 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[10] ) );
  dff_sg \shifter_0/reg_w_0_reg[11]  ( .D(\shifter_0/n10550 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[11] ) );
  dff_sg \shifter_0/reg_w_0_reg[12]  ( .D(\shifter_0/n10549 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[12] ) );
  dff_sg \shifter_0/reg_w_0_reg[13]  ( .D(\shifter_0/n10548 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[13] ) );
  dff_sg \shifter_0/reg_w_0_reg[14]  ( .D(\shifter_0/n10547 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[14] ) );
  dff_sg \shifter_0/reg_w_0_reg[15]  ( .D(\shifter_0/n10546 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[15] ) );
  dff_sg \shifter_0/reg_w_0_reg[16]  ( .D(\shifter_0/n10545 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[16] ) );
  dff_sg \shifter_0/reg_w_0_reg[17]  ( .D(\shifter_0/n10544 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[17] ) );
  dff_sg \shifter_0/reg_w_0_reg[18]  ( .D(\shifter_0/n10543 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[18] ) );
  dff_sg \shifter_0/reg_w_0_reg[19]  ( .D(\shifter_0/n10542 ), .CP(clk), .Q(
        \shifter_0/reg_w_0[19] ) );
  dff_sg \shifter_0/reg_w_1_reg[0]  ( .D(\shifter_0/n10541 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[0] ) );
  dff_sg \shifter_0/reg_w_1_reg[1]  ( .D(\shifter_0/n10540 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[1] ) );
  dff_sg \shifter_0/reg_w_1_reg[2]  ( .D(\shifter_0/n10539 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[2] ) );
  dff_sg \shifter_0/reg_w_1_reg[3]  ( .D(\shifter_0/n10538 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[3] ) );
  dff_sg \shifter_0/reg_w_1_reg[4]  ( .D(\shifter_0/n10537 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[4] ) );
  dff_sg \shifter_0/reg_w_1_reg[5]  ( .D(\shifter_0/n10536 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[5] ) );
  dff_sg \shifter_0/reg_w_1_reg[6]  ( .D(\shifter_0/n10535 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[6] ) );
  dff_sg \shifter_0/reg_w_1_reg[7]  ( .D(\shifter_0/n10534 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[7] ) );
  dff_sg \shifter_0/reg_w_1_reg[8]  ( .D(\shifter_0/n10533 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[8] ) );
  dff_sg \shifter_0/reg_w_1_reg[9]  ( .D(\shifter_0/n10532 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[9] ) );
  dff_sg \shifter_0/reg_w_1_reg[10]  ( .D(\shifter_0/n10531 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[10] ) );
  dff_sg \shifter_0/reg_w_1_reg[11]  ( .D(\shifter_0/n10530 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[11] ) );
  dff_sg \shifter_0/reg_w_1_reg[12]  ( .D(\shifter_0/n10529 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[12] ) );
  dff_sg \shifter_0/reg_w_1_reg[13]  ( .D(\shifter_0/n10528 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[13] ) );
  dff_sg \shifter_0/reg_w_1_reg[14]  ( .D(\shifter_0/n10527 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[14] ) );
  dff_sg \shifter_0/reg_w_1_reg[15]  ( .D(\shifter_0/n10526 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[15] ) );
  dff_sg \shifter_0/reg_w_1_reg[16]  ( .D(\shifter_0/n10525 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[16] ) );
  dff_sg \shifter_0/reg_w_1_reg[17]  ( .D(\shifter_0/n10524 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[17] ) );
  dff_sg \shifter_0/reg_w_1_reg[18]  ( .D(\shifter_0/n10523 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[18] ) );
  dff_sg \shifter_0/reg_w_1_reg[19]  ( .D(\shifter_0/n10522 ), .CP(clk), .Q(
        \shifter_0/reg_w_1[19] ) );
  dff_sg \shifter_0/reg_w_2_reg[0]  ( .D(\shifter_0/n10521 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[0] ) );
  dff_sg \shifter_0/reg_w_2_reg[1]  ( .D(\shifter_0/n10520 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[1] ) );
  dff_sg \shifter_0/reg_w_2_reg[2]  ( .D(\shifter_0/n10519 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[2] ) );
  dff_sg \shifter_0/reg_w_2_reg[3]  ( .D(\shifter_0/n10518 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[3] ) );
  dff_sg \shifter_0/reg_w_2_reg[4]  ( .D(\shifter_0/n10517 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[4] ) );
  dff_sg \shifter_0/reg_w_2_reg[5]  ( .D(\shifter_0/n10516 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[5] ) );
  dff_sg \shifter_0/reg_w_2_reg[6]  ( .D(\shifter_0/n10515 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[6] ) );
  dff_sg \shifter_0/reg_w_2_reg[7]  ( .D(\shifter_0/n10514 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[7] ) );
  dff_sg \shifter_0/reg_w_2_reg[8]  ( .D(\shifter_0/n10513 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[8] ) );
  dff_sg \shifter_0/reg_w_2_reg[9]  ( .D(\shifter_0/n10512 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[9] ) );
  dff_sg \shifter_0/reg_w_2_reg[10]  ( .D(\shifter_0/n10511 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[10] ) );
  dff_sg \shifter_0/reg_w_2_reg[11]  ( .D(\shifter_0/n10510 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[11] ) );
  dff_sg \shifter_0/reg_w_2_reg[12]  ( .D(\shifter_0/n10509 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[12] ) );
  dff_sg \shifter_0/reg_w_2_reg[13]  ( .D(\shifter_0/n10508 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[13] ) );
  dff_sg \shifter_0/reg_w_2_reg[14]  ( .D(\shifter_0/n10507 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[14] ) );
  dff_sg \shifter_0/reg_w_2_reg[15]  ( .D(\shifter_0/n10506 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[15] ) );
  dff_sg \shifter_0/reg_w_2_reg[16]  ( .D(\shifter_0/n10505 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[16] ) );
  dff_sg \shifter_0/reg_w_2_reg[17]  ( .D(\shifter_0/n10504 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[17] ) );
  dff_sg \shifter_0/reg_w_2_reg[18]  ( .D(\shifter_0/n10503 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[18] ) );
  dff_sg \shifter_0/reg_w_2_reg[19]  ( .D(\shifter_0/n10502 ), .CP(clk), .Q(
        \shifter_0/reg_w_2[19] ) );
  dff_sg \shifter_0/reg_w_3_reg[0]  ( .D(\shifter_0/n10501 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[0] ) );
  dff_sg \shifter_0/reg_w_3_reg[1]  ( .D(\shifter_0/n10500 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[1] ) );
  dff_sg \shifter_0/reg_w_3_reg[2]  ( .D(\shifter_0/n10499 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[2] ) );
  dff_sg \shifter_0/reg_w_3_reg[3]  ( .D(\shifter_0/n10498 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[3] ) );
  dff_sg \shifter_0/reg_w_3_reg[4]  ( .D(\shifter_0/n10497 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[4] ) );
  dff_sg \shifter_0/reg_w_3_reg[5]  ( .D(\shifter_0/n10496 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[5] ) );
  dff_sg \shifter_0/reg_w_3_reg[6]  ( .D(\shifter_0/n10495 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[6] ) );
  dff_sg \shifter_0/reg_w_3_reg[7]  ( .D(\shifter_0/n10494 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[7] ) );
  dff_sg \shifter_0/reg_w_3_reg[8]  ( .D(\shifter_0/n10493 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[8] ) );
  dff_sg \shifter_0/reg_w_3_reg[9]  ( .D(\shifter_0/n10492 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[9] ) );
  dff_sg \shifter_0/reg_w_3_reg[10]  ( .D(\shifter_0/n10491 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[10] ) );
  dff_sg \shifter_0/reg_w_3_reg[11]  ( .D(\shifter_0/n10490 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[11] ) );
  dff_sg \shifter_0/reg_w_3_reg[12]  ( .D(\shifter_0/n10489 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[12] ) );
  dff_sg \shifter_0/reg_w_3_reg[13]  ( .D(\shifter_0/n10488 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[13] ) );
  dff_sg \shifter_0/reg_w_3_reg[14]  ( .D(\shifter_0/n10487 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[14] ) );
  dff_sg \shifter_0/reg_w_3_reg[15]  ( .D(\shifter_0/n10486 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[15] ) );
  dff_sg \shifter_0/reg_w_3_reg[16]  ( .D(\shifter_0/n10485 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[16] ) );
  dff_sg \shifter_0/reg_w_3_reg[17]  ( .D(\shifter_0/n10484 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[17] ) );
  dff_sg \shifter_0/reg_w_3_reg[18]  ( .D(\shifter_0/n10483 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[18] ) );
  dff_sg \shifter_0/reg_w_3_reg[19]  ( .D(\shifter_0/n10482 ), .CP(clk), .Q(
        \shifter_0/reg_w_3[19] ) );
  dff_sg \shifter_0/reg_w_4_reg[0]  ( .D(\shifter_0/n10481 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[0] ) );
  dff_sg \shifter_0/reg_w_4_reg[1]  ( .D(\shifter_0/n10480 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[1] ) );
  dff_sg \shifter_0/reg_w_4_reg[2]  ( .D(\shifter_0/n10479 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[2] ) );
  dff_sg \shifter_0/reg_w_4_reg[3]  ( .D(\shifter_0/n10478 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[3] ) );
  dff_sg \shifter_0/reg_w_4_reg[4]  ( .D(\shifter_0/n10477 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[4] ) );
  dff_sg \shifter_0/reg_w_4_reg[5]  ( .D(\shifter_0/n10476 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[5] ) );
  dff_sg \shifter_0/reg_w_4_reg[6]  ( .D(\shifter_0/n10475 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[6] ) );
  dff_sg \shifter_0/reg_w_4_reg[7]  ( .D(\shifter_0/n10474 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[7] ) );
  dff_sg \shifter_0/reg_w_4_reg[8]  ( .D(\shifter_0/n10473 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[8] ) );
  dff_sg \shifter_0/reg_w_4_reg[9]  ( .D(\shifter_0/n10472 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[9] ) );
  dff_sg \shifter_0/reg_w_4_reg[10]  ( .D(\shifter_0/n10471 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[10] ) );
  dff_sg \shifter_0/reg_w_4_reg[11]  ( .D(\shifter_0/n10470 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[11] ) );
  dff_sg \shifter_0/reg_w_4_reg[12]  ( .D(\shifter_0/n10469 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[12] ) );
  dff_sg \shifter_0/reg_w_4_reg[13]  ( .D(\shifter_0/n10468 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[13] ) );
  dff_sg \shifter_0/reg_w_4_reg[14]  ( .D(\shifter_0/n10467 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[14] ) );
  dff_sg \shifter_0/reg_w_4_reg[15]  ( .D(\shifter_0/n10466 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[15] ) );
  dff_sg \shifter_0/reg_w_4_reg[16]  ( .D(\shifter_0/n10465 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[16] ) );
  dff_sg \shifter_0/reg_w_4_reg[17]  ( .D(\shifter_0/n10464 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[17] ) );
  dff_sg \shifter_0/reg_w_4_reg[18]  ( .D(\shifter_0/n10463 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[18] ) );
  dff_sg \shifter_0/reg_w_4_reg[19]  ( .D(\shifter_0/n10462 ), .CP(clk), .Q(
        \shifter_0/reg_w_4[19] ) );
  dff_sg \shifter_0/reg_w_5_reg[0]  ( .D(\shifter_0/n10461 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[0] ) );
  dff_sg \shifter_0/reg_w_5_reg[1]  ( .D(\shifter_0/n10460 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[1] ) );
  dff_sg \shifter_0/reg_w_5_reg[2]  ( .D(\shifter_0/n10459 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[2] ) );
  dff_sg \shifter_0/reg_w_5_reg[3]  ( .D(\shifter_0/n10458 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[3] ) );
  dff_sg \shifter_0/reg_w_5_reg[4]  ( .D(\shifter_0/n10457 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[4] ) );
  dff_sg \shifter_0/reg_w_5_reg[5]  ( .D(\shifter_0/n10456 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[5] ) );
  dff_sg \shifter_0/reg_w_5_reg[6]  ( .D(\shifter_0/n10455 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[6] ) );
  dff_sg \shifter_0/reg_w_5_reg[7]  ( .D(\shifter_0/n10454 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[7] ) );
  dff_sg \shifter_0/reg_w_5_reg[8]  ( .D(\shifter_0/n10453 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[8] ) );
  dff_sg \shifter_0/reg_w_5_reg[9]  ( .D(\shifter_0/n10452 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[9] ) );
  dff_sg \shifter_0/reg_w_5_reg[10]  ( .D(\shifter_0/n10451 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[10] ) );
  dff_sg \shifter_0/reg_w_5_reg[11]  ( .D(\shifter_0/n10450 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[11] ) );
  dff_sg \shifter_0/reg_w_5_reg[12]  ( .D(\shifter_0/n10449 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[12] ) );
  dff_sg \shifter_0/reg_w_5_reg[13]  ( .D(\shifter_0/n10448 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[13] ) );
  dff_sg \shifter_0/reg_w_5_reg[14]  ( .D(\shifter_0/n10447 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[14] ) );
  dff_sg \shifter_0/reg_w_5_reg[15]  ( .D(\shifter_0/n10446 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[15] ) );
  dff_sg \shifter_0/reg_w_5_reg[16]  ( .D(\shifter_0/n10445 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[16] ) );
  dff_sg \shifter_0/reg_w_5_reg[17]  ( .D(\shifter_0/n10444 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[17] ) );
  dff_sg \shifter_0/reg_w_5_reg[18]  ( .D(\shifter_0/n10443 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[18] ) );
  dff_sg \shifter_0/reg_w_5_reg[19]  ( .D(\shifter_0/n10442 ), .CP(clk), .Q(
        \shifter_0/reg_w_5[19] ) );
  dff_sg \shifter_0/reg_w_6_reg[0]  ( .D(\shifter_0/n10441 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[0] ) );
  dff_sg \shifter_0/reg_w_6_reg[1]  ( .D(\shifter_0/n10440 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[1] ) );
  dff_sg \shifter_0/reg_w_6_reg[2]  ( .D(\shifter_0/n10439 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[2] ) );
  dff_sg \shifter_0/reg_w_6_reg[3]  ( .D(\shifter_0/n10438 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[3] ) );
  dff_sg \shifter_0/reg_w_6_reg[4]  ( .D(\shifter_0/n10437 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[4] ) );
  dff_sg \shifter_0/reg_w_6_reg[5]  ( .D(\shifter_0/n10436 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[5] ) );
  dff_sg \shifter_0/reg_w_6_reg[6]  ( .D(\shifter_0/n10435 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[6] ) );
  dff_sg \shifter_0/reg_w_6_reg[7]  ( .D(\shifter_0/n10434 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[7] ) );
  dff_sg \shifter_0/reg_w_6_reg[8]  ( .D(\shifter_0/n10433 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[8] ) );
  dff_sg \shifter_0/reg_w_6_reg[9]  ( .D(\shifter_0/n10432 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[9] ) );
  dff_sg \shifter_0/reg_w_6_reg[10]  ( .D(\shifter_0/n10431 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[10] ) );
  dff_sg \shifter_0/reg_w_6_reg[11]  ( .D(\shifter_0/n10430 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[11] ) );
  dff_sg \shifter_0/reg_w_6_reg[12]  ( .D(\shifter_0/n10429 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[12] ) );
  dff_sg \shifter_0/reg_w_6_reg[13]  ( .D(\shifter_0/n10428 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[13] ) );
  dff_sg \shifter_0/reg_w_6_reg[14]  ( .D(\shifter_0/n10427 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[14] ) );
  dff_sg \shifter_0/reg_w_6_reg[15]  ( .D(\shifter_0/n10426 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[15] ) );
  dff_sg \shifter_0/reg_w_6_reg[16]  ( .D(\shifter_0/n10425 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[16] ) );
  dff_sg \shifter_0/reg_w_6_reg[17]  ( .D(\shifter_0/n10424 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[17] ) );
  dff_sg \shifter_0/reg_w_6_reg[18]  ( .D(\shifter_0/n10423 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[18] ) );
  dff_sg \shifter_0/reg_w_6_reg[19]  ( .D(\shifter_0/n10422 ), .CP(clk), .Q(
        \shifter_0/reg_w_6[19] ) );
  dff_sg \shifter_0/reg_w_7_reg[0]  ( .D(\shifter_0/n10421 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[0] ) );
  dff_sg \shifter_0/reg_w_7_reg[1]  ( .D(\shifter_0/n10420 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[1] ) );
  dff_sg \shifter_0/reg_w_7_reg[2]  ( .D(\shifter_0/n10419 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[2] ) );
  dff_sg \shifter_0/reg_w_7_reg[3]  ( .D(\shifter_0/n10418 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[3] ) );
  dff_sg \shifter_0/reg_w_7_reg[4]  ( .D(\shifter_0/n10417 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[4] ) );
  dff_sg \shifter_0/reg_w_7_reg[5]  ( .D(\shifter_0/n10416 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[5] ) );
  dff_sg \shifter_0/reg_w_7_reg[6]  ( .D(\shifter_0/n10415 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[6] ) );
  dff_sg \shifter_0/reg_w_7_reg[7]  ( .D(\shifter_0/n10414 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[7] ) );
  dff_sg \shifter_0/reg_w_7_reg[8]  ( .D(\shifter_0/n10413 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[8] ) );
  dff_sg \shifter_0/reg_w_7_reg[9]  ( .D(\shifter_0/n10412 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[9] ) );
  dff_sg \shifter_0/reg_w_7_reg[10]  ( .D(\shifter_0/n10411 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[10] ) );
  dff_sg \shifter_0/reg_w_7_reg[11]  ( .D(\shifter_0/n10410 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[11] ) );
  dff_sg \shifter_0/reg_w_7_reg[12]  ( .D(\shifter_0/n10409 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[12] ) );
  dff_sg \shifter_0/reg_w_7_reg[13]  ( .D(\shifter_0/n10408 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[13] ) );
  dff_sg \shifter_0/reg_w_7_reg[14]  ( .D(\shifter_0/n10407 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[14] ) );
  dff_sg \shifter_0/reg_w_7_reg[15]  ( .D(\shifter_0/n10406 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[15] ) );
  dff_sg \shifter_0/reg_w_7_reg[16]  ( .D(\shifter_0/n10405 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[16] ) );
  dff_sg \shifter_0/reg_w_7_reg[17]  ( .D(\shifter_0/n10404 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[17] ) );
  dff_sg \shifter_0/reg_w_7_reg[18]  ( .D(\shifter_0/n10403 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[18] ) );
  dff_sg \shifter_0/reg_w_7_reg[19]  ( .D(\shifter_0/n10402 ), .CP(clk), .Q(
        \shifter_0/reg_w_7[19] ) );
  dff_sg \shifter_0/reg_w_8_reg[0]  ( .D(\shifter_0/n10401 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[0] ) );
  dff_sg \shifter_0/reg_w_8_reg[1]  ( .D(\shifter_0/n10400 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[1] ) );
  dff_sg \shifter_0/reg_w_8_reg[2]  ( .D(\shifter_0/n10399 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[2] ) );
  dff_sg \shifter_0/reg_w_8_reg[3]  ( .D(\shifter_0/n10398 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[3] ) );
  dff_sg \shifter_0/reg_w_8_reg[4]  ( .D(\shifter_0/n10397 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[4] ) );
  dff_sg \shifter_0/reg_w_8_reg[5]  ( .D(\shifter_0/n10396 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[5] ) );
  dff_sg \shifter_0/reg_w_8_reg[6]  ( .D(\shifter_0/n10395 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[6] ) );
  dff_sg \shifter_0/reg_w_8_reg[7]  ( .D(\shifter_0/n10394 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[7] ) );
  dff_sg \shifter_0/reg_w_8_reg[8]  ( .D(\shifter_0/n10393 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[8] ) );
  dff_sg \shifter_0/reg_w_8_reg[9]  ( .D(\shifter_0/n10392 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[9] ) );
  dff_sg \shifter_0/reg_w_8_reg[10]  ( .D(\shifter_0/n10391 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[10] ) );
  dff_sg \shifter_0/reg_w_8_reg[11]  ( .D(\shifter_0/n10390 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[11] ) );
  dff_sg \shifter_0/reg_w_8_reg[12]  ( .D(\shifter_0/n10389 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[12] ) );
  dff_sg \shifter_0/reg_w_8_reg[13]  ( .D(\shifter_0/n10388 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[13] ) );
  dff_sg \shifter_0/reg_w_8_reg[14]  ( .D(\shifter_0/n10387 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[14] ) );
  dff_sg \shifter_0/reg_w_8_reg[15]  ( .D(\shifter_0/n10386 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[15] ) );
  dff_sg \shifter_0/reg_w_8_reg[16]  ( .D(\shifter_0/n10385 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[16] ) );
  dff_sg \shifter_0/reg_w_8_reg[17]  ( .D(\shifter_0/n10384 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[17] ) );
  dff_sg \shifter_0/reg_w_8_reg[18]  ( .D(\shifter_0/n10383 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[18] ) );
  dff_sg \shifter_0/reg_w_8_reg[19]  ( .D(\shifter_0/n10382 ), .CP(clk), .Q(
        \shifter_0/reg_w_8[19] ) );
  dff_sg \shifter_0/reg_w_9_reg[0]  ( .D(\shifter_0/n10381 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[0] ) );
  dff_sg \shifter_0/reg_w_9_reg[1]  ( .D(\shifter_0/n10380 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[1] ) );
  dff_sg \shifter_0/reg_w_9_reg[2]  ( .D(\shifter_0/n10379 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[2] ) );
  dff_sg \shifter_0/reg_w_9_reg[3]  ( .D(\shifter_0/n10378 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[3] ) );
  dff_sg \shifter_0/reg_w_9_reg[4]  ( .D(\shifter_0/n10377 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[4] ) );
  dff_sg \shifter_0/reg_w_9_reg[5]  ( .D(\shifter_0/n10376 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[5] ) );
  dff_sg \shifter_0/reg_w_9_reg[6]  ( .D(\shifter_0/n10375 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[6] ) );
  dff_sg \shifter_0/reg_w_9_reg[7]  ( .D(\shifter_0/n10374 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[7] ) );
  dff_sg \shifter_0/reg_w_9_reg[8]  ( .D(\shifter_0/n10373 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[8] ) );
  dff_sg \shifter_0/reg_w_9_reg[9]  ( .D(\shifter_0/n10372 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[9] ) );
  dff_sg \shifter_0/reg_w_9_reg[10]  ( .D(\shifter_0/n10371 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[10] ) );
  dff_sg \shifter_0/reg_w_9_reg[11]  ( .D(\shifter_0/n10370 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[11] ) );
  dff_sg \shifter_0/reg_w_9_reg[12]  ( .D(\shifter_0/n10369 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[12] ) );
  dff_sg \shifter_0/reg_w_9_reg[13]  ( .D(\shifter_0/n10368 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[13] ) );
  dff_sg \shifter_0/reg_w_9_reg[14]  ( .D(\shifter_0/n10367 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[14] ) );
  dff_sg \shifter_0/reg_w_9_reg[15]  ( .D(\shifter_0/n10366 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[15] ) );
  dff_sg \shifter_0/reg_w_9_reg[16]  ( .D(\shifter_0/n10365 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[16] ) );
  dff_sg \shifter_0/reg_w_9_reg[17]  ( .D(\shifter_0/n10364 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[17] ) );
  dff_sg \shifter_0/reg_w_9_reg[18]  ( .D(\shifter_0/n10363 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[18] ) );
  dff_sg \shifter_0/reg_w_9_reg[19]  ( .D(\shifter_0/n10362 ), .CP(clk), .Q(
        \shifter_0/reg_w_9[19] ) );
  dff_sg \shifter_0/reg_w_10_reg[0]  ( .D(\shifter_0/n10361 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[0] ) );
  dff_sg \shifter_0/reg_w_10_reg[1]  ( .D(\shifter_0/n10360 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[1] ) );
  dff_sg \shifter_0/reg_w_10_reg[2]  ( .D(\shifter_0/n10359 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[2] ) );
  dff_sg \shifter_0/reg_w_10_reg[3]  ( .D(\shifter_0/n10358 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[3] ) );
  dff_sg \shifter_0/reg_w_10_reg[4]  ( .D(\shifter_0/n10357 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[4] ) );
  dff_sg \shifter_0/reg_w_10_reg[5]  ( .D(\shifter_0/n10356 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[5] ) );
  dff_sg \shifter_0/reg_w_10_reg[6]  ( .D(\shifter_0/n10355 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[6] ) );
  dff_sg \shifter_0/reg_w_10_reg[7]  ( .D(\shifter_0/n10354 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[7] ) );
  dff_sg \shifter_0/reg_w_10_reg[8]  ( .D(\shifter_0/n10353 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[8] ) );
  dff_sg \shifter_0/reg_w_10_reg[9]  ( .D(\shifter_0/n10352 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[9] ) );
  dff_sg \shifter_0/reg_w_10_reg[10]  ( .D(\shifter_0/n10351 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[10] ) );
  dff_sg \shifter_0/reg_w_10_reg[11]  ( .D(\shifter_0/n10350 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[11] ) );
  dff_sg \shifter_0/reg_w_10_reg[12]  ( .D(\shifter_0/n10349 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[12] ) );
  dff_sg \shifter_0/reg_w_10_reg[13]  ( .D(\shifter_0/n10348 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[13] ) );
  dff_sg \shifter_0/reg_w_10_reg[14]  ( .D(\shifter_0/n10347 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[14] ) );
  dff_sg \shifter_0/reg_w_10_reg[15]  ( .D(\shifter_0/n10346 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[15] ) );
  dff_sg \shifter_0/reg_w_10_reg[16]  ( .D(\shifter_0/n10345 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[16] ) );
  dff_sg \shifter_0/reg_w_10_reg[17]  ( .D(\shifter_0/n10344 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[17] ) );
  dff_sg \shifter_0/reg_w_10_reg[18]  ( .D(\shifter_0/n10343 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[18] ) );
  dff_sg \shifter_0/reg_w_10_reg[19]  ( .D(\shifter_0/n10342 ), .CP(clk), .Q(
        \shifter_0/reg_w_10[19] ) );
  dff_sg \shifter_0/reg_w_11_reg[0]  ( .D(\shifter_0/n10341 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[0] ) );
  dff_sg \shifter_0/reg_w_11_reg[1]  ( .D(\shifter_0/n10340 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[1] ) );
  dff_sg \shifter_0/reg_w_11_reg[2]  ( .D(\shifter_0/n10339 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[2] ) );
  dff_sg \shifter_0/reg_w_11_reg[3]  ( .D(\shifter_0/n10338 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[3] ) );
  dff_sg \shifter_0/reg_w_11_reg[4]  ( .D(\shifter_0/n10337 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[4] ) );
  dff_sg \shifter_0/reg_w_11_reg[5]  ( .D(\shifter_0/n10336 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[5] ) );
  dff_sg \shifter_0/reg_w_11_reg[6]  ( .D(\shifter_0/n10335 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[6] ) );
  dff_sg \shifter_0/reg_w_11_reg[7]  ( .D(\shifter_0/n10334 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[7] ) );
  dff_sg \shifter_0/reg_w_11_reg[8]  ( .D(\shifter_0/n10333 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[8] ) );
  dff_sg \shifter_0/reg_w_11_reg[9]  ( .D(\shifter_0/n10332 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[9] ) );
  dff_sg \shifter_0/reg_w_11_reg[10]  ( .D(\shifter_0/n10331 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[10] ) );
  dff_sg \shifter_0/reg_w_11_reg[11]  ( .D(\shifter_0/n10330 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[11] ) );
  dff_sg \shifter_0/reg_w_11_reg[12]  ( .D(\shifter_0/n10329 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[12] ) );
  dff_sg \shifter_0/reg_w_11_reg[13]  ( .D(\shifter_0/n10328 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[13] ) );
  dff_sg \shifter_0/reg_w_11_reg[14]  ( .D(\shifter_0/n10327 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[14] ) );
  dff_sg \shifter_0/reg_w_11_reg[15]  ( .D(\shifter_0/n10326 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[15] ) );
  dff_sg \shifter_0/reg_w_11_reg[16]  ( .D(\shifter_0/n10325 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[16] ) );
  dff_sg \shifter_0/reg_w_11_reg[17]  ( .D(\shifter_0/n10324 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[17] ) );
  dff_sg \shifter_0/reg_w_11_reg[18]  ( .D(\shifter_0/n10323 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[18] ) );
  dff_sg \shifter_0/reg_w_11_reg[19]  ( .D(\shifter_0/n10322 ), .CP(clk), .Q(
        \shifter_0/reg_w_11[19] ) );
  dff_sg \shifter_0/reg_w_12_reg[0]  ( .D(\shifter_0/n10321 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[0] ) );
  dff_sg \shifter_0/reg_w_12_reg[1]  ( .D(\shifter_0/n10320 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[1] ) );
  dff_sg \shifter_0/reg_w_12_reg[2]  ( .D(\shifter_0/n10319 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[2] ) );
  dff_sg \shifter_0/reg_w_12_reg[3]  ( .D(\shifter_0/n10318 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[3] ) );
  dff_sg \shifter_0/reg_w_12_reg[4]  ( .D(\shifter_0/n10317 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[4] ) );
  dff_sg \shifter_0/reg_w_12_reg[5]  ( .D(\shifter_0/n10316 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[5] ) );
  dff_sg \shifter_0/reg_w_12_reg[6]  ( .D(\shifter_0/n10315 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[6] ) );
  dff_sg \shifter_0/reg_w_12_reg[7]  ( .D(\shifter_0/n10314 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[7] ) );
  dff_sg \shifter_0/reg_w_12_reg[8]  ( .D(\shifter_0/n10313 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[8] ) );
  dff_sg \shifter_0/reg_w_12_reg[9]  ( .D(\shifter_0/n10312 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[9] ) );
  dff_sg \shifter_0/reg_w_12_reg[10]  ( .D(\shifter_0/n10311 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[10] ) );
  dff_sg \shifter_0/reg_w_12_reg[11]  ( .D(\shifter_0/n10310 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[11] ) );
  dff_sg \shifter_0/reg_w_12_reg[12]  ( .D(\shifter_0/n10309 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[12] ) );
  dff_sg \shifter_0/reg_w_12_reg[13]  ( .D(\shifter_0/n10308 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[13] ) );
  dff_sg \shifter_0/reg_w_12_reg[14]  ( .D(\shifter_0/n10307 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[14] ) );
  dff_sg \shifter_0/reg_w_12_reg[15]  ( .D(\shifter_0/n10306 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[15] ) );
  dff_sg \shifter_0/reg_w_12_reg[16]  ( .D(\shifter_0/n10305 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[16] ) );
  dff_sg \shifter_0/reg_w_12_reg[17]  ( .D(\shifter_0/n10304 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[17] ) );
  dff_sg \shifter_0/reg_w_12_reg[18]  ( .D(\shifter_0/n10303 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[18] ) );
  dff_sg \shifter_0/reg_w_12_reg[19]  ( .D(\shifter_0/n10302 ), .CP(clk), .Q(
        \shifter_0/reg_w_12[19] ) );
  dff_sg \shifter_0/reg_w_13_reg[0]  ( .D(\shifter_0/n10301 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[0] ) );
  dff_sg \shifter_0/reg_w_13_reg[1]  ( .D(\shifter_0/n10300 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[1] ) );
  dff_sg \shifter_0/reg_w_13_reg[2]  ( .D(\shifter_0/n10299 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[2] ) );
  dff_sg \shifter_0/reg_w_13_reg[3]  ( .D(\shifter_0/n10298 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[3] ) );
  dff_sg \shifter_0/reg_w_13_reg[4]  ( .D(\shifter_0/n10297 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[4] ) );
  dff_sg \shifter_0/reg_w_13_reg[5]  ( .D(\shifter_0/n10296 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[5] ) );
  dff_sg \shifter_0/reg_w_13_reg[6]  ( .D(\shifter_0/n10295 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[6] ) );
  dff_sg \shifter_0/reg_w_13_reg[7]  ( .D(\shifter_0/n10294 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[7] ) );
  dff_sg \shifter_0/reg_w_13_reg[8]  ( .D(\shifter_0/n10293 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[8] ) );
  dff_sg \shifter_0/reg_w_13_reg[9]  ( .D(\shifter_0/n10292 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[9] ) );
  dff_sg \shifter_0/reg_w_13_reg[10]  ( .D(\shifter_0/n10291 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[10] ) );
  dff_sg \shifter_0/reg_w_13_reg[11]  ( .D(\shifter_0/n10290 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[11] ) );
  dff_sg \shifter_0/reg_w_13_reg[12]  ( .D(\shifter_0/n10289 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[12] ) );
  dff_sg \shifter_0/reg_w_13_reg[13]  ( .D(\shifter_0/n10288 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[13] ) );
  dff_sg \shifter_0/reg_w_13_reg[14]  ( .D(\shifter_0/n10287 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[14] ) );
  dff_sg \shifter_0/reg_w_13_reg[15]  ( .D(\shifter_0/n10286 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[15] ) );
  dff_sg \shifter_0/reg_w_13_reg[16]  ( .D(\shifter_0/n10285 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[16] ) );
  dff_sg \shifter_0/reg_w_13_reg[17]  ( .D(\shifter_0/n10284 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[17] ) );
  dff_sg \shifter_0/reg_w_13_reg[18]  ( .D(\shifter_0/n10283 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[18] ) );
  dff_sg \shifter_0/reg_w_13_reg[19]  ( .D(\shifter_0/n10282 ), .CP(clk), .Q(
        \shifter_0/reg_w_13[19] ) );
  dff_sg \shifter_0/reg_w_14_reg[0]  ( .D(\shifter_0/n10281 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[0] ) );
  dff_sg \shifter_0/reg_w_14_reg[1]  ( .D(\shifter_0/n10280 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[1] ) );
  dff_sg \shifter_0/reg_w_14_reg[2]  ( .D(\shifter_0/n10279 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[2] ) );
  dff_sg \shifter_0/reg_w_14_reg[3]  ( .D(\shifter_0/n10278 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[3] ) );
  dff_sg \shifter_0/reg_w_14_reg[4]  ( .D(\shifter_0/n10277 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[4] ) );
  dff_sg \shifter_0/reg_w_14_reg[5]  ( .D(\shifter_0/n10276 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[5] ) );
  dff_sg \shifter_0/reg_w_14_reg[6]  ( .D(\shifter_0/n10275 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[6] ) );
  dff_sg \shifter_0/reg_w_14_reg[7]  ( .D(\shifter_0/n10274 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[7] ) );
  dff_sg \shifter_0/reg_w_14_reg[8]  ( .D(\shifter_0/n10273 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[8] ) );
  dff_sg \shifter_0/reg_w_14_reg[9]  ( .D(\shifter_0/n10272 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[9] ) );
  dff_sg \shifter_0/reg_w_14_reg[10]  ( .D(\shifter_0/n10271 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[10] ) );
  dff_sg \shifter_0/reg_w_14_reg[11]  ( .D(\shifter_0/n10270 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[11] ) );
  dff_sg \shifter_0/reg_w_14_reg[12]  ( .D(\shifter_0/n10269 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[12] ) );
  dff_sg \shifter_0/reg_w_14_reg[13]  ( .D(\shifter_0/n10268 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[13] ) );
  dff_sg \shifter_0/reg_w_14_reg[14]  ( .D(\shifter_0/n10267 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[14] ) );
  dff_sg \shifter_0/reg_w_14_reg[15]  ( .D(\shifter_0/n10266 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[15] ) );
  dff_sg \shifter_0/reg_w_14_reg[16]  ( .D(\shifter_0/n10265 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[16] ) );
  dff_sg \shifter_0/reg_w_14_reg[17]  ( .D(\shifter_0/n10264 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[17] ) );
  dff_sg \shifter_0/reg_w_14_reg[18]  ( .D(\shifter_0/n10263 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[18] ) );
  dff_sg \shifter_0/reg_w_14_reg[19]  ( .D(\shifter_0/n10262 ), .CP(clk), .Q(
        \shifter_0/reg_w_14[19] ) );
  dff_sg \shifter_0/reg_w_15_reg[0]  ( .D(\shifter_0/n10261 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[0] ) );
  dff_sg \shifter_0/reg_w_15_reg[1]  ( .D(\shifter_0/n10260 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[1] ) );
  dff_sg \shifter_0/reg_w_15_reg[2]  ( .D(\shifter_0/n10259 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[2] ) );
  dff_sg \shifter_0/reg_w_15_reg[3]  ( .D(\shifter_0/n10258 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[3] ) );
  dff_sg \shifter_0/reg_w_15_reg[4]  ( .D(\shifter_0/n10257 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[4] ) );
  dff_sg \shifter_0/reg_w_15_reg[5]  ( .D(\shifter_0/n10256 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[5] ) );
  dff_sg \shifter_0/reg_w_15_reg[6]  ( .D(\shifter_0/n10255 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[6] ) );
  dff_sg \shifter_0/reg_w_15_reg[7]  ( .D(\shifter_0/n10254 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[7] ) );
  dff_sg \shifter_0/reg_w_15_reg[8]  ( .D(\shifter_0/n10253 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[8] ) );
  dff_sg \shifter_0/reg_w_15_reg[9]  ( .D(\shifter_0/n10252 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[9] ) );
  dff_sg \shifter_0/reg_w_15_reg[10]  ( .D(\shifter_0/n10251 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[10] ) );
  dff_sg \shifter_0/reg_w_15_reg[11]  ( .D(\shifter_0/n10250 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[11] ) );
  dff_sg \shifter_0/reg_w_15_reg[12]  ( .D(\shifter_0/n10249 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[12] ) );
  dff_sg \shifter_0/reg_w_15_reg[13]  ( .D(\shifter_0/n10248 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[13] ) );
  dff_sg \shifter_0/reg_w_15_reg[14]  ( .D(\shifter_0/n10247 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[14] ) );
  dff_sg \shifter_0/reg_w_15_reg[15]  ( .D(\shifter_0/n10246 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[15] ) );
  dff_sg \shifter_0/reg_w_15_reg[16]  ( .D(\shifter_0/n10245 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[16] ) );
  dff_sg \shifter_0/reg_w_15_reg[17]  ( .D(\shifter_0/n10244 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[17] ) );
  dff_sg \shifter_0/reg_w_15_reg[18]  ( .D(\shifter_0/n10243 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[18] ) );
  dff_sg \shifter_0/reg_w_15_reg[19]  ( .D(\shifter_0/n10242 ), .CP(clk), .Q(
        \shifter_0/reg_w_15[19] ) );
  dff_sg \shifter_0/state_reg[0]  ( .D(\shifter_0/n10883 ), .CP(clk), .Q(
        shifter_state[0]) );
  dff_sg \shifter_0/state_reg[1]  ( .D(\shifter_0/n10884 ), .CP(clk), .Q(
        shifter_state[1]) );
  dff_sg \shifter_0/pointer_reg[0]  ( .D(\shifter_0/n10886 ), .CP(clk), .Q(
        \shifter_0/pointer[0] ) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n4984 ), 
        .force_10(\filter_0/n4985 ), .force_11(1'b0), .Q(\filter_0/n8243 ) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n4988 ), 
        .force_10(\filter_0/n4989 ), .force_11(1'b0), .Q(\filter_0/n8242 ) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n4992 ), 
        .force_10(\filter_0/n4993 ), .force_11(1'b0), .Q(\filter_0/n8241 ) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n4996 ), 
        .force_10(\filter_0/n4997 ), .force_11(1'b0), .Q(\filter_0/n8240 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5000 ), .force_10(\filter_0/n5001 ), 
        .force_11(1'b0), .Q(\filter_0/n8239 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5004 ), .force_10(\filter_0/n5005 ), 
        .force_11(1'b0), .Q(\filter_0/n8238 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5008 ), .force_10(\filter_0/n5009 ), 
        .force_11(1'b0), .Q(\filter_0/n8237 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5012 ), .force_10(\filter_0/n5013 ), 
        .force_11(1'b0), .Q(\filter_0/n8236 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5016 ), .force_10(\filter_0/n5017 ), 
        .force_11(1'b0), .Q(\filter_0/n8235 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5020 ), .force_10(\filter_0/n5021 ), 
        .force_11(1'b0), .Q(\filter_0/n8234 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5024 ), .force_10(\filter_0/n5025 ), 
        .force_11(1'b0), .Q(\filter_0/n8233 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5028 ), .force_10(\filter_0/n5029 ), 
        .force_11(1'b0), .Q(\filter_0/n8232 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5032 ), .force_10(\filter_0/n5033 ), 
        .force_11(1'b0), .Q(\filter_0/n8231 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5036 ), .force_10(\filter_0/n5037 ), 
        .force_11(1'b0), .Q(\filter_0/n8230 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5040 ), .force_10(
        \filter_0/n5041 ), .force_11(1'b0), .Q(\filter_0/n8229 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5044 ), .force_10(
        \filter_0/n5045 ), .force_11(1'b0), .Q(\filter_0/n8228 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5048 ), .force_10(
        \filter_0/n5049 ), .force_11(1'b0), .Q(\filter_0/n8227 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5052 ), .force_10(
        \filter_0/n5053 ), .force_11(1'b0), .Q(\filter_0/n8226 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5056 ), .force_10(
        \filter_0/n5057 ), .force_11(1'b0), .Q(\filter_0/n8225 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5060 ), .force_10(
        \filter_0/n5061 ), .force_11(1'b0), .Q(\filter_0/n8224 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5064 ), .force_10(
        \filter_0/n5065 ), .force_11(1'b0), .Q(\filter_0/n8223 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5068 ), .force_10(
        \filter_0/n5069 ), .force_11(1'b0), .Q(\filter_0/n8222 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5072 ), .force_10(
        \filter_0/n5073 ), .force_11(1'b0), .Q(\filter_0/n8221 ) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5076 ), .force_10(
        \filter_0/n5077 ), .force_11(1'b0), .Q(\filter_0/n8220 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5080 ), .force_10(\filter_0/n5081 ), 
        .force_11(1'b0), .Q(\filter_0/n8219 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5084 ), .force_10(\filter_0/n5085 ), 
        .force_11(1'b0), .Q(\filter_0/n8218 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5088 ), .force_10(\filter_0/n5089 ), 
        .force_11(1'b0), .Q(\filter_0/n8217 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5092 ), .force_10(\filter_0/n5093 ), 
        .force_11(1'b0), .Q(\filter_0/n8216 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5096 ), .force_10(\filter_0/n5097 ), 
        .force_11(1'b0), .Q(\filter_0/n8215 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5100 ), .force_10(\filter_0/n5101 ), 
        .force_11(1'b0), .Q(\filter_0/n8214 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5104 ), .force_10(\filter_0/n5105 ), 
        .force_11(1'b0), .Q(\filter_0/n8213 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5108 ), .force_10(\filter_0/n5109 ), 
        .force_11(1'b0), .Q(\filter_0/n8212 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5112 ), .force_10(\filter_0/n5113 ), 
        .force_11(1'b0), .Q(\filter_0/n8211 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5116 ), .force_10(\filter_0/n5117 ), 
        .force_11(1'b0), .Q(\filter_0/n8210 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5120 ), .force_10(
        \filter_0/n5121 ), .force_11(1'b0), .Q(\filter_0/n8209 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5124 ), .force_10(
        \filter_0/n5125 ), .force_11(1'b0), .Q(\filter_0/n8208 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5128 ), .force_10(
        \filter_0/n5129 ), .force_11(1'b0), .Q(\filter_0/n8207 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5132 ), .force_10(
        \filter_0/n5133 ), .force_11(1'b0), .Q(\filter_0/n8206 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5136 ), .force_10(
        \filter_0/n5137 ), .force_11(1'b0), .Q(\filter_0/n8205 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5140 ), .force_10(
        \filter_0/n5141 ), .force_11(1'b0), .Q(\filter_0/n8204 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5144 ), .force_10(
        \filter_0/n5145 ), .force_11(1'b0), .Q(\filter_0/n8203 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5148 ), .force_10(
        \filter_0/n5149 ), .force_11(1'b0), .Q(\filter_0/n8202 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5152 ), .force_10(
        \filter_0/n5153 ), .force_11(1'b0), .Q(\filter_0/n8201 ) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5156 ), .force_10(
        \filter_0/n5157 ), .force_11(1'b0), .Q(\filter_0/n8200 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5160 ), .force_10(\filter_0/n5161 ), 
        .force_11(1'b0), .Q(\filter_0/n8199 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5164 ), .force_10(\filter_0/n5165 ), 
        .force_11(1'b0), .Q(\filter_0/n8198 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5168 ), .force_10(\filter_0/n5169 ), 
        .force_11(1'b0), .Q(\filter_0/n8197 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5172 ), .force_10(\filter_0/n5173 ), 
        .force_11(1'b0), .Q(\filter_0/n8196 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5176 ), .force_10(\filter_0/n5177 ), 
        .force_11(1'b0), .Q(\filter_0/n8195 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5180 ), .force_10(\filter_0/n5181 ), 
        .force_11(1'b0), .Q(\filter_0/n8194 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5184 ), .force_10(\filter_0/n5185 ), 
        .force_11(1'b0), .Q(\filter_0/n8193 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5188 ), .force_10(\filter_0/n5189 ), 
        .force_11(1'b0), .Q(\filter_0/n8192 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5192 ), .force_10(\filter_0/n5193 ), 
        .force_11(1'b0), .Q(\filter_0/n8191 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5196 ), .force_10(\filter_0/n5197 ), 
        .force_11(1'b0), .Q(\filter_0/n8190 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5200 ), .force_10(
        \filter_0/n5201 ), .force_11(1'b0), .Q(\filter_0/n8189 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5204 ), .force_10(
        \filter_0/n5205 ), .force_11(1'b0), .Q(\filter_0/n8188 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5208 ), .force_10(
        \filter_0/n5209 ), .force_11(1'b0), .Q(\filter_0/n8187 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5212 ), .force_10(
        \filter_0/n5213 ), .force_11(1'b0), .Q(\filter_0/n8186 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5216 ), .force_10(
        \filter_0/n5217 ), .force_11(1'b0), .Q(\filter_0/n8185 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5220 ), .force_10(
        \filter_0/n5221 ), .force_11(1'b0), .Q(\filter_0/n8184 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5224 ), .force_10(
        \filter_0/n5225 ), .force_11(1'b0), .Q(\filter_0/n8183 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5228 ), .force_10(
        \filter_0/n5229 ), .force_11(1'b0), .Q(\filter_0/n8182 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5232 ), .force_10(
        \filter_0/n5233 ), .force_11(1'b0), .Q(\filter_0/n8181 ) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5236 ), .force_10(
        \filter_0/n5237 ), .force_11(1'b0), .Q(\filter_0/n8180 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5240 ), .force_10(\filter_0/n5241 ), 
        .force_11(1'b0), .Q(\filter_0/n8179 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5244 ), .force_10(\filter_0/n5245 ), 
        .force_11(1'b0), .Q(\filter_0/n8178 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5248 ), .force_10(\filter_0/n5249 ), 
        .force_11(1'b0), .Q(\filter_0/n8177 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5252 ), .force_10(\filter_0/n5253 ), 
        .force_11(1'b0), .Q(\filter_0/n8176 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5256 ), .force_10(\filter_0/n5257 ), 
        .force_11(1'b0), .Q(\filter_0/n8175 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5260 ), .force_10(\filter_0/n5261 ), 
        .force_11(1'b0), .Q(\filter_0/n8174 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5264 ), .force_10(\filter_0/n5265 ), 
        .force_11(1'b0), .Q(\filter_0/n8173 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5268 ), .force_10(\filter_0/n5269 ), 
        .force_11(1'b0), .Q(\filter_0/n8172 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5272 ), .force_10(\filter_0/n5273 ), 
        .force_11(1'b0), .Q(\filter_0/n8171 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5276 ), .force_10(\filter_0/n5277 ), 
        .force_11(1'b0), .Q(\filter_0/n8170 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5280 ), .force_10(
        \filter_0/n5281 ), .force_11(1'b0), .Q(\filter_0/n8169 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5284 ), .force_10(
        \filter_0/n5285 ), .force_11(1'b0), .Q(\filter_0/n8168 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5288 ), .force_10(
        \filter_0/n5289 ), .force_11(1'b0), .Q(\filter_0/n8167 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5292 ), .force_10(
        \filter_0/n5293 ), .force_11(1'b0), .Q(\filter_0/n8166 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5296 ), .force_10(
        \filter_0/n5297 ), .force_11(1'b0), .Q(\filter_0/n8165 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5300 ), .force_10(
        \filter_0/n5301 ), .force_11(1'b0), .Q(\filter_0/n8164 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5304 ), .force_10(
        \filter_0/n5305 ), .force_11(1'b0), .Q(\filter_0/n8163 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5308 ), .force_10(
        \filter_0/n5309 ), .force_11(1'b0), .Q(\filter_0/n8162 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5312 ), .force_10(
        \filter_0/n5313 ), .force_11(1'b0), .Q(\filter_0/n8161 ) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5316 ), .force_10(
        \filter_0/n5317 ), .force_11(1'b0), .Q(\filter_0/n8160 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5320 ), .force_10(\filter_0/n5321 ), 
        .force_11(1'b0), .Q(\filter_0/n8159 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5324 ), .force_10(\filter_0/n5325 ), 
        .force_11(1'b0), .Q(\filter_0/n8158 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5328 ), .force_10(\filter_0/n5329 ), 
        .force_11(1'b0), .Q(\filter_0/n8157 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5332 ), .force_10(\filter_0/n5333 ), 
        .force_11(1'b0), .Q(\filter_0/n8156 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5336 ), .force_10(\filter_0/n5337 ), 
        .force_11(1'b0), .Q(\filter_0/n8155 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5340 ), .force_10(\filter_0/n5341 ), 
        .force_11(1'b0), .Q(\filter_0/n8154 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5344 ), .force_10(\filter_0/n5345 ), 
        .force_11(1'b0), .Q(\filter_0/n8153 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5348 ), .force_10(\filter_0/n5349 ), 
        .force_11(1'b0), .Q(\filter_0/n8152 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5352 ), .force_10(\filter_0/n5353 ), 
        .force_11(1'b0), .Q(\filter_0/n8151 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5356 ), .force_10(\filter_0/n5357 ), 
        .force_11(1'b0), .Q(\filter_0/n8150 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5360 ), .force_10(
        \filter_0/n5361 ), .force_11(1'b0), .Q(\filter_0/n8149 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5364 ), .force_10(
        \filter_0/n5365 ), .force_11(1'b0), .Q(\filter_0/n8148 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5368 ), .force_10(
        \filter_0/n5369 ), .force_11(1'b0), .Q(\filter_0/n8147 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5372 ), .force_10(
        \filter_0/n5373 ), .force_11(1'b0), .Q(\filter_0/n8146 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5376 ), .force_10(
        \filter_0/n5377 ), .force_11(1'b0), .Q(\filter_0/n8145 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5380 ), .force_10(
        \filter_0/n5381 ), .force_11(1'b0), .Q(\filter_0/n8144 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5384 ), .force_10(
        \filter_0/n5385 ), .force_11(1'b0), .Q(\filter_0/n8143 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5388 ), .force_10(
        \filter_0/n5389 ), .force_11(1'b0), .Q(\filter_0/n8142 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5392 ), .force_10(
        \filter_0/n5393 ), .force_11(1'b0), .Q(\filter_0/n8141 ) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5396 ), .force_10(
        \filter_0/n5397 ), .force_11(1'b0), .Q(\filter_0/n8140 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5400 ), .force_10(\filter_0/n5401 ), 
        .force_11(1'b0), .Q(\filter_0/n8139 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5404 ), .force_10(\filter_0/n5405 ), 
        .force_11(1'b0), .Q(\filter_0/n8138 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5408 ), .force_10(\filter_0/n5409 ), 
        .force_11(1'b0), .Q(\filter_0/n8137 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5412 ), .force_10(\filter_0/n5413 ), 
        .force_11(1'b0), .Q(\filter_0/n8136 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5416 ), .force_10(\filter_0/n5417 ), 
        .force_11(1'b0), .Q(\filter_0/n8135 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5420 ), .force_10(\filter_0/n5421 ), 
        .force_11(1'b0), .Q(\filter_0/n8134 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5424 ), .force_10(\filter_0/n5425 ), 
        .force_11(1'b0), .Q(\filter_0/n8133 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5428 ), .force_10(\filter_0/n5429 ), 
        .force_11(1'b0), .Q(\filter_0/n8132 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5432 ), .force_10(\filter_0/n5433 ), 
        .force_11(1'b0), .Q(\filter_0/n8131 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5436 ), .force_10(\filter_0/n5437 ), 
        .force_11(1'b0), .Q(\filter_0/n8130 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5440 ), .force_10(
        \filter_0/n5441 ), .force_11(1'b0), .Q(\filter_0/n8129 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5444 ), .force_10(
        \filter_0/n5445 ), .force_11(1'b0), .Q(\filter_0/n8128 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5448 ), .force_10(
        \filter_0/n5449 ), .force_11(1'b0), .Q(\filter_0/n8127 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5452 ), .force_10(
        \filter_0/n5453 ), .force_11(1'b0), .Q(\filter_0/n8126 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5456 ), .force_10(
        \filter_0/n5457 ), .force_11(1'b0), .Q(\filter_0/n8125 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5460 ), .force_10(
        \filter_0/n5461 ), .force_11(1'b0), .Q(\filter_0/n8124 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5464 ), .force_10(
        \filter_0/n5465 ), .force_11(1'b0), .Q(\filter_0/n8123 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5468 ), .force_10(
        \filter_0/n5469 ), .force_11(1'b0), .Q(\filter_0/n8122 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5472 ), .force_10(
        \filter_0/n5473 ), .force_11(1'b0), .Q(\filter_0/n8121 ) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5476 ), .force_10(
        \filter_0/n5477 ), .force_11(1'b0), .Q(\filter_0/n8120 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5480 ), .force_10(\filter_0/n5481 ), 
        .force_11(1'b0), .Q(\filter_0/n8119 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5484 ), .force_10(\filter_0/n5485 ), 
        .force_11(1'b0), .Q(\filter_0/n8118 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5488 ), .force_10(\filter_0/n5489 ), 
        .force_11(1'b0), .Q(\filter_0/n8117 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5492 ), .force_10(\filter_0/n5493 ), 
        .force_11(1'b0), .Q(\filter_0/n8116 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5496 ), .force_10(\filter_0/n5497 ), 
        .force_11(1'b0), .Q(\filter_0/n8115 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5500 ), .force_10(\filter_0/n5501 ), 
        .force_11(1'b0), .Q(\filter_0/n8114 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5504 ), .force_10(\filter_0/n5505 ), 
        .force_11(1'b0), .Q(\filter_0/n8113 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5508 ), .force_10(\filter_0/n5509 ), 
        .force_11(1'b0), .Q(\filter_0/n8112 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5512 ), .force_10(\filter_0/n5513 ), 
        .force_11(1'b0), .Q(\filter_0/n8111 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5516 ), .force_10(\filter_0/n5517 ), 
        .force_11(1'b0), .Q(\filter_0/n8110 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5520 ), .force_10(
        \filter_0/n5521 ), .force_11(1'b0), .Q(\filter_0/n8109 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5524 ), .force_10(
        \filter_0/n5525 ), .force_11(1'b0), .Q(\filter_0/n8108 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5528 ), .force_10(
        \filter_0/n5529 ), .force_11(1'b0), .Q(\filter_0/n8107 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5532 ), .force_10(
        \filter_0/n5533 ), .force_11(1'b0), .Q(\filter_0/n8106 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5536 ), .force_10(
        \filter_0/n5537 ), .force_11(1'b0), .Q(\filter_0/n8105 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5540 ), .force_10(
        \filter_0/n5541 ), .force_11(1'b0), .Q(\filter_0/n8104 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5544 ), .force_10(
        \filter_0/n5545 ), .force_11(1'b0), .Q(\filter_0/n8103 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5548 ), .force_10(
        \filter_0/n5549 ), .force_11(1'b0), .Q(\filter_0/n8102 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5552 ), .force_10(
        \filter_0/n5553 ), .force_11(1'b0), .Q(\filter_0/n8101 ) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5556 ), .force_10(
        \filter_0/n5557 ), .force_11(1'b0), .Q(\filter_0/n8100 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5560 ), .force_10(\filter_0/n5561 ), 
        .force_11(1'b0), .Q(\filter_0/n8099 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5564 ), .force_10(\filter_0/n5565 ), 
        .force_11(1'b0), .Q(\filter_0/n8098 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5568 ), .force_10(\filter_0/n5569 ), 
        .force_11(1'b0), .Q(\filter_0/n8097 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5572 ), .force_10(\filter_0/n5573 ), 
        .force_11(1'b0), .Q(\filter_0/n8096 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5576 ), .force_10(\filter_0/n5577 ), 
        .force_11(1'b0), .Q(\filter_0/n8095 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5580 ), .force_10(\filter_0/n5581 ), 
        .force_11(1'b0), .Q(\filter_0/n8094 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5584 ), .force_10(\filter_0/n5585 ), 
        .force_11(1'b0), .Q(\filter_0/n8093 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5588 ), .force_10(\filter_0/n5589 ), 
        .force_11(1'b0), .Q(\filter_0/n8092 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5592 ), .force_10(\filter_0/n5593 ), 
        .force_11(1'b0), .Q(\filter_0/n8091 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n5596 ), .force_10(\filter_0/n5597 ), 
        .force_11(1'b0), .Q(\filter_0/n8090 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5600 ), .force_10(
        \filter_0/n5601 ), .force_11(1'b0), .Q(\filter_0/n8089 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5604 ), .force_10(
        \filter_0/n5605 ), .force_11(1'b0), .Q(\filter_0/n8088 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5608 ), .force_10(
        \filter_0/n5609 ), .force_11(1'b0), .Q(\filter_0/n8087 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5612 ), .force_10(
        \filter_0/n5613 ), .force_11(1'b0), .Q(\filter_0/n8086 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5616 ), .force_10(
        \filter_0/n5617 ), .force_11(1'b0), .Q(\filter_0/n8085 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5620 ), .force_10(
        \filter_0/n5621 ), .force_11(1'b0), .Q(\filter_0/n8084 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5624 ), .force_10(
        \filter_0/n5625 ), .force_11(1'b0), .Q(\filter_0/n8083 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5628 ), .force_10(
        \filter_0/n5629 ), .force_11(1'b0), .Q(\filter_0/n8082 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5632 ), .force_10(
        \filter_0/n5633 ), .force_11(1'b0), .Q(\filter_0/n8081 ) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5636 ), .force_10(
        \filter_0/n5637 ), .force_11(1'b0), .Q(\filter_0/n8080 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5640 ), .force_10(
        \filter_0/n5641 ), .force_11(1'b0), .Q(\filter_0/n8079 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5644 ), .force_10(
        \filter_0/n5645 ), .force_11(1'b0), .Q(\filter_0/n8078 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5648 ), .force_10(
        \filter_0/n5649 ), .force_11(1'b0), .Q(\filter_0/n8077 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5652 ), .force_10(
        \filter_0/n5653 ), .force_11(1'b0), .Q(\filter_0/n8076 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5656 ), .force_10(
        \filter_0/n5657 ), .force_11(1'b0), .Q(\filter_0/n8075 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5660 ), .force_10(
        \filter_0/n5661 ), .force_11(1'b0), .Q(\filter_0/n8074 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5664 ), .force_10(
        \filter_0/n5665 ), .force_11(1'b0), .Q(\filter_0/n8073 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5668 ), .force_10(
        \filter_0/n5669 ), .force_11(1'b0), .Q(\filter_0/n8072 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5672 ), .force_10(
        \filter_0/n5673 ), .force_11(1'b0), .Q(\filter_0/n8071 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5676 ), .force_10(
        \filter_0/n5677 ), .force_11(1'b0), .Q(\filter_0/n8070 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5680 ), .force_10(
        \filter_0/n5681 ), .force_11(1'b0), .Q(\filter_0/n8069 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5684 ), .force_10(
        \filter_0/n5685 ), .force_11(1'b0), .Q(\filter_0/n8068 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5688 ), .force_10(
        \filter_0/n5689 ), .force_11(1'b0), .Q(\filter_0/n8067 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5692 ), .force_10(
        \filter_0/n5693 ), .force_11(1'b0), .Q(\filter_0/n8066 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5696 ), .force_10(
        \filter_0/n5697 ), .force_11(1'b0), .Q(\filter_0/n8065 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5700 ), .force_10(
        \filter_0/n5701 ), .force_11(1'b0), .Q(\filter_0/n8064 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5704 ), .force_10(
        \filter_0/n5705 ), .force_11(1'b0), .Q(\filter_0/n8063 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5708 ), .force_10(
        \filter_0/n5709 ), .force_11(1'b0), .Q(\filter_0/n8062 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5712 ), .force_10(
        \filter_0/n5713 ), .force_11(1'b0), .Q(\filter_0/n8061 ) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5716 ), .force_10(
        \filter_0/n5717 ), .force_11(1'b0), .Q(\filter_0/n8060 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5720 ), .force_10(
        \filter_0/n5721 ), .force_11(1'b0), .Q(\filter_0/n8059 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5724 ), .force_10(
        \filter_0/n5725 ), .force_11(1'b0), .Q(\filter_0/n8058 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5728 ), .force_10(
        \filter_0/n5729 ), .force_11(1'b0), .Q(\filter_0/n8057 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5732 ), .force_10(
        \filter_0/n5733 ), .force_11(1'b0), .Q(\filter_0/n8056 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5736 ), .force_10(
        \filter_0/n5737 ), .force_11(1'b0), .Q(\filter_0/n8055 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5740 ), .force_10(
        \filter_0/n5741 ), .force_11(1'b0), .Q(\filter_0/n8054 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5744 ), .force_10(
        \filter_0/n5745 ), .force_11(1'b0), .Q(\filter_0/n8053 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5748 ), .force_10(
        \filter_0/n5749 ), .force_11(1'b0), .Q(\filter_0/n8052 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5752 ), .force_10(
        \filter_0/n5753 ), .force_11(1'b0), .Q(\filter_0/n8051 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5756 ), .force_10(
        \filter_0/n5757 ), .force_11(1'b0), .Q(\filter_0/n8050 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5760 ), .force_10(
        \filter_0/n5761 ), .force_11(1'b0), .Q(\filter_0/n8049 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5764 ), .force_10(
        \filter_0/n5765 ), .force_11(1'b0), .Q(\filter_0/n8048 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5768 ), .force_10(
        \filter_0/n5769 ), .force_11(1'b0), .Q(\filter_0/n8047 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5772 ), .force_10(
        \filter_0/n5773 ), .force_11(1'b0), .Q(\filter_0/n8046 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5776 ), .force_10(
        \filter_0/n5777 ), .force_11(1'b0), .Q(\filter_0/n8045 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5780 ), .force_10(
        \filter_0/n5781 ), .force_11(1'b0), .Q(\filter_0/n8044 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5784 ), .force_10(
        \filter_0/n5785 ), .force_11(1'b0), .Q(\filter_0/n8043 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5788 ), .force_10(
        \filter_0/n5789 ), .force_11(1'b0), .Q(\filter_0/n8042 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5792 ), .force_10(
        \filter_0/n5793 ), .force_11(1'b0), .Q(\filter_0/n8041 ) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5796 ), .force_10(
        \filter_0/n5797 ), .force_11(1'b0), .Q(\filter_0/n8040 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5800 ), .force_10(
        \filter_0/n5801 ), .force_11(1'b0), .Q(\filter_0/n8039 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5804 ), .force_10(
        \filter_0/n5805 ), .force_11(1'b0), .Q(\filter_0/n8038 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5808 ), .force_10(
        \filter_0/n5809 ), .force_11(1'b0), .Q(\filter_0/n8037 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5812 ), .force_10(
        \filter_0/n5813 ), .force_11(1'b0), .Q(\filter_0/n8036 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5816 ), .force_10(
        \filter_0/n5817 ), .force_11(1'b0), .Q(\filter_0/n8035 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5820 ), .force_10(
        \filter_0/n5821 ), .force_11(1'b0), .Q(\filter_0/n8034 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5824 ), .force_10(
        \filter_0/n5825 ), .force_11(1'b0), .Q(\filter_0/n8033 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5828 ), .force_10(
        \filter_0/n5829 ), .force_11(1'b0), .Q(\filter_0/n8032 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5832 ), .force_10(
        \filter_0/n5833 ), .force_11(1'b0), .Q(\filter_0/n8031 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5836 ), .force_10(
        \filter_0/n5837 ), .force_11(1'b0), .Q(\filter_0/n8030 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5840 ), .force_10(
        \filter_0/n5841 ), .force_11(1'b0), .Q(\filter_0/n8029 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5844 ), .force_10(
        \filter_0/n5845 ), .force_11(1'b0), .Q(\filter_0/n8028 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5848 ), .force_10(
        \filter_0/n5849 ), .force_11(1'b0), .Q(\filter_0/n8027 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5852 ), .force_10(
        \filter_0/n5853 ), .force_11(1'b0), .Q(\filter_0/n8026 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5856 ), .force_10(
        \filter_0/n5857 ), .force_11(1'b0), .Q(\filter_0/n8025 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5860 ), .force_10(
        \filter_0/n5861 ), .force_11(1'b0), .Q(\filter_0/n8024 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5864 ), .force_10(
        \filter_0/n5865 ), .force_11(1'b0), .Q(\filter_0/n8023 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5868 ), .force_10(
        \filter_0/n5869 ), .force_11(1'b0), .Q(\filter_0/n8022 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5872 ), .force_10(
        \filter_0/n5873 ), .force_11(1'b0), .Q(\filter_0/n8021 ) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5876 ), .force_10(
        \filter_0/n5877 ), .force_11(1'b0), .Q(\filter_0/n8020 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5880 ), .force_10(
        \filter_0/n5881 ), .force_11(1'b0), .Q(\filter_0/n8019 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5884 ), .force_10(
        \filter_0/n5885 ), .force_11(1'b0), .Q(\filter_0/n8018 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5888 ), .force_10(
        \filter_0/n5889 ), .force_11(1'b0), .Q(\filter_0/n8017 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5892 ), .force_10(
        \filter_0/n5893 ), .force_11(1'b0), .Q(\filter_0/n8016 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5896 ), .force_10(
        \filter_0/n5897 ), .force_11(1'b0), .Q(\filter_0/n8015 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5900 ), .force_10(
        \filter_0/n5901 ), .force_11(1'b0), .Q(\filter_0/n8014 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5904 ), .force_10(
        \filter_0/n5905 ), .force_11(1'b0), .Q(\filter_0/n8013 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5908 ), .force_10(
        \filter_0/n5909 ), .force_11(1'b0), .Q(\filter_0/n8012 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5912 ), .force_10(
        \filter_0/n5913 ), .force_11(1'b0), .Q(\filter_0/n8011 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5916 ), .force_10(
        \filter_0/n5917 ), .force_11(1'b0), .Q(\filter_0/n8010 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5920 ), .force_10(
        \filter_0/n5921 ), .force_11(1'b0), .Q(\filter_0/n8009 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5924 ), .force_10(
        \filter_0/n5925 ), .force_11(1'b0), .Q(\filter_0/n8008 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5928 ), .force_10(
        \filter_0/n5929 ), .force_11(1'b0), .Q(\filter_0/n8007 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5932 ), .force_10(
        \filter_0/n5933 ), .force_11(1'b0), .Q(\filter_0/n8006 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5936 ), .force_10(
        \filter_0/n5937 ), .force_11(1'b0), .Q(\filter_0/n8005 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5940 ), .force_10(
        \filter_0/n5941 ), .force_11(1'b0), .Q(\filter_0/n8004 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5944 ), .force_10(
        \filter_0/n5945 ), .force_11(1'b0), .Q(\filter_0/n8003 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5948 ), .force_10(
        \filter_0/n5949 ), .force_11(1'b0), .Q(\filter_0/n8002 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5952 ), .force_10(
        \filter_0/n5953 ), .force_11(1'b0), .Q(\filter_0/n8001 ) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5956 ), .force_10(
        \filter_0/n5957 ), .force_11(1'b0), .Q(\filter_0/n8000 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5960 ), .force_10(
        \filter_0/n5961 ), .force_11(1'b0), .Q(\filter_0/n7999 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5964 ), .force_10(
        \filter_0/n5965 ), .force_11(1'b0), .Q(\filter_0/n7998 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5968 ), .force_10(
        \filter_0/n5969 ), .force_11(1'b0), .Q(\filter_0/n7997 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5972 ), .force_10(
        \filter_0/n5973 ), .force_11(1'b0), .Q(\filter_0/n7996 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5976 ), .force_10(
        \filter_0/n5977 ), .force_11(1'b0), .Q(\filter_0/n7995 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5980 ), .force_10(
        \filter_0/n5981 ), .force_11(1'b0), .Q(\filter_0/n7994 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5984 ), .force_10(
        \filter_0/n5985 ), .force_11(1'b0), .Q(\filter_0/n7993 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5988 ), .force_10(
        \filter_0/n5989 ), .force_11(1'b0), .Q(\filter_0/n7992 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5992 ), .force_10(
        \filter_0/n5993 ), .force_11(1'b0), .Q(\filter_0/n7991 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n5996 ), .force_10(
        \filter_0/n5997 ), .force_11(1'b0), .Q(\filter_0/n7990 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6000 ), .force_10(
        \filter_0/n6001 ), .force_11(1'b0), .Q(\filter_0/n7989 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6004 ), .force_10(
        \filter_0/n6005 ), .force_11(1'b0), .Q(\filter_0/n7988 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6008 ), .force_10(
        \filter_0/n6009 ), .force_11(1'b0), .Q(\filter_0/n7987 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6012 ), .force_10(
        \filter_0/n6013 ), .force_11(1'b0), .Q(\filter_0/n7986 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6016 ), .force_10(
        \filter_0/n6017 ), .force_11(1'b0), .Q(\filter_0/n7985 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6020 ), .force_10(
        \filter_0/n6021 ), .force_11(1'b0), .Q(\filter_0/n7984 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6024 ), .force_10(
        \filter_0/n6025 ), .force_11(1'b0), .Q(\filter_0/n7983 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6028 ), .force_10(
        \filter_0/n6029 ), .force_11(1'b0), .Q(\filter_0/n7982 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6032 ), .force_10(
        \filter_0/n6033 ), .force_11(1'b0), .Q(\filter_0/n7981 ) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6036 ), .force_10(
        \filter_0/n6037 ), .force_11(1'b0), .Q(\filter_0/n7980 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6040 ), .force_10(
        \filter_0/n6041 ), .force_11(1'b0), .Q(\filter_0/n7979 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6044 ), .force_10(
        \filter_0/n6045 ), .force_11(1'b0), .Q(\filter_0/n7978 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6048 ), .force_10(
        \filter_0/n6049 ), .force_11(1'b0), .Q(\filter_0/n7977 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6052 ), .force_10(
        \filter_0/n6053 ), .force_11(1'b0), .Q(\filter_0/n7976 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6056 ), .force_10(
        \filter_0/n6057 ), .force_11(1'b0), .Q(\filter_0/n7975 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6060 ), .force_10(
        \filter_0/n6061 ), .force_11(1'b0), .Q(\filter_0/n7974 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6064 ), .force_10(
        \filter_0/n6065 ), .force_11(1'b0), .Q(\filter_0/n7973 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6068 ), .force_10(
        \filter_0/n6069 ), .force_11(1'b0), .Q(\filter_0/n7972 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6072 ), .force_10(
        \filter_0/n6073 ), .force_11(1'b0), .Q(\filter_0/n7971 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6076 ), .force_10(
        \filter_0/n6077 ), .force_11(1'b0), .Q(\filter_0/n7970 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6080 ), .force_10(
        \filter_0/n6081 ), .force_11(1'b0), .Q(\filter_0/n7969 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6084 ), .force_10(
        \filter_0/n6085 ), .force_11(1'b0), .Q(\filter_0/n7968 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6088 ), .force_10(
        \filter_0/n6089 ), .force_11(1'b0), .Q(\filter_0/n7967 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6092 ), .force_10(
        \filter_0/n6093 ), .force_11(1'b0), .Q(\filter_0/n7966 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6096 ), .force_10(
        \filter_0/n6097 ), .force_11(1'b0), .Q(\filter_0/n7965 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6100 ), .force_10(
        \filter_0/n6101 ), .force_11(1'b0), .Q(\filter_0/n7964 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6104 ), .force_10(
        \filter_0/n6105 ), .force_11(1'b0), .Q(\filter_0/n7963 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6108 ), .force_10(
        \filter_0/n6109 ), .force_11(1'b0), .Q(\filter_0/n7962 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6112 ), .force_10(
        \filter_0/n6113 ), .force_11(1'b0), .Q(\filter_0/n7961 ) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6116 ), .force_10(
        \filter_0/n6117 ), .force_11(1'b0), .Q(\filter_0/n7960 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6120 ), .force_10(\filter_0/n6121 ), 
        .force_11(1'b0), .Q(\filter_0/n7959 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6124 ), .force_10(\filter_0/n6125 ), 
        .force_11(1'b0), .Q(\filter_0/n7958 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6128 ), .force_10(\filter_0/n6129 ), 
        .force_11(1'b0), .Q(\filter_0/n7957 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6132 ), .force_10(\filter_0/n6133 ), 
        .force_11(1'b0), .Q(\filter_0/n7956 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6136 ), .force_10(\filter_0/n6137 ), 
        .force_11(1'b0), .Q(\filter_0/n7955 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6140 ), .force_10(\filter_0/n6141 ), 
        .force_11(1'b0), .Q(\filter_0/n7954 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6144 ), .force_10(\filter_0/n6145 ), 
        .force_11(1'b0), .Q(\filter_0/n7953 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6148 ), .force_10(\filter_0/n6149 ), 
        .force_11(1'b0), .Q(\filter_0/n7952 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6152 ), .force_10(\filter_0/n6153 ), 
        .force_11(1'b0), .Q(\filter_0/n7951 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6156 ), .force_10(\filter_0/n6157 ), 
        .force_11(1'b0), .Q(\filter_0/n7950 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6160 ), .force_10(
        \filter_0/n6161 ), .force_11(1'b0), .Q(\filter_0/n7949 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6164 ), .force_10(
        \filter_0/n6165 ), .force_11(1'b0), .Q(\filter_0/n7948 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6168 ), .force_10(
        \filter_0/n6169 ), .force_11(1'b0), .Q(\filter_0/n7947 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6172 ), .force_10(
        \filter_0/n6173 ), .force_11(1'b0), .Q(\filter_0/n7946 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6176 ), .force_10(
        \filter_0/n6177 ), .force_11(1'b0), .Q(\filter_0/n7945 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6180 ), .force_10(
        \filter_0/n6181 ), .force_11(1'b0), .Q(\filter_0/n7944 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6184 ), .force_10(
        \filter_0/n6185 ), .force_11(1'b0), .Q(\filter_0/n7943 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6188 ), .force_10(
        \filter_0/n6189 ), .force_11(1'b0), .Q(\filter_0/n7942 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6192 ), .force_10(
        \filter_0/n6193 ), .force_11(1'b0), .Q(\filter_0/n7941 ) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6196 ), .force_10(
        \filter_0/n6197 ), .force_11(1'b0), .Q(\filter_0/n7940 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6200 ), .force_10(\filter_0/n6201 ), 
        .force_11(1'b0), .Q(\filter_0/n7939 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6204 ), .force_10(\filter_0/n6205 ), 
        .force_11(1'b0), .Q(\filter_0/n7938 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6208 ), .force_10(\filter_0/n6209 ), 
        .force_11(1'b0), .Q(\filter_0/n7937 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6212 ), .force_10(\filter_0/n6213 ), 
        .force_11(1'b0), .Q(\filter_0/n7936 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6216 ), .force_10(\filter_0/n6217 ), 
        .force_11(1'b0), .Q(\filter_0/n7935 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6220 ), .force_10(\filter_0/n6221 ), 
        .force_11(1'b0), .Q(\filter_0/n7934 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6224 ), .force_10(\filter_0/n6225 ), 
        .force_11(1'b0), .Q(\filter_0/n7933 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6228 ), .force_10(\filter_0/n6229 ), 
        .force_11(1'b0), .Q(\filter_0/n7932 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6232 ), .force_10(\filter_0/n6233 ), 
        .force_11(1'b0), .Q(\filter_0/n7931 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6236 ), .force_10(\filter_0/n6237 ), 
        .force_11(1'b0), .Q(\filter_0/n7930 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6240 ), .force_10(
        \filter_0/n6241 ), .force_11(1'b0), .Q(\filter_0/n7929 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6244 ), .force_10(
        \filter_0/n6245 ), .force_11(1'b0), .Q(\filter_0/n7928 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6248 ), .force_10(
        \filter_0/n6249 ), .force_11(1'b0), .Q(\filter_0/n7927 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6252 ), .force_10(
        \filter_0/n6253 ), .force_11(1'b0), .Q(\filter_0/n7926 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6256 ), .force_10(
        \filter_0/n6257 ), .force_11(1'b0), .Q(\filter_0/n7925 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6260 ), .force_10(
        \filter_0/n6261 ), .force_11(1'b0), .Q(\filter_0/n7924 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6264 ), .force_10(
        \filter_0/n6265 ), .force_11(1'b0), .Q(\filter_0/n7923 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6268 ), .force_10(
        \filter_0/n6269 ), .force_11(1'b0), .Q(\filter_0/n7922 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6272 ), .force_10(
        \filter_0/n6273 ), .force_11(1'b0), .Q(\filter_0/n7921 ) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6276 ), .force_10(
        \filter_0/n6277 ), .force_11(1'b0), .Q(\filter_0/n7920 ) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6280 ), 
        .force_10(\filter_0/n6281 ), .force_11(1'b0), .Q(\filter_0/n7919 ) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6284 ), 
        .force_10(\filter_0/n6285 ), .force_11(1'b0), .Q(\filter_0/n7918 ) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6288 ), 
        .force_10(\filter_0/n6289 ), .force_11(1'b0), .Q(\filter_0/n7917 ) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6292 ), 
        .force_10(\filter_0/n6293 ), .force_11(1'b0), .Q(\filter_0/n7916 ) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6296 ), 
        .force_10(\filter_0/n6297 ), .force_11(1'b0), .Q(\filter_0/n7915 ) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6300 ), 
        .force_10(\filter_0/n6301 ), .force_11(1'b0), .Q(\filter_0/n7914 ) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6304 ), 
        .force_10(\filter_0/n6305 ), .force_11(1'b0), .Q(\filter_0/n7913 ) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6308 ), 
        .force_10(\filter_0/n6309 ), .force_11(1'b0), .Q(\filter_0/n7912 ) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6312 ), 
        .force_10(\filter_0/n6313 ), .force_11(1'b0), .Q(\filter_0/n7911 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6316 ), .force_10(\filter_0/n6317 ), 
        .force_11(1'b0), .Q(\filter_0/n7910 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6320 ), .force_10(\filter_0/n6321 ), 
        .force_11(1'b0), .Q(\filter_0/n7909 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6324 ), .force_10(\filter_0/n6325 ), 
        .force_11(1'b0), .Q(\filter_0/n7908 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6328 ), .force_10(\filter_0/n6329 ), 
        .force_11(1'b0), .Q(\filter_0/n7907 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6332 ), .force_10(\filter_0/n6333 ), 
        .force_11(1'b0), .Q(\filter_0/n7906 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6336 ), .force_10(\filter_0/n6337 ), 
        .force_11(1'b0), .Q(\filter_0/n7905 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6340 ), .force_10(\filter_0/n6341 ), 
        .force_11(1'b0), .Q(\filter_0/n7904 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6344 ), .force_10(\filter_0/n6345 ), 
        .force_11(1'b0), .Q(\filter_0/n7903 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6348 ), .force_10(\filter_0/n6349 ), 
        .force_11(1'b0), .Q(\filter_0/n7902 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6352 ), .force_10(\filter_0/n6353 ), 
        .force_11(1'b0), .Q(\filter_0/n7901 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6356 ), .force_10(
        \filter_0/n6357 ), .force_11(1'b0), .Q(\filter_0/n7900 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6360 ), .force_10(
        \filter_0/n6361 ), .force_11(1'b0), .Q(\filter_0/n7899 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6364 ), .force_10(
        \filter_0/n6365 ), .force_11(1'b0), .Q(\filter_0/n7898 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6368 ), .force_10(
        \filter_0/n6369 ), .force_11(1'b0), .Q(\filter_0/n7897 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6372 ), .force_10(
        \filter_0/n6373 ), .force_11(1'b0), .Q(\filter_0/n7896 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6376 ), .force_10(
        \filter_0/n6377 ), .force_11(1'b0), .Q(\filter_0/n7895 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6380 ), .force_10(
        \filter_0/n6381 ), .force_11(1'b0), .Q(\filter_0/n7894 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6384 ), .force_10(
        \filter_0/n6385 ), .force_11(1'b0), .Q(\filter_0/n7893 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6388 ), .force_10(
        \filter_0/n6389 ), .force_11(1'b0), .Q(\filter_0/n7892 ) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6392 ), .force_10(
        \filter_0/n6393 ), .force_11(1'b0), .Q(\filter_0/n7891 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6396 ), .force_10(\filter_0/n6397 ), 
        .force_11(1'b0), .Q(\filter_0/n7890 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6400 ), .force_10(\filter_0/n6401 ), 
        .force_11(1'b0), .Q(\filter_0/n7889 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6404 ), .force_10(\filter_0/n6405 ), 
        .force_11(1'b0), .Q(\filter_0/n7888 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6408 ), .force_10(\filter_0/n6409 ), 
        .force_11(1'b0), .Q(\filter_0/n7887 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6412 ), .force_10(\filter_0/n6413 ), 
        .force_11(1'b0), .Q(\filter_0/n7886 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6416 ), .force_10(\filter_0/n6417 ), 
        .force_11(1'b0), .Q(\filter_0/n7885 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6420 ), .force_10(\filter_0/n6421 ), 
        .force_11(1'b0), .Q(\filter_0/n7884 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6424 ), .force_10(\filter_0/n6425 ), 
        .force_11(1'b0), .Q(\filter_0/n7883 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6428 ), .force_10(\filter_0/n6429 ), 
        .force_11(1'b0), .Q(\filter_0/n7882 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6432 ), .force_10(\filter_0/n6433 ), 
        .force_11(1'b0), .Q(\filter_0/n7881 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6436 ), .force_10(
        \filter_0/n6437 ), .force_11(1'b0), .Q(\filter_0/n7880 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6440 ), .force_10(
        \filter_0/n6441 ), .force_11(1'b0), .Q(\filter_0/n7879 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6444 ), .force_10(
        \filter_0/n6445 ), .force_11(1'b0), .Q(\filter_0/n7878 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6448 ), .force_10(
        \filter_0/n6449 ), .force_11(1'b0), .Q(\filter_0/n7877 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6452 ), .force_10(
        \filter_0/n6453 ), .force_11(1'b0), .Q(\filter_0/n7876 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6456 ), .force_10(
        \filter_0/n6457 ), .force_11(1'b0), .Q(\filter_0/n7875 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6460 ), .force_10(
        \filter_0/n6461 ), .force_11(1'b0), .Q(\filter_0/n7874 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6464 ), .force_10(
        \filter_0/n6465 ), .force_11(1'b0), .Q(\filter_0/n7873 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6468 ), .force_10(
        \filter_0/n6469 ), .force_11(1'b0), .Q(\filter_0/n7872 ) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6472 ), .force_10(
        \filter_0/n6473 ), .force_11(1'b0), .Q(\filter_0/n7871 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6476 ), .force_10(\filter_0/n6477 ), 
        .force_11(1'b0), .Q(\filter_0/n7870 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6480 ), .force_10(\filter_0/n6481 ), 
        .force_11(1'b0), .Q(\filter_0/n7869 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6484 ), .force_10(\filter_0/n6485 ), 
        .force_11(1'b0), .Q(\filter_0/n7868 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6488 ), .force_10(\filter_0/n6489 ), 
        .force_11(1'b0), .Q(\filter_0/n7867 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6492 ), .force_10(\filter_0/n6493 ), 
        .force_11(1'b0), .Q(\filter_0/n7866 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6496 ), .force_10(\filter_0/n6497 ), 
        .force_11(1'b0), .Q(\filter_0/n7865 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6500 ), .force_10(\filter_0/n6501 ), 
        .force_11(1'b0), .Q(\filter_0/n7864 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6504 ), .force_10(\filter_0/n6505 ), 
        .force_11(1'b0), .Q(\filter_0/n7863 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6508 ), .force_10(\filter_0/n6509 ), 
        .force_11(1'b0), .Q(\filter_0/n7862 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6512 ), .force_10(\filter_0/n6513 ), 
        .force_11(1'b0), .Q(\filter_0/n7861 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6516 ), .force_10(
        \filter_0/n6517 ), .force_11(1'b0), .Q(\filter_0/n7860 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6520 ), .force_10(
        \filter_0/n6521 ), .force_11(1'b0), .Q(\filter_0/n7859 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6524 ), .force_10(
        \filter_0/n6525 ), .force_11(1'b0), .Q(\filter_0/n7858 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6528 ), .force_10(
        \filter_0/n6529 ), .force_11(1'b0), .Q(\filter_0/n7857 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6532 ), .force_10(
        \filter_0/n6533 ), .force_11(1'b0), .Q(\filter_0/n7856 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6536 ), .force_10(
        \filter_0/n6537 ), .force_11(1'b0), .Q(\filter_0/n7855 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6540 ), .force_10(
        \filter_0/n6541 ), .force_11(1'b0), .Q(\filter_0/n7854 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6544 ), .force_10(
        \filter_0/n6545 ), .force_11(1'b0), .Q(\filter_0/n7853 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6548 ), .force_10(
        \filter_0/n6549 ), .force_11(1'b0), .Q(\filter_0/n7852 ) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6552 ), .force_10(
        \filter_0/n6553 ), .force_11(1'b0), .Q(\filter_0/n7851 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6556 ), .force_10(\filter_0/n6557 ), 
        .force_11(1'b0), .Q(\filter_0/n7850 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6560 ), .force_10(\filter_0/n6561 ), 
        .force_11(1'b0), .Q(\filter_0/n7849 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6564 ), .force_10(\filter_0/n6565 ), 
        .force_11(1'b0), .Q(\filter_0/n7848 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6568 ), .force_10(\filter_0/n6569 ), 
        .force_11(1'b0), .Q(\filter_0/n7847 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6572 ), .force_10(\filter_0/n6573 ), 
        .force_11(1'b0), .Q(\filter_0/n7846 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6576 ), .force_10(\filter_0/n6577 ), 
        .force_11(1'b0), .Q(\filter_0/n7845 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6580 ), .force_10(\filter_0/n6581 ), 
        .force_11(1'b0), .Q(\filter_0/n7844 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6584 ), .force_10(\filter_0/n6585 ), 
        .force_11(1'b0), .Q(\filter_0/n7843 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6588 ), .force_10(\filter_0/n6589 ), 
        .force_11(1'b0), .Q(\filter_0/n7842 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6592 ), .force_10(\filter_0/n6593 ), 
        .force_11(1'b0), .Q(\filter_0/n7841 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6596 ), .force_10(
        \filter_0/n6597 ), .force_11(1'b0), .Q(\filter_0/n7840 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6600 ), .force_10(
        \filter_0/n6601 ), .force_11(1'b0), .Q(\filter_0/n7839 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6604 ), .force_10(
        \filter_0/n6605 ), .force_11(1'b0), .Q(\filter_0/n7838 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6608 ), .force_10(
        \filter_0/n6609 ), .force_11(1'b0), .Q(\filter_0/n7837 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6612 ), .force_10(
        \filter_0/n6613 ), .force_11(1'b0), .Q(\filter_0/n7836 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6616 ), .force_10(
        \filter_0/n6617 ), .force_11(1'b0), .Q(\filter_0/n7835 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6620 ), .force_10(
        \filter_0/n6621 ), .force_11(1'b0), .Q(\filter_0/n7834 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6624 ), .force_10(
        \filter_0/n6625 ), .force_11(1'b0), .Q(\filter_0/n7833 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6628 ), .force_10(
        \filter_0/n6629 ), .force_11(1'b0), .Q(\filter_0/n7832 ) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6632 ), .force_10(
        \filter_0/n6633 ), .force_11(1'b0), .Q(\filter_0/n7831 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6636 ), .force_10(\filter_0/n6637 ), 
        .force_11(1'b0), .Q(\filter_0/n7830 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6640 ), .force_10(\filter_0/n6641 ), 
        .force_11(1'b0), .Q(\filter_0/n7829 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6644 ), .force_10(\filter_0/n6645 ), 
        .force_11(1'b0), .Q(\filter_0/n7828 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6648 ), .force_10(\filter_0/n6649 ), 
        .force_11(1'b0), .Q(\filter_0/n7827 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6652 ), .force_10(\filter_0/n6653 ), 
        .force_11(1'b0), .Q(\filter_0/n7826 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6656 ), .force_10(\filter_0/n6657 ), 
        .force_11(1'b0), .Q(\filter_0/n7825 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6660 ), .force_10(\filter_0/n6661 ), 
        .force_11(1'b0), .Q(\filter_0/n7824 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6664 ), .force_10(\filter_0/n6665 ), 
        .force_11(1'b0), .Q(\filter_0/n7823 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6668 ), .force_10(\filter_0/n6669 ), 
        .force_11(1'b0), .Q(\filter_0/n7822 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6672 ), .force_10(\filter_0/n6673 ), 
        .force_11(1'b0), .Q(\filter_0/n7821 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6676 ), .force_10(
        \filter_0/n6677 ), .force_11(1'b0), .Q(\filter_0/n7820 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6680 ), .force_10(
        \filter_0/n6681 ), .force_11(1'b0), .Q(\filter_0/n7819 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6684 ), .force_10(
        \filter_0/n6685 ), .force_11(1'b0), .Q(\filter_0/n7818 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6688 ), .force_10(
        \filter_0/n6689 ), .force_11(1'b0), .Q(\filter_0/n7817 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6692 ), .force_10(
        \filter_0/n6693 ), .force_11(1'b0), .Q(\filter_0/n7816 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6696 ), .force_10(
        \filter_0/n6697 ), .force_11(1'b0), .Q(\filter_0/n7815 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6700 ), .force_10(
        \filter_0/n6701 ), .force_11(1'b0), .Q(\filter_0/n7814 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6704 ), .force_10(
        \filter_0/n6705 ), .force_11(1'b0), .Q(\filter_0/n7813 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6708 ), .force_10(
        \filter_0/n6709 ), .force_11(1'b0), .Q(\filter_0/n7812 ) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6712 ), .force_10(
        \filter_0/n6713 ), .force_11(1'b0), .Q(\filter_0/n7811 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6716 ), .force_10(\filter_0/n6717 ), 
        .force_11(1'b0), .Q(\filter_0/n7810 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6720 ), .force_10(\filter_0/n6721 ), 
        .force_11(1'b0), .Q(\filter_0/n7809 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6724 ), .force_10(\filter_0/n6725 ), 
        .force_11(1'b0), .Q(\filter_0/n7808 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6728 ), .force_10(\filter_0/n6729 ), 
        .force_11(1'b0), .Q(\filter_0/n7807 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6732 ), .force_10(\filter_0/n6733 ), 
        .force_11(1'b0), .Q(\filter_0/n7806 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6736 ), .force_10(\filter_0/n6737 ), 
        .force_11(1'b0), .Q(\filter_0/n7805 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6740 ), .force_10(\filter_0/n6741 ), 
        .force_11(1'b0), .Q(\filter_0/n7804 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6744 ), .force_10(\filter_0/n6745 ), 
        .force_11(1'b0), .Q(\filter_0/n7803 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6748 ), .force_10(\filter_0/n6749 ), 
        .force_11(1'b0), .Q(\filter_0/n7802 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6752 ), .force_10(\filter_0/n6753 ), 
        .force_11(1'b0), .Q(\filter_0/n7801 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6756 ), .force_10(
        \filter_0/n6757 ), .force_11(1'b0), .Q(\filter_0/n7800 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6760 ), .force_10(
        \filter_0/n6761 ), .force_11(1'b0), .Q(\filter_0/n7799 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6764 ), .force_10(
        \filter_0/n6765 ), .force_11(1'b0), .Q(\filter_0/n7798 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6768 ), .force_10(
        \filter_0/n6769 ), .force_11(1'b0), .Q(\filter_0/n7797 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6772 ), .force_10(
        \filter_0/n6773 ), .force_11(1'b0), .Q(\filter_0/n7796 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6776 ), .force_10(
        \filter_0/n6777 ), .force_11(1'b0), .Q(\filter_0/n7795 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6780 ), .force_10(
        \filter_0/n6781 ), .force_11(1'b0), .Q(\filter_0/n7794 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6784 ), .force_10(
        \filter_0/n6785 ), .force_11(1'b0), .Q(\filter_0/n7793 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6788 ), .force_10(
        \filter_0/n6789 ), .force_11(1'b0), .Q(\filter_0/n7792 ) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6792 ), .force_10(
        \filter_0/n6793 ), .force_11(1'b0), .Q(\filter_0/n7791 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6796 ), .force_10(\filter_0/n6797 ), 
        .force_11(1'b0), .Q(\filter_0/n7790 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6800 ), .force_10(\filter_0/n6801 ), 
        .force_11(1'b0), .Q(\filter_0/n7789 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6804 ), .force_10(\filter_0/n6805 ), 
        .force_11(1'b0), .Q(\filter_0/n7788 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6808 ), .force_10(\filter_0/n6809 ), 
        .force_11(1'b0), .Q(\filter_0/n7787 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6812 ), .force_10(\filter_0/n6813 ), 
        .force_11(1'b0), .Q(\filter_0/n7786 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6816 ), .force_10(\filter_0/n6817 ), 
        .force_11(1'b0), .Q(\filter_0/n7785 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6820 ), .force_10(\filter_0/n6821 ), 
        .force_11(1'b0), .Q(\filter_0/n7784 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6824 ), .force_10(\filter_0/n6825 ), 
        .force_11(1'b0), .Q(\filter_0/n7783 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6828 ), .force_10(\filter_0/n6829 ), 
        .force_11(1'b0), .Q(\filter_0/n7782 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6832 ), .force_10(\filter_0/n6833 ), 
        .force_11(1'b0), .Q(\filter_0/n7781 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6836 ), .force_10(
        \filter_0/n6837 ), .force_11(1'b0), .Q(\filter_0/n7780 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6840 ), .force_10(
        \filter_0/n6841 ), .force_11(1'b0), .Q(\filter_0/n7779 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6844 ), .force_10(
        \filter_0/n6845 ), .force_11(1'b0), .Q(\filter_0/n7778 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6848 ), .force_10(
        \filter_0/n6849 ), .force_11(1'b0), .Q(\filter_0/n7777 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6852 ), .force_10(
        \filter_0/n6853 ), .force_11(1'b0), .Q(\filter_0/n7776 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6856 ), .force_10(
        \filter_0/n6857 ), .force_11(1'b0), .Q(\filter_0/n7775 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6860 ), .force_10(
        \filter_0/n6861 ), .force_11(1'b0), .Q(\filter_0/n7774 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6864 ), .force_10(
        \filter_0/n6865 ), .force_11(1'b0), .Q(\filter_0/n7773 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6868 ), .force_10(
        \filter_0/n6869 ), .force_11(1'b0), .Q(\filter_0/n7772 ) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6872 ), .force_10(
        \filter_0/n6873 ), .force_11(1'b0), .Q(\filter_0/n7771 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6876 ), .force_10(\filter_0/n6877 ), 
        .force_11(1'b0), .Q(\filter_0/n7770 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6880 ), .force_10(\filter_0/n6881 ), 
        .force_11(1'b0), .Q(\filter_0/n7769 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6884 ), .force_10(\filter_0/n6885 ), 
        .force_11(1'b0), .Q(\filter_0/n7768 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6888 ), .force_10(\filter_0/n6889 ), 
        .force_11(1'b0), .Q(\filter_0/n7767 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6892 ), .force_10(\filter_0/n6893 ), 
        .force_11(1'b0), .Q(\filter_0/n7766 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6896 ), .force_10(\filter_0/n6897 ), 
        .force_11(1'b0), .Q(\filter_0/n7765 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6900 ), .force_10(\filter_0/n6901 ), 
        .force_11(1'b0), .Q(\filter_0/n7764 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6904 ), .force_10(\filter_0/n6905 ), 
        .force_11(1'b0), .Q(\filter_0/n7763 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6908 ), .force_10(\filter_0/n6909 ), 
        .force_11(1'b0), .Q(\filter_0/n7762 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n6912 ), .force_10(\filter_0/n6913 ), 
        .force_11(1'b0), .Q(\filter_0/n7761 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6916 ), .force_10(
        \filter_0/n6917 ), .force_11(1'b0), .Q(\filter_0/n7760 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6920 ), .force_10(
        \filter_0/n6921 ), .force_11(1'b0), .Q(\filter_0/n7759 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6924 ), .force_10(
        \filter_0/n6925 ), .force_11(1'b0), .Q(\filter_0/n7758 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6928 ), .force_10(
        \filter_0/n6929 ), .force_11(1'b0), .Q(\filter_0/n7757 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6932 ), .force_10(
        \filter_0/n6933 ), .force_11(1'b0), .Q(\filter_0/n7756 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6936 ), .force_10(
        \filter_0/n6937 ), .force_11(1'b0), .Q(\filter_0/n7755 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6940 ), .force_10(
        \filter_0/n6941 ), .force_11(1'b0), .Q(\filter_0/n7754 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6944 ), .force_10(
        \filter_0/n6945 ), .force_11(1'b0), .Q(\filter_0/n7753 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6948 ), .force_10(
        \filter_0/n6949 ), .force_11(1'b0), .Q(\filter_0/n7752 ) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6952 ), .force_10(
        \filter_0/n6953 ), .force_11(1'b0), .Q(\filter_0/n7751 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6956 ), .force_10(
        \filter_0/n6957 ), .force_11(1'b0), .Q(\filter_0/n7750 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6960 ), .force_10(
        \filter_0/n6961 ), .force_11(1'b0), .Q(\filter_0/n7749 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6964 ), .force_10(
        \filter_0/n6965 ), .force_11(1'b0), .Q(\filter_0/n7748 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6968 ), .force_10(
        \filter_0/n6969 ), .force_11(1'b0), .Q(\filter_0/n7747 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6972 ), .force_10(
        \filter_0/n6973 ), .force_11(1'b0), .Q(\filter_0/n7746 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6976 ), .force_10(
        \filter_0/n6977 ), .force_11(1'b0), .Q(\filter_0/n7745 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6980 ), .force_10(
        \filter_0/n6981 ), .force_11(1'b0), .Q(\filter_0/n7744 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6984 ), .force_10(
        \filter_0/n6985 ), .force_11(1'b0), .Q(\filter_0/n7743 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6988 ), .force_10(
        \filter_0/n6989 ), .force_11(1'b0), .Q(\filter_0/n7742 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6992 ), .force_10(
        \filter_0/n6993 ), .force_11(1'b0), .Q(\filter_0/n7741 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n6996 ), .force_10(
        \filter_0/n6997 ), .force_11(1'b0), .Q(\filter_0/n7740 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7000 ), .force_10(
        \filter_0/n7001 ), .force_11(1'b0), .Q(\filter_0/n7739 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7004 ), .force_10(
        \filter_0/n7005 ), .force_11(1'b0), .Q(\filter_0/n7738 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7008 ), .force_10(
        \filter_0/n7009 ), .force_11(1'b0), .Q(\filter_0/n7737 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7012 ), .force_10(
        \filter_0/n7013 ), .force_11(1'b0), .Q(\filter_0/n7736 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7016 ), .force_10(
        \filter_0/n7017 ), .force_11(1'b0), .Q(\filter_0/n7735 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7020 ), .force_10(
        \filter_0/n7021 ), .force_11(1'b0), .Q(\filter_0/n7734 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7024 ), .force_10(
        \filter_0/n7025 ), .force_11(1'b0), .Q(\filter_0/n7733 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7028 ), .force_10(
        \filter_0/n7029 ), .force_11(1'b0), .Q(\filter_0/n7732 ) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7032 ), .force_10(
        \filter_0/n7033 ), .force_11(1'b0), .Q(\filter_0/n7731 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7036 ), .force_10(
        \filter_0/n7037 ), .force_11(1'b0), .Q(\filter_0/n7730 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7040 ), .force_10(
        \filter_0/n7041 ), .force_11(1'b0), .Q(\filter_0/n7729 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7044 ), .force_10(
        \filter_0/n7045 ), .force_11(1'b0), .Q(\filter_0/n7728 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7048 ), .force_10(
        \filter_0/n7049 ), .force_11(1'b0), .Q(\filter_0/n7727 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7052 ), .force_10(
        \filter_0/n7053 ), .force_11(1'b0), .Q(\filter_0/n7726 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7056 ), .force_10(
        \filter_0/n7057 ), .force_11(1'b0), .Q(\filter_0/n7725 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7060 ), .force_10(
        \filter_0/n7061 ), .force_11(1'b0), .Q(\filter_0/n7724 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7064 ), .force_10(
        \filter_0/n7065 ), .force_11(1'b0), .Q(\filter_0/n7723 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7068 ), .force_10(
        \filter_0/n7069 ), .force_11(1'b0), .Q(\filter_0/n7722 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7072 ), .force_10(
        \filter_0/n7073 ), .force_11(1'b0), .Q(\filter_0/n7721 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7076 ), .force_10(
        \filter_0/n7077 ), .force_11(1'b0), .Q(\filter_0/n7720 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7080 ), .force_10(
        \filter_0/n7081 ), .force_11(1'b0), .Q(\filter_0/n7719 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7084 ), .force_10(
        \filter_0/n7085 ), .force_11(1'b0), .Q(\filter_0/n7718 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7088 ), .force_10(
        \filter_0/n7089 ), .force_11(1'b0), .Q(\filter_0/n7717 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7092 ), .force_10(
        \filter_0/n7093 ), .force_11(1'b0), .Q(\filter_0/n7716 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7096 ), .force_10(
        \filter_0/n7097 ), .force_11(1'b0), .Q(\filter_0/n7715 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7100 ), .force_10(
        \filter_0/n7101 ), .force_11(1'b0), .Q(\filter_0/n7714 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7104 ), .force_10(
        \filter_0/n7105 ), .force_11(1'b0), .Q(\filter_0/n7713 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7108 ), .force_10(
        \filter_0/n7109 ), .force_11(1'b0), .Q(\filter_0/n7712 ) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7112 ), .force_10(
        \filter_0/n7113 ), .force_11(1'b0), .Q(\filter_0/n7711 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7116 ), .force_10(
        \filter_0/n7117 ), .force_11(1'b0), .Q(\filter_0/n7710 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7120 ), .force_10(
        \filter_0/n7121 ), .force_11(1'b0), .Q(\filter_0/n7709 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7124 ), .force_10(
        \filter_0/n7125 ), .force_11(1'b0), .Q(\filter_0/n7708 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7128 ), .force_10(
        \filter_0/n7129 ), .force_11(1'b0), .Q(\filter_0/n7707 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7132 ), .force_10(
        \filter_0/n7133 ), .force_11(1'b0), .Q(\filter_0/n7706 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7136 ), .force_10(
        \filter_0/n7137 ), .force_11(1'b0), .Q(\filter_0/n7705 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7140 ), .force_10(
        \filter_0/n7141 ), .force_11(1'b0), .Q(\filter_0/n7704 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7144 ), .force_10(
        \filter_0/n7145 ), .force_11(1'b0), .Q(\filter_0/n7703 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7148 ), .force_10(
        \filter_0/n7149 ), .force_11(1'b0), .Q(\filter_0/n7702 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7152 ), .force_10(
        \filter_0/n7153 ), .force_11(1'b0), .Q(\filter_0/n7701 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7156 ), .force_10(
        \filter_0/n7157 ), .force_11(1'b0), .Q(\filter_0/n7700 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7160 ), .force_10(
        \filter_0/n7161 ), .force_11(1'b0), .Q(\filter_0/n7699 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7164 ), .force_10(
        \filter_0/n7165 ), .force_11(1'b0), .Q(\filter_0/n7698 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7168 ), .force_10(
        \filter_0/n7169 ), .force_11(1'b0), .Q(\filter_0/n7697 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7172 ), .force_10(
        \filter_0/n7173 ), .force_11(1'b0), .Q(\filter_0/n7696 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7176 ), .force_10(
        \filter_0/n7177 ), .force_11(1'b0), .Q(\filter_0/n7695 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7180 ), .force_10(
        \filter_0/n7181 ), .force_11(1'b0), .Q(\filter_0/n7694 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7184 ), .force_10(
        \filter_0/n7185 ), .force_11(1'b0), .Q(\filter_0/n7693 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7188 ), .force_10(
        \filter_0/n7189 ), .force_11(1'b0), .Q(\filter_0/n7692 ) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7192 ), .force_10(
        \filter_0/n7193 ), .force_11(1'b0), .Q(\filter_0/n7691 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7196 ), .force_10(
        \filter_0/n7197 ), .force_11(1'b0), .Q(\filter_0/n7690 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7200 ), .force_10(
        \filter_0/n7201 ), .force_11(1'b0), .Q(\filter_0/n7689 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7204 ), .force_10(
        \filter_0/n7205 ), .force_11(1'b0), .Q(\filter_0/n7688 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7208 ), .force_10(
        \filter_0/n7209 ), .force_11(1'b0), .Q(\filter_0/n7687 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7212 ), .force_10(
        \filter_0/n7213 ), .force_11(1'b0), .Q(\filter_0/n7686 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7216 ), .force_10(
        \filter_0/n7217 ), .force_11(1'b0), .Q(\filter_0/n7685 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7220 ), .force_10(
        \filter_0/n7221 ), .force_11(1'b0), .Q(\filter_0/n7684 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7224 ), .force_10(
        \filter_0/n7225 ), .force_11(1'b0), .Q(\filter_0/n7683 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7228 ), .force_10(
        \filter_0/n7229 ), .force_11(1'b0), .Q(\filter_0/n7682 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7232 ), .force_10(
        \filter_0/n7233 ), .force_11(1'b0), .Q(\filter_0/n7681 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7236 ), .force_10(
        \filter_0/n7237 ), .force_11(1'b0), .Q(\filter_0/n7680 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7240 ), .force_10(
        \filter_0/n7241 ), .force_11(1'b0), .Q(\filter_0/n7679 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7244 ), .force_10(
        \filter_0/n7245 ), .force_11(1'b0), .Q(\filter_0/n7678 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7248 ), .force_10(
        \filter_0/n7249 ), .force_11(1'b0), .Q(\filter_0/n7677 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7252 ), .force_10(
        \filter_0/n7253 ), .force_11(1'b0), .Q(\filter_0/n7676 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7256 ), .force_10(
        \filter_0/n7257 ), .force_11(1'b0), .Q(\filter_0/n7675 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7260 ), .force_10(
        \filter_0/n7261 ), .force_11(1'b0), .Q(\filter_0/n7674 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7264 ), .force_10(
        \filter_0/n7265 ), .force_11(1'b0), .Q(\filter_0/n7673 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7268 ), .force_10(
        \filter_0/n7269 ), .force_11(1'b0), .Q(\filter_0/n7672 ) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7272 ), .force_10(
        \filter_0/n7273 ), .force_11(1'b0), .Q(\filter_0/n7671 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7276 ), .force_10(
        \filter_0/n7277 ), .force_11(1'b0), .Q(\filter_0/n7670 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7280 ), .force_10(
        \filter_0/n7281 ), .force_11(1'b0), .Q(\filter_0/n7669 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7284 ), .force_10(
        \filter_0/n7285 ), .force_11(1'b0), .Q(\filter_0/n7668 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7288 ), .force_10(
        \filter_0/n7289 ), .force_11(1'b0), .Q(\filter_0/n7667 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7292 ), .force_10(
        \filter_0/n7293 ), .force_11(1'b0), .Q(\filter_0/n7666 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7296 ), .force_10(
        \filter_0/n7297 ), .force_11(1'b0), .Q(\filter_0/n7665 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7300 ), .force_10(
        \filter_0/n7301 ), .force_11(1'b0), .Q(\filter_0/n7664 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7304 ), .force_10(
        \filter_0/n7305 ), .force_11(1'b0), .Q(\filter_0/n7663 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7308 ), .force_10(
        \filter_0/n7309 ), .force_11(1'b0), .Q(\filter_0/n7662 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7312 ), .force_10(
        \filter_0/n7313 ), .force_11(1'b0), .Q(\filter_0/n7661 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7316 ), .force_10(
        \filter_0/n7317 ), .force_11(1'b0), .Q(\filter_0/n7660 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7320 ), .force_10(
        \filter_0/n7321 ), .force_11(1'b0), .Q(\filter_0/n7659 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7324 ), .force_10(
        \filter_0/n7325 ), .force_11(1'b0), .Q(\filter_0/n7658 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7328 ), .force_10(
        \filter_0/n7329 ), .force_11(1'b0), .Q(\filter_0/n7657 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7332 ), .force_10(
        \filter_0/n7333 ), .force_11(1'b0), .Q(\filter_0/n7656 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7336 ), .force_10(
        \filter_0/n7337 ), .force_11(1'b0), .Q(\filter_0/n7655 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7340 ), .force_10(
        \filter_0/n7341 ), .force_11(1'b0), .Q(\filter_0/n7654 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7344 ), .force_10(
        \filter_0/n7345 ), .force_11(1'b0), .Q(\filter_0/n7653 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7348 ), .force_10(
        \filter_0/n7349 ), .force_11(1'b0), .Q(\filter_0/n7652 ) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7352 ), .force_10(
        \filter_0/n7353 ), .force_11(1'b0), .Q(\filter_0/n7651 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7356 ), .force_10(
        \filter_0/n7357 ), .force_11(1'b0), .Q(\filter_0/n7650 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7360 ), .force_10(
        \filter_0/n7361 ), .force_11(1'b0), .Q(\filter_0/n7649 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7364 ), .force_10(
        \filter_0/n7365 ), .force_11(1'b0), .Q(\filter_0/n7648 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7368 ), .force_10(
        \filter_0/n7369 ), .force_11(1'b0), .Q(\filter_0/n7647 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7372 ), .force_10(
        \filter_0/n7373 ), .force_11(1'b0), .Q(\filter_0/n7646 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7376 ), .force_10(
        \filter_0/n7377 ), .force_11(1'b0), .Q(\filter_0/n7645 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7380 ), .force_10(
        \filter_0/n7381 ), .force_11(1'b0), .Q(\filter_0/n7644 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7384 ), .force_10(
        \filter_0/n7385 ), .force_11(1'b0), .Q(\filter_0/n7643 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7388 ), .force_10(
        \filter_0/n7389 ), .force_11(1'b0), .Q(\filter_0/n7642 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7392 ), .force_10(
        \filter_0/n7393 ), .force_11(1'b0), .Q(\filter_0/n7641 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7396 ), .force_10(
        \filter_0/n7397 ), .force_11(1'b0), .Q(\filter_0/n7640 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7400 ), .force_10(
        \filter_0/n7401 ), .force_11(1'b0), .Q(\filter_0/n7639 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7404 ), .force_10(
        \filter_0/n7405 ), .force_11(1'b0), .Q(\filter_0/n7638 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7408 ), .force_10(
        \filter_0/n7409 ), .force_11(1'b0), .Q(\filter_0/n7637 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7412 ), .force_10(
        \filter_0/n7413 ), .force_11(1'b0), .Q(\filter_0/n7636 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7416 ), .force_10(
        \filter_0/n7417 ), .force_11(1'b0), .Q(\filter_0/n7635 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7420 ), .force_10(
        \filter_0/n7421 ), .force_11(1'b0), .Q(\filter_0/n7634 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7424 ), .force_10(
        \filter_0/n7425 ), .force_11(1'b0), .Q(\filter_0/n7633 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7428 ), .force_10(
        \filter_0/n7429 ), .force_11(1'b0), .Q(\filter_0/n7632 ) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7432 ), .force_10(
        \filter_0/n7433 ), .force_11(1'b0), .Q(\filter_0/n7631 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7436 ), .force_10(\filter_0/n7437 ), 
        .force_11(1'b0), .Q(\filter_0/n7630 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7440 ), .force_10(\filter_0/n7441 ), 
        .force_11(1'b0), .Q(\filter_0/n7629 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7444 ), .force_10(\filter_0/n7445 ), 
        .force_11(1'b0), .Q(\filter_0/n7628 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7448 ), .force_10(\filter_0/n7449 ), 
        .force_11(1'b0), .Q(\filter_0/n7627 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7452 ), .force_10(\filter_0/n7453 ), 
        .force_11(1'b0), .Q(\filter_0/n7626 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7456 ), .force_10(\filter_0/n7457 ), 
        .force_11(1'b0), .Q(\filter_0/n7625 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7460 ), .force_10(\filter_0/n7461 ), 
        .force_11(1'b0), .Q(\filter_0/n7624 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7464 ), .force_10(\filter_0/n7465 ), 
        .force_11(1'b0), .Q(\filter_0/n7623 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7468 ), .force_10(\filter_0/n7469 ), 
        .force_11(1'b0), .Q(\filter_0/n7622 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7472 ), .force_10(\filter_0/n7473 ), 
        .force_11(1'b0), .Q(\filter_0/n7621 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7476 ), .force_10(
        \filter_0/n7477 ), .force_11(1'b0), .Q(\filter_0/n7620 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7480 ), .force_10(
        \filter_0/n7481 ), .force_11(1'b0), .Q(\filter_0/n7619 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7484 ), .force_10(
        \filter_0/n7485 ), .force_11(1'b0), .Q(\filter_0/n7618 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7488 ), .force_10(
        \filter_0/n7489 ), .force_11(1'b0), .Q(\filter_0/n7617 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7492 ), .force_10(
        \filter_0/n7493 ), .force_11(1'b0), .Q(\filter_0/n7616 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7496 ), .force_10(
        \filter_0/n7497 ), .force_11(1'b0), .Q(\filter_0/n7615 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7500 ), .force_10(
        \filter_0/n7501 ), .force_11(1'b0), .Q(\filter_0/n7614 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7504 ), .force_10(
        \filter_0/n7505 ), .force_11(1'b0), .Q(\filter_0/n7613 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7508 ), .force_10(
        \filter_0/n7509 ), .force_11(1'b0), .Q(\filter_0/n7612 ) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7512 ), .force_10(
        \filter_0/n7513 ), .force_11(1'b0), .Q(\filter_0/n7611 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7516 ), .force_10(\filter_0/n7517 ), 
        .force_11(1'b0), .Q(\filter_0/n7610 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7520 ), .force_10(\filter_0/n7521 ), 
        .force_11(1'b0), .Q(\filter_0/n7609 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7524 ), .force_10(\filter_0/n7525 ), 
        .force_11(1'b0), .Q(\filter_0/n7608 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7528 ), .force_10(\filter_0/n7529 ), 
        .force_11(1'b0), .Q(\filter_0/n7607 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7532 ), .force_10(\filter_0/n7533 ), 
        .force_11(1'b0), .Q(\filter_0/n7606 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7536 ), .force_10(\filter_0/n7537 ), 
        .force_11(1'b0), .Q(\filter_0/n7605 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7540 ), .force_10(\filter_0/n7541 ), 
        .force_11(1'b0), .Q(\filter_0/n7604 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7544 ), .force_10(\filter_0/n7545 ), 
        .force_11(1'b0), .Q(\filter_0/n7603 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7548 ), .force_10(\filter_0/n7549 ), 
        .force_11(1'b0), .Q(\filter_0/n7602 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n7552 ), .force_10(\filter_0/n7553 ), 
        .force_11(1'b0), .Q(\filter_0/n7601 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7556 ), .force_10(
        \filter_0/n7557 ), .force_11(1'b0), .Q(\filter_0/n7600 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7560 ), .force_10(
        \filter_0/n7561 ), .force_11(1'b0), .Q(\filter_0/n7599 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7564 ), .force_10(
        \filter_0/n7565 ), .force_11(1'b0), .Q(\filter_0/n7598 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7568 ), .force_10(
        \filter_0/n7569 ), .force_11(1'b0), .Q(\filter_0/n7597 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7572 ), .force_10(
        \filter_0/n7573 ), .force_11(1'b0), .Q(\filter_0/n7596 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7576 ), .force_10(
        \filter_0/n7577 ), .force_11(1'b0), .Q(\filter_0/n7595 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7580 ), .force_10(
        \filter_0/n7581 ), .force_11(1'b0), .Q(\filter_0/n7594 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7584 ), .force_10(
        \filter_0/n7585 ), .force_11(1'b0), .Q(\filter_0/n7593 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n7588 ), .force_10(
        \filter_0/n7589 ), .force_11(1'b0), .Q(\filter_0/n7592 ) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n4980 ), .force_10(
        \filter_0/n4981 ), .force_11(1'b0), .Q(\filter_0/n7591 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6397 ), .force_10(
        \shifter_0/n6398 ), .force_11(1'b0), .Q(\shifter_0/n9591 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6401 ), .force_10(
        \shifter_0/n6402 ), .force_11(1'b0), .Q(\shifter_0/n9590 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6405 ), .force_10(
        \shifter_0/n6406 ), .force_11(1'b0), .Q(\shifter_0/n9589 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6409 ), .force_10(
        \shifter_0/n6410 ), .force_11(1'b0), .Q(\shifter_0/n9588 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6413 ), .force_10(
        \shifter_0/n6414 ), .force_11(1'b0), .Q(\shifter_0/n9587 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6417 ), .force_10(
        \shifter_0/n6418 ), .force_11(1'b0), .Q(\shifter_0/n9586 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6421 ), .force_10(
        \shifter_0/n6422 ), .force_11(1'b0), .Q(\shifter_0/n9585 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6425 ), .force_10(
        \shifter_0/n6426 ), .force_11(1'b0), .Q(\shifter_0/n9584 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6429 ), .force_10(
        \shifter_0/n6430 ), .force_11(1'b0), .Q(\shifter_0/n9583 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6433 ), .force_10(
        \shifter_0/n6434 ), .force_11(1'b0), .Q(\shifter_0/n9582 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6437 ), .force_10(
        \shifter_0/n6438 ), .force_11(1'b0), .Q(\shifter_0/n9581 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6441 ), .force_10(
        \shifter_0/n6442 ), .force_11(1'b0), .Q(\shifter_0/n9580 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6445 ), .force_10(
        \shifter_0/n6446 ), .force_11(1'b0), .Q(\shifter_0/n9579 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6449 ), .force_10(
        \shifter_0/n6450 ), .force_11(1'b0), .Q(\shifter_0/n9578 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6453 ), .force_10(
        \shifter_0/n6454 ), .force_11(1'b0), .Q(\shifter_0/n9577 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6457 ), .force_10(
        \shifter_0/n6458 ), .force_11(1'b0), .Q(\shifter_0/n9576 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6461 ), .force_10(
        \shifter_0/n6462 ), .force_11(1'b0), .Q(\shifter_0/n9575 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6465 ), .force_10(
        \shifter_0/n6466 ), .force_11(1'b0), .Q(\shifter_0/n9574 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6469 ), .force_10(
        \shifter_0/n6470 ), .force_11(1'b0), .Q(\shifter_0/n9573 ) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6473 ), .force_10(
        \shifter_0/n6474 ), .force_11(1'b0), .Q(\shifter_0/n9572 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6477 ), .force_10(n41624), .force_11(1'b0), .Q(\shifter_0/n9571 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6481 ), .force_10(n41623), .force_11(1'b0), .Q(\shifter_0/n9570 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6485 ), .force_10(n41622), .force_11(1'b0), .Q(\shifter_0/n9569 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6489 ), .force_10(n41621), .force_11(1'b0), .Q(\shifter_0/n9568 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6493 ), .force_10(n41620), .force_11(1'b0), .Q(\shifter_0/n9567 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6497 ), .force_10(n41619), .force_11(1'b0), .Q(\shifter_0/n9566 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6501 ), .force_10(n41618), .force_11(1'b0), .Q(\shifter_0/n9565 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6505 ), .force_10(n41617), .force_11(1'b0), .Q(\shifter_0/n9564 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6509 ), .force_10(n41616), .force_11(1'b0), .Q(\shifter_0/n9563 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6513 ), .force_10(n41615), .force_11(1'b0), .Q(\shifter_0/n9562 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6517 ), .force_10(n41614), .force_11(1'b0), .Q(\shifter_0/n9561 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6521 ), .force_10(n41613), .force_11(1'b0), .Q(\shifter_0/n9560 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6525 ), .force_10(n41612), .force_11(1'b0), .Q(\shifter_0/n9559 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6529 ), .force_10(n41611), .force_11(1'b0), .Q(\shifter_0/n9558 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6533 ), .force_10(n41610), .force_11(1'b0), .Q(\shifter_0/n9557 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6537 ), .force_10(n41609), .force_11(1'b0), .Q(\shifter_0/n9556 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6541 ), .force_10(n41608), .force_11(1'b0), .Q(\shifter_0/n9555 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6545 ), .force_10(n41607), .force_11(1'b0), .Q(\shifter_0/n9554 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6549 ), .force_10(n41606), .force_11(1'b0), .Q(\shifter_0/n9553 ) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6553 ), .force_10(n41605), .force_11(1'b0), .Q(\shifter_0/n9552 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6557 ), .force_10(n41341), .force_11(1'b0), .Q(\shifter_0/n9551 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6561 ), .force_10(n41345), .force_11(1'b0), .Q(\shifter_0/n9550 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6565 ), .force_10(n41349), .force_11(1'b0), .Q(\shifter_0/n9549 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6569 ), .force_10(n41353), .force_11(1'b0), .Q(\shifter_0/n9548 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6573 ), .force_10(n41357), .force_11(1'b0), .Q(\shifter_0/n9547 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6577 ), .force_10(n41361), .force_11(1'b0), .Q(\shifter_0/n9546 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6581 ), .force_10(n41365), .force_11(1'b0), .Q(\shifter_0/n9545 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6585 ), .force_10(n41369), .force_11(1'b0), .Q(\shifter_0/n9544 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6589 ), .force_10(n41373), .force_11(1'b0), .Q(\shifter_0/n9543 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6593 ), .force_10(n41377), .force_11(1'b0), .Q(\shifter_0/n9542 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6597 ), .force_10(n41381), .force_11(1'b0), .Q(\shifter_0/n9541 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6601 ), .force_10(n41385), .force_11(1'b0), .Q(\shifter_0/n9540 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6605 ), .force_10(n41389), .force_11(1'b0), .Q(\shifter_0/n9539 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6609 ), .force_10(n41393), .force_11(1'b0), .Q(\shifter_0/n9538 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6613 ), .force_10(n41397), .force_11(1'b0), .Q(\shifter_0/n9537 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6617 ), .force_10(n41401), .force_11(1'b0), .Q(\shifter_0/n9536 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6621 ), .force_10(n41405), .force_11(1'b0), .Q(\shifter_0/n9535 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6625 ), .force_10(n41409), .force_11(1'b0), .Q(\shifter_0/n9534 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6629 ), .force_10(n41413), .force_11(1'b0), .Q(\shifter_0/n9533 ) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6633 ), .force_10(n41417), .force_11(1'b0), .Q(\shifter_0/n9532 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6637 ), .force_10(n41644), .force_11(1'b0), .Q(\shifter_0/n9531 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6641 ), .force_10(n41643), .force_11(1'b0), .Q(\shifter_0/n9530 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6645 ), .force_10(n41642), .force_11(1'b0), .Q(\shifter_0/n9529 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6649 ), .force_10(n41641), .force_11(1'b0), .Q(\shifter_0/n9528 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6653 ), .force_10(n41640), .force_11(1'b0), .Q(\shifter_0/n9527 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6657 ), .force_10(n41639), .force_11(1'b0), .Q(\shifter_0/n9526 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6661 ), .force_10(n41638), .force_11(1'b0), .Q(\shifter_0/n9525 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6665 ), .force_10(n41637), .force_11(1'b0), .Q(\shifter_0/n9524 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6669 ), .force_10(n41636), .force_11(1'b0), .Q(\shifter_0/n9523 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6673 ), .force_10(n41635), .force_11(1'b0), .Q(\shifter_0/n9522 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6677 ), .force_10(n41634), .force_11(1'b0), .Q(\shifter_0/n9521 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6681 ), .force_10(n41633), .force_11(1'b0), .Q(\shifter_0/n9520 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6685 ), .force_10(n41632), .force_11(1'b0), .Q(\shifter_0/n9519 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6689 ), .force_10(n41631), .force_11(1'b0), .Q(\shifter_0/n9518 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6693 ), .force_10(n41630), .force_11(1'b0), .Q(\shifter_0/n9517 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6697 ), .force_10(n41629), .force_11(1'b0), .Q(\shifter_0/n9516 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6701 ), .force_10(n41628), .force_11(1'b0), .Q(\shifter_0/n9515 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6705 ), .force_10(n41627), .force_11(1'b0), .Q(\shifter_0/n9514 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6709 ), .force_10(n41626), .force_11(1'b0), .Q(\shifter_0/n9513 ) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6713 ), .force_10(n41625), .force_11(1'b0), .Q(\shifter_0/n9512 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6717 ), .force_10(n41340), .force_11(1'b0), .Q(\shifter_0/n9511 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6721 ), .force_10(n41344), .force_11(1'b0), .Q(\shifter_0/n9510 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6725 ), .force_10(n41348), .force_11(1'b0), .Q(\shifter_0/n9509 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6729 ), .force_10(n41352), .force_11(1'b0), .Q(\shifter_0/n9508 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6733 ), .force_10(n41356), .force_11(1'b0), .Q(\shifter_0/n9507 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6737 ), .force_10(n41360), .force_11(1'b0), .Q(\shifter_0/n9506 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6741 ), .force_10(n41364), .force_11(1'b0), .Q(\shifter_0/n9505 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6745 ), .force_10(n41368), .force_11(1'b0), .Q(\shifter_0/n9504 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6749 ), .force_10(n41372), .force_11(1'b0), .Q(\shifter_0/n9503 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6753 ), .force_10(n41376), .force_11(1'b0), .Q(\shifter_0/n9502 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6757 ), .force_10(n41380), .force_11(1'b0), .Q(\shifter_0/n9501 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6761 ), .force_10(n41384), .force_11(1'b0), .Q(\shifter_0/n9500 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6765 ), .force_10(n41388), .force_11(1'b0), .Q(\shifter_0/n9499 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6769 ), .force_10(n41392), .force_11(1'b0), .Q(\shifter_0/n9498 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6773 ), .force_10(n41396), .force_11(1'b0), .Q(\shifter_0/n9497 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6777 ), .force_10(n41400), .force_11(1'b0), .Q(\shifter_0/n9496 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6781 ), .force_10(n41404), .force_11(1'b0), .Q(\shifter_0/n9495 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6785 ), .force_10(n41408), .force_11(1'b0), .Q(\shifter_0/n9494 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6789 ), .force_10(n41412), .force_11(1'b0), .Q(\shifter_0/n9493 ) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6793 ), .force_10(n41416), .force_11(1'b0), .Q(\shifter_0/n9492 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6797 ), .force_10(n41704), .force_11(1'b0), .Q(\shifter_0/n9491 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6801 ), .force_10(n41703), .force_11(1'b0), .Q(\shifter_0/n9490 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6805 ), .force_10(n41702), .force_11(1'b0), .Q(\shifter_0/n9489 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6809 ), .force_10(n41701), .force_11(1'b0), .Q(\shifter_0/n9488 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6813 ), .force_10(n41700), .force_11(1'b0), .Q(\shifter_0/n9487 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6817 ), .force_10(n41699), .force_11(1'b0), .Q(\shifter_0/n9486 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6821 ), .force_10(n41698), .force_11(1'b0), .Q(\shifter_0/n9485 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6825 ), .force_10(n41697), .force_11(1'b0), .Q(\shifter_0/n9484 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6829 ), .force_10(n41696), .force_11(1'b0), .Q(\shifter_0/n9483 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6833 ), .force_10(n41695), .force_11(1'b0), .Q(\shifter_0/n9482 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6837 ), .force_10(n41694), .force_11(1'b0), .Q(\shifter_0/n9481 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6841 ), .force_10(n41693), .force_11(1'b0), .Q(\shifter_0/n9480 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6845 ), .force_10(n41692), .force_11(1'b0), .Q(\shifter_0/n9479 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6849 ), .force_10(n41691), .force_11(1'b0), .Q(\shifter_0/n9478 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6853 ), .force_10(n41690), .force_11(1'b0), .Q(\shifter_0/n9477 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6857 ), .force_10(n41689), .force_11(1'b0), .Q(\shifter_0/n9476 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6861 ), .force_10(n41688), .force_11(1'b0), .Q(\shifter_0/n9475 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6865 ), .force_10(n41687), .force_11(1'b0), .Q(\shifter_0/n9474 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6869 ), .force_10(n41686), .force_11(1'b0), .Q(\shifter_0/n9473 ) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6873 ), .force_10(n41685), .force_11(1'b0), .Q(\shifter_0/n9472 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6877 ), .force_10(n41543), .force_11(1'b0), .Q(\shifter_0/n9471 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6881 ), .force_10(n41542), .force_11(1'b0), .Q(\shifter_0/n9470 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6885 ), .force_10(n41541), .force_11(1'b0), .Q(\shifter_0/n9469 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6889 ), .force_10(n41540), .force_11(1'b0), .Q(\shifter_0/n9468 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6893 ), .force_10(n41539), .force_11(1'b0), .Q(\shifter_0/n9467 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6897 ), .force_10(n41538), .force_11(1'b0), .Q(\shifter_0/n9466 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6901 ), .force_10(n41537), .force_11(1'b0), .Q(\shifter_0/n9465 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6905 ), .force_10(n41536), .force_11(1'b0), .Q(\shifter_0/n9464 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6909 ), .force_10(n41535), .force_11(1'b0), .Q(\shifter_0/n9463 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6913 ), .force_10(n41534), .force_11(1'b0), .Q(\shifter_0/n9462 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6917 ), .force_10(n41533), .force_11(1'b0), .Q(\shifter_0/n9461 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6921 ), .force_10(n41532), .force_11(1'b0), .Q(\shifter_0/n9460 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6925 ), .force_10(n41531), .force_11(1'b0), .Q(\shifter_0/n9459 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6929 ), .force_10(n41530), .force_11(1'b0), .Q(\shifter_0/n9458 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6933 ), .force_10(n41529), .force_11(1'b0), .Q(\shifter_0/n9457 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6937 ), .force_10(n41528), .force_11(1'b0), .Q(\shifter_0/n9456 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6941 ), .force_10(n41527), .force_11(1'b0), .Q(\shifter_0/n9455 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6945 ), .force_10(n41526), .force_11(1'b0), .Q(\shifter_0/n9454 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6949 ), .force_10(n41525), .force_11(1'b0), .Q(\shifter_0/n9453 ) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6953 ), .force_10(n41524), .force_11(1'b0), .Q(\shifter_0/n9452 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6957 ), .force_10(n41725), .force_11(1'b0), .Q(\shifter_0/n9451 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6961 ), .force_10(n41724), .force_11(1'b0), .Q(\shifter_0/n9450 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6965 ), .force_10(n41723), .force_11(1'b0), .Q(\shifter_0/n9449 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6969 ), .force_10(n41722), .force_11(1'b0), .Q(\shifter_0/n9448 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6973 ), .force_10(n41721), .force_11(1'b0), .Q(\shifter_0/n9447 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6977 ), .force_10(n41720), .force_11(1'b0), .Q(\shifter_0/n9446 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6981 ), .force_10(n41719), .force_11(1'b0), .Q(\shifter_0/n9445 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6985 ), .force_10(n41718), .force_11(1'b0), .Q(\shifter_0/n9444 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6989 ), .force_10(n41717), .force_11(1'b0), .Q(\shifter_0/n9443 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6993 ), .force_10(n41716), .force_11(1'b0), .Q(\shifter_0/n9442 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6997 ), .force_10(n41715), .force_11(1'b0), .Q(\shifter_0/n9441 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7001 ), .force_10(n41714), .force_11(1'b0), .Q(\shifter_0/n9440 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7005 ), .force_10(n41713), .force_11(1'b0), .Q(\shifter_0/n9439 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7009 ), .force_10(n41712), .force_11(1'b0), .Q(\shifter_0/n9438 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7013 ), .force_10(n41711), .force_11(1'b0), .Q(\shifter_0/n9437 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7017 ), .force_10(n41710), .force_11(1'b0), .Q(\shifter_0/n9436 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7021 ), .force_10(n41709), .force_11(1'b0), .Q(\shifter_0/n9435 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7025 ), .force_10(n41708), .force_11(1'b0), .Q(\shifter_0/n9434 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7029 ), .force_10(n41707), .force_11(1'b0), .Q(\shifter_0/n9433 ) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7033 ), .force_10(n41706), .force_11(1'b0), .Q(\shifter_0/n9432 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7037 ), .force_10(n41339), .force_11(1'b0), .Q(\shifter_0/n9431 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7041 ), .force_10(n41343), .force_11(1'b0), .Q(\shifter_0/n9430 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7045 ), .force_10(n41347), .force_11(1'b0), .Q(\shifter_0/n9429 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7049 ), .force_10(n41351), .force_11(1'b0), .Q(\shifter_0/n9428 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7053 ), .force_10(n41355), .force_11(1'b0), .Q(\shifter_0/n9427 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7057 ), .force_10(n41359), .force_11(1'b0), .Q(\shifter_0/n9426 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7061 ), .force_10(n41363), .force_11(1'b0), .Q(\shifter_0/n9425 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7065 ), .force_10(n41367), .force_11(1'b0), .Q(\shifter_0/n9424 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7069 ), .force_10(n41371), .force_11(1'b0), .Q(\shifter_0/n9423 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7073 ), .force_10(n41375), .force_11(1'b0), .Q(\shifter_0/n9422 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7077 ), .force_10(n41379), .force_11(1'b0), .Q(\shifter_0/n9421 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7081 ), .force_10(n41383), .force_11(1'b0), .Q(\shifter_0/n9420 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7085 ), .force_10(n41387), .force_11(1'b0), .Q(\shifter_0/n9419 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7089 ), .force_10(n41391), .force_11(1'b0), .Q(\shifter_0/n9418 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7093 ), .force_10(n41395), .force_11(1'b0), .Q(\shifter_0/n9417 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7097 ), .force_10(n41399), .force_11(1'b0), .Q(\shifter_0/n9416 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7101 ), .force_10(n41403), .force_11(1'b0), .Q(\shifter_0/n9415 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7105 ), .force_10(n41407), .force_11(1'b0), .Q(\shifter_0/n9414 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7109 ), .force_10(n41411), .force_11(1'b0), .Q(\shifter_0/n9413 ) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7113 ), .force_10(n41415), .force_11(1'b0), .Q(\shifter_0/n9412 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7117 ), .force_10(
        \shifter_0/n7118 ), .force_11(1'b0), .Q(\shifter_0/n9411 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7121 ), .force_10(
        \shifter_0/n7122 ), .force_11(1'b0), .Q(\shifter_0/n9410 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7125 ), .force_10(
        \shifter_0/n7126 ), .force_11(1'b0), .Q(\shifter_0/n9409 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7129 ), .force_10(
        \shifter_0/n7130 ), .force_11(1'b0), .Q(\shifter_0/n9408 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7133 ), .force_10(
        \shifter_0/n7134 ), .force_11(1'b0), .Q(\shifter_0/n9407 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7137 ), .force_10(
        \shifter_0/n7138 ), .force_11(1'b0), .Q(\shifter_0/n9406 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7141 ), .force_10(
        \shifter_0/n7142 ), .force_11(1'b0), .Q(\shifter_0/n9405 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7145 ), .force_10(
        \shifter_0/n7146 ), .force_11(1'b0), .Q(\shifter_0/n9404 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7149 ), .force_10(
        \shifter_0/n7150 ), .force_11(1'b0), .Q(\shifter_0/n9403 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7153 ), .force_10(
        \shifter_0/n7154 ), .force_11(1'b0), .Q(\shifter_0/n9402 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7157 ), .force_10(
        \shifter_0/n7158 ), .force_11(1'b0), .Q(\shifter_0/n9401 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7161 ), .force_10(
        \shifter_0/n7162 ), .force_11(1'b0), .Q(\shifter_0/n9400 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7165 ), .force_10(
        \shifter_0/n7166 ), .force_11(1'b0), .Q(\shifter_0/n9399 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7169 ), .force_10(
        \shifter_0/n7170 ), .force_11(1'b0), .Q(\shifter_0/n9398 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7173 ), .force_10(
        \shifter_0/n7174 ), .force_11(1'b0), .Q(\shifter_0/n9397 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7177 ), .force_10(
        \shifter_0/n7178 ), .force_11(1'b0), .Q(\shifter_0/n9396 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7181 ), .force_10(
        \shifter_0/n7182 ), .force_11(1'b0), .Q(\shifter_0/n9395 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7185 ), .force_10(
        \shifter_0/n7186 ), .force_11(1'b0), .Q(\shifter_0/n9394 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7189 ), .force_10(
        \shifter_0/n7190 ), .force_11(1'b0), .Q(\shifter_0/n9393 ) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7193 ), .force_10(
        \shifter_0/n7194 ), .force_11(1'b0), .Q(\shifter_0/n9392 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7197 ), .force_10(
        \shifter_0/n7198 ), .force_11(1'b0), .Q(\shifter_0/n9391 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7201 ), .force_10(
        \shifter_0/n7202 ), .force_11(1'b0), .Q(\shifter_0/n9390 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7205 ), .force_10(
        \shifter_0/n7206 ), .force_11(1'b0), .Q(\shifter_0/n9389 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7209 ), .force_10(
        \shifter_0/n7210 ), .force_11(1'b0), .Q(\shifter_0/n9388 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7213 ), .force_10(
        \shifter_0/n7214 ), .force_11(1'b0), .Q(\shifter_0/n9387 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7217 ), .force_10(
        \shifter_0/n7218 ), .force_11(1'b0), .Q(\shifter_0/n9386 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7221 ), .force_10(
        \shifter_0/n7222 ), .force_11(1'b0), .Q(\shifter_0/n9385 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7225 ), .force_10(
        \shifter_0/n7226 ), .force_11(1'b0), .Q(\shifter_0/n9384 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7229 ), .force_10(
        \shifter_0/n7230 ), .force_11(1'b0), .Q(\shifter_0/n9383 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7233 ), .force_10(
        \shifter_0/n7234 ), .force_11(1'b0), .Q(\shifter_0/n9382 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7237 ), .force_10(
        \shifter_0/n7238 ), .force_11(1'b0), .Q(\shifter_0/n9381 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7241 ), .force_10(
        \shifter_0/n7242 ), .force_11(1'b0), .Q(\shifter_0/n9380 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7245 ), .force_10(
        \shifter_0/n7246 ), .force_11(1'b0), .Q(\shifter_0/n9379 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7249 ), .force_10(
        \shifter_0/n7250 ), .force_11(1'b0), .Q(\shifter_0/n9378 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7253 ), .force_10(
        \shifter_0/n7254 ), .force_11(1'b0), .Q(\shifter_0/n9377 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7257 ), .force_10(
        \shifter_0/n7258 ), .force_11(1'b0), .Q(\shifter_0/n9376 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7261 ), .force_10(
        \shifter_0/n7262 ), .force_11(1'b0), .Q(\shifter_0/n9375 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7265 ), .force_10(
        \shifter_0/n7266 ), .force_11(1'b0), .Q(\shifter_0/n9374 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7269 ), .force_10(
        \shifter_0/n7270 ), .force_11(1'b0), .Q(\shifter_0/n9373 ) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7273 ), .force_10(
        \shifter_0/n7274 ), .force_11(1'b0), .Q(\shifter_0/n9372 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7277 ), .force_10(n41684), .force_11(1'b0), .Q(\shifter_0/n9371 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7281 ), .force_10(n41683), .force_11(1'b0), .Q(\shifter_0/n9370 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7285 ), .force_10(n41682), .force_11(1'b0), .Q(\shifter_0/n9369 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7289 ), .force_10(n41681), .force_11(1'b0), .Q(\shifter_0/n9368 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7293 ), .force_10(n41680), .force_11(1'b0), .Q(\shifter_0/n9367 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7297 ), .force_10(n41679), .force_11(1'b0), .Q(\shifter_0/n9366 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7301 ), .force_10(n41678), .force_11(1'b0), .Q(\shifter_0/n9365 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7305 ), .force_10(n41677), .force_11(1'b0), .Q(\shifter_0/n9364 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7309 ), .force_10(n41676), .force_11(1'b0), .Q(\shifter_0/n9363 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7313 ), .force_10(n41675), .force_11(1'b0), .Q(\shifter_0/n9362 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7317 ), .force_10(n41674), .force_11(1'b0), .Q(\shifter_0/n9361 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7321 ), .force_10(n41673), .force_11(1'b0), .Q(\shifter_0/n9360 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7325 ), .force_10(n41672), .force_11(1'b0), .Q(\shifter_0/n9359 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7329 ), .force_10(n41671), .force_11(1'b0), .Q(\shifter_0/n9358 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7333 ), .force_10(n41670), .force_11(1'b0), .Q(\shifter_0/n9357 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7337 ), .force_10(n41669), .force_11(1'b0), .Q(\shifter_0/n9356 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7341 ), .force_10(n41668), .force_11(1'b0), .Q(\shifter_0/n9355 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7345 ), .force_10(n41667), .force_11(1'b0), .Q(\shifter_0/n9354 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7349 ), .force_10(n41666), .force_11(1'b0), .Q(\shifter_0/n9353 ) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7353 ), .force_10(n41665), .force_11(1'b0), .Q(\shifter_0/n9352 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7357 ), .force_10(n41544), .force_11(1'b0), .Q(\shifter_0/n9351 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7361 ), .force_10(n41545), .force_11(1'b0), .Q(\shifter_0/n9350 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7365 ), .force_10(n41546), .force_11(1'b0), .Q(\shifter_0/n9349 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7369 ), .force_10(n41547), .force_11(1'b0), .Q(\shifter_0/n9348 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7373 ), .force_10(n41548), .force_11(1'b0), .Q(\shifter_0/n9347 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7377 ), .force_10(n41549), .force_11(1'b0), .Q(\shifter_0/n9346 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7381 ), .force_10(n41550), .force_11(1'b0), .Q(\shifter_0/n9345 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7385 ), .force_10(n41551), .force_11(1'b0), .Q(\shifter_0/n9344 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7389 ), .force_10(n41552), .force_11(1'b0), .Q(\shifter_0/n9343 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7393 ), .force_10(n41553), .force_11(1'b0), .Q(\shifter_0/n9342 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7397 ), .force_10(n41554), .force_11(1'b0), .Q(\shifter_0/n9341 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7401 ), .force_10(n41555), .force_11(1'b0), .Q(\shifter_0/n9340 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7405 ), .force_10(n41556), .force_11(1'b0), .Q(\shifter_0/n9339 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7409 ), .force_10(n41557), .force_11(1'b0), .Q(\shifter_0/n9338 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7413 ), .force_10(n41558), .force_11(1'b0), .Q(\shifter_0/n9337 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7417 ), .force_10(n41559), .force_11(1'b0), .Q(\shifter_0/n9336 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7421 ), .force_10(n41560), .force_11(1'b0), .Q(\shifter_0/n9335 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7425 ), .force_10(n41561), .force_11(1'b0), .Q(\shifter_0/n9334 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7429 ), .force_10(n41562), .force_11(1'b0), .Q(\shifter_0/n9333 ) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7433 ), .force_10(n41563), .force_11(1'b0), .Q(\shifter_0/n9332 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7437 ), .force_10(
        \shifter_0/n7438 ), .force_11(1'b0), .Q(\shifter_0/n9331 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7441 ), .force_10(
        \shifter_0/n7442 ), .force_11(1'b0), .Q(\shifter_0/n9330 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7445 ), .force_10(
        \shifter_0/n7446 ), .force_11(1'b0), .Q(\shifter_0/n9329 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7449 ), .force_10(
        \shifter_0/n7450 ), .force_11(1'b0), .Q(\shifter_0/n9328 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7453 ), .force_10(
        \shifter_0/n7454 ), .force_11(1'b0), .Q(\shifter_0/n9327 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7457 ), .force_10(
        \shifter_0/n7458 ), .force_11(1'b0), .Q(\shifter_0/n9326 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7461 ), .force_10(
        \shifter_0/n7462 ), .force_11(1'b0), .Q(\shifter_0/n9325 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7465 ), .force_10(
        \shifter_0/n7466 ), .force_11(1'b0), .Q(\shifter_0/n9324 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7469 ), .force_10(
        \shifter_0/n7470 ), .force_11(1'b0), .Q(\shifter_0/n9323 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7473 ), .force_10(
        \shifter_0/n7474 ), .force_11(1'b0), .Q(\shifter_0/n9322 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7477 ), .force_10(
        \shifter_0/n7478 ), .force_11(1'b0), .Q(\shifter_0/n9321 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7481 ), .force_10(
        \shifter_0/n7482 ), .force_11(1'b0), .Q(\shifter_0/n9320 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7485 ), .force_10(
        \shifter_0/n7486 ), .force_11(1'b0), .Q(\shifter_0/n9319 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7489 ), .force_10(
        \shifter_0/n7490 ), .force_11(1'b0), .Q(\shifter_0/n9318 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7493 ), .force_10(
        \shifter_0/n7494 ), .force_11(1'b0), .Q(\shifter_0/n9317 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7497 ), .force_10(
        \shifter_0/n7498 ), .force_11(1'b0), .Q(\shifter_0/n9316 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7501 ), .force_10(
        \shifter_0/n7502 ), .force_11(1'b0), .Q(\shifter_0/n9315 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7505 ), .force_10(
        \shifter_0/n7506 ), .force_11(1'b0), .Q(\shifter_0/n9314 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7509 ), .force_10(
        \shifter_0/n7510 ), .force_11(1'b0), .Q(\shifter_0/n9313 ) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7513 ), .force_10(
        \shifter_0/n7514 ), .force_11(1'b0), .Q(\shifter_0/n9312 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7517 ), .force_10(
        \shifter_0/n7518 ), .force_11(1'b0), .Q(\shifter_0/n9311 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7521 ), .force_10(
        \shifter_0/n7522 ), .force_11(1'b0), .Q(\shifter_0/n9310 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7525 ), .force_10(
        \shifter_0/n7526 ), .force_11(1'b0), .Q(\shifter_0/n9309 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7529 ), .force_10(
        \shifter_0/n7530 ), .force_11(1'b0), .Q(\shifter_0/n9308 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7533 ), .force_10(
        \shifter_0/n7534 ), .force_11(1'b0), .Q(\shifter_0/n9307 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7537 ), .force_10(
        \shifter_0/n7538 ), .force_11(1'b0), .Q(\shifter_0/n9306 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7541 ), .force_10(
        \shifter_0/n7542 ), .force_11(1'b0), .Q(\shifter_0/n9305 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7545 ), .force_10(
        \shifter_0/n7546 ), .force_11(1'b0), .Q(\shifter_0/n9304 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7549 ), .force_10(
        \shifter_0/n7550 ), .force_11(1'b0), .Q(\shifter_0/n9303 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7553 ), .force_10(
        \shifter_0/n7554 ), .force_11(1'b0), .Q(\shifter_0/n9302 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7557 ), .force_10(
        \shifter_0/n7558 ), .force_11(1'b0), .Q(\shifter_0/n9301 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7561 ), .force_10(
        \shifter_0/n7562 ), .force_11(1'b0), .Q(\shifter_0/n9300 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7565 ), .force_10(
        \shifter_0/n7566 ), .force_11(1'b0), .Q(\shifter_0/n9299 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7569 ), .force_10(
        \shifter_0/n7570 ), .force_11(1'b0), .Q(\shifter_0/n9298 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7573 ), .force_10(
        \shifter_0/n7574 ), .force_11(1'b0), .Q(\shifter_0/n9297 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7577 ), .force_10(
        \shifter_0/n7578 ), .force_11(1'b0), .Q(\shifter_0/n9296 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7581 ), .force_10(
        \shifter_0/n7582 ), .force_11(1'b0), .Q(\shifter_0/n9295 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7585 ), .force_10(
        \shifter_0/n7586 ), .force_11(1'b0), .Q(\shifter_0/n9294 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7589 ), .force_10(
        \shifter_0/n7590 ), .force_11(1'b0), .Q(\shifter_0/n9293 ) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7593 ), .force_10(
        \shifter_0/n7594 ), .force_11(1'b0), .Q(\shifter_0/n9292 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7597 ), .force_10(
        \shifter_0/n7598 ), .force_11(1'b0), .Q(\shifter_0/n9291 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7601 ), .force_10(
        \shifter_0/n7602 ), .force_11(1'b0), .Q(\shifter_0/n9290 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7605 ), .force_10(
        \shifter_0/n7606 ), .force_11(1'b0), .Q(\shifter_0/n9289 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7609 ), .force_10(
        \shifter_0/n7610 ), .force_11(1'b0), .Q(\shifter_0/n9288 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7613 ), .force_10(
        \shifter_0/n7614 ), .force_11(1'b0), .Q(\shifter_0/n9287 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7617 ), .force_10(
        \shifter_0/n7618 ), .force_11(1'b0), .Q(\shifter_0/n9286 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7621 ), .force_10(
        \shifter_0/n7622 ), .force_11(1'b0), .Q(\shifter_0/n9285 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7625 ), .force_10(
        \shifter_0/n7626 ), .force_11(1'b0), .Q(\shifter_0/n9284 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7629 ), .force_10(
        \shifter_0/n7630 ), .force_11(1'b0), .Q(\shifter_0/n9283 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7633 ), .force_10(
        \shifter_0/n7634 ), .force_11(1'b0), .Q(\shifter_0/n9282 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7637 ), .force_10(
        \shifter_0/n7638 ), .force_11(1'b0), .Q(\shifter_0/n9281 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7641 ), .force_10(
        \shifter_0/n7642 ), .force_11(1'b0), .Q(\shifter_0/n9280 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7645 ), .force_10(
        \shifter_0/n7646 ), .force_11(1'b0), .Q(\shifter_0/n9279 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7649 ), .force_10(
        \shifter_0/n7650 ), .force_11(1'b0), .Q(\shifter_0/n9278 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7653 ), .force_10(
        \shifter_0/n7654 ), .force_11(1'b0), .Q(\shifter_0/n9277 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7657 ), .force_10(
        \shifter_0/n7658 ), .force_11(1'b0), .Q(\shifter_0/n9276 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7661 ), .force_10(
        \shifter_0/n7662 ), .force_11(1'b0), .Q(\shifter_0/n9275 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7665 ), .force_10(
        \shifter_0/n7666 ), .force_11(1'b0), .Q(\shifter_0/n9274 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7669 ), .force_10(
        \shifter_0/n7670 ), .force_11(1'b0), .Q(\shifter_0/n9273 ) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7673 ), .force_10(
        \shifter_0/n7674 ), .force_11(1'b0), .Q(\shifter_0/n9272 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7677 ), .force_10(
        \shifter_0/n7678 ), .force_11(1'b0), .Q(\shifter_0/n9271 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7681 ), .force_10(
        \shifter_0/n7682 ), .force_11(1'b0), .Q(\shifter_0/n9270 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7685 ), .force_10(
        \shifter_0/n7686 ), .force_11(1'b0), .Q(\shifter_0/n9269 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7689 ), .force_10(
        \shifter_0/n7690 ), .force_11(1'b0), .Q(\shifter_0/n9268 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7693 ), .force_10(
        \shifter_0/n7694 ), .force_11(1'b0), .Q(\shifter_0/n9267 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7697 ), .force_10(
        \shifter_0/n7698 ), .force_11(1'b0), .Q(\shifter_0/n9266 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7701 ), .force_10(
        \shifter_0/n7702 ), .force_11(1'b0), .Q(\shifter_0/n9265 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7705 ), .force_10(
        \shifter_0/n7706 ), .force_11(1'b0), .Q(\shifter_0/n9264 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7709 ), .force_10(
        \shifter_0/n7710 ), .force_11(1'b0), .Q(\shifter_0/n9263 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7713 ), .force_10(
        \shifter_0/n7714 ), .force_11(1'b0), .Q(\shifter_0/n9262 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7717 ), .force_10(
        \shifter_0/n7718 ), .force_11(1'b0), .Q(\shifter_0/n9261 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7721 ), .force_10(
        \shifter_0/n7722 ), .force_11(1'b0), .Q(\shifter_0/n9260 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7725 ), .force_10(
        \shifter_0/n7726 ), .force_11(1'b0), .Q(\shifter_0/n9259 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7729 ), .force_10(
        \shifter_0/n7730 ), .force_11(1'b0), .Q(\shifter_0/n9258 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7733 ), .force_10(
        \shifter_0/n7734 ), .force_11(1'b0), .Q(\shifter_0/n9257 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7737 ), .force_10(
        \shifter_0/n7738 ), .force_11(1'b0), .Q(\shifter_0/n9256 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7741 ), .force_10(
        \shifter_0/n7742 ), .force_11(1'b0), .Q(\shifter_0/n9255 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7745 ), .force_10(
        \shifter_0/n7746 ), .force_11(1'b0), .Q(\shifter_0/n9254 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7749 ), .force_10(
        \shifter_0/n7750 ), .force_11(1'b0), .Q(\shifter_0/n9253 ) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7753 ), .force_10(
        \shifter_0/n7754 ), .force_11(1'b0), .Q(\shifter_0/n9252 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7757 ), .force_10(
        \shifter_0/n7758 ), .force_11(1'b0), .Q(\shifter_0/n9251 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7761 ), .force_10(
        \shifter_0/n7762 ), .force_11(1'b0), .Q(\shifter_0/n9250 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7765 ), .force_10(
        \shifter_0/n7766 ), .force_11(1'b0), .Q(\shifter_0/n9249 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7769 ), .force_10(
        \shifter_0/n7770 ), .force_11(1'b0), .Q(\shifter_0/n9248 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7773 ), .force_10(
        \shifter_0/n7774 ), .force_11(1'b0), .Q(\shifter_0/n9247 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7777 ), .force_10(
        \shifter_0/n7778 ), .force_11(1'b0), .Q(\shifter_0/n9246 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7781 ), .force_10(
        \shifter_0/n7782 ), .force_11(1'b0), .Q(\shifter_0/n9245 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7785 ), .force_10(
        \shifter_0/n7786 ), .force_11(1'b0), .Q(\shifter_0/n9244 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7789 ), .force_10(
        \shifter_0/n7790 ), .force_11(1'b0), .Q(\shifter_0/n9243 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7793 ), .force_10(
        \shifter_0/n7794 ), .force_11(1'b0), .Q(\shifter_0/n9242 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7797 ), .force_10(
        \shifter_0/n7798 ), .force_11(1'b0), .Q(\shifter_0/n9241 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7801 ), .force_10(
        \shifter_0/n7802 ), .force_11(1'b0), .Q(\shifter_0/n9240 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7805 ), .force_10(
        \shifter_0/n7806 ), .force_11(1'b0), .Q(\shifter_0/n9239 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7809 ), .force_10(
        \shifter_0/n7810 ), .force_11(1'b0), .Q(\shifter_0/n9238 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7813 ), .force_10(
        \shifter_0/n7814 ), .force_11(1'b0), .Q(\shifter_0/n9237 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7817 ), .force_10(
        \shifter_0/n7818 ), .force_11(1'b0), .Q(\shifter_0/n9236 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7821 ), .force_10(
        \shifter_0/n7822 ), .force_11(1'b0), .Q(\shifter_0/n9235 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7825 ), .force_10(
        \shifter_0/n7826 ), .force_11(1'b0), .Q(\shifter_0/n9234 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7829 ), .force_10(
        \shifter_0/n7830 ), .force_11(1'b0), .Q(\shifter_0/n9233 ) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7833 ), .force_10(
        \shifter_0/n7834 ), .force_11(1'b0), .Q(\shifter_0/n9232 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7837 ), .force_10(
        \shifter_0/n7838 ), .force_11(1'b0), .Q(\shifter_0/n9231 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7841 ), .force_10(
        \shifter_0/n7842 ), .force_11(1'b0), .Q(\shifter_0/n9230 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7845 ), .force_10(
        \shifter_0/n7846 ), .force_11(1'b0), .Q(\shifter_0/n9229 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7849 ), .force_10(
        \shifter_0/n7850 ), .force_11(1'b0), .Q(\shifter_0/n9228 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7853 ), .force_10(
        \shifter_0/n7854 ), .force_11(1'b0), .Q(\shifter_0/n9227 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7857 ), .force_10(
        \shifter_0/n7858 ), .force_11(1'b0), .Q(\shifter_0/n9226 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7861 ), .force_10(
        \shifter_0/n7862 ), .force_11(1'b0), .Q(\shifter_0/n9225 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7865 ), .force_10(
        \shifter_0/n7866 ), .force_11(1'b0), .Q(\shifter_0/n9224 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7869 ), .force_10(
        \shifter_0/n7870 ), .force_11(1'b0), .Q(\shifter_0/n9223 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7873 ), .force_10(
        \shifter_0/n7874 ), .force_11(1'b0), .Q(\shifter_0/n9222 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7877 ), .force_10(
        \shifter_0/n7878 ), .force_11(1'b0), .Q(\shifter_0/n9221 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7881 ), .force_10(
        \shifter_0/n7882 ), .force_11(1'b0), .Q(\shifter_0/n9220 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7885 ), .force_10(
        \shifter_0/n7886 ), .force_11(1'b0), .Q(\shifter_0/n9219 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7889 ), .force_10(
        \shifter_0/n7890 ), .force_11(1'b0), .Q(\shifter_0/n9218 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7893 ), .force_10(
        \shifter_0/n7894 ), .force_11(1'b0), .Q(\shifter_0/n9217 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7897 ), .force_10(
        \shifter_0/n7898 ), .force_11(1'b0), .Q(\shifter_0/n9216 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7901 ), .force_10(
        \shifter_0/n7902 ), .force_11(1'b0), .Q(\shifter_0/n9215 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7905 ), .force_10(
        \shifter_0/n7906 ), .force_11(1'b0), .Q(\shifter_0/n9214 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7909 ), .force_10(
        \shifter_0/n7910 ), .force_11(1'b0), .Q(\shifter_0/n9213 ) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7913 ), .force_10(
        \shifter_0/n7914 ), .force_11(1'b0), .Q(\shifter_0/n9212 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7917 ), .force_10(n41664), .force_11(1'b0), .Q(\shifter_0/n9211 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7921 ), .force_10(n41663), .force_11(1'b0), .Q(\shifter_0/n9210 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7925 ), .force_10(n41662), .force_11(1'b0), .Q(\shifter_0/n9209 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7929 ), .force_10(n41661), .force_11(1'b0), .Q(\shifter_0/n9208 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7933 ), .force_10(n41660), .force_11(1'b0), .Q(\shifter_0/n9207 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7937 ), .force_10(n41659), .force_11(1'b0), .Q(\shifter_0/n9206 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7941 ), .force_10(n41658), .force_11(1'b0), .Q(\shifter_0/n9205 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7945 ), .force_10(n41657), .force_11(1'b0), .Q(\shifter_0/n9204 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7949 ), .force_10(n41656), .force_11(1'b0), .Q(\shifter_0/n9203 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7953 ), .force_10(n41655), .force_11(1'b0), .Q(\shifter_0/n9202 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7957 ), .force_10(n41654), .force_11(1'b0), .Q(\shifter_0/n9201 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7961 ), .force_10(n41653), .force_11(1'b0), .Q(\shifter_0/n9200 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7965 ), .force_10(n41652), .force_11(1'b0), .Q(\shifter_0/n9199 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7969 ), .force_10(n41651), .force_11(1'b0), .Q(\shifter_0/n9198 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7973 ), .force_10(n41650), .force_11(1'b0), .Q(\shifter_0/n9197 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7977 ), .force_10(n41649), .force_11(1'b0), .Q(\shifter_0/n9196 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7981 ), .force_10(n41648), .force_11(1'b0), .Q(\shifter_0/n9195 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7985 ), .force_10(n41647), .force_11(1'b0), .Q(\shifter_0/n9194 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7989 ), .force_10(n41646), .force_11(1'b0), .Q(\shifter_0/n9193 ) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7993 ), .force_10(n41645), .force_11(1'b0), .Q(\shifter_0/n9192 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n7997 ), .force_10(n41519), .force_11(1'b0), .Q(\shifter_0/n9191 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8001 ), .force_10(n41518), .force_11(1'b0), .Q(\shifter_0/n9190 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8005 ), .force_10(n41517), .force_11(1'b0), .Q(\shifter_0/n9189 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8009 ), .force_10(n41516), .force_11(1'b0), .Q(\shifter_0/n9188 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8013 ), .force_10(n41515), .force_11(1'b0), .Q(\shifter_0/n9187 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8017 ), .force_10(n41514), .force_11(1'b0), .Q(\shifter_0/n9186 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8021 ), .force_10(n41513), .force_11(1'b0), .Q(\shifter_0/n9185 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8025 ), .force_10(n41512), .force_11(1'b0), .Q(\shifter_0/n9184 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8029 ), .force_10(n41511), .force_11(1'b0), .Q(\shifter_0/n9183 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8033 ), .force_10(n41510), .force_11(1'b0), .Q(\shifter_0/n9182 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8037 ), .force_10(n41509), .force_11(1'b0), .Q(\shifter_0/n9181 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8041 ), .force_10(n41508), .force_11(1'b0), .Q(\shifter_0/n9180 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8045 ), .force_10(n41507), .force_11(1'b0), .Q(\shifter_0/n9179 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8049 ), .force_10(n41506), .force_11(1'b0), .Q(\shifter_0/n9178 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8053 ), .force_10(n41505), .force_11(1'b0), .Q(\shifter_0/n9177 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8057 ), .force_10(n41504), .force_11(1'b0), .Q(\shifter_0/n9176 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8061 ), .force_10(n41503), .force_11(1'b0), .Q(\shifter_0/n9175 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8065 ), .force_10(n41502), .force_11(1'b0), .Q(\shifter_0/n9174 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8069 ), .force_10(n41501), .force_11(1'b0), .Q(\shifter_0/n9173 ) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8073 ), .force_10(n41500), .force_11(1'b0), .Q(\shifter_0/n9172 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8077 ), .force_10(
        \shifter_0/n8078 ), .force_11(1'b0), .Q(\shifter_0/n9171 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8081 ), .force_10(
        \shifter_0/n8082 ), .force_11(1'b0), .Q(\shifter_0/n9170 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8085 ), .force_10(
        \shifter_0/n8086 ), .force_11(1'b0), .Q(\shifter_0/n9169 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8089 ), .force_10(
        \shifter_0/n8090 ), .force_11(1'b0), .Q(\shifter_0/n9168 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8093 ), .force_10(
        \shifter_0/n8094 ), .force_11(1'b0), .Q(\shifter_0/n9167 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8097 ), .force_10(
        \shifter_0/n8098 ), .force_11(1'b0), .Q(\shifter_0/n9166 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8101 ), .force_10(
        \shifter_0/n8102 ), .force_11(1'b0), .Q(\shifter_0/n9165 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8105 ), .force_10(
        \shifter_0/n8106 ), .force_11(1'b0), .Q(\shifter_0/n9164 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8109 ), .force_10(
        \shifter_0/n8110 ), .force_11(1'b0), .Q(\shifter_0/n9163 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8113 ), .force_10(
        \shifter_0/n8114 ), .force_11(1'b0), .Q(\shifter_0/n9162 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8117 ), .force_10(
        \shifter_0/n8118 ), .force_11(1'b0), .Q(\shifter_0/n9161 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8121 ), .force_10(
        \shifter_0/n8122 ), .force_11(1'b0), .Q(\shifter_0/n9160 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8125 ), .force_10(
        \shifter_0/n8126 ), .force_11(1'b0), .Q(\shifter_0/n9159 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8129 ), .force_10(
        \shifter_0/n8130 ), .force_11(1'b0), .Q(\shifter_0/n9158 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8133 ), .force_10(
        \shifter_0/n8134 ), .force_11(1'b0), .Q(\shifter_0/n9157 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8137 ), .force_10(
        \shifter_0/n8138 ), .force_11(1'b0), .Q(\shifter_0/n9156 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8141 ), .force_10(
        \shifter_0/n8142 ), .force_11(1'b0), .Q(\shifter_0/n9155 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8145 ), .force_10(
        \shifter_0/n8146 ), .force_11(1'b0), .Q(\shifter_0/n9154 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8149 ), .force_10(
        \shifter_0/n8150 ), .force_11(1'b0), .Q(\shifter_0/n9153 ) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8153 ), .force_10(
        \shifter_0/n8154 ), .force_11(1'b0), .Q(\shifter_0/n9152 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8157 ), .force_10(
        \shifter_0/n8158 ), .force_11(1'b0), .Q(\shifter_0/n9151 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8161 ), .force_10(
        \shifter_0/n8162 ), .force_11(1'b0), .Q(\shifter_0/n9150 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8165 ), .force_10(
        \shifter_0/n8166 ), .force_11(1'b0), .Q(\shifter_0/n9149 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8169 ), .force_10(
        \shifter_0/n8170 ), .force_11(1'b0), .Q(\shifter_0/n9148 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8173 ), .force_10(
        \shifter_0/n8174 ), .force_11(1'b0), .Q(\shifter_0/n9147 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8177 ), .force_10(
        \shifter_0/n8178 ), .force_11(1'b0), .Q(\shifter_0/n9146 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8181 ), .force_10(
        \shifter_0/n8182 ), .force_11(1'b0), .Q(\shifter_0/n9145 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8185 ), .force_10(
        \shifter_0/n8186 ), .force_11(1'b0), .Q(\shifter_0/n9144 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8189 ), .force_10(
        \shifter_0/n8190 ), .force_11(1'b0), .Q(\shifter_0/n9143 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8193 ), .force_10(
        \shifter_0/n8194 ), .force_11(1'b0), .Q(\shifter_0/n9142 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8197 ), .force_10(
        \shifter_0/n8198 ), .force_11(1'b0), .Q(\shifter_0/n9141 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8201 ), .force_10(
        \shifter_0/n8202 ), .force_11(1'b0), .Q(\shifter_0/n9140 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8205 ), .force_10(
        \shifter_0/n8206 ), .force_11(1'b0), .Q(\shifter_0/n9139 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8209 ), .force_10(
        \shifter_0/n8210 ), .force_11(1'b0), .Q(\shifter_0/n9138 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8213 ), .force_10(
        \shifter_0/n8214 ), .force_11(1'b0), .Q(\shifter_0/n9137 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8217 ), .force_10(
        \shifter_0/n8218 ), .force_11(1'b0), .Q(\shifter_0/n9136 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8221 ), .force_10(
        \shifter_0/n8222 ), .force_11(1'b0), .Q(\shifter_0/n9135 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8225 ), .force_10(
        \shifter_0/n8226 ), .force_11(1'b0), .Q(\shifter_0/n9134 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8229 ), .force_10(
        \shifter_0/n8230 ), .force_11(1'b0), .Q(\shifter_0/n9133 ) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8233 ), .force_10(
        \shifter_0/n8234 ), .force_11(1'b0), .Q(\shifter_0/n9132 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8237 ), .force_10(
        \shifter_0/n8238 ), .force_11(1'b0), .Q(\shifter_0/n9131 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8241 ), .force_10(
        \shifter_0/n8242 ), .force_11(1'b0), .Q(\shifter_0/n9130 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8245 ), .force_10(
        \shifter_0/n8246 ), .force_11(1'b0), .Q(\shifter_0/n9129 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8249 ), .force_10(
        \shifter_0/n8250 ), .force_11(1'b0), .Q(\shifter_0/n9128 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8253 ), .force_10(
        \shifter_0/n8254 ), .force_11(1'b0), .Q(\shifter_0/n9127 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8257 ), .force_10(
        \shifter_0/n8258 ), .force_11(1'b0), .Q(\shifter_0/n9126 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8261 ), .force_10(
        \shifter_0/n8262 ), .force_11(1'b0), .Q(\shifter_0/n9125 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8265 ), .force_10(
        \shifter_0/n8266 ), .force_11(1'b0), .Q(\shifter_0/n9124 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8269 ), .force_10(
        \shifter_0/n8270 ), .force_11(1'b0), .Q(\shifter_0/n9123 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8273 ), .force_10(
        \shifter_0/n8274 ), .force_11(1'b0), .Q(\shifter_0/n9122 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8277 ), .force_10(
        \shifter_0/n8278 ), .force_11(1'b0), .Q(\shifter_0/n9121 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8281 ), .force_10(
        \shifter_0/n8282 ), .force_11(1'b0), .Q(\shifter_0/n9120 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8285 ), .force_10(
        \shifter_0/n8286 ), .force_11(1'b0), .Q(\shifter_0/n9119 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8289 ), .force_10(
        \shifter_0/n8290 ), .force_11(1'b0), .Q(\shifter_0/n9118 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8293 ), .force_10(
        \shifter_0/n8294 ), .force_11(1'b0), .Q(\shifter_0/n9117 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8297 ), .force_10(
        \shifter_0/n8298 ), .force_11(1'b0), .Q(\shifter_0/n9116 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8301 ), .force_10(
        \shifter_0/n8302 ), .force_11(1'b0), .Q(\shifter_0/n9115 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8305 ), .force_10(
        \shifter_0/n8306 ), .force_11(1'b0), .Q(\shifter_0/n9114 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8309 ), .force_10(
        \shifter_0/n8310 ), .force_11(1'b0), .Q(\shifter_0/n9113 ) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8313 ), .force_10(
        \shifter_0/n8314 ), .force_11(1'b0), .Q(\shifter_0/n9112 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8317 ), .force_10(
        \shifter_0/n8318 ), .force_11(1'b0), .Q(\shifter_0/n9111 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8321 ), .force_10(
        \shifter_0/n8322 ), .force_11(1'b0), .Q(\shifter_0/n9110 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8325 ), .force_10(
        \shifter_0/n8326 ), .force_11(1'b0), .Q(\shifter_0/n9109 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8329 ), .force_10(
        \shifter_0/n8330 ), .force_11(1'b0), .Q(\shifter_0/n9108 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8333 ), .force_10(
        \shifter_0/n8334 ), .force_11(1'b0), .Q(\shifter_0/n9107 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8337 ), .force_10(
        \shifter_0/n8338 ), .force_11(1'b0), .Q(\shifter_0/n9106 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8341 ), .force_10(
        \shifter_0/n8342 ), .force_11(1'b0), .Q(\shifter_0/n9105 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8345 ), .force_10(
        \shifter_0/n8346 ), .force_11(1'b0), .Q(\shifter_0/n9104 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8349 ), .force_10(
        \shifter_0/n8350 ), .force_11(1'b0), .Q(\shifter_0/n9103 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8353 ), .force_10(
        \shifter_0/n8354 ), .force_11(1'b0), .Q(\shifter_0/n9102 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8357 ), .force_10(
        \shifter_0/n8358 ), .force_11(1'b0), .Q(\shifter_0/n9101 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8361 ), .force_10(
        \shifter_0/n8362 ), .force_11(1'b0), .Q(\shifter_0/n9100 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8365 ), .force_10(
        \shifter_0/n8366 ), .force_11(1'b0), .Q(\shifter_0/n9099 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8369 ), .force_10(
        \shifter_0/n8370 ), .force_11(1'b0), .Q(\shifter_0/n9098 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8373 ), .force_10(
        \shifter_0/n8374 ), .force_11(1'b0), .Q(\shifter_0/n9097 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8377 ), .force_10(
        \shifter_0/n8378 ), .force_11(1'b0), .Q(\shifter_0/n9096 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8381 ), .force_10(
        \shifter_0/n8382 ), .force_11(1'b0), .Q(\shifter_0/n9095 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8385 ), .force_10(
        \shifter_0/n8386 ), .force_11(1'b0), .Q(\shifter_0/n9094 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8389 ), .force_10(
        \shifter_0/n8390 ), .force_11(1'b0), .Q(\shifter_0/n9093 ) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8393 ), .force_10(
        \shifter_0/n8394 ), .force_11(1'b0), .Q(\shifter_0/n9092 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8397 ), .force_10(
        \shifter_0/n8398 ), .force_11(1'b0), .Q(\shifter_0/n9091 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8401 ), .force_10(
        \shifter_0/n8402 ), .force_11(1'b0), .Q(\shifter_0/n9090 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8405 ), .force_10(
        \shifter_0/n8406 ), .force_11(1'b0), .Q(\shifter_0/n9089 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8409 ), .force_10(
        \shifter_0/n8410 ), .force_11(1'b0), .Q(\shifter_0/n9088 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8413 ), .force_10(
        \shifter_0/n8414 ), .force_11(1'b0), .Q(\shifter_0/n9087 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8417 ), .force_10(
        \shifter_0/n8418 ), .force_11(1'b0), .Q(\shifter_0/n9086 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8421 ), .force_10(
        \shifter_0/n8422 ), .force_11(1'b0), .Q(\shifter_0/n9085 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8425 ), .force_10(
        \shifter_0/n8426 ), .force_11(1'b0), .Q(\shifter_0/n9084 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8429 ), .force_10(
        \shifter_0/n8430 ), .force_11(1'b0), .Q(\shifter_0/n9083 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8433 ), .force_10(
        \shifter_0/n8434 ), .force_11(1'b0), .Q(\shifter_0/n9082 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8437 ), .force_10(
        \shifter_0/n8438 ), .force_11(1'b0), .Q(\shifter_0/n9081 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8441 ), .force_10(
        \shifter_0/n8442 ), .force_11(1'b0), .Q(\shifter_0/n9080 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8445 ), .force_10(
        \shifter_0/n8446 ), .force_11(1'b0), .Q(\shifter_0/n9079 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8449 ), .force_10(
        \shifter_0/n8450 ), .force_11(1'b0), .Q(\shifter_0/n9078 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8453 ), .force_10(
        \shifter_0/n8454 ), .force_11(1'b0), .Q(\shifter_0/n9077 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8457 ), .force_10(
        \shifter_0/n8458 ), .force_11(1'b0), .Q(\shifter_0/n9076 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8461 ), .force_10(
        \shifter_0/n8462 ), .force_11(1'b0), .Q(\shifter_0/n9075 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8465 ), .force_10(
        \shifter_0/n8466 ), .force_11(1'b0), .Q(\shifter_0/n9074 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8469 ), .force_10(
        \shifter_0/n8470 ), .force_11(1'b0), .Q(\shifter_0/n9073 ) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8473 ), .force_10(
        \shifter_0/n8474 ), .force_11(1'b0), .Q(\shifter_0/n9072 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8477 ), .force_10(
        \shifter_0/n8478 ), .force_11(1'b0), .Q(\shifter_0/n9071 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8481 ), .force_10(
        \shifter_0/n8482 ), .force_11(1'b0), .Q(\shifter_0/n9070 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8485 ), .force_10(
        \shifter_0/n8486 ), .force_11(1'b0), .Q(\shifter_0/n9069 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8489 ), .force_10(
        \shifter_0/n8490 ), .force_11(1'b0), .Q(\shifter_0/n9068 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8493 ), .force_10(
        \shifter_0/n8494 ), .force_11(1'b0), .Q(\shifter_0/n9067 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8497 ), .force_10(
        \shifter_0/n8498 ), .force_11(1'b0), .Q(\shifter_0/n9066 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8501 ), .force_10(
        \shifter_0/n8502 ), .force_11(1'b0), .Q(\shifter_0/n9065 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8505 ), .force_10(
        \shifter_0/n8506 ), .force_11(1'b0), .Q(\shifter_0/n9064 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8509 ), .force_10(
        \shifter_0/n8510 ), .force_11(1'b0), .Q(\shifter_0/n9063 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8513 ), .force_10(
        \shifter_0/n8514 ), .force_11(1'b0), .Q(\shifter_0/n9062 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8517 ), .force_10(
        \shifter_0/n8518 ), .force_11(1'b0), .Q(\shifter_0/n9061 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8521 ), .force_10(
        \shifter_0/n8522 ), .force_11(1'b0), .Q(\shifter_0/n9060 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8525 ), .force_10(
        \shifter_0/n8526 ), .force_11(1'b0), .Q(\shifter_0/n9059 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8529 ), .force_10(
        \shifter_0/n8530 ), .force_11(1'b0), .Q(\shifter_0/n9058 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8533 ), .force_10(
        \shifter_0/n8534 ), .force_11(1'b0), .Q(\shifter_0/n9057 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8537 ), .force_10(
        \shifter_0/n8538 ), .force_11(1'b0), .Q(\shifter_0/n9056 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8541 ), .force_10(
        \shifter_0/n8542 ), .force_11(1'b0), .Q(\shifter_0/n9055 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8545 ), .force_10(
        \shifter_0/n8546 ), .force_11(1'b0), .Q(\shifter_0/n9054 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8549 ), .force_10(
        \shifter_0/n8550 ), .force_11(1'b0), .Q(\shifter_0/n9053 ) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8553 ), .force_10(
        \shifter_0/n8554 ), .force_11(1'b0), .Q(\shifter_0/n9052 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8557 ), .force_10(
        \shifter_0/n8558 ), .force_11(1'b0), .Q(\shifter_0/n9051 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8561 ), .force_10(
        \shifter_0/n8562 ), .force_11(1'b0), .Q(\shifter_0/n9050 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8565 ), .force_10(
        \shifter_0/n8566 ), .force_11(1'b0), .Q(\shifter_0/n9049 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8569 ), .force_10(
        \shifter_0/n8570 ), .force_11(1'b0), .Q(\shifter_0/n9048 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8573 ), .force_10(
        \shifter_0/n8574 ), .force_11(1'b0), .Q(\shifter_0/n9047 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8577 ), .force_10(
        \shifter_0/n8578 ), .force_11(1'b0), .Q(\shifter_0/n9046 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8581 ), .force_10(
        \shifter_0/n8582 ), .force_11(1'b0), .Q(\shifter_0/n9045 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8585 ), .force_10(
        \shifter_0/n8586 ), .force_11(1'b0), .Q(\shifter_0/n9044 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8589 ), .force_10(
        \shifter_0/n8590 ), .force_11(1'b0), .Q(\shifter_0/n9043 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8593 ), .force_10(
        \shifter_0/n8594 ), .force_11(1'b0), .Q(\shifter_0/n9042 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8597 ), .force_10(
        \shifter_0/n8598 ), .force_11(1'b0), .Q(\shifter_0/n9041 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8601 ), .force_10(
        \shifter_0/n8602 ), .force_11(1'b0), .Q(\shifter_0/n9040 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8605 ), .force_10(
        \shifter_0/n8606 ), .force_11(1'b0), .Q(\shifter_0/n9039 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8609 ), .force_10(
        \shifter_0/n8610 ), .force_11(1'b0), .Q(\shifter_0/n9038 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8613 ), .force_10(
        \shifter_0/n8614 ), .force_11(1'b0), .Q(\shifter_0/n9037 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8617 ), .force_10(
        \shifter_0/n8618 ), .force_11(1'b0), .Q(\shifter_0/n9036 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8621 ), .force_10(
        \shifter_0/n8622 ), .force_11(1'b0), .Q(\shifter_0/n9035 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8625 ), .force_10(
        \shifter_0/n8626 ), .force_11(1'b0), .Q(\shifter_0/n9034 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8629 ), .force_10(
        \shifter_0/n8630 ), .force_11(1'b0), .Q(\shifter_0/n9033 ) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8633 ), .force_10(
        \shifter_0/n8634 ), .force_11(1'b0), .Q(\shifter_0/n9032 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8637 ), .force_10(
        \shifter_0/n8638 ), .force_11(1'b0), .Q(\shifter_0/n9031 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8641 ), .force_10(
        \shifter_0/n8642 ), .force_11(1'b0), .Q(\shifter_0/n9030 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8645 ), .force_10(
        \shifter_0/n8646 ), .force_11(1'b0), .Q(\shifter_0/n9029 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8649 ), .force_10(
        \shifter_0/n8650 ), .force_11(1'b0), .Q(\shifter_0/n9028 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8653 ), .force_10(
        \shifter_0/n8654 ), .force_11(1'b0), .Q(\shifter_0/n9027 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8657 ), .force_10(
        \shifter_0/n8658 ), .force_11(1'b0), .Q(\shifter_0/n9026 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8661 ), .force_10(
        \shifter_0/n8662 ), .force_11(1'b0), .Q(\shifter_0/n9025 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8665 ), .force_10(
        \shifter_0/n8666 ), .force_11(1'b0), .Q(\shifter_0/n9024 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8669 ), .force_10(
        \shifter_0/n8670 ), .force_11(1'b0), .Q(\shifter_0/n9023 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8673 ), .force_10(
        \shifter_0/n8674 ), .force_11(1'b0), .Q(\shifter_0/n9022 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8677 ), .force_10(
        \shifter_0/n8678 ), .force_11(1'b0), .Q(\shifter_0/n9021 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8681 ), .force_10(
        \shifter_0/n8682 ), .force_11(1'b0), .Q(\shifter_0/n9020 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8685 ), .force_10(
        \shifter_0/n8686 ), .force_11(1'b0), .Q(\shifter_0/n9019 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8689 ), .force_10(
        \shifter_0/n8690 ), .force_11(1'b0), .Q(\shifter_0/n9018 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8693 ), .force_10(
        \shifter_0/n8694 ), .force_11(1'b0), .Q(\shifter_0/n9017 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8697 ), .force_10(
        \shifter_0/n8698 ), .force_11(1'b0), .Q(\shifter_0/n9016 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8701 ), .force_10(
        \shifter_0/n8702 ), .force_11(1'b0), .Q(\shifter_0/n9015 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8705 ), .force_10(
        \shifter_0/n8706 ), .force_11(1'b0), .Q(\shifter_0/n9014 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8709 ), .force_10(
        \shifter_0/n8710 ), .force_11(1'b0), .Q(\shifter_0/n9013 ) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8713 ), .force_10(
        \shifter_0/n8714 ), .force_11(1'b0), .Q(\shifter_0/n9012 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8717 ), .force_10(
        \shifter_0/n8718 ), .force_11(1'b0), .Q(\shifter_0/n9011 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8721 ), .force_10(
        \shifter_0/n8722 ), .force_11(1'b0), .Q(\shifter_0/n9010 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8725 ), .force_10(
        \shifter_0/n8726 ), .force_11(1'b0), .Q(\shifter_0/n9009 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8729 ), .force_10(
        \shifter_0/n8730 ), .force_11(1'b0), .Q(\shifter_0/n9008 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8733 ), .force_10(
        \shifter_0/n8734 ), .force_11(1'b0), .Q(\shifter_0/n9007 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8737 ), .force_10(
        \shifter_0/n8738 ), .force_11(1'b0), .Q(\shifter_0/n9006 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8741 ), .force_10(
        \shifter_0/n8742 ), .force_11(1'b0), .Q(\shifter_0/n9005 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8745 ), .force_10(
        \shifter_0/n8746 ), .force_11(1'b0), .Q(\shifter_0/n9004 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8749 ), .force_10(
        \shifter_0/n8750 ), .force_11(1'b0), .Q(\shifter_0/n9003 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8753 ), .force_10(
        \shifter_0/n8754 ), .force_11(1'b0), .Q(\shifter_0/n9002 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8757 ), .force_10(
        \shifter_0/n8758 ), .force_11(1'b0), .Q(\shifter_0/n9001 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8761 ), .force_10(
        \shifter_0/n8762 ), .force_11(1'b0), .Q(\shifter_0/n9000 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8765 ), .force_10(
        \shifter_0/n8766 ), .force_11(1'b0), .Q(\shifter_0/n8999 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8769 ), .force_10(
        \shifter_0/n8770 ), .force_11(1'b0), .Q(\shifter_0/n8998 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8773 ), .force_10(
        \shifter_0/n8774 ), .force_11(1'b0), .Q(\shifter_0/n8997 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8777 ), .force_10(
        \shifter_0/n8778 ), .force_11(1'b0), .Q(\shifter_0/n8996 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8781 ), .force_10(
        \shifter_0/n8782 ), .force_11(1'b0), .Q(\shifter_0/n8995 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8785 ), .force_10(
        \shifter_0/n8786 ), .force_11(1'b0), .Q(\shifter_0/n8994 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8789 ), .force_10(
        \shifter_0/n8790 ), .force_11(1'b0), .Q(\shifter_0/n8993 ) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8793 ), .force_10(
        \shifter_0/n8794 ), .force_11(1'b0), .Q(\shifter_0/n8992 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8797 ), .force_10(
        \shifter_0/n8798 ), .force_11(1'b0), .Q(\shifter_0/n8991 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8801 ), .force_10(
        \shifter_0/n8802 ), .force_11(1'b0), .Q(\shifter_0/n8990 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8805 ), .force_10(
        \shifter_0/n8806 ), .force_11(1'b0), .Q(\shifter_0/n8989 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8809 ), .force_10(
        \shifter_0/n8810 ), .force_11(1'b0), .Q(\shifter_0/n8988 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8813 ), .force_10(
        \shifter_0/n8814 ), .force_11(1'b0), .Q(\shifter_0/n8987 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8817 ), .force_10(
        \shifter_0/n8818 ), .force_11(1'b0), .Q(\shifter_0/n8986 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8821 ), .force_10(
        \shifter_0/n8822 ), .force_11(1'b0), .Q(\shifter_0/n8985 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8825 ), .force_10(
        \shifter_0/n8826 ), .force_11(1'b0), .Q(\shifter_0/n8984 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8829 ), .force_10(
        \shifter_0/n8830 ), .force_11(1'b0), .Q(\shifter_0/n8983 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8833 ), .force_10(
        \shifter_0/n8834 ), .force_11(1'b0), .Q(\shifter_0/n8982 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8837 ), .force_10(
        \shifter_0/n8838 ), .force_11(1'b0), .Q(\shifter_0/n8981 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8841 ), .force_10(
        \shifter_0/n8842 ), .force_11(1'b0), .Q(\shifter_0/n8980 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8845 ), .force_10(
        \shifter_0/n8846 ), .force_11(1'b0), .Q(\shifter_0/n8979 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8849 ), .force_10(
        \shifter_0/n8850 ), .force_11(1'b0), .Q(\shifter_0/n8978 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8853 ), .force_10(
        \shifter_0/n8854 ), .force_11(1'b0), .Q(\shifter_0/n8977 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8857 ), .force_10(
        \shifter_0/n8858 ), .force_11(1'b0), .Q(\shifter_0/n8976 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8861 ), .force_10(
        \shifter_0/n8862 ), .force_11(1'b0), .Q(\shifter_0/n8975 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8865 ), .force_10(
        \shifter_0/n8866 ), .force_11(1'b0), .Q(\shifter_0/n8974 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8869 ), .force_10(
        \shifter_0/n8870 ), .force_11(1'b0), .Q(\shifter_0/n8973 ) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8873 ), .force_10(
        \shifter_0/n8874 ), .force_11(1'b0), .Q(\shifter_0/n8972 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8877 ), .force_10(
        \shifter_0/n8878 ), .force_11(1'b0), .Q(\shifter_0/n8971 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8881 ), .force_10(
        \shifter_0/n8882 ), .force_11(1'b0), .Q(\shifter_0/n8970 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8885 ), .force_10(
        \shifter_0/n8886 ), .force_11(1'b0), .Q(\shifter_0/n8969 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8889 ), .force_10(
        \shifter_0/n8890 ), .force_11(1'b0), .Q(\shifter_0/n8968 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8893 ), .force_10(
        \shifter_0/n8894 ), .force_11(1'b0), .Q(\shifter_0/n8967 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8897 ), .force_10(
        \shifter_0/n8898 ), .force_11(1'b0), .Q(\shifter_0/n8966 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8901 ), .force_10(
        \shifter_0/n8902 ), .force_11(1'b0), .Q(\shifter_0/n8965 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8905 ), .force_10(
        \shifter_0/n8906 ), .force_11(1'b0), .Q(\shifter_0/n8964 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8909 ), .force_10(
        \shifter_0/n8910 ), .force_11(1'b0), .Q(\shifter_0/n8963 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8913 ), .force_10(
        \shifter_0/n8914 ), .force_11(1'b0), .Q(\shifter_0/n8962 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8917 ), .force_10(
        \shifter_0/n8918 ), .force_11(1'b0), .Q(\shifter_0/n8961 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8921 ), .force_10(
        \shifter_0/n8922 ), .force_11(1'b0), .Q(\shifter_0/n8960 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8925 ), .force_10(
        \shifter_0/n8926 ), .force_11(1'b0), .Q(\shifter_0/n8959 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8929 ), .force_10(
        \shifter_0/n8930 ), .force_11(1'b0), .Q(\shifter_0/n8958 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8933 ), .force_10(
        \shifter_0/n8934 ), .force_11(1'b0), .Q(\shifter_0/n8957 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8937 ), .force_10(
        \shifter_0/n8938 ), .force_11(1'b0), .Q(\shifter_0/n8956 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8941 ), .force_10(
        \shifter_0/n8942 ), .force_11(1'b0), .Q(\shifter_0/n8955 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8945 ), .force_10(
        \shifter_0/n8946 ), .force_11(1'b0), .Q(\shifter_0/n8954 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n8949 ), .force_10(
        \shifter_0/n8950 ), .force_11(1'b0), .Q(\shifter_0/n8953 ) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n6393 ), .force_10(
        \shifter_0/n6394 ), .force_11(1'b0), .Q(\shifter_0/n8952 ) );
  nand_x1_sg U35199 ( .A(n11840), .B(n11841), .X(n35654) );
  nand_x1_sg U35200 ( .A(n11842), .B(n11612), .X(n11841) );
  nand_x1_sg U35201 ( .A(n13091), .B(n13092), .X(n35643) );
  nand_x1_sg U35202 ( .A(n11888), .B(n11889), .X(n35652) );
  nand_x1_sg U35203 ( .A(n12962), .B(n12963), .X(n12842) );
  inv_x1_sg U35204 ( .A(n12448), .X(n41139) );
  inv_x1_sg U35205 ( .A(n12457), .X(n41140) );
  inv_x1_sg U35206 ( .A(n12510), .X(n41141) );
  inv_x1_sg U35207 ( .A(n12515), .X(n41142) );
  nand_x1_sg U35208 ( .A(n13287), .B(n13288), .X(n35639) );
  nand_x1_sg U35209 ( .A(n13483), .B(n13484), .X(n35620) );
  nand_x1_sg U35210 ( .A(n13696), .B(n13697), .X(n35637) );
  nand_x1_sg U35211 ( .A(n13778), .B(n13779), .X(n35636) );
  nand_x1_sg U35212 ( .A(n35463), .B(n21370), .X(n21326) );
  nand_x2_sg U35213 ( .A(n15299), .B(n15300), .X(n15298) );
  nand_x1_sg U35214 ( .A(n21189), .B(n21190), .X(n20988) );
  nand_x1_sg U35215 ( .A(n21229), .B(n21230), .X(n20997) );
  nand_x1_sg U35216 ( .A(n21247), .B(n21248), .X(n20998) );
  nand_x1_sg U35217 ( .A(n21285), .B(n21286), .X(n21002) );
  nand_x1_sg U35218 ( .A(n21091), .B(n21092), .X(n20977) );
  nand_x1_sg U35219 ( .A(n21109), .B(n21110), .X(n20978) );
  nand_x1_sg U35220 ( .A(n21147), .B(n21148), .X(n20982) );
  nand_x1_sg U35221 ( .A(n21012), .B(n21013), .X(n20966) );
  nand_x1_sg U35222 ( .A(n21030), .B(n21031), .X(n20967) );
  nand_x1_sg U35223 ( .A(n21068), .B(n21069), .X(n20972) );
  nand_x1_sg U35224 ( .A(n21689), .B(n21690), .X(n21662) );
  nand_x1_sg U35225 ( .A(n21600), .B(n21601), .X(n21571) );
  nand_x1_sg U35226 ( .A(n21582), .B(n21583), .X(n21570) );
  nand_x1_sg U35227 ( .A(n21638), .B(n21639), .X(n21575) );
  nand_x1_sg U35228 ( .A(n21413), .B(n21414), .X(n21384) );
  nand_x1_sg U35229 ( .A(n21395), .B(n21396), .X(n21383) );
  nand_x1_sg U35230 ( .A(n21451), .B(n21452), .X(n21388) );
  nand_x1_sg U35231 ( .A(n21505), .B(n21506), .X(n21477) );
  nand_x1_sg U35232 ( .A(n21487), .B(n21488), .X(n21476) );
  nand_x1_sg U35233 ( .A(n21543), .B(n21544), .X(n21481) );
  nand_x2_sg U35234 ( .A(n15315), .B(n15316), .X(n15314) );
  nand_x1_sg U35235 ( .A(n21168), .B(n21169), .X(n20991) );
  nand_x1_sg U35236 ( .A(n21207), .B(n21208), .X(n20992) );
  nand_x1_sg U35237 ( .A(n20988), .B(n31695), .X(n20987) );
  nand_x1_sg U35238 ( .A(n21267), .B(n21268), .X(n21001) );
  nand_x1_sg U35239 ( .A(n21050), .B(n21051), .X(n20971) );
  nand_x1_sg U35240 ( .A(n21129), .B(n21130), .X(n20981) );
  nand_x1_sg U35241 ( .A(n21668), .B(n21669), .X(n21665) );
  nand_x1_sg U35242 ( .A(n21707), .B(n21708), .X(n21666) );
  nand_x1_sg U35243 ( .A(n21620), .B(n21621), .X(n21574) );
  nand_x1_sg U35244 ( .A(n21433), .B(n21434), .X(n21387) );
  nand_x1_sg U35245 ( .A(n21525), .B(n21526), .X(n21480) );
  nand_x1_sg U35246 ( .A(n15285), .B(n15286), .X(n29667) );
  nand_x1_sg U35247 ( .A(n15287), .B(n31874), .X(n15286) );
  nor_x1_sg U35248 ( .A(n15254), .B(n15255), .X(n15253) );
  inv_x1_sg U35249 ( .A(n21086), .X(n42543) );
  inv_x1_sg U35250 ( .A(n21007), .X(n42544) );
  inv_x1_sg U35251 ( .A(n21577), .X(n42539) );
  inv_x1_sg U35252 ( .A(n21390), .X(n42541) );
  inv_x1_sg U35253 ( .A(n21482), .X(n42540) );
  nand_x1_sg U35254 ( .A(n34449), .B(n11845), .X(n11840) );
  nand_x1_sg U35255 ( .A(n12117), .B(n35560), .X(n35624) );
  nand_x1_sg U35256 ( .A(n12119), .B(n11609), .X(n35560) );
  nand_x1_sg U35257 ( .A(n12344), .B(n12345), .X(n35623) );
  nand_x1_sg U35258 ( .A(n12346), .B(n11639), .X(n12345) );
  nand_x1_sg U35259 ( .A(n12430), .B(n12431), .X(n35649) );
  nand_x1_sg U35260 ( .A(n19579), .B(n12432), .X(n12431) );
  nand_x1_sg U35261 ( .A(n13093), .B(n13094), .X(n13092) );
  nand_x1_sg U35262 ( .A(n12977), .B(n13791), .X(n13364) );
  nand_x1_sg U35263 ( .A(n12983), .B(n13828), .X(n13372) );
  nand_x1_sg U35264 ( .A(n12989), .B(n13859), .X(n13378) );
  nand_x1_sg U35265 ( .A(n12995), .B(n13890), .X(n13384) );
  nand_x1_sg U35266 ( .A(n13001), .B(n13921), .X(n13390) );
  nand_x1_sg U35267 ( .A(n13007), .B(n13952), .X(n13396) );
  nand_x1_sg U35268 ( .A(n13013), .B(n13983), .X(n13402) );
  nand_x1_sg U35269 ( .A(n13019), .B(n14014), .X(n13408) );
  nand_x1_sg U35270 ( .A(n13025), .B(n14045), .X(n13414) );
  nand_x1_sg U35271 ( .A(n13031), .B(n14076), .X(n13420) );
  nand_x1_sg U35272 ( .A(n13037), .B(n14107), .X(n13426) );
  nand_x1_sg U35273 ( .A(n13043), .B(n14138), .X(n13432) );
  nand_x1_sg U35274 ( .A(n13049), .B(n14169), .X(n13438) );
  nand_x1_sg U35275 ( .A(n13055), .B(n14200), .X(n13444) );
  nand_x1_sg U35276 ( .A(n13061), .B(n14231), .X(n13450) );
  nand_x1_sg U35277 ( .A(n13067), .B(n14262), .X(n13456) );
  nand_x1_sg U35278 ( .A(n13073), .B(n14293), .X(n13462) );
  nand_x1_sg U35279 ( .A(n13079), .B(n14324), .X(n13468) );
  nand_x1_sg U35280 ( .A(n13085), .B(n14355), .X(n13474) );
  nand_x1_sg U35281 ( .A(n13099), .B(n14386), .X(n13480) );
  nand_x1_sg U35282 ( .A(n13108), .B(n14418), .X(n13493) );
  nand_x1_sg U35283 ( .A(n13114), .B(n14449), .X(n13499) );
  nand_x1_sg U35284 ( .A(n13125), .B(n14513), .X(n13510) );
  nand_x1_sg U35285 ( .A(n13136), .B(n14575), .X(n13521) );
  nand_x1_sg U35286 ( .A(n13142), .B(n14606), .X(n13527) );
  nand_x1_sg U35287 ( .A(n13148), .B(n14637), .X(n13533) );
  nand_x1_sg U35288 ( .A(n13154), .B(n14668), .X(n13539) );
  nand_x1_sg U35289 ( .A(n13160), .B(n14699), .X(n13545) );
  nand_x1_sg U35290 ( .A(n13166), .B(n14730), .X(n13551) );
  nand_x1_sg U35291 ( .A(n13172), .B(n14761), .X(n13557) );
  nand_x1_sg U35292 ( .A(n13178), .B(n14792), .X(n13563) );
  nand_x1_sg U35293 ( .A(n13184), .B(n14823), .X(n13569) );
  nand_x1_sg U35294 ( .A(n13190), .B(n14854), .X(n13575) );
  nand_x1_sg U35295 ( .A(n13196), .B(n14885), .X(n13581) );
  nand_x1_sg U35296 ( .A(n13202), .B(n14916), .X(n13587) );
  nand_x1_sg U35297 ( .A(n13225), .B(n15009), .X(n13603) );
  nand_x1_sg U35298 ( .A(n28967), .B(n31662), .X(n15284) );
  nor_x1_sg U35299 ( .A(n15125), .B(n15126), .X(n15124) );
  nand_x1_sg U35300 ( .A(n29666), .B(n31661), .X(n15183) );
  nand_x1_sg U35301 ( .A(n21725), .B(n21726), .X(n21370) );
  nand_x1_sg U35302 ( .A(n28255), .B(n28256), .X(n35485) );
  nand_x1_sg U35303 ( .A(n28255), .B(n28256), .X(n32008) );
  inv_x1_sg U35304 ( .A(n34389), .X(n33880) );
  inv_x1_sg U35305 ( .A(n33879), .X(n33886) );
  inv_x1_sg U35306 ( .A(n33879), .X(n33883) );
  nand_x1_sg U35307 ( .A(n11890), .B(n19581), .X(n11889) );
  nand_x1_sg U35308 ( .A(n41459), .B(n11898), .X(n11800) );
  nand_x1_sg U35309 ( .A(n41460), .B(n11910), .X(n11803) );
  nand_x1_sg U35310 ( .A(n41461), .B(n11921), .X(n11805) );
  nand_x1_sg U35311 ( .A(n41462), .B(n11932), .X(n11807) );
  nand_x1_sg U35312 ( .A(n41463), .B(n11943), .X(n11809) );
  nand_x1_sg U35313 ( .A(n41464), .B(n11954), .X(n11811) );
  nand_x1_sg U35314 ( .A(n41465), .B(n11965), .X(n11813) );
  nand_x1_sg U35315 ( .A(n41466), .B(n11976), .X(n11815) );
  nand_x1_sg U35316 ( .A(n41467), .B(n11987), .X(n11817) );
  nand_x1_sg U35317 ( .A(n41468), .B(n11998), .X(n11819) );
  nand_x1_sg U35318 ( .A(n41469), .B(n12009), .X(n11821) );
  nand_x1_sg U35319 ( .A(n41470), .B(n12020), .X(n11823) );
  nand_x1_sg U35320 ( .A(n41471), .B(n12031), .X(n11825) );
  nand_x1_sg U35321 ( .A(n41472), .B(n12042), .X(n11827) );
  nand_x1_sg U35322 ( .A(n41473), .B(n12053), .X(n11829) );
  nand_x1_sg U35323 ( .A(n41474), .B(n12064), .X(n11831) );
  nand_x1_sg U35324 ( .A(n41475), .B(n12075), .X(n11833) );
  nand_x1_sg U35325 ( .A(n41476), .B(n12086), .X(n11835) );
  nand_x1_sg U35326 ( .A(n41477), .B(n12097), .X(n11837) );
  nand_x1_sg U35327 ( .A(n41478), .B(n12108), .X(n11839) );
  nand_x1_sg U35328 ( .A(n41479), .B(n12126), .X(n11848) );
  nand_x1_sg U35329 ( .A(n41480), .B(n12138), .X(n11851) );
  nand_x1_sg U35330 ( .A(n41481), .B(n12149), .X(n11853) );
  nand_x1_sg U35331 ( .A(n41482), .B(n12160), .X(n11855) );
  nand_x1_sg U35332 ( .A(n41483), .B(n12171), .X(n11857) );
  nand_x1_sg U35333 ( .A(n41484), .B(n12182), .X(n11859) );
  nand_x1_sg U35334 ( .A(n41485), .B(n12193), .X(n11861) );
  nand_x1_sg U35335 ( .A(n41486), .B(n12204), .X(n11863) );
  nand_x1_sg U35336 ( .A(n41487), .B(n12215), .X(n11865) );
  nand_x1_sg U35337 ( .A(n41488), .B(n12226), .X(n11867) );
  nand_x1_sg U35338 ( .A(n41489), .B(n12237), .X(n11869) );
  nand_x1_sg U35339 ( .A(n41490), .B(n12248), .X(n11871) );
  nand_x1_sg U35340 ( .A(n41491), .B(n12259), .X(n11873) );
  nand_x1_sg U35341 ( .A(n41492), .B(n12270), .X(n11875) );
  nand_x1_sg U35342 ( .A(n41493), .B(n12281), .X(n11877) );
  nand_x1_sg U35343 ( .A(n41494), .B(n12292), .X(n11879) );
  nand_x1_sg U35344 ( .A(n41495), .B(n12303), .X(n11881) );
  nand_x1_sg U35345 ( .A(n41496), .B(n12314), .X(n11883) );
  nand_x1_sg U35346 ( .A(n41497), .B(n12325), .X(n11885) );
  nand_x1_sg U35347 ( .A(n41498), .B(n12336), .X(n11887) );
  nand_x1_sg U35348 ( .A(n12834), .B(n12964), .X(n12963) );
  nand_x1_sg U35349 ( .A(n11637), .B(n12966), .X(n12962) );
  nand_x1_sg U35350 ( .A(n14488), .B(n14489), .X(n12448) );
  inv_x1_sg U35351 ( .A(n13117), .X(n41135) );
  nand_x1_sg U35352 ( .A(n14552), .B(n14553), .X(n12457) );
  inv_x1_sg U35353 ( .A(n35453), .X(n41136) );
  nand_x1_sg U35354 ( .A(n14955), .B(n14956), .X(n12510) );
  inv_x1_sg U35355 ( .A(n13205), .X(n41137) );
  nand_x1_sg U35356 ( .A(n14986), .B(n14987), .X(n12515) );
  inv_x1_sg U35357 ( .A(n13210), .X(n41138) );
  nand_x1_sg U35358 ( .A(n13289), .B(n31200), .X(n13288) );
  nand_x1_sg U35359 ( .A(n13291), .B(n35102), .X(n13357) );
  nand_x1_sg U35360 ( .A(n13485), .B(n30134), .X(n13484) );
  nand_x1_sg U35361 ( .A(n13487), .B(n13098), .X(n13483) );
  nand_x1_sg U35362 ( .A(n13698), .B(n13098), .X(n13697) );
  nand_x1_sg U35363 ( .A(n13780), .B(n13222), .X(n13779) );
  nor_x1_sg U35364 ( .A(n22210), .B(reset), .X(n19606) );
  nand_x1_sg U35365 ( .A(n20938), .B(n20954), .X(n20953) );
  nand_x1_sg U35366 ( .A(n20955), .B(n20956), .X(n20954) );
  nand_x1_sg U35367 ( .A(n35484), .B(n21332), .X(n21330) );
  nand_x1_sg U35368 ( .A(n21333), .B(n21334), .X(n21332) );
  nand_x1_sg U35369 ( .A(n28255), .B(n28256), .X(n32007) );
  nand_x1_sg U35370 ( .A(n33716), .B(n12731), .X(n12730) );
  nand_x1_sg U35371 ( .A(n33796), .B(n12861), .X(n12860) );
  nand_x1_sg U35372 ( .A(n33733), .B(n13237), .X(n13236) );
  nand_x1_sg U35373 ( .A(n33635), .B(n13304), .X(n13303) );
  nand_x1_sg U35374 ( .A(n33741), .B(n13382), .X(n13381) );
  nand_x1_sg U35375 ( .A(n33720), .B(n13508), .X(n13507) );
  nand_x1_sg U35376 ( .A(n33737), .B(n13629), .X(n13628) );
  nand_x1_sg U35377 ( .A(n33724), .B(n13714), .X(n13713) );
  nand_x1_sg U35378 ( .A(n33523), .B(n14474), .X(n14473) );
  nand_x4_sg U35379 ( .A(n26574), .B(n35527), .X(n31201) );
  inv_x1_sg U35380 ( .A(n35012), .X(n29671) );
  inv_x1_sg U35381 ( .A(n30693), .X(n29672) );
  inv_x1_sg U35382 ( .A(n32485), .X(n29673) );
  inv_x1_sg U35383 ( .A(n30778), .X(n29674) );
  inv_x1_sg U35384 ( .A(n29674), .X(n29675) );
  inv_x1_sg U35385 ( .A(n19589), .X(n29676) );
  inv_x1_sg U35386 ( .A(n31061), .X(n29677) );
  inv_x1_sg U35387 ( .A(n31066), .X(n29678) );
  inv_x1_sg U35388 ( .A(n31228), .X(n29679) );
  inv_x1_sg U35389 ( .A(n31239), .X(n29680) );
  inv_x1_sg U35390 ( .A(n31244), .X(n29681) );
  inv_x1_sg U35391 ( .A(n31477), .X(n29682) );
  inv_x1_sg U35392 ( .A(n29800), .X(n29683) );
  inv_x1_sg U35393 ( .A(n35685), .X(n29684) );
  inv_x1_sg U35394 ( .A(n31103), .X(n29685) );
  inv_x1_sg U35395 ( .A(n31616), .X(n29686) );
  inv_x1_sg U35396 ( .A(n31098), .X(n29687) );
  inv_x1_sg U35397 ( .A(n30912), .X(n29688) );
  inv_x1_sg U35398 ( .A(n29675), .X(n29689) );
  inv_x1_sg U35399 ( .A(n29675), .X(n29690) );
  inv_x1_sg U35400 ( .A(n31679), .X(n29691) );
  inv_x1_sg U35401 ( .A(n29691), .X(n29692) );
  inv_x1_sg U35402 ( .A(n31680), .X(n29693) );
  inv_x1_sg U35403 ( .A(n29693), .X(n29694) );
  inv_x1_sg U35404 ( .A(n31681), .X(n29695) );
  inv_x1_sg U35405 ( .A(n29695), .X(n29696) );
  inv_x1_sg U35406 ( .A(n31682), .X(n29697) );
  inv_x1_sg U35407 ( .A(n29697), .X(n29698) );
  inv_x1_sg U35408 ( .A(n31683), .X(n29699) );
  inv_x1_sg U35409 ( .A(n29699), .X(n29700) );
  inv_x1_sg U35410 ( .A(n31684), .X(n29701) );
  inv_x1_sg U35411 ( .A(n29701), .X(n29702) );
  inv_x1_sg U35412 ( .A(n30533), .X(n29703) );
  inv_x1_sg U35413 ( .A(n30531), .X(n29704) );
  inv_x1_sg U35414 ( .A(n31304), .X(n29705) );
  inv_x1_sg U35415 ( .A(n31307), .X(n29706) );
  inv_x1_sg U35416 ( .A(n31310), .X(n29707) );
  inv_x1_sg U35417 ( .A(n31313), .X(n29708) );
  inv_x1_sg U35418 ( .A(n31316), .X(n29709) );
  inv_x1_sg U35419 ( .A(n31319), .X(n29710) );
  inv_x1_sg U35420 ( .A(n31322), .X(n29711) );
  inv_x1_sg U35421 ( .A(n31325), .X(n29712) );
  inv_x1_sg U35422 ( .A(n31328), .X(n29713) );
  inv_x1_sg U35423 ( .A(n31331), .X(n29714) );
  inv_x1_sg U35424 ( .A(n31334), .X(n29715) );
  inv_x1_sg U35425 ( .A(n31337), .X(n29716) );
  inv_x1_sg U35426 ( .A(n31340), .X(n29717) );
  inv_x1_sg U35427 ( .A(n31343), .X(n29718) );
  inv_x1_sg U35428 ( .A(n31346), .X(n29719) );
  inv_x1_sg U35429 ( .A(n31349), .X(n29720) );
  inv_x1_sg U35430 ( .A(n31352), .X(n29721) );
  inv_x1_sg U35431 ( .A(n31355), .X(n29722) );
  inv_x1_sg U35432 ( .A(n31358), .X(n29723) );
  inv_x1_sg U35433 ( .A(n31361), .X(n29724) );
  inv_x1_sg U35434 ( .A(n31364), .X(n29725) );
  inv_x1_sg U35435 ( .A(n31367), .X(n29726) );
  inv_x1_sg U35436 ( .A(n31370), .X(n29727) );
  inv_x1_sg U35437 ( .A(n31385), .X(n29728) );
  inv_x1_sg U35438 ( .A(n31388), .X(n29729) );
  inv_x1_sg U35439 ( .A(n31391), .X(n29730) );
  inv_x1_sg U35440 ( .A(n31394), .X(n29731) );
  inv_x1_sg U35441 ( .A(n31397), .X(n29732) );
  inv_x1_sg U35442 ( .A(n31406), .X(n29733) );
  inv_x1_sg U35443 ( .A(n31409), .X(n29734) );
  inv_x1_sg U35444 ( .A(n31415), .X(n29735) );
  inv_x1_sg U35445 ( .A(n31418), .X(n29736) );
  inv_x1_sg U35446 ( .A(n31421), .X(n29737) );
  inv_x1_sg U35447 ( .A(n31424), .X(n29738) );
  inv_x1_sg U35448 ( .A(n31427), .X(n29739) );
  inv_x1_sg U35449 ( .A(n31430), .X(n29740) );
  inv_x1_sg U35450 ( .A(n31433), .X(n29741) );
  inv_x1_sg U35451 ( .A(n31436), .X(n29742) );
  inv_x1_sg U35452 ( .A(n31439), .X(n29743) );
  inv_x1_sg U35453 ( .A(n31442), .X(n29744) );
  inv_x1_sg U35454 ( .A(n31445), .X(n29745) );
  inv_x1_sg U35455 ( .A(n31448), .X(n29746) );
  inv_x1_sg U35456 ( .A(n31451), .X(n29747) );
  inv_x1_sg U35457 ( .A(n31454), .X(n29748) );
  inv_x1_sg U35458 ( .A(n32053), .X(n29749) );
  inv_x1_sg U35459 ( .A(n29749), .X(n29750) );
  inv_x1_sg U35460 ( .A(n29753), .X(n29751) );
  inv_x1_sg U35461 ( .A(n29753), .X(n29752) );
  inv_x1_sg U35462 ( .A(n32083), .X(n29753) );
  inv_x1_sg U35463 ( .A(n29753), .X(n29754) );
  inv_x1_sg U35464 ( .A(n30139), .X(n29755) );
  inv_x1_sg U35465 ( .A(n30139), .X(n29756) );
  inv_x1_sg U35466 ( .A(n30862), .X(n29757) );
  inv_x1_sg U35467 ( .A(n30721), .X(n29758) );
  inv_x1_sg U35468 ( .A(n34654), .X(n29759) );
  inv_x1_sg U35469 ( .A(n35316), .X(n29760) );
  inv_x1_sg U35470 ( .A(n29672), .X(n29761) );
  inv_x1_sg U35471 ( .A(n30710), .X(n29762) );
  inv_x1_sg U35472 ( .A(n30710), .X(n29763) );
  inv_x1_sg U35473 ( .A(n29766), .X(n29764) );
  inv_x1_sg U35474 ( .A(n29766), .X(n29765) );
  inv_x1_sg U35475 ( .A(n32745), .X(n29766) );
  inv_x1_sg U35476 ( .A(n29766), .X(n29767) );
  inv_x1_sg U35477 ( .A(n30728), .X(n29768) );
  inv_x1_sg U35478 ( .A(n31024), .X(n29769) );
  inv_x1_sg U35479 ( .A(n32896), .X(n29770) );
  inv_x1_sg U35480 ( .A(n29770), .X(n29771) );
  inv_x1_sg U35481 ( .A(n30042), .X(n29772) );
  inv_x1_sg U35482 ( .A(n32916), .X(n29773) );
  inv_x1_sg U35483 ( .A(n29773), .X(n29774) );
  inv_x1_sg U35484 ( .A(n32921), .X(n29775) );
  inv_x1_sg U35485 ( .A(n29775), .X(n29776) );
  inv_x1_sg U35486 ( .A(n32952), .X(n29777) );
  inv_x1_sg U35487 ( .A(n29777), .X(n29778) );
  inv_x1_sg U35488 ( .A(n32953), .X(n29779) );
  inv_x1_sg U35489 ( .A(n29779), .X(n29780) );
  inv_x1_sg U35490 ( .A(n32954), .X(n29781) );
  inv_x1_sg U35491 ( .A(n29781), .X(n29782) );
  inv_x1_sg U35492 ( .A(n32959), .X(n29783) );
  inv_x1_sg U35493 ( .A(n29783), .X(n29784) );
  inv_x1_sg U35494 ( .A(n32960), .X(n29785) );
  inv_x1_sg U35495 ( .A(n29785), .X(n29786) );
  inv_x1_sg U35496 ( .A(n32961), .X(n29787) );
  inv_x1_sg U35497 ( .A(n29787), .X(n29788) );
  inv_x1_sg U35498 ( .A(n32966), .X(n29789) );
  inv_x1_sg U35499 ( .A(n29789), .X(n29790) );
  inv_x1_sg U35500 ( .A(n32967), .X(n29791) );
  inv_x1_sg U35501 ( .A(n29791), .X(n29792) );
  inv_x1_sg U35502 ( .A(n32968), .X(n29793) );
  inv_x1_sg U35503 ( .A(n29793), .X(n29794) );
  inv_x1_sg U35504 ( .A(n30129), .X(n29795) );
  inv_x1_sg U35505 ( .A(n32972), .X(n29796) );
  inv_x1_sg U35506 ( .A(n32084), .X(n29797) );
  inv_x1_sg U35507 ( .A(n29797), .X(n29798) );
  inv_x1_sg U35508 ( .A(n29800), .X(n29799) );
  inv_x1_sg U35509 ( .A(n31212), .X(n29800) );
  inv_x1_sg U35510 ( .A(n29800), .X(n29801) );
  inv_x1_sg U35511 ( .A(n33055), .X(n29802) );
  inv_x1_sg U35512 ( .A(n29802), .X(n29803) );
  inv_x1_sg U35513 ( .A(n33055), .X(n29804) );
  inv_x1_sg U35514 ( .A(n33060), .X(n29805) );
  inv_x1_sg U35515 ( .A(n29805), .X(n29806) );
  inv_x1_sg U35516 ( .A(n33060), .X(n29807) );
  inv_x1_sg U35517 ( .A(n33067), .X(n29808) );
  inv_x1_sg U35518 ( .A(n29808), .X(n29809) );
  inv_x1_sg U35519 ( .A(n33067), .X(n29810) );
  inv_x1_sg U35520 ( .A(n33072), .X(n29811) );
  inv_x1_sg U35521 ( .A(n29811), .X(n29812) );
  inv_x1_sg U35522 ( .A(n33072), .X(n29813) );
  inv_x1_sg U35523 ( .A(n33077), .X(n29814) );
  inv_x1_sg U35524 ( .A(n29814), .X(n29815) );
  inv_x1_sg U35525 ( .A(n33079), .X(n29816) );
  inv_x1_sg U35526 ( .A(n29816), .X(n29817) );
  inv_x1_sg U35527 ( .A(n33079), .X(n29818) );
  inv_x1_sg U35528 ( .A(n33084), .X(n29819) );
  inv_x1_sg U35529 ( .A(n29819), .X(n29820) );
  inv_x1_sg U35530 ( .A(n33084), .X(n29821) );
  inv_x1_sg U35531 ( .A(n30242), .X(n29822) );
  inv_x1_sg U35532 ( .A(n30244), .X(n29823) );
  inv_x1_sg U35533 ( .A(n33096), .X(n29824) );
  inv_x1_sg U35534 ( .A(n29828), .X(n29825) );
  inv_x1_sg U35535 ( .A(n29828), .X(n29826) );
  inv_x1_sg U35536 ( .A(n33108), .X(n29827) );
  inv_x1_sg U35537 ( .A(n33113), .X(n29828) );
  inv_x1_sg U35538 ( .A(n29828), .X(n29829) );
  inv_x1_sg U35539 ( .A(n33115), .X(n29830) );
  inv_x1_sg U35540 ( .A(n29832), .X(n29831) );
  inv_x1_sg U35541 ( .A(n33126), .X(n29832) );
  inv_x1_sg U35542 ( .A(n29832), .X(n29833) );
  inv_x1_sg U35543 ( .A(n33127), .X(n29834) );
  inv_x1_sg U35544 ( .A(n29834), .X(n29835) );
  inv_x1_sg U35545 ( .A(n33127), .X(n29836) );
  inv_x1_sg U35546 ( .A(n33134), .X(n29837) );
  inv_x1_sg U35547 ( .A(n29837), .X(n29838) );
  inv_x1_sg U35548 ( .A(n29838), .X(n29839) );
  inv_x1_sg U35549 ( .A(n33139), .X(n29840) );
  inv_x1_sg U35550 ( .A(n29840), .X(n29841) );
  inv_x1_sg U35551 ( .A(n29841), .X(n29842) );
  inv_x1_sg U35552 ( .A(n30218), .X(n29843) );
  inv_x1_sg U35553 ( .A(n30237), .X(n29844) );
  inv_x1_sg U35554 ( .A(n33151), .X(n29845) );
  inv_x1_sg U35555 ( .A(n33158), .X(n29846) );
  inv_x1_sg U35556 ( .A(n29848), .X(n29847) );
  inv_x1_sg U35557 ( .A(n33167), .X(n29848) );
  inv_x1_sg U35558 ( .A(n29848), .X(n29849) );
  inv_x1_sg U35559 ( .A(n33174), .X(n29850) );
  inv_x1_sg U35560 ( .A(n30229), .X(n29851) );
  inv_x1_sg U35561 ( .A(n30228), .X(n29852) );
  inv_x1_sg U35562 ( .A(n33181), .X(n29853) );
  inv_x1_sg U35563 ( .A(n33186), .X(n29854) );
  inv_x1_sg U35564 ( .A(n29854), .X(n29855) );
  inv_x1_sg U35565 ( .A(n29855), .X(n29856) );
  inv_x1_sg U35566 ( .A(n33193), .X(n29857) );
  inv_x1_sg U35567 ( .A(n33198), .X(n29858) );
  inv_x1_sg U35568 ( .A(n29858), .X(n29859) );
  inv_x1_sg U35569 ( .A(n29859), .X(n29860) );
  inv_x1_sg U35570 ( .A(n33205), .X(n29861) );
  inv_x1_sg U35571 ( .A(n29861), .X(n29862) );
  inv_x1_sg U35572 ( .A(n29862), .X(n29863) );
  inv_x1_sg U35573 ( .A(n33210), .X(n29864) );
  inv_x1_sg U35574 ( .A(n33217), .X(n29865) );
  inv_x1_sg U35575 ( .A(n29865), .X(n29866) );
  inv_x1_sg U35576 ( .A(n33217), .X(n29867) );
  inv_x1_sg U35577 ( .A(n33222), .X(n29868) );
  inv_x1_sg U35578 ( .A(n29868), .X(n29869) );
  inv_x1_sg U35579 ( .A(n33223), .X(n29870) );
  inv_x1_sg U35580 ( .A(n29870), .X(n29871) );
  inv_x1_sg U35581 ( .A(n29896), .X(n29872) );
  inv_x1_sg U35582 ( .A(n29868), .X(n29873) );
  inv_x1_sg U35583 ( .A(n29868), .X(n29874) );
  inv_x1_sg U35584 ( .A(n29868), .X(n29875) );
  inv_x1_sg U35585 ( .A(n33229), .X(n29876) );
  inv_x1_sg U35586 ( .A(n29876), .X(n29877) );
  inv_x1_sg U35587 ( .A(n33230), .X(n29878) );
  inv_x1_sg U35588 ( .A(n29878), .X(n29879) );
  inv_x1_sg U35589 ( .A(n33232), .X(n29880) );
  inv_x1_sg U35590 ( .A(n29880), .X(n29881) );
  inv_x1_sg U35591 ( .A(n33233), .X(n29882) );
  inv_x1_sg U35592 ( .A(n29882), .X(n29883) );
  inv_x1_sg U35593 ( .A(n33234), .X(n29884) );
  inv_x1_sg U35594 ( .A(n29884), .X(n29885) );
  inv_x1_sg U35595 ( .A(n33235), .X(n29886) );
  inv_x1_sg U35596 ( .A(n29886), .X(n29887) );
  inv_x1_sg U35597 ( .A(n33237), .X(n29888) );
  inv_x1_sg U35598 ( .A(n29888), .X(n29889) );
  inv_x1_sg U35599 ( .A(n33238), .X(n29890) );
  inv_x1_sg U35600 ( .A(n29890), .X(n29891) );
  inv_x1_sg U35601 ( .A(n33239), .X(n29892) );
  inv_x1_sg U35602 ( .A(n29892), .X(n29893) );
  inv_x1_sg U35603 ( .A(n33240), .X(n29894) );
  inv_x1_sg U35604 ( .A(n29894), .X(n29895) );
  inv_x1_sg U35605 ( .A(n34843), .X(n29896) );
  inv_x1_sg U35606 ( .A(n29896), .X(n29897) );
  inv_x1_sg U35607 ( .A(n29870), .X(n29898) );
  inv_x1_sg U35608 ( .A(n34831), .X(n29899) );
  inv_x1_sg U35609 ( .A(n29899), .X(n29900) );
  inv_x1_sg U35610 ( .A(n29900), .X(n29901) );
  inv_x1_sg U35611 ( .A(n35055), .X(n29902) );
  inv_x1_sg U35612 ( .A(n33254), .X(n29903) );
  inv_x1_sg U35613 ( .A(n30212), .X(n29904) );
  inv_x1_sg U35614 ( .A(n33259), .X(n29905) );
  inv_x1_sg U35615 ( .A(n30119), .X(n29906) );
  inv_x1_sg U35616 ( .A(n30119), .X(n29907) );
  inv_x1_sg U35617 ( .A(n35642), .X(n29908) );
  inv_x1_sg U35618 ( .A(n33274), .X(n29909) );
  inv_x1_sg U35619 ( .A(n35648), .X(n29910) );
  inv_x1_sg U35620 ( .A(n33279), .X(n29911) );
  inv_x1_sg U35621 ( .A(n12976), .X(n29912) );
  inv_x1_sg U35622 ( .A(n33284), .X(n29913) );
  inv_x1_sg U35623 ( .A(n12353), .X(n29914) );
  inv_x1_sg U35624 ( .A(n33289), .X(n29915) );
  inv_x1_sg U35625 ( .A(n35659), .X(n29916) );
  inv_x1_sg U35626 ( .A(n29916), .X(n29917) );
  inv_x1_sg U35627 ( .A(n29492), .X(n29918) );
  inv_x1_sg U35628 ( .A(n29918), .X(n29919) );
  inv_x1_sg U35629 ( .A(n28978), .X(n29920) );
  inv_x1_sg U35630 ( .A(n29920), .X(n29921) );
  inv_x1_sg U35631 ( .A(n35662), .X(n29922) );
  inv_x1_sg U35632 ( .A(n29922), .X(n29923) );
  inv_x1_sg U35633 ( .A(n35668), .X(n29924) );
  inv_x1_sg U35634 ( .A(n29924), .X(n29925) );
  inv_x1_sg U35635 ( .A(n35670), .X(n29926) );
  inv_x1_sg U35636 ( .A(n29926), .X(n29927) );
  inv_x1_sg U35637 ( .A(n35658), .X(n29928) );
  inv_x1_sg U35638 ( .A(n29928), .X(n29929) );
  inv_x1_sg U35639 ( .A(n35660), .X(n29930) );
  inv_x1_sg U35640 ( .A(n29930), .X(n29931) );
  inv_x1_sg U35641 ( .A(n35671), .X(n29932) );
  inv_x1_sg U35642 ( .A(n29932), .X(n29933) );
  inv_x1_sg U35643 ( .A(n35674), .X(n29934) );
  inv_x1_sg U35644 ( .A(n29934), .X(n29935) );
  inv_x1_sg U35645 ( .A(n28452), .X(n29936) );
  inv_x1_sg U35646 ( .A(n29936), .X(n29937) );
  inv_x1_sg U35647 ( .A(n35681), .X(n29938) );
  inv_x1_sg U35648 ( .A(n29938), .X(n29939) );
  inv_x1_sg U35649 ( .A(n35672), .X(n29940) );
  inv_x1_sg U35650 ( .A(n29940), .X(n29941) );
  inv_x1_sg U35651 ( .A(n28621), .X(n29942) );
  inv_x1_sg U35652 ( .A(n29942), .X(n29943) );
  inv_x1_sg U35653 ( .A(n35680), .X(n29944) );
  inv_x1_sg U35654 ( .A(n29944), .X(n29945) );
  inv_x1_sg U35655 ( .A(n28705), .X(n29946) );
  inv_x1_sg U35656 ( .A(n29946), .X(n29947) );
  inv_x1_sg U35657 ( .A(n35673), .X(n29948) );
  inv_x1_sg U35658 ( .A(n29948), .X(n29949) );
  inv_x1_sg U35659 ( .A(n35675), .X(n29950) );
  inv_x1_sg U35660 ( .A(n29950), .X(n29951) );
  inv_x1_sg U35661 ( .A(n35678), .X(n29952) );
  inv_x1_sg U35662 ( .A(n29952), .X(n29953) );
  inv_x1_sg U35663 ( .A(n29623), .X(n29954) );
  inv_x1_sg U35664 ( .A(n29954), .X(n29955) );
  inv_x1_sg U35665 ( .A(n35664), .X(n29956) );
  inv_x1_sg U35666 ( .A(n29956), .X(n29957) );
  inv_x1_sg U35667 ( .A(n29447), .X(n29958) );
  inv_x1_sg U35668 ( .A(n29958), .X(n29959) );
  inv_x1_sg U35669 ( .A(n35663), .X(n29960) );
  inv_x1_sg U35670 ( .A(n29960), .X(n29961) );
  inv_x1_sg U35671 ( .A(n12134), .X(n29962) );
  inv_x1_sg U35672 ( .A(n33409), .X(n29963) );
  inv_x1_sg U35673 ( .A(n11906), .X(n29964) );
  inv_x1_sg U35674 ( .A(n33414), .X(n29965) );
  inv_x1_sg U35675 ( .A(n11895), .X(n29966) );
  inv_x1_sg U35676 ( .A(n33419), .X(n29967) );
  inv_x1_sg U35677 ( .A(n35651), .X(n29968) );
  inv_x1_sg U35678 ( .A(n33424), .X(n29969) );
  inv_x1_sg U35679 ( .A(n35676), .X(n29970) );
  inv_x1_sg U35680 ( .A(n29970), .X(n29971) );
  inv_x1_sg U35681 ( .A(n35665), .X(n29972) );
  inv_x1_sg U35682 ( .A(n29972), .X(n29973) );
  inv_x1_sg U35683 ( .A(n35661), .X(n29974) );
  inv_x1_sg U35684 ( .A(n29974), .X(n29975) );
  inv_x1_sg U35685 ( .A(n35679), .X(n29976) );
  inv_x1_sg U35686 ( .A(n29976), .X(n29977) );
  inv_x1_sg U35687 ( .A(n35669), .X(n29978) );
  inv_x1_sg U35688 ( .A(n29978), .X(n29979) );
  inv_x1_sg U35689 ( .A(n35667), .X(n29980) );
  inv_x1_sg U35690 ( .A(n29980), .X(n29981) );
  inv_x1_sg U35691 ( .A(n35666), .X(n29982) );
  inv_x1_sg U35692 ( .A(n29982), .X(n29983) );
  inv_x1_sg U35693 ( .A(n29064), .X(n29984) );
  inv_x1_sg U35694 ( .A(n29984), .X(n29985) );
  inv_x1_sg U35695 ( .A(n35677), .X(n29986) );
  inv_x1_sg U35696 ( .A(n29986), .X(n29987) );
  inv_x1_sg U35697 ( .A(n33523), .X(n29988) );
  inv_x1_sg U35698 ( .A(n29988), .X(n29989) );
  inv_x1_sg U35699 ( .A(n33631), .X(n29990) );
  inv_x1_sg U35700 ( .A(n29990), .X(n29991) );
  nand_x2_sg U35701 ( .A(n13357), .B(n13358), .X(n35621) );
  inv_x1_sg U35702 ( .A(n33635), .X(n29992) );
  inv_x1_sg U35703 ( .A(n29992), .X(n29993) );
  inv_x1_sg U35704 ( .A(n33716), .X(n29994) );
  inv_x1_sg U35705 ( .A(n29994), .X(n29995) );
  inv_x1_sg U35706 ( .A(n33720), .X(n29996) );
  inv_x1_sg U35707 ( .A(n29996), .X(n29997) );
  inv_x1_sg U35708 ( .A(n33724), .X(n29998) );
  inv_x1_sg U35709 ( .A(n29998), .X(n29999) );
  inv_x1_sg U35710 ( .A(n33733), .X(n30000) );
  inv_x1_sg U35711 ( .A(n30000), .X(n30001) );
  inv_x1_sg U35712 ( .A(n33737), .X(n30002) );
  inv_x1_sg U35713 ( .A(n30002), .X(n30003) );
  inv_x1_sg U35714 ( .A(n33741), .X(n30004) );
  inv_x1_sg U35715 ( .A(n30004), .X(n30005) );
  inv_x1_sg U35716 ( .A(n33750), .X(n30006) );
  inv_x1_sg U35717 ( .A(n30006), .X(n30007) );
  inv_x1_sg U35718 ( .A(n35654), .X(n30008) );
  inv_x2_sg U35719 ( .A(n35654), .X(n33753) );
  inv_x1_sg U35720 ( .A(n33755), .X(n30009) );
  inv_x1_sg U35721 ( .A(n30009), .X(n30010) );
  inv_x1_sg U35722 ( .A(n35643), .X(n30011) );
  inv_x2_sg U35723 ( .A(n35643), .X(n33758) );
  inv_x1_sg U35724 ( .A(n33796), .X(n30012) );
  inv_x1_sg U35725 ( .A(n30012), .X(n30013) );
  inv_x1_sg U35726 ( .A(n30139), .X(n30014) );
  inv_x1_sg U35727 ( .A(n35314), .X(n30015) );
  inv_x1_sg U35728 ( .A(n30912), .X(n30016) );
  inv_x1_sg U35729 ( .A(n30911), .X(n30017) );
  inv_x1_sg U35730 ( .A(n33963), .X(n30018) );
  inv_x1_sg U35731 ( .A(n33986), .X(n30019) );
  inv_x1_sg U35732 ( .A(n30019), .X(n30020) );
  inv_x1_sg U35733 ( .A(n30531), .X(n30021) );
  inv_x1_sg U35734 ( .A(n30533), .X(n30022) );
  inv_x1_sg U35735 ( .A(n31026), .X(n30023) );
  inv_x1_sg U35736 ( .A(n30871), .X(n30024) );
  inv_x1_sg U35737 ( .A(n31063), .X(n30025) );
  inv_x1_sg U35738 ( .A(n29677), .X(n30026) );
  inv_x1_sg U35739 ( .A(n31068), .X(n30027) );
  inv_x1_sg U35740 ( .A(n29678), .X(n30028) );
  inv_x1_sg U35741 ( .A(n30930), .X(n30029) );
  inv_x1_sg U35742 ( .A(n30928), .X(n30030) );
  inv_x1_sg U35743 ( .A(n30938), .X(n30031) );
  inv_x1_sg U35744 ( .A(n30924), .X(n30032) );
  inv_x1_sg U35745 ( .A(n30936), .X(n30033) );
  inv_x1_sg U35746 ( .A(n30932), .X(n30034) );
  inv_x1_sg U35747 ( .A(n30922), .X(n30035) );
  inv_x1_sg U35748 ( .A(n30934), .X(n30036) );
  inv_x1_sg U35749 ( .A(n30873), .X(n30037) );
  inv_x1_sg U35750 ( .A(n13221), .X(n30038) );
  inv_x1_sg U35751 ( .A(n31493), .X(n30039) );
  inv_x1_sg U35752 ( .A(n30038), .X(n30040) );
  inv_x1_sg U35753 ( .A(n34100), .X(n30041) );
  inv_x1_sg U35754 ( .A(n30041), .X(n30042) );
  inv_x1_sg U35755 ( .A(n31484), .X(n30043) );
  inv_x1_sg U35756 ( .A(n31483), .X(n30044) );
  inv_x1_sg U35757 ( .A(n31474), .X(n30045) );
  inv_x1_sg U35758 ( .A(n30181), .X(n30046) );
  inv_x1_sg U35759 ( .A(n35606), .X(n30047) );
  inv_x1_sg U35760 ( .A(n30047), .X(n30048) );
  inv_x1_sg U35761 ( .A(n35600), .X(n30049) );
  inv_x1_sg U35762 ( .A(n35464), .X(n30050) );
  inv_x1_sg U35763 ( .A(n30050), .X(n30051) );
  inv_x1_sg U35764 ( .A(n11737), .X(n30052) );
  inv_x1_sg U35765 ( .A(n35462), .X(n30053) );
  inv_x1_sg U35766 ( .A(n30053), .X(n30054) );
  inv_x1_sg U35767 ( .A(n11791), .X(n30055) );
  inv_x1_sg U35768 ( .A(n35461), .X(n30056) );
  inv_x1_sg U35769 ( .A(n30056), .X(n30057) );
  inv_x1_sg U35770 ( .A(n11710), .X(n30058) );
  inv_x1_sg U35771 ( .A(n15171), .X(n30059) );
  inv_x1_sg U35772 ( .A(n30059), .X(n30060) );
  inv_x1_sg U35773 ( .A(n34128), .X(n30061) );
  inv_x1_sg U35774 ( .A(n34133), .X(n30062) );
  inv_x1_sg U35775 ( .A(n34138), .X(n30063) );
  inv_x1_sg U35776 ( .A(n34143), .X(n30064) );
  inv_x1_sg U35777 ( .A(n34148), .X(n30065) );
  inv_x1_sg U35778 ( .A(n34153), .X(n30066) );
  inv_x1_sg U35779 ( .A(n34158), .X(n30067) );
  inv_x1_sg U35780 ( .A(n34163), .X(n30068) );
  inv_x1_sg U35781 ( .A(n34168), .X(n30069) );
  inv_x1_sg U35782 ( .A(n34173), .X(n30070) );
  inv_x1_sg U35783 ( .A(n34178), .X(n30071) );
  inv_x1_sg U35784 ( .A(n34183), .X(n30072) );
  inv_x1_sg U35785 ( .A(n34188), .X(n30073) );
  inv_x1_sg U35786 ( .A(n34193), .X(n30074) );
  inv_x1_sg U35787 ( .A(n34198), .X(n30075) );
  inv_x1_sg U35788 ( .A(n34203), .X(n30076) );
  inv_x1_sg U35789 ( .A(n34208), .X(n30077) );
  inv_x1_sg U35790 ( .A(n34213), .X(n30078) );
  inv_x1_sg U35791 ( .A(n34218), .X(n30079) );
  inv_x1_sg U35792 ( .A(n34223), .X(n30080) );
  inv_x1_sg U35793 ( .A(n34228), .X(n30081) );
  inv_x1_sg U35794 ( .A(n34233), .X(n30082) );
  inv_x1_sg U35795 ( .A(n34238), .X(n30083) );
  inv_x1_sg U35796 ( .A(n34243), .X(n30084) );
  inv_x1_sg U35797 ( .A(n34248), .X(n30085) );
  inv_x1_sg U35798 ( .A(n34253), .X(n30086) );
  inv_x1_sg U35799 ( .A(n34258), .X(n30087) );
  inv_x1_sg U35800 ( .A(n34263), .X(n30088) );
  inv_x1_sg U35801 ( .A(n34268), .X(n30089) );
  inv_x1_sg U35802 ( .A(n34273), .X(n30090) );
  inv_x1_sg U35803 ( .A(n34278), .X(n30091) );
  inv_x1_sg U35804 ( .A(n34283), .X(n30092) );
  inv_x1_sg U35805 ( .A(n34288), .X(n30093) );
  inv_x1_sg U35806 ( .A(n34293), .X(n30094) );
  inv_x1_sg U35807 ( .A(n34298), .X(n30095) );
  inv_x1_sg U35808 ( .A(n34303), .X(n30096) );
  inv_x1_sg U35809 ( .A(n34308), .X(n30097) );
  inv_x1_sg U35810 ( .A(n34313), .X(n30098) );
  inv_x1_sg U35811 ( .A(n34318), .X(n30099) );
  inv_x1_sg U35812 ( .A(n34323), .X(n30100) );
  inv_x1_sg U35813 ( .A(n34328), .X(n30101) );
  inv_x1_sg U35814 ( .A(n34333), .X(n30102) );
  inv_x1_sg U35815 ( .A(n34338), .X(n30103) );
  inv_x1_sg U35816 ( .A(n34343), .X(n30104) );
  inv_x1_sg U35817 ( .A(n34348), .X(n30105) );
  inv_x1_sg U35818 ( .A(n34353), .X(n30106) );
  inv_x1_sg U35819 ( .A(n34358), .X(n30107) );
  inv_x1_sg U35820 ( .A(n34363), .X(n30108) );
  inv_x1_sg U35821 ( .A(n34368), .X(n30109) );
  inv_x1_sg U35822 ( .A(n34373), .X(n30110) );
  inv_x1_sg U35823 ( .A(n34378), .X(n30111) );
  inv_x1_sg U35824 ( .A(n34383), .X(n30112) );
  inv_x1_sg U35825 ( .A(n30858), .X(n30113) );
  inv_x1_sg U35826 ( .A(n30856), .X(n30114) );
  inv_x1_sg U35827 ( .A(n30852), .X(n30115) );
  inv_x1_sg U35828 ( .A(n34421), .X(n30116) );
  inv_x1_sg U35829 ( .A(n34426), .X(n30117) );
  inv_x1_sg U35830 ( .A(n30829), .X(n30118) );
  inv_x1_sg U35831 ( .A(n30133), .X(n30119) );
  inv_x1_sg U35832 ( .A(n33224), .X(n30120) );
  inv_x1_sg U35833 ( .A(n33225), .X(n30121) );
  inv_x1_sg U35834 ( .A(n29687), .X(n30122) );
  inv_x1_sg U35835 ( .A(n34494), .X(n30123) );
  inv_x1_sg U35836 ( .A(n30123), .X(n30124) );
  inv_x1_sg U35837 ( .A(n30123), .X(n30125) );
  inv_x1_sg U35838 ( .A(n30813), .X(n30126) );
  inv_x1_sg U35839 ( .A(n30794), .X(n30127) );
  inv_x1_sg U35840 ( .A(n30131), .X(n30128) );
  inv_x1_sg U35841 ( .A(n31004), .X(n30129) );
  inv_x1_sg U35842 ( .A(n31479), .X(n30130) );
  inv_x1_sg U35843 ( .A(n30211), .X(n30131) );
  inv_x1_sg U35844 ( .A(n30211), .X(n30132) );
  inv_x1_sg U35845 ( .A(n30211), .X(n30133) );
  inv_x1_sg U35846 ( .A(n31705), .X(n30134) );
  inv_x1_sg U35847 ( .A(n29676), .X(n30135) );
  inv_x1_sg U35848 ( .A(n32055), .X(n30136) );
  inv_x1_sg U35849 ( .A(n34543), .X(n30137) );
  inv_x1_sg U35850 ( .A(n31298), .X(n30138) );
  inv_x1_sg U35851 ( .A(n34553), .X(n30139) );
  inv_x1_sg U35852 ( .A(n30139), .X(n30140) );
  inv_x1_sg U35853 ( .A(n34562), .X(n30141) );
  inv_x1_sg U35854 ( .A(n30141), .X(n30142) );
  inv_x1_sg U35855 ( .A(n32168), .X(n30143) );
  inv_x1_sg U35856 ( .A(n30154), .X(n30144) );
  inv_x1_sg U35857 ( .A(n30152), .X(n30145) );
  inv_x1_sg U35858 ( .A(n34567), .X(n30146) );
  inv_x1_sg U35859 ( .A(n30146), .X(n30147) );
  inv_x1_sg U35860 ( .A(n34568), .X(n30148) );
  inv_x1_sg U35861 ( .A(n30148), .X(n30149) );
  inv_x1_sg U35862 ( .A(n34576), .X(n30150) );
  inv_x1_sg U35863 ( .A(n30150), .X(n30151) );
  inv_x1_sg U35864 ( .A(n34577), .X(n30152) );
  inv_x1_sg U35865 ( .A(n30152), .X(n30153) );
  inv_x1_sg U35866 ( .A(n34578), .X(n30154) );
  inv_x1_sg U35867 ( .A(n30154), .X(n30155) );
  inv_x1_sg U35868 ( .A(n34581), .X(n30156) );
  inv_x1_sg U35869 ( .A(n30156), .X(n30157) );
  inv_x1_sg U35870 ( .A(n29675), .X(n30158) );
  inv_x1_sg U35871 ( .A(n30776), .X(n30159) );
  inv_x1_sg U35872 ( .A(n30163), .X(n30160) );
  inv_x1_sg U35873 ( .A(n30163), .X(n30161) );
  inv_x1_sg U35874 ( .A(n34627), .X(n30162) );
  inv_x1_sg U35875 ( .A(n30162), .X(n30163) );
  inv_x1_sg U35876 ( .A(n30769), .X(n30164) );
  inv_x1_sg U35877 ( .A(n34637), .X(n30165) );
  inv_x1_sg U35878 ( .A(n30165), .X(n30166) );
  inv_x1_sg U35879 ( .A(n30247), .X(n30167) );
  inv_x1_sg U35880 ( .A(n30759), .X(n30168) );
  inv_x1_sg U35881 ( .A(n30756), .X(n30169) );
  inv_x1_sg U35882 ( .A(n34649), .X(n30170) );
  inv_x1_sg U35883 ( .A(n35394), .X(n30171) );
  inv_x1_sg U35884 ( .A(n35238), .X(n30172) );
  inv_x1_sg U35885 ( .A(n30706), .X(n30173) );
  inv_x1_sg U35886 ( .A(n30708), .X(n30174) );
  inv_x1_sg U35887 ( .A(n30731), .X(n30175) );
  inv_x1_sg U35888 ( .A(n34694), .X(n30176) );
  inv_x1_sg U35889 ( .A(n35378), .X(n30177) );
  inv_x1_sg U35890 ( .A(n35331), .X(n30178) );
  inv_x1_sg U35891 ( .A(n35331), .X(n30179) );
  inv_x1_sg U35892 ( .A(n35360), .X(n30180) );
  inv_x1_sg U35893 ( .A(n34956), .X(n30181) );
  inv_x1_sg U35894 ( .A(n30216), .X(n30182) );
  inv_x1_sg U35895 ( .A(n34755), .X(n30183) );
  inv_x1_sg U35896 ( .A(n30183), .X(n30184) );
  inv_x1_sg U35897 ( .A(n30648), .X(n30185) );
  inv_x1_sg U35898 ( .A(n30652), .X(n30186) );
  inv_x1_sg U35899 ( .A(n34797), .X(n30187) );
  inv_x1_sg U35900 ( .A(n30187), .X(n30188) );
  inv_x1_sg U35901 ( .A(n30215), .X(n30189) );
  inv_x1_sg U35902 ( .A(n31274), .X(n30190) );
  inv_x1_sg U35903 ( .A(n31275), .X(n30191) );
  inv_x1_sg U35904 ( .A(n31270), .X(n30192) );
  inv_x1_sg U35905 ( .A(n31265), .X(n30193) );
  inv_x1_sg U35906 ( .A(n31256), .X(n30194) );
  inv_x1_sg U35907 ( .A(n30150), .X(n30195) );
  inv_x1_sg U35908 ( .A(n30150), .X(n30196) );
  inv_x1_sg U35909 ( .A(n30150), .X(n30197) );
  inv_x1_sg U35910 ( .A(n30637), .X(n30198) );
  inv_x1_sg U35911 ( .A(n34854), .X(n30199) );
  inv_x1_sg U35912 ( .A(n30199), .X(n30200) );
  inv_x1_sg U35913 ( .A(n34862), .X(n30201) );
  inv_x1_sg U35914 ( .A(n34867), .X(n30202) );
  inv_x1_sg U35915 ( .A(n30631), .X(n30203) );
  inv_x1_sg U35916 ( .A(n30926), .X(n30204) );
  inv_x1_sg U35917 ( .A(n30626), .X(n30205) );
  inv_x1_sg U35918 ( .A(n34896), .X(n30206) );
  inv_x1_sg U35919 ( .A(n30206), .X(n30207) );
  inv_x1_sg U35920 ( .A(n32051), .X(n30208) );
  inv_x1_sg U35921 ( .A(n29681), .X(n30209) );
  inv_x1_sg U35922 ( .A(n31241), .X(n30210) );
  inv_x1_sg U35923 ( .A(n34915), .X(n30211) );
  inv_x1_sg U35924 ( .A(n30211), .X(n30212) );
  inv_x1_sg U35925 ( .A(n30154), .X(n30213) );
  inv_x1_sg U35926 ( .A(n30675), .X(n30214) );
  inv_x1_sg U35927 ( .A(n31107), .X(n30215) );
  inv_x1_sg U35928 ( .A(n31609), .X(n30216) );
  inv_x1_sg U35929 ( .A(n29679), .X(n30217) );
  inv_x1_sg U35930 ( .A(n34974), .X(n30218) );
  inv_x1_sg U35931 ( .A(n30218), .X(n30219) );
  inv_x1_sg U35932 ( .A(n30218), .X(n30220) );
  inv_x1_sg U35933 ( .A(n34978), .X(n30221) );
  inv_x1_sg U35934 ( .A(n30221), .X(n30222) );
  inv_x1_sg U35935 ( .A(n31231), .X(n30223) );
  inv_x1_sg U35936 ( .A(n31230), .X(n30224) );
  inv_x1_sg U35937 ( .A(n34983), .X(n30225) );
  inv_x1_sg U35938 ( .A(n30225), .X(n30226) );
  inv_x1_sg U35939 ( .A(n34971), .X(n30227) );
  inv_x1_sg U35940 ( .A(n30229), .X(n30228) );
  inv_x1_sg U35941 ( .A(n34994), .X(n30229) );
  inv_x1_sg U35942 ( .A(n30229), .X(n30230) );
  inv_x1_sg U35943 ( .A(n31113), .X(n30231) );
  inv_x1_sg U35944 ( .A(n34999), .X(n30232) );
  inv_x1_sg U35945 ( .A(n30232), .X(n30233) );
  inv_x1_sg U35946 ( .A(n30218), .X(n30234) );
  inv_x1_sg U35947 ( .A(n35002), .X(n30235) );
  inv_x1_sg U35948 ( .A(n30235), .X(n30236) );
  inv_x1_sg U35949 ( .A(n35003), .X(n30237) );
  inv_x1_sg U35950 ( .A(n30237), .X(n30238) );
  inv_x1_sg U35951 ( .A(n35594), .X(n30239) );
  inv_x1_sg U35952 ( .A(n31217), .X(n30240) );
  inv_x1_sg U35953 ( .A(n35034), .X(n30241) );
  inv_x1_sg U35954 ( .A(n35027), .X(n30242) );
  inv_x1_sg U35955 ( .A(n30242), .X(n30243) );
  inv_x1_sg U35956 ( .A(n30245), .X(n30244) );
  inv_x1_sg U35957 ( .A(n30974), .X(n30245) );
  inv_x1_sg U35958 ( .A(n35033), .X(n30246) );
  nand_x4_sg U35959 ( .A(n22215), .B(n23631), .X(n35455) );
  inv_x1_sg U35960 ( .A(n31109), .X(n30247) );
  inv_x1_sg U35961 ( .A(n30763), .X(n30248) );
  inv_x1_sg U35962 ( .A(n30746), .X(n30249) );
  inv_x1_sg U35963 ( .A(n30774), .X(n30250) );
  inv_x1_sg U35964 ( .A(n30771), .X(n30251) );
  inv_x1_sg U35965 ( .A(n30766), .X(n30252) );
  inv_x1_sg U35966 ( .A(n29620), .X(n30253) );
  inv_x1_sg U35967 ( .A(n28921), .X(n30254) );
  inv_x1_sg U35968 ( .A(shifter_state[0]), .X(n30255) );
  inv_x1_sg U35969 ( .A(n30628), .X(n30256) );
  inv_x1_sg U35970 ( .A(n30258), .X(n30257) );
  inv_x1_sg U35971 ( .A(n15181), .X(n30258) );
  inv_x1_sg U35972 ( .A(n30260), .X(n30259) );
  inv_x1_sg U35973 ( .A(n15180), .X(n30260) );
  inv_x1_sg U35974 ( .A(n30262), .X(n30261) );
  inv_x1_sg U35975 ( .A(n15177), .X(n30262) );
  inv_x1_sg U35976 ( .A(n30264), .X(n30263) );
  inv_x1_sg U35977 ( .A(n15048), .X(n30264) );
  inv_x1_sg U35978 ( .A(n30266), .X(n30265) );
  inv_x1_sg U35979 ( .A(n15044), .X(n30266) );
  inv_x1_sg U35980 ( .A(n30268), .X(n30267) );
  inv_x1_sg U35981 ( .A(n15190), .X(n30268) );
  inv_x1_sg U35982 ( .A(n30270), .X(n30269) );
  inv_x1_sg U35983 ( .A(n15182), .X(n30270) );
  inv_x1_sg U35984 ( .A(n30272), .X(n30271) );
  inv_x1_sg U35985 ( .A(n15055), .X(n30272) );
  inv_x1_sg U35986 ( .A(n30274), .X(n30273) );
  inv_x1_sg U35987 ( .A(n15049), .X(n30274) );
  inv_x1_sg U35988 ( .A(n30276), .X(n30275) );
  inv_x1_sg U35989 ( .A(n15172), .X(n30276) );
  inv_x1_sg U35990 ( .A(n30278), .X(n30277) );
  inv_x1_sg U35991 ( .A(n15170), .X(n30278) );
  inv_x1_sg U35992 ( .A(n30280), .X(n30279) );
  inv_x1_sg U35993 ( .A(n15039), .X(n30280) );
  inv_x1_sg U35994 ( .A(n30282), .X(n30281) );
  inv_x1_sg U35995 ( .A(n15038), .X(n30282) );
  inv_x1_sg U35996 ( .A(n30284), .X(n30283) );
  inv_x1_sg U35997 ( .A(n15037), .X(n30284) );
  inv_x1_sg U35998 ( .A(n30286), .X(n30285) );
  inv_x1_sg U35999 ( .A(n13808), .X(n30286) );
  inv_x1_sg U36000 ( .A(n31412), .X(n30287) );
  inv_x1_sg U36001 ( .A(n30289), .X(n30288) );
  inv_x1_sg U36002 ( .A(n35644), .X(n30289) );
  inv_x1_sg U36003 ( .A(n30291), .X(n30290) );
  inv_x1_sg U36004 ( .A(n35645), .X(n30291) );
  inv_x1_sg U36005 ( .A(n30293), .X(n30292) );
  inv_x1_sg U36006 ( .A(n13787), .X(n30293) );
  inv_x1_sg U36007 ( .A(n31403), .X(n30294) );
  inv_x1_sg U36008 ( .A(n30296), .X(n30295) );
  inv_x1_sg U36009 ( .A(n12531), .X(n30296) );
  inv_x1_sg U36010 ( .A(n31400), .X(n30297) );
  inv_x1_sg U36011 ( .A(n30299), .X(n30298) );
  inv_x1_sg U36012 ( .A(n35633), .X(n30299) );
  inv_x1_sg U36013 ( .A(n30301), .X(n30300) );
  inv_x1_sg U36014 ( .A(n12533), .X(n30301) );
  inv_x1_sg U36015 ( .A(n30303), .X(n30302) );
  inv_x1_sg U36016 ( .A(n35629), .X(n30303) );
  inv_x1_sg U36017 ( .A(n30305), .X(n30304) );
  inv_x1_sg U36018 ( .A(n35630), .X(n30305) );
  inv_x1_sg U36019 ( .A(n30307), .X(n30306) );
  inv_x1_sg U36020 ( .A(n35632), .X(n30307) );
  inv_x1_sg U36021 ( .A(n30309), .X(n30308) );
  inv_x1_sg U36022 ( .A(n35650), .X(n30309) );
  inv_x1_sg U36023 ( .A(n31382), .X(n30310) );
  inv_x1_sg U36024 ( .A(n30312), .X(n30311) );
  inv_x1_sg U36025 ( .A(n13816), .X(n30312) );
  inv_x1_sg U36026 ( .A(n31379), .X(n30313) );
  inv_x1_sg U36027 ( .A(n30315), .X(n30314) );
  inv_x1_sg U36028 ( .A(n13805), .X(n30315) );
  inv_x1_sg U36029 ( .A(n31376), .X(n30316) );
  inv_x1_sg U36030 ( .A(n30318), .X(n30317) );
  inv_x1_sg U36031 ( .A(n13804), .X(n30318) );
  inv_x1_sg U36032 ( .A(n31373), .X(n30319) );
  inv_x1_sg U36033 ( .A(n30321), .X(n30320) );
  inv_x1_sg U36034 ( .A(n13367), .X(n30321) );
  inv_x1_sg U36035 ( .A(n30323), .X(n30322) );
  inv_x1_sg U36036 ( .A(n11667), .X(n30323) );
  inv_x1_sg U36037 ( .A(n30325), .X(n30324) );
  inv_x1_sg U36038 ( .A(n11535), .X(n30325) );
  inv_x1_sg U36039 ( .A(n30327), .X(n30326) );
  inv_x1_sg U36040 ( .A(n15184), .X(n30327) );
  inv_x1_sg U36041 ( .A(n30329), .X(n30328) );
  inv_x1_sg U36042 ( .A(n15179), .X(n30329) );
  inv_x1_sg U36043 ( .A(n30331), .X(n30330) );
  inv_x1_sg U36044 ( .A(n15050), .X(n30331) );
  inv_x1_sg U36045 ( .A(n30333), .X(n30332) );
  inv_x1_sg U36046 ( .A(n15046), .X(n30333) );
  inv_x1_sg U36047 ( .A(n30335), .X(n30334) );
  inv_x1_sg U36048 ( .A(n35599), .X(n30335) );
  inv_x1_sg U36049 ( .A(n30337), .X(n30336) );
  inv_x1_sg U36050 ( .A(n35598), .X(n30337) );
  inv_x1_sg U36051 ( .A(n30339), .X(n30338) );
  inv_x1_sg U36052 ( .A(n35597), .X(n30339) );
  inv_x1_sg U36053 ( .A(n30341), .X(n30340) );
  inv_x1_sg U36054 ( .A(n35596), .X(n30341) );
  inv_x1_sg U36055 ( .A(n30343), .X(n30342) );
  inv_x1_sg U36056 ( .A(n35595), .X(n30343) );
  inv_x1_sg U36057 ( .A(n30345), .X(n30344) );
  inv_x1_sg U36058 ( .A(n15047), .X(n30345) );
  inv_x1_sg U36059 ( .A(n30347), .X(n30346) );
  inv_x1_sg U36060 ( .A(n15187), .X(n30347) );
  inv_x1_sg U36061 ( .A(n30349), .X(n30348) );
  inv_x1_sg U36062 ( .A(n13368), .X(n30349) );
  inv_x1_sg U36063 ( .A(n30351), .X(n30350) );
  inv_x1_sg U36064 ( .A(n35631), .X(n30351) );
  inv_x1_sg U36065 ( .A(n30353), .X(n30352) );
  inv_x1_sg U36066 ( .A(n11562), .X(n30353) );
  inv_x1_sg U36067 ( .A(n30355), .X(n30354) );
  inv_x1_sg U36068 ( .A(n11586), .X(n30355) );
  inv_x1_sg U36069 ( .A(n30357), .X(n30356) );
  inv_x1_sg U36070 ( .A(n11536), .X(n30357) );
  inv_x1_sg U36071 ( .A(n30359), .X(n30358) );
  inv_x1_sg U36072 ( .A(n11641), .X(n30359) );
  inv_x1_sg U36073 ( .A(n30361), .X(n30360) );
  inv_x1_sg U36074 ( .A(n35458), .X(n30361) );
  inv_x1_sg U36075 ( .A(n30363), .X(n30362) );
  inv_x1_sg U36076 ( .A(n35483), .X(n30363) );
  inv_x1_sg U36077 ( .A(n30365), .X(n30364) );
  inv_x1_sg U36078 ( .A(n15053), .X(n30365) );
  inv_x1_sg U36079 ( .A(n31287), .X(n30366) );
  inv_x1_sg U36080 ( .A(n30366), .X(n30367) );
  inv_x1_sg U36081 ( .A(n30366), .X(n30368) );
  inv_x1_sg U36082 ( .A(n34926), .X(n30369) );
  inv_x1_sg U36083 ( .A(n30369), .X(n30370) );
  inv_x1_sg U36084 ( .A(n30369), .X(n30371) );
  inv_x1_sg U36085 ( .A(n31278), .X(n30372) );
  inv_x1_sg U36086 ( .A(n30372), .X(n30373) );
  inv_x1_sg U36087 ( .A(n30376), .X(n30374) );
  inv_x1_sg U36088 ( .A(n30372), .X(n30375) );
  inv_x1_sg U36089 ( .A(n30377), .X(n30376) );
  inv_x1_sg U36090 ( .A(n31273), .X(n30377) );
  inv_x1_sg U36091 ( .A(n30377), .X(n30378) );
  inv_x1_sg U36092 ( .A(n30380), .X(n30379) );
  inv_x1_sg U36093 ( .A(n31268), .X(n30380) );
  inv_x1_sg U36094 ( .A(n30380), .X(n30381) );
  inv_x1_sg U36095 ( .A(n31264), .X(n30382) );
  inv_x1_sg U36096 ( .A(n31260), .X(n30383) );
  inv_x1_sg U36097 ( .A(n31261), .X(n30384) );
  inv_x1_sg U36098 ( .A(n31255), .X(n30385) );
  inv_x1_sg U36099 ( .A(n29681), .X(n30386) );
  inv_x1_sg U36100 ( .A(n31241), .X(n30387) );
  inv_x1_sg U36101 ( .A(\filter_0/N13 ), .X(n30388) );
  inv_x1_sg U36102 ( .A(n30388), .X(n30389) );
  inv_x1_sg U36103 ( .A(n35153), .X(n30390) );
  inv_x1_sg U36104 ( .A(n35152), .X(n30391) );
  inv_x1_sg U36105 ( .A(n35151), .X(n30392) );
  inv_x1_sg U36106 ( .A(n35150), .X(n30393) );
  inv_x1_sg U36107 ( .A(n35149), .X(n30394) );
  inv_x1_sg U36108 ( .A(n35148), .X(n30395) );
  inv_x1_sg U36109 ( .A(n35147), .X(n30396) );
  inv_x1_sg U36110 ( .A(n35146), .X(n30397) );
  inv_x1_sg U36111 ( .A(n35145), .X(n30398) );
  inv_x1_sg U36112 ( .A(n35144), .X(n30399) );
  inv_x1_sg U36113 ( .A(n35143), .X(n30400) );
  inv_x1_sg U36114 ( .A(n35142), .X(n30401) );
  inv_x1_sg U36115 ( .A(n35141), .X(n30402) );
  inv_x1_sg U36116 ( .A(n35140), .X(n30403) );
  inv_x1_sg U36117 ( .A(n35139), .X(n30404) );
  inv_x1_sg U36118 ( .A(\shifter_0/reg_i_8[0] ), .X(n30405) );
  inv_x1_sg U36119 ( .A(n30405), .X(n30406) );
  inv_x1_sg U36120 ( .A(\shifter_0/reg_i_8[1] ), .X(n30407) );
  inv_x1_sg U36121 ( .A(n30407), .X(n30408) );
  inv_x1_sg U36122 ( .A(\shifter_0/reg_i_8[2] ), .X(n30409) );
  inv_x1_sg U36123 ( .A(n30409), .X(n30410) );
  inv_x1_sg U36124 ( .A(\shifter_0/reg_i_8[3] ), .X(n30411) );
  inv_x1_sg U36125 ( .A(n30411), .X(n30412) );
  inv_x1_sg U36126 ( .A(\shifter_0/reg_i_8[4] ), .X(n30413) );
  inv_x1_sg U36127 ( .A(n30413), .X(n30414) );
  inv_x1_sg U36128 ( .A(\shifter_0/reg_i_8[5] ), .X(n30415) );
  inv_x1_sg U36129 ( .A(n30415), .X(n30416) );
  inv_x1_sg U36130 ( .A(\shifter_0/reg_i_8[6] ), .X(n30417) );
  inv_x1_sg U36131 ( .A(n30417), .X(n30418) );
  inv_x1_sg U36132 ( .A(\shifter_0/reg_i_8[7] ), .X(n30419) );
  inv_x1_sg U36133 ( .A(n30419), .X(n30420) );
  inv_x1_sg U36134 ( .A(\shifter_0/reg_i_8[8] ), .X(n30421) );
  inv_x1_sg U36135 ( .A(n30421), .X(n30422) );
  inv_x1_sg U36136 ( .A(\shifter_0/reg_i_8[9] ), .X(n30423) );
  inv_x1_sg U36137 ( .A(n30423), .X(n30424) );
  inv_x1_sg U36138 ( .A(\shifter_0/reg_i_8[10] ), .X(n30425) );
  inv_x1_sg U36139 ( .A(n30425), .X(n30426) );
  inv_x1_sg U36140 ( .A(\shifter_0/reg_i_8[11] ), .X(n30427) );
  inv_x1_sg U36141 ( .A(n30427), .X(n30428) );
  inv_x1_sg U36142 ( .A(\shifter_0/reg_i_8[12] ), .X(n30429) );
  inv_x1_sg U36143 ( .A(n30429), .X(n30430) );
  inv_x1_sg U36144 ( .A(\shifter_0/reg_i_8[13] ), .X(n30431) );
  inv_x1_sg U36145 ( .A(n30431), .X(n30432) );
  inv_x1_sg U36146 ( .A(\shifter_0/reg_i_8[14] ), .X(n30433) );
  inv_x1_sg U36147 ( .A(n30433), .X(n30434) );
  inv_x1_sg U36148 ( .A(\shifter_0/reg_i_8[15] ), .X(n30435) );
  inv_x1_sg U36149 ( .A(n30435), .X(n30436) );
  inv_x1_sg U36150 ( .A(\shifter_0/reg_i_8[16] ), .X(n30437) );
  inv_x1_sg U36151 ( .A(n30437), .X(n30438) );
  inv_x1_sg U36152 ( .A(\shifter_0/reg_i_8[17] ), .X(n30439) );
  inv_x1_sg U36153 ( .A(n30439), .X(n30440) );
  inv_x1_sg U36154 ( .A(\shifter_0/reg_i_8[18] ), .X(n30441) );
  inv_x1_sg U36155 ( .A(n30441), .X(n30442) );
  inv_x1_sg U36156 ( .A(\shifter_0/reg_i_8[19] ), .X(n30443) );
  inv_x1_sg U36157 ( .A(n30443), .X(n30444) );
  inv_x1_sg U36158 ( .A(n35138), .X(n30445) );
  inv_x1_sg U36159 ( .A(n35137), .X(n30446) );
  inv_x1_sg U36160 ( .A(n35136), .X(n30447) );
  inv_x1_sg U36161 ( .A(n35135), .X(n30448) );
  inv_x1_sg U36162 ( .A(n35134), .X(n30449) );
  inv_x1_sg U36163 ( .A(n35133), .X(n30450) );
  inv_x1_sg U36164 ( .A(n35132), .X(n30451) );
  inv_x1_sg U36165 ( .A(n35131), .X(n30452) );
  inv_x1_sg U36166 ( .A(n35130), .X(n30453) );
  inv_x1_sg U36167 ( .A(n35129), .X(n30454) );
  inv_x1_sg U36168 ( .A(n35128), .X(n30455) );
  inv_x1_sg U36169 ( .A(n35127), .X(n30456) );
  inv_x1_sg U36170 ( .A(n35126), .X(n30457) );
  inv_x1_sg U36171 ( .A(n35125), .X(n30458) );
  inv_x1_sg U36172 ( .A(n35124), .X(n30459) );
  inv_x1_sg U36173 ( .A(n35123), .X(n30460) );
  inv_x1_sg U36174 ( .A(n35122), .X(n30461) );
  inv_x1_sg U36175 ( .A(n35121), .X(n30462) );
  inv_x1_sg U36176 ( .A(n35120), .X(n30463) );
  inv_x1_sg U36177 ( .A(n35119), .X(n30464) );
  inv_x1_sg U36178 ( .A(n35118), .X(n30465) );
  inv_x1_sg U36179 ( .A(n35117), .X(n30466) );
  inv_x1_sg U36180 ( .A(\shifter_0/reg_w_8[0] ), .X(n30467) );
  inv_x1_sg U36181 ( .A(n30467), .X(n30468) );
  inv_x1_sg U36182 ( .A(\shifter_0/reg_w_8[1] ), .X(n30469) );
  inv_x1_sg U36183 ( .A(n30469), .X(n30470) );
  inv_x1_sg U36184 ( .A(\shifter_0/reg_w_8[2] ), .X(n30471) );
  inv_x1_sg U36185 ( .A(n30471), .X(n30472) );
  inv_x1_sg U36186 ( .A(\shifter_0/reg_w_8[3] ), .X(n30473) );
  inv_x1_sg U36187 ( .A(n30473), .X(n30474) );
  inv_x1_sg U36188 ( .A(\shifter_0/reg_w_8[4] ), .X(n30475) );
  inv_x1_sg U36189 ( .A(n30475), .X(n30476) );
  inv_x1_sg U36190 ( .A(\shifter_0/reg_w_8[5] ), .X(n30477) );
  inv_x1_sg U36191 ( .A(n30477), .X(n30478) );
  inv_x1_sg U36192 ( .A(\shifter_0/reg_w_8[6] ), .X(n30479) );
  inv_x1_sg U36193 ( .A(n30479), .X(n30480) );
  inv_x1_sg U36194 ( .A(\shifter_0/reg_w_8[7] ), .X(n30481) );
  inv_x1_sg U36195 ( .A(n30481), .X(n30482) );
  inv_x1_sg U36196 ( .A(\shifter_0/reg_w_8[8] ), .X(n30483) );
  inv_x1_sg U36197 ( .A(n30483), .X(n30484) );
  inv_x1_sg U36198 ( .A(\shifter_0/reg_w_8[9] ), .X(n30485) );
  inv_x1_sg U36199 ( .A(n30485), .X(n30486) );
  inv_x1_sg U36200 ( .A(\shifter_0/reg_w_8[10] ), .X(n30487) );
  inv_x1_sg U36201 ( .A(n30487), .X(n30488) );
  inv_x1_sg U36202 ( .A(\shifter_0/reg_w_8[11] ), .X(n30489) );
  inv_x1_sg U36203 ( .A(n30489), .X(n30490) );
  inv_x1_sg U36204 ( .A(\shifter_0/reg_w_8[12] ), .X(n30491) );
  inv_x1_sg U36205 ( .A(n30491), .X(n30492) );
  inv_x1_sg U36206 ( .A(\shifter_0/reg_w_8[13] ), .X(n30493) );
  inv_x1_sg U36207 ( .A(n30493), .X(n30494) );
  inv_x1_sg U36208 ( .A(\shifter_0/reg_w_8[14] ), .X(n30495) );
  inv_x1_sg U36209 ( .A(n30495), .X(n30496) );
  inv_x1_sg U36210 ( .A(\shifter_0/reg_w_8[15] ), .X(n30497) );
  inv_x1_sg U36211 ( .A(n30497), .X(n30498) );
  inv_x1_sg U36212 ( .A(\shifter_0/reg_w_8[16] ), .X(n30499) );
  inv_x1_sg U36213 ( .A(n30499), .X(n30500) );
  inv_x1_sg U36214 ( .A(\shifter_0/reg_w_8[17] ), .X(n30501) );
  inv_x1_sg U36215 ( .A(n30501), .X(n30502) );
  inv_x1_sg U36216 ( .A(\shifter_0/reg_w_8[18] ), .X(n30503) );
  inv_x1_sg U36217 ( .A(n30503), .X(n30504) );
  inv_x1_sg U36218 ( .A(\shifter_0/reg_w_8[19] ), .X(n30505) );
  inv_x1_sg U36219 ( .A(n30505), .X(n30506) );
  inv_x1_sg U36220 ( .A(n35116), .X(n30507) );
  inv_x1_sg U36221 ( .A(n35115), .X(n30508) );
  inv_x1_sg U36222 ( .A(n35114), .X(n30509) );
  inv_x1_sg U36223 ( .A(n35113), .X(n30510) );
  inv_x1_sg U36224 ( .A(n35112), .X(n30511) );
  inv_x1_sg U36225 ( .A(n35111), .X(n30512) );
  inv_x1_sg U36226 ( .A(n35110), .X(n30513) );
  inv_x1_sg U36227 ( .A(n35109), .X(n30514) );
  inv_x1_sg U36228 ( .A(n35108), .X(n30515) );
  inv_x1_sg U36229 ( .A(n35107), .X(n30516) );
  inv_x1_sg U36230 ( .A(n35106), .X(n30517) );
  inv_x1_sg U36231 ( .A(n35105), .X(n30518) );
  inv_x1_sg U36232 ( .A(n29664), .X(n30519) );
  inv_x1_sg U36233 ( .A(n30519), .X(n30520) );
  inv_x1_sg U36234 ( .A(n28965), .X(n30521) );
  inv_x1_sg U36235 ( .A(n30521), .X(n30522) );
  inv_x1_sg U36236 ( .A(n35104), .X(n30523) );
  inv_x1_sg U36237 ( .A(n35103), .X(n30524) );
  inv_x1_sg U36238 ( .A(n35102), .X(n30525) );
  inv_x1_sg U36239 ( .A(n19579), .X(n30526) );
  inv_x1_sg U36240 ( .A(n30526), .X(n30527) );
  inv_x1_sg U36241 ( .A(n19580), .X(n30528) );
  inv_x1_sg U36242 ( .A(n30528), .X(n30529) );
  inv_x1_sg U36243 ( .A(n14497), .X(n30530) );
  inv_x1_sg U36244 ( .A(n30530), .X(n30531) );
  inv_x1_sg U36245 ( .A(n14496), .X(n30532) );
  inv_x1_sg U36246 ( .A(n30532), .X(n30533) );
  inv_x1_sg U36247 ( .A(n35099), .X(n30534) );
  inv_x1_sg U36248 ( .A(n35098), .X(n30535) );
  inv_x1_sg U36249 ( .A(n19585), .X(n30536) );
  inv_x1_sg U36250 ( .A(n30536), .X(n30537) );
  inv_x1_sg U36251 ( .A(n11664), .X(n30538) );
  inv_x1_sg U36252 ( .A(n30538), .X(n30539) );
  nand_x2_sg U36253 ( .A(n35463), .B(n21304), .X(n30540) );
  nand_x2_sg U36254 ( .A(n35463), .B(n21304), .X(n35605) );
  inv_x1_sg U36255 ( .A(n42407), .X(n30541) );
  nor_x1_sg U36256 ( .A(n26195), .B(reset), .X(n22215) );
  inv_x1_sg U36257 ( .A(n35097), .X(n30542) );
  nand_x1_sg U36258 ( .A(n35582), .B(n15215), .X(n30543) );
  inv_x1_sg U36259 ( .A(n31216), .X(n30544) );
  inv_x1_sg U36260 ( .A(n31574), .X(n30545) );
  inv_x1_sg U36261 ( .A(n13007), .X(n30546) );
  nand_x4_sg U36262 ( .A(n13959), .B(n13960), .X(n13007) );
  inv_x1_sg U36263 ( .A(n13019), .X(n30547) );
  nand_x4_sg U36264 ( .A(n14021), .B(n14022), .X(n13019) );
  inv_x1_sg U36265 ( .A(n13031), .X(n30548) );
  nand_x4_sg U36266 ( .A(n14083), .B(n14084), .X(n13031) );
  inv_x1_sg U36267 ( .A(n13043), .X(n30549) );
  nand_x4_sg U36268 ( .A(n14145), .B(n14146), .X(n13043) );
  inv_x1_sg U36269 ( .A(n13055), .X(n30550) );
  nand_x4_sg U36270 ( .A(n14207), .B(n14208), .X(n13055) );
  inv_x1_sg U36271 ( .A(n12977), .X(n30551) );
  nand_x4_sg U36272 ( .A(n13798), .B(n13799), .X(n12977) );
  inv_x1_sg U36273 ( .A(n12989), .X(n30552) );
  nand_x4_sg U36274 ( .A(n13866), .B(n13867), .X(n12989) );
  inv_x1_sg U36275 ( .A(n13025), .X(n30553) );
  nand_x4_sg U36276 ( .A(n14052), .B(n14053), .X(n13025) );
  inv_x1_sg U36277 ( .A(n13049), .X(n30554) );
  nand_x4_sg U36278 ( .A(n14176), .B(n14177), .X(n13049) );
  inv_x1_sg U36279 ( .A(n13061), .X(n30555) );
  nand_x4_sg U36280 ( .A(n14238), .B(n14239), .X(n13061) );
  inv_x1_sg U36281 ( .A(n13067), .X(n30556) );
  nand_x4_sg U36282 ( .A(n14269), .B(n14270), .X(n13067) );
  inv_x1_sg U36283 ( .A(n13079), .X(n30557) );
  nand_x4_sg U36284 ( .A(n14331), .B(n14332), .X(n13079) );
  inv_x1_sg U36285 ( .A(n13085), .X(n30558) );
  nand_x4_sg U36286 ( .A(n14362), .B(n14363), .X(n13085) );
  inv_x1_sg U36287 ( .A(n13001), .X(n30559) );
  nand_x4_sg U36288 ( .A(n13928), .B(n13929), .X(n13001) );
  inv_x1_sg U36289 ( .A(n13099), .X(n30560) );
  nand_x4_sg U36290 ( .A(n14393), .B(n14394), .X(n13099) );
  inv_x1_sg U36291 ( .A(n13037), .X(n30561) );
  nand_x4_sg U36292 ( .A(n14114), .B(n14115), .X(n13037) );
  inv_x1_sg U36293 ( .A(n13073), .X(n30562) );
  nand_x4_sg U36294 ( .A(n14300), .B(n14301), .X(n13073) );
  inv_x1_sg U36295 ( .A(n35465), .X(n30563) );
  inv_x1_sg U36296 ( .A(n30563), .X(n30564) );
  inv_x1_sg U36297 ( .A(n13114), .X(n30565) );
  nand_x4_sg U36298 ( .A(n14456), .B(n14457), .X(n13114) );
  inv_x1_sg U36299 ( .A(n13114), .X(n35593) );
  inv_x1_sg U36300 ( .A(n12983), .X(n30566) );
  nand_x4_sg U36301 ( .A(n13835), .B(n13836), .X(n12983) );
  inv_x1_sg U36302 ( .A(n12983), .X(n35561) );
  inv_x1_sg U36303 ( .A(n13148), .X(n30567) );
  nand_x4_sg U36304 ( .A(n14644), .B(n14645), .X(n13148) );
  inv_x1_sg U36305 ( .A(n13148), .X(n35506) );
  inv_x1_sg U36306 ( .A(n13225), .X(n30568) );
  nand_x4_sg U36307 ( .A(n15016), .B(n15017), .X(n13225) );
  inv_x1_sg U36308 ( .A(n13225), .X(n35583) );
  inv_x1_sg U36309 ( .A(n13108), .X(n30569) );
  nand_x4_sg U36310 ( .A(n14425), .B(n14426), .X(n13108) );
  inv_x1_sg U36311 ( .A(n13108), .X(n35503) );
  inv_x1_sg U36312 ( .A(n13202), .X(n30570) );
  nand_x4_sg U36313 ( .A(n14923), .B(n14924), .X(n13202) );
  inv_x1_sg U36314 ( .A(n13202), .X(n35512) );
  inv_x1_sg U36315 ( .A(n12995), .X(n30571) );
  nand_x4_sg U36316 ( .A(n13897), .B(n13898), .X(n12995) );
  inv_x1_sg U36317 ( .A(n12995), .X(n35509) );
  inv_x1_sg U36318 ( .A(n13013), .X(n30572) );
  nand_x4_sg U36319 ( .A(n13990), .B(n13991), .X(n13013) );
  inv_x1_sg U36320 ( .A(n13013), .X(n35514) );
  inv_x1_sg U36321 ( .A(n13166), .X(n30573) );
  nand_x4_sg U36322 ( .A(n14737), .B(n14738), .X(n13166) );
  inv_x1_sg U36323 ( .A(n13166), .X(n35513) );
  inv_x1_sg U36324 ( .A(n13184), .X(n30574) );
  nand_x4_sg U36325 ( .A(n14830), .B(n14831), .X(n13184) );
  inv_x1_sg U36326 ( .A(n13184), .X(n35505) );
  inv_x1_sg U36327 ( .A(n13196), .X(n30575) );
  nand_x4_sg U36328 ( .A(n14892), .B(n14893), .X(n13196) );
  inv_x1_sg U36329 ( .A(n13196), .X(n35584) );
  inv_x1_sg U36330 ( .A(n13190), .X(n30576) );
  nand_x4_sg U36331 ( .A(n14861), .B(n14862), .X(n13190) );
  inv_x1_sg U36332 ( .A(n13190), .X(n35585) );
  inv_x1_sg U36333 ( .A(n13178), .X(n30577) );
  nand_x4_sg U36334 ( .A(n14799), .B(n14800), .X(n13178) );
  inv_x1_sg U36335 ( .A(n13178), .X(n35586) );
  inv_x1_sg U36336 ( .A(n13172), .X(n30578) );
  nand_x4_sg U36337 ( .A(n14768), .B(n14769), .X(n13172) );
  inv_x1_sg U36338 ( .A(n13172), .X(n35587) );
  inv_x1_sg U36339 ( .A(n13160), .X(n30579) );
  nand_x4_sg U36340 ( .A(n14706), .B(n14707), .X(n13160) );
  inv_x1_sg U36341 ( .A(n13160), .X(n35588) );
  inv_x1_sg U36342 ( .A(n13154), .X(n30580) );
  nand_x4_sg U36343 ( .A(n14675), .B(n14676), .X(n13154) );
  inv_x1_sg U36344 ( .A(n13154), .X(n35589) );
  inv_x1_sg U36345 ( .A(n13142), .X(n30581) );
  nand_x4_sg U36346 ( .A(n14613), .B(n14614), .X(n13142) );
  inv_x1_sg U36347 ( .A(n13142), .X(n35590) );
  inv_x1_sg U36348 ( .A(n13136), .X(n30582) );
  nand_x4_sg U36349 ( .A(n14582), .B(n14583), .X(n13136) );
  inv_x1_sg U36350 ( .A(n13136), .X(n35591) );
  inv_x1_sg U36351 ( .A(n13125), .X(n30583) );
  nand_x4_sg U36352 ( .A(n14520), .B(n14521), .X(n13125) );
  inv_x1_sg U36353 ( .A(n13125), .X(n35592) );
  inv_x1_sg U36354 ( .A(\filter_0/w_pointer[0] ), .X(n30584) );
  inv_x1_sg U36355 ( .A(n21303), .X(n30585) );
  inv_x1_sg U36356 ( .A(n30590), .X(n30586) );
  inv_x1_sg U36357 ( .A(n35180), .X(n30587) );
  inv_x1_sg U36358 ( .A(n30715), .X(n30588) );
  inv_x1_sg U36359 ( .A(n30715), .X(n30589) );
  inv_x1_sg U36360 ( .A(n35086), .X(n30590) );
  inv_x1_sg U36361 ( .A(n30590), .X(n30591) );
  inv_x1_sg U36362 ( .A(n35365), .X(n30592) );
  inv_x1_sg U36363 ( .A(n35170), .X(n30593) );
  inv_x1_sg U36364 ( .A(n35174), .X(n30594) );
  inv_x1_sg U36365 ( .A(n35188), .X(n30595) );
  inv_x1_sg U36366 ( .A(n30598), .X(n30596) );
  inv_x1_sg U36367 ( .A(n30598), .X(n30597) );
  inv_x1_sg U36368 ( .A(n34937), .X(n30598) );
  inv_x1_sg U36369 ( .A(n30598), .X(n30599) );
  inv_x1_sg U36370 ( .A(n30617), .X(n30600) );
  inv_x1_sg U36371 ( .A(n30545), .X(n30601) );
  inv_x1_sg U36372 ( .A(n30604), .X(n30602) );
  inv_x1_sg U36373 ( .A(n33054), .X(n30603) );
  inv_x1_sg U36374 ( .A(n35010), .X(n30604) );
  inv_x1_sg U36375 ( .A(n35031), .X(n30605) );
  inv_x1_sg U36376 ( .A(n35040), .X(n30606) );
  inv_x1_sg U36377 ( .A(n31219), .X(n30607) );
  inv_x1_sg U36378 ( .A(n34944), .X(n30608) );
  inv_x1_sg U36379 ( .A(n34943), .X(n30609) );
  inv_x1_sg U36380 ( .A(n30609), .X(n30610) );
  inv_x1_sg U36381 ( .A(n30152), .X(n30611) );
  inv_x1_sg U36382 ( .A(n31612), .X(n30612) );
  inv_x1_sg U36383 ( .A(n29682), .X(n30613) );
  inv_x1_sg U36384 ( .A(n31479), .X(n30614) );
  inv_x1_sg U36385 ( .A(n31617), .X(n30615) );
  inv_x1_sg U36386 ( .A(n30600), .X(n30616) );
  inv_x1_sg U36387 ( .A(n35051), .X(n30617) );
  inv_x1_sg U36388 ( .A(n30620), .X(n30618) );
  inv_x1_sg U36389 ( .A(n30618), .X(n30619) );
  inv_x1_sg U36390 ( .A(n31608), .X(n30620) );
  inv_x1_sg U36391 ( .A(n30152), .X(n30621) );
  inv_x1_sg U36392 ( .A(n30624), .X(n30622) );
  inv_x1_sg U36393 ( .A(n34892), .X(n30623) );
  inv_x1_sg U36394 ( .A(n34939), .X(n30624) );
  inv_x1_sg U36395 ( .A(n34887), .X(n30625) );
  inv_x1_sg U36396 ( .A(n34890), .X(n30626) );
  inv_x1_sg U36397 ( .A(n34882), .X(n30627) );
  inv_x1_sg U36398 ( .A(n30627), .X(n30628) );
  inv_x1_sg U36399 ( .A(n34877), .X(n30629) );
  inv_x1_sg U36400 ( .A(n30629), .X(n30630) );
  inv_x1_sg U36401 ( .A(n26350), .X(n30631) );
  inv_x1_sg U36402 ( .A(n30202), .X(n30632) );
  inv_x1_sg U36403 ( .A(n31620), .X(n30633) );
  inv_x1_sg U36404 ( .A(n26352), .X(n30634) );
  inv_x1_sg U36405 ( .A(n35417), .X(n30635) );
  inv_x1_sg U36406 ( .A(n34853), .X(n30636) );
  inv_x1_sg U36407 ( .A(n29756), .X(n30637) );
  inv_x1_sg U36408 ( .A(n34805), .X(n30638) );
  inv_x1_sg U36409 ( .A(n33828), .X(n30639) );
  inv_x1_sg U36410 ( .A(n30643), .X(n30640) );
  inv_x1_sg U36411 ( .A(n34800), .X(n30641) );
  inv_x1_sg U36412 ( .A(n34800), .X(n30642) );
  inv_x1_sg U36413 ( .A(n30642), .X(n30643) );
  inv_x1_sg U36414 ( .A(n34795), .X(n30644) );
  inv_x1_sg U36415 ( .A(n30646), .X(n30645) );
  inv_x1_sg U36416 ( .A(n26219), .X(n30646) );
  inv_x1_sg U36417 ( .A(n30650), .X(n30647) );
  inv_x1_sg U36418 ( .A(n34790), .X(n30648) );
  inv_x1_sg U36419 ( .A(n30672), .X(n30649) );
  inv_x1_sg U36420 ( .A(n30649), .X(n30650) );
  inv_x1_sg U36421 ( .A(n30654), .X(n30651) );
  inv_x1_sg U36422 ( .A(n34785), .X(n30652) );
  inv_x1_sg U36423 ( .A(n32097), .X(n30653) );
  inv_x1_sg U36424 ( .A(n30653), .X(n30654) );
  inv_x1_sg U36425 ( .A(n30658), .X(n30655) );
  inv_x1_sg U36426 ( .A(n34780), .X(n30656) );
  inv_x1_sg U36427 ( .A(n30186), .X(n30657) );
  inv_x1_sg U36428 ( .A(n30657), .X(n30658) );
  inv_x1_sg U36429 ( .A(n30662), .X(n30659) );
  inv_x1_sg U36430 ( .A(n34775), .X(n30660) );
  inv_x1_sg U36431 ( .A(n30185), .X(n30661) );
  inv_x1_sg U36432 ( .A(n30661), .X(n30662) );
  inv_x1_sg U36433 ( .A(n30666), .X(n30663) );
  inv_x1_sg U36434 ( .A(n34770), .X(n30664) );
  inv_x1_sg U36435 ( .A(n32093), .X(n30665) );
  inv_x1_sg U36436 ( .A(n30665), .X(n30666) );
  inv_x1_sg U36437 ( .A(n30670), .X(n30667) );
  inv_x1_sg U36438 ( .A(n34765), .X(n30668) );
  inv_x1_sg U36439 ( .A(n30123), .X(n30669) );
  inv_x1_sg U36440 ( .A(n30669), .X(n30670) );
  inv_x1_sg U36441 ( .A(n34760), .X(n30671) );
  inv_x1_sg U36442 ( .A(n30671), .X(n30672) );
  inv_x1_sg U36443 ( .A(n30672), .X(n30673) );
  inv_x1_sg U36444 ( .A(n34760), .X(n30674) );
  inv_x1_sg U36445 ( .A(n30677), .X(n30675) );
  inv_x1_sg U36446 ( .A(n30679), .X(n30676) );
  inv_x1_sg U36447 ( .A(n34755), .X(n30677) );
  inv_x1_sg U36448 ( .A(n34755), .X(n30678) );
  inv_x1_sg U36449 ( .A(n30678), .X(n30679) );
  inv_x1_sg U36450 ( .A(n29672), .X(n30680) );
  inv_x1_sg U36451 ( .A(n34750), .X(n30681) );
  inv_x1_sg U36452 ( .A(n30189), .X(n30682) );
  inv_x1_sg U36453 ( .A(n30682), .X(n30683) );
  inv_x1_sg U36454 ( .A(n30687), .X(n30684) );
  inv_x1_sg U36455 ( .A(n34745), .X(n30685) );
  inv_x1_sg U36456 ( .A(n30182), .X(n30686) );
  inv_x1_sg U36457 ( .A(n30686), .X(n30687) );
  inv_x1_sg U36458 ( .A(n30691), .X(n30688) );
  inv_x1_sg U36459 ( .A(n34740), .X(n30689) );
  inv_x1_sg U36460 ( .A(n34740), .X(n30690) );
  inv_x1_sg U36461 ( .A(n30690), .X(n30691) );
  inv_x1_sg U36462 ( .A(n30695), .X(n30692) );
  inv_x1_sg U36463 ( .A(n30181), .X(n30693) );
  inv_x1_sg U36464 ( .A(n34735), .X(n30694) );
  inv_x1_sg U36465 ( .A(n30694), .X(n30695) );
  inv_x1_sg U36466 ( .A(n30699), .X(n30696) );
  inv_x1_sg U36467 ( .A(n30683), .X(n30697) );
  inv_x1_sg U36468 ( .A(n30703), .X(n30698) );
  inv_x1_sg U36469 ( .A(n30698), .X(n30699) );
  inv_x1_sg U36470 ( .A(n34962), .X(n30700) );
  inv_x1_sg U36471 ( .A(n30700), .X(n30701) );
  inv_x1_sg U36472 ( .A(n30700), .X(n30702) );
  inv_x1_sg U36473 ( .A(n31236), .X(n30703) );
  inv_x1_sg U36474 ( .A(n34723), .X(n30704) );
  inv_x1_sg U36475 ( .A(n30704), .X(n30705) );
  inv_x1_sg U36476 ( .A(n34722), .X(n30706) );
  inv_x1_sg U36477 ( .A(n30706), .X(n30707) );
  inv_x1_sg U36478 ( .A(n34721), .X(n30708) );
  inv_x1_sg U36479 ( .A(n30708), .X(n30709) );
  inv_x1_sg U36480 ( .A(n31093), .X(n30710) );
  inv_x1_sg U36481 ( .A(n30706), .X(n30711) );
  inv_x1_sg U36482 ( .A(n30708), .X(n30712) );
  inv_x1_sg U36483 ( .A(n30590), .X(n30713) );
  inv_x1_sg U36484 ( .A(n30718), .X(n30714) );
  inv_x1_sg U36485 ( .A(n34711), .X(n30715) );
  inv_x1_sg U36486 ( .A(n30715), .X(n30716) );
  inv_x1_sg U36487 ( .A(n35383), .X(n30717) );
  inv_x1_sg U36488 ( .A(n35343), .X(n30718) );
  inv_x1_sg U36489 ( .A(n34707), .X(n30719) );
  inv_x1_sg U36490 ( .A(n30719), .X(n30720) );
  inv_x1_sg U36491 ( .A(n34706), .X(n30721) );
  inv_x1_sg U36492 ( .A(n30721), .X(n30722) );
  inv_x1_sg U36493 ( .A(n34705), .X(n30723) );
  inv_x1_sg U36494 ( .A(n30723), .X(n30724) );
  inv_x1_sg U36495 ( .A(n35192), .X(n30725) );
  inv_x1_sg U36496 ( .A(n35176), .X(n30726) );
  inv_x1_sg U36497 ( .A(n35190), .X(n30727) );
  inv_x1_sg U36498 ( .A(n30178), .X(n30728) );
  inv_x1_sg U36499 ( .A(n35166), .X(n30729) );
  inv_x1_sg U36500 ( .A(n30780), .X(n30730) );
  inv_x1_sg U36501 ( .A(n34942), .X(n30731) );
  inv_x1_sg U36502 ( .A(n30734), .X(n30732) );
  inv_x1_sg U36503 ( .A(n34689), .X(n30733) );
  inv_x1_sg U36504 ( .A(n35064), .X(n30734) );
  inv_x1_sg U36505 ( .A(n34684), .X(n30735) );
  inv_x1_sg U36506 ( .A(n30737), .X(n30736) );
  inv_x1_sg U36507 ( .A(n35065), .X(n30737) );
  inv_x1_sg U36508 ( .A(n34679), .X(n30738) );
  inv_x1_sg U36509 ( .A(n30740), .X(n30739) );
  inv_x1_sg U36510 ( .A(n35061), .X(n30740) );
  inv_x1_sg U36511 ( .A(n34674), .X(n30741) );
  inv_x1_sg U36512 ( .A(n30743), .X(n30742) );
  inv_x1_sg U36513 ( .A(n35065), .X(n30743) );
  inv_x1_sg U36514 ( .A(n34669), .X(n30744) );
  inv_x1_sg U36515 ( .A(n34669), .X(n30745) );
  inv_x1_sg U36516 ( .A(n30745), .X(n30746) );
  inv_x1_sg U36517 ( .A(n30714), .X(n30747) );
  inv_x1_sg U36518 ( .A(n30880), .X(n30748) );
  inv_x1_sg U36519 ( .A(n34664), .X(n30749) );
  inv_x1_sg U36520 ( .A(n30749), .X(n30750) );
  inv_x1_sg U36521 ( .A(n35393), .X(n30751) );
  inv_x1_sg U36522 ( .A(n30753), .X(n30752) );
  inv_x1_sg U36523 ( .A(n35683), .X(n30753) );
  inv_x1_sg U36524 ( .A(n30779), .X(n30754) );
  inv_x1_sg U36525 ( .A(n30783), .X(n30755) );
  inv_x1_sg U36526 ( .A(n34941), .X(n30756) );
  inv_x1_sg U36527 ( .A(n34644), .X(n30757) );
  inv_x1_sg U36528 ( .A(n30167), .X(n30758) );
  inv_x1_sg U36529 ( .A(n30758), .X(n30759) );
  inv_x1_sg U36530 ( .A(n30166), .X(n30760) );
  inv_x1_sg U36531 ( .A(n30760), .X(n30761) );
  inv_x1_sg U36532 ( .A(n30760), .X(n30762) );
  inv_x1_sg U36533 ( .A(n31922), .X(n30763) );
  inv_x1_sg U36534 ( .A(n34632), .X(n30764) );
  inv_x1_sg U36535 ( .A(n34632), .X(n30765) );
  inv_x1_sg U36536 ( .A(n30765), .X(n30766) );
  inv_x1_sg U36537 ( .A(n30163), .X(n30767) );
  inv_x1_sg U36538 ( .A(n34627), .X(n30768) );
  inv_x1_sg U36539 ( .A(n30768), .X(n30769) );
  inv_x1_sg U36540 ( .A(n34622), .X(n30770) );
  inv_x1_sg U36541 ( .A(n30770), .X(n30771) );
  inv_x1_sg U36542 ( .A(n30771), .X(n30772) );
  inv_x1_sg U36543 ( .A(n30771), .X(n30773) );
  inv_x1_sg U36544 ( .A(n31916), .X(n30774) );
  inv_x1_sg U36545 ( .A(n34605), .X(n30775) );
  inv_x1_sg U36546 ( .A(n34607), .X(n30776) );
  inv_x1_sg U36547 ( .A(n34600), .X(n30777) );
  inv_x1_sg U36548 ( .A(n30777), .X(n30778) );
  inv_x1_sg U36549 ( .A(n32288), .X(n30779) );
  inv_x1_sg U36550 ( .A(n32282), .X(n30780) );
  inv_x1_sg U36551 ( .A(n32283), .X(n30781) );
  inv_x1_sg U36552 ( .A(n34564), .X(n30782) );
  inv_x1_sg U36553 ( .A(n30782), .X(n30783) );
  inv_x1_sg U36554 ( .A(n35263), .X(n30784) );
  inv_x1_sg U36555 ( .A(n34512), .X(n30785) );
  inv_x1_sg U36556 ( .A(n30787), .X(n30786) );
  inv_x1_sg U36557 ( .A(n11716), .X(n30787) );
  inv_x1_sg U36558 ( .A(n30791), .X(n30788) );
  inv_x1_sg U36559 ( .A(n30128), .X(n30789) );
  inv_x1_sg U36560 ( .A(n34507), .X(n30790) );
  inv_x1_sg U36561 ( .A(n30790), .X(n30791) );
  inv_x1_sg U36562 ( .A(n30126), .X(n30792) );
  inv_x1_sg U36563 ( .A(n34502), .X(n30793) );
  inv_x1_sg U36564 ( .A(n30793), .X(n30794) );
  inv_x1_sg U36565 ( .A(n30797), .X(n30795) );
  inv_x1_sg U36566 ( .A(n34497), .X(n30796) );
  inv_x1_sg U36567 ( .A(n30610), .X(n30797) );
  inv_x1_sg U36568 ( .A(n30800), .X(n30798) );
  inv_x1_sg U36569 ( .A(n34492), .X(n30799) );
  inv_x1_sg U36570 ( .A(n30608), .X(n30800) );
  inv_x1_sg U36571 ( .A(n30804), .X(n30801) );
  inv_x1_sg U36572 ( .A(n30122), .X(n30802) );
  inv_x1_sg U36573 ( .A(n34487), .X(n30803) );
  inv_x1_sg U36574 ( .A(n30803), .X(n30804) );
  inv_x1_sg U36575 ( .A(n30808), .X(n30805) );
  inv_x1_sg U36576 ( .A(n30121), .X(n30806) );
  inv_x1_sg U36577 ( .A(n34482), .X(n30807) );
  inv_x1_sg U36578 ( .A(n30807), .X(n30808) );
  inv_x1_sg U36579 ( .A(n30812), .X(n30809) );
  inv_x1_sg U36580 ( .A(n30120), .X(n30810) );
  inv_x1_sg U36581 ( .A(n34477), .X(n30811) );
  inv_x1_sg U36582 ( .A(n30811), .X(n30812) );
  inv_x1_sg U36583 ( .A(n31617), .X(n30813) );
  inv_x1_sg U36584 ( .A(n30817), .X(n30814) );
  inv_x1_sg U36585 ( .A(n34470), .X(n30815) );
  inv_x1_sg U36586 ( .A(n30128), .X(n30816) );
  inv_x1_sg U36587 ( .A(n30816), .X(n30817) );
  inv_x1_sg U36588 ( .A(n30821), .X(n30818) );
  inv_x1_sg U36589 ( .A(n30119), .X(n30819) );
  inv_x1_sg U36590 ( .A(n34465), .X(n30820) );
  inv_x1_sg U36591 ( .A(n30820), .X(n30821) );
  inv_x1_sg U36592 ( .A(n31614), .X(n30822) );
  inv_x1_sg U36593 ( .A(n31615), .X(n30823) );
  inv_x1_sg U36594 ( .A(n30827), .X(n30824) );
  inv_x1_sg U36595 ( .A(n30118), .X(n30825) );
  inv_x1_sg U36596 ( .A(n34458), .X(n30826) );
  inv_x1_sg U36597 ( .A(n30826), .X(n30827) );
  inv_x1_sg U36598 ( .A(n30831), .X(n30828) );
  inv_x1_sg U36599 ( .A(n29902), .X(n30829) );
  inv_x1_sg U36600 ( .A(n34453), .X(n30830) );
  inv_x1_sg U36601 ( .A(n30830), .X(n30831) );
  inv_x1_sg U36602 ( .A(n30120), .X(n30832) );
  inv_x1_sg U36603 ( .A(n35653), .X(n30833) );
  inv_x1_sg U36604 ( .A(n30833), .X(n30834) );
  inv_x1_sg U36605 ( .A(n34446), .X(n30835) );
  inv_x1_sg U36606 ( .A(n11561), .X(n30836) );
  inv_x1_sg U36607 ( .A(n30836), .X(n30837) );
  inv_x1_sg U36608 ( .A(n34441), .X(n30838) );
  inv_x1_sg U36609 ( .A(n30841), .X(n30839) );
  inv_x1_sg U36610 ( .A(n34436), .X(n30840) );
  inv_x1_sg U36611 ( .A(n19582), .X(n30841) );
  inv_x1_sg U36612 ( .A(n35657), .X(n30842) );
  inv_x1_sg U36613 ( .A(n30842), .X(n30843) );
  inv_x1_sg U36614 ( .A(n34431), .X(n30844) );
  inv_x1_sg U36615 ( .A(n30846), .X(n30845) );
  inv_x1_sg U36616 ( .A(n13619), .X(n30846) );
  inv_x1_sg U36617 ( .A(n30848), .X(n30847) );
  inv_x1_sg U36618 ( .A(n11611), .X(n30848) );
  inv_x1_sg U36619 ( .A(n35634), .X(n30849) );
  inv_x1_sg U36620 ( .A(n30849), .X(n30850) );
  inv_x1_sg U36621 ( .A(n34416), .X(n30851) );
  inv_x1_sg U36622 ( .A(n31984), .X(n30852) );
  inv_x1_sg U36623 ( .A(n34107), .X(n30853) );
  inv_x1_sg U36624 ( .A(n30042), .X(n30854) );
  inv_x1_sg U36625 ( .A(n34407), .X(n30855) );
  inv_x1_sg U36626 ( .A(n19591), .X(n30856) );
  inv_x1_sg U36627 ( .A(n34402), .X(n30857) );
  inv_x1_sg U36628 ( .A(n31998), .X(n30858) );
  inv_x1_sg U36629 ( .A(n35389), .X(n30859) );
  inv_x1_sg U36630 ( .A(n35213), .X(n30860) );
  inv_x1_sg U36631 ( .A(n35400), .X(n30861) );
  inv_x1_sg U36632 ( .A(n34084), .X(n30862) );
  inv_x1_sg U36633 ( .A(n30862), .X(n30863) );
  inv_x1_sg U36634 ( .A(n35178), .X(n30864) );
  inv_x1_sg U36635 ( .A(n30862), .X(n30865) );
  inv_x1_sg U36636 ( .A(n30721), .X(n30866) );
  inv_x1_sg U36637 ( .A(n30704), .X(n30867) );
  inv_x1_sg U36638 ( .A(n30704), .X(n30868) );
  inv_x1_sg U36639 ( .A(n29766), .X(n30869) );
  inv_x1_sg U36640 ( .A(n30706), .X(n30870) );
  inv_x1_sg U36641 ( .A(n34074), .X(n30871) );
  inv_x1_sg U36642 ( .A(n30871), .X(n30872) );
  inv_x1_sg U36643 ( .A(n34073), .X(n30873) );
  inv_x1_sg U36644 ( .A(n30873), .X(n30874) );
  inv_x1_sg U36645 ( .A(n30708), .X(n30875) );
  inv_x1_sg U36646 ( .A(n30723), .X(n30876) );
  inv_x1_sg U36647 ( .A(n35352), .X(n30877) );
  inv_x1_sg U36648 ( .A(n35402), .X(n30878) );
  inv_x1_sg U36649 ( .A(n30719), .X(n30879) );
  inv_x1_sg U36650 ( .A(n31489), .X(n30880) );
  inv_x1_sg U36651 ( .A(n30873), .X(n30881) );
  inv_x1_sg U36652 ( .A(n30871), .X(n30882) );
  inv_x1_sg U36653 ( .A(n31026), .X(n30883) );
  inv_x1_sg U36654 ( .A(n31024), .X(n30884) );
  inv_x1_sg U36655 ( .A(n31490), .X(n30885) );
  inv_x1_sg U36656 ( .A(n34048), .X(n30886) );
  inv_x1_sg U36657 ( .A(n30886), .X(n30887) );
  inv_x1_sg U36658 ( .A(n34047), .X(n30888) );
  inv_x1_sg U36659 ( .A(n30888), .X(n30889) );
  inv_x1_sg U36660 ( .A(n34046), .X(n30890) );
  inv_x1_sg U36661 ( .A(n30890), .X(n30891) );
  inv_x1_sg U36662 ( .A(n30893), .X(n30892) );
  inv_x1_sg U36663 ( .A(n31492), .X(n30893) );
  inv_x1_sg U36664 ( .A(n34007), .X(n30894) );
  inv_x1_sg U36665 ( .A(n30894), .X(n30895) );
  inv_x1_sg U36666 ( .A(n34006), .X(n30896) );
  inv_x1_sg U36667 ( .A(n30896), .X(n30897) );
  inv_x1_sg U36668 ( .A(n30900), .X(n30898) );
  inv_x1_sg U36669 ( .A(n30900), .X(n30899) );
  inv_x1_sg U36670 ( .A(n31094), .X(n30900) );
  inv_x1_sg U36671 ( .A(n34002), .X(n30901) );
  inv_x1_sg U36672 ( .A(n30901), .X(n30902) );
  inv_x1_sg U36673 ( .A(n30907), .X(n30903) );
  inv_x1_sg U36674 ( .A(n34000), .X(n30904) );
  inv_x1_sg U36675 ( .A(n30904), .X(n30905) );
  inv_x1_sg U36676 ( .A(n30907), .X(n30906) );
  inv_x1_sg U36677 ( .A(n35227), .X(n30907) );
  inv_x1_sg U36678 ( .A(n30910), .X(n30908) );
  inv_x1_sg U36679 ( .A(n33983), .X(n30909) );
  inv_x1_sg U36680 ( .A(n19590), .X(n30910) );
  inv_x1_sg U36681 ( .A(n26587), .X(n30911) );
  inv_x1_sg U36682 ( .A(n35274), .X(n30912) );
  inv_x1_sg U36683 ( .A(n13699), .X(n30913) );
  inv_x1_sg U36684 ( .A(n34569), .X(n30914) );
  inv_x1_sg U36685 ( .A(n33952), .X(n30915) );
  inv_x1_sg U36686 ( .A(n30915), .X(n30916) );
  inv_x1_sg U36687 ( .A(n33948), .X(n30917) );
  inv_x1_sg U36688 ( .A(n30917), .X(n30918) );
  inv_x1_sg U36689 ( .A(n33947), .X(n30919) );
  inv_x1_sg U36690 ( .A(n30919), .X(n30920) );
  inv_x1_sg U36691 ( .A(n33937), .X(n30921) );
  inv_x1_sg U36692 ( .A(n30921), .X(n30922) );
  inv_x1_sg U36693 ( .A(n33932), .X(n30923) );
  inv_x1_sg U36694 ( .A(n30923), .X(n30924) );
  inv_x1_sg U36695 ( .A(n33927), .X(n30925) );
  inv_x1_sg U36696 ( .A(n30925), .X(n30926) );
  inv_x1_sg U36697 ( .A(n33922), .X(n30927) );
  inv_x1_sg U36698 ( .A(n30927), .X(n30928) );
  inv_x1_sg U36699 ( .A(n33917), .X(n30929) );
  inv_x1_sg U36700 ( .A(n30929), .X(n30930) );
  inv_x1_sg U36701 ( .A(n33910), .X(n30931) );
  inv_x1_sg U36702 ( .A(n30931), .X(n30932) );
  inv_x1_sg U36703 ( .A(n33905), .X(n30933) );
  inv_x1_sg U36704 ( .A(n30933), .X(n30934) );
  inv_x1_sg U36705 ( .A(n33898), .X(n30935) );
  inv_x1_sg U36706 ( .A(n30935), .X(n30936) );
  inv_x1_sg U36707 ( .A(n33891), .X(n30937) );
  inv_x1_sg U36708 ( .A(n30937), .X(n30938) );
  inv_x1_sg U36709 ( .A(n35647), .X(n30939) );
  inv_x1_sg U36710 ( .A(n30939), .X(n30940) );
  inv_x1_sg U36711 ( .A(n33874), .X(n30941) );
  inv_x1_sg U36712 ( .A(n35641), .X(n30942) );
  inv_x1_sg U36713 ( .A(n30942), .X(n30943) );
  inv_x1_sg U36714 ( .A(n33869), .X(n30944) );
  inv_x1_sg U36715 ( .A(n35640), .X(n30945) );
  inv_x1_sg U36716 ( .A(n30945), .X(n30946) );
  inv_x1_sg U36717 ( .A(n33864), .X(n30947) );
  inv_x1_sg U36718 ( .A(n35646), .X(n30948) );
  inv_x1_sg U36719 ( .A(n30948), .X(n30949) );
  inv_x1_sg U36720 ( .A(n33859), .X(n30950) );
  inv_x1_sg U36721 ( .A(n34866), .X(n30951) );
  inv_x1_sg U36722 ( .A(n33854), .X(n30952) );
  inv_x1_sg U36723 ( .A(n33854), .X(n30953) );
  inv_x1_sg U36724 ( .A(n33849), .X(n30954) );
  inv_x1_sg U36725 ( .A(n30954), .X(n30955) );
  inv_x1_sg U36726 ( .A(n33849), .X(n30956) );
  inv_x1_sg U36727 ( .A(n33849), .X(n30957) );
  inv_x1_sg U36728 ( .A(n33844), .X(n30958) );
  inv_x1_sg U36729 ( .A(n30958), .X(n30959) );
  inv_x1_sg U36730 ( .A(n33844), .X(n30960) );
  inv_x1_sg U36731 ( .A(n33844), .X(n30961) );
  inv_x1_sg U36732 ( .A(n30968), .X(n30962) );
  inv_x1_sg U36733 ( .A(n33835), .X(n30963) );
  inv_x1_sg U36734 ( .A(n33835), .X(n30964) );
  inv_x1_sg U36735 ( .A(n33830), .X(n30965) );
  inv_x1_sg U36736 ( .A(n30965), .X(n30966) );
  inv_x1_sg U36737 ( .A(n33830), .X(n30967) );
  inv_x1_sg U36738 ( .A(n33830), .X(n30968) );
  inv_x1_sg U36739 ( .A(n31220), .X(n30969) );
  inv_x1_sg U36740 ( .A(n30969), .X(n30970) );
  inv_x1_sg U36741 ( .A(n30969), .X(n30971) );
  inv_x1_sg U36742 ( .A(n29825), .X(n30972) );
  inv_x1_sg U36743 ( .A(n30972), .X(n30973) );
  inv_x1_sg U36744 ( .A(n30972), .X(n30974) );
  inv_x1_sg U36745 ( .A(n35259), .X(n30975) );
  inv_x1_sg U36746 ( .A(n30975), .X(n30976) );
  inv_x1_sg U36747 ( .A(n33813), .X(n30977) );
  inv_x1_sg U36748 ( .A(n35260), .X(n30978) );
  inv_x1_sg U36749 ( .A(n30978), .X(n30979) );
  inv_x1_sg U36750 ( .A(n33808), .X(n30980) );
  inv_x1_sg U36751 ( .A(n35261), .X(n30981) );
  inv_x1_sg U36752 ( .A(n30981), .X(n30982) );
  inv_x1_sg U36753 ( .A(n33803), .X(n30983) );
  inv_x1_sg U36754 ( .A(n35410), .X(n30984) );
  inv_x1_sg U36755 ( .A(n30984), .X(n30985) );
  inv_x1_sg U36756 ( .A(n33799), .X(n30986) );
  inv_x1_sg U36757 ( .A(n33795), .X(n30987) );
  inv_x1_sg U36758 ( .A(n33758), .X(n30988) );
  inv_x1_sg U36759 ( .A(n33753), .X(n30989) );
  inv_x1_sg U36760 ( .A(n33749), .X(n30990) );
  inv_x1_sg U36761 ( .A(n30980), .X(n30991) );
  inv_x1_sg U36762 ( .A(n33740), .X(n30992) );
  inv_x1_sg U36763 ( .A(n33736), .X(n30993) );
  inv_x1_sg U36764 ( .A(n33732), .X(n30994) );
  inv_x1_sg U36765 ( .A(n30983), .X(n30995) );
  inv_x1_sg U36766 ( .A(n33723), .X(n30996) );
  inv_x1_sg U36767 ( .A(n33719), .X(n30997) );
  inv_x1_sg U36768 ( .A(n33715), .X(n30998) );
  inv_x1_sg U36769 ( .A(n30977), .X(n30999) );
  inv_x1_sg U36770 ( .A(n33634), .X(n31000) );
  inv_x1_sg U36771 ( .A(n33630), .X(n31001) );
  inv_x1_sg U36772 ( .A(n33522), .X(n31002) );
  inv_x1_sg U36773 ( .A(n31101), .X(n31003) );
  inv_x1_sg U36774 ( .A(n31003), .X(n31004) );
  inv_x1_sg U36775 ( .A(n31626), .X(n31005) );
  inv_x1_sg U36776 ( .A(n31004), .X(n31006) );
  inv_x1_sg U36777 ( .A(n31005), .X(n31007) );
  inv_x1_sg U36778 ( .A(n32073), .X(n31008) );
  inv_x1_sg U36779 ( .A(n31008), .X(n31009) );
  inv_x1_sg U36780 ( .A(n31008), .X(n31010) );
  inv_x1_sg U36781 ( .A(n31009), .X(n31011) );
  inv_x1_sg U36782 ( .A(n31010), .X(n31012) );
  inv_x1_sg U36783 ( .A(n29753), .X(n31013) );
  inv_x1_sg U36784 ( .A(n31013), .X(n31014) );
  inv_x1_sg U36785 ( .A(n31013), .X(n31015) );
  inv_x1_sg U36786 ( .A(n31014), .X(n31016) );
  inv_x1_sg U36787 ( .A(n31015), .X(n31017) );
  inv_x1_sg U36788 ( .A(n13224), .X(n31018) );
  inv_x1_sg U36789 ( .A(n34533), .X(n31019) );
  inv_x1_sg U36790 ( .A(n31018), .X(n31020) );
  inv_x1_sg U36791 ( .A(n19589), .X(n31021) );
  inv_x1_sg U36792 ( .A(n31021), .X(n31022) );
  inv_x1_sg U36793 ( .A(n34538), .X(n31023) );
  inv_x1_sg U36794 ( .A(n31873), .X(n31024) );
  inv_x1_sg U36795 ( .A(n31024), .X(n31025) );
  inv_x1_sg U36796 ( .A(n31872), .X(n31026) );
  inv_x1_sg U36797 ( .A(n31026), .X(n31027) );
  inv_x1_sg U36798 ( .A(n31871), .X(n31028) );
  inv_x1_sg U36799 ( .A(n31028), .X(n31029) );
  inv_x1_sg U36800 ( .A(n31870), .X(n31030) );
  inv_x1_sg U36801 ( .A(n31030), .X(n31031) );
  inv_x1_sg U36802 ( .A(n31869), .X(n31032) );
  inv_x1_sg U36803 ( .A(n31032), .X(n31033) );
  inv_x1_sg U36804 ( .A(n31868), .X(n31034) );
  inv_x1_sg U36805 ( .A(n31034), .X(n31035) );
  inv_x1_sg U36806 ( .A(n31865), .X(n31036) );
  inv_x1_sg U36807 ( .A(n31036), .X(n31037) );
  inv_x1_sg U36808 ( .A(n31864), .X(n31038) );
  inv_x1_sg U36809 ( .A(n31038), .X(n31039) );
  inv_x1_sg U36810 ( .A(n31863), .X(n31040) );
  inv_x1_sg U36811 ( .A(n31040), .X(n31041) );
  inv_x1_sg U36812 ( .A(n31862), .X(n31042) );
  inv_x1_sg U36813 ( .A(n31042), .X(n31043) );
  inv_x1_sg U36814 ( .A(n31620), .X(n31044) );
  inv_x1_sg U36815 ( .A(n34868), .X(n31045) );
  inv_x1_sg U36816 ( .A(n31619), .X(n31046) );
  inv_x1_sg U36817 ( .A(n35414), .X(n31047) );
  inv_x1_sg U36818 ( .A(n31047), .X(n31048) );
  inv_x1_sg U36819 ( .A(n33988), .X(n31049) );
  inv_x1_sg U36820 ( .A(n35413), .X(n31050) );
  inv_x1_sg U36821 ( .A(n31050), .X(n31051) );
  inv_x1_sg U36822 ( .A(n33992), .X(n31052) );
  inv_x1_sg U36823 ( .A(n31692), .X(n31053) );
  inv_x1_sg U36824 ( .A(n31053), .X(n31054) );
  inv_x1_sg U36825 ( .A(n31691), .X(n31055) );
  inv_x1_sg U36826 ( .A(n31055), .X(n31056) );
  inv_x1_sg U36827 ( .A(n31690), .X(n31057) );
  inv_x1_sg U36828 ( .A(n31057), .X(n31058) );
  inv_x1_sg U36829 ( .A(n31689), .X(n31059) );
  inv_x1_sg U36830 ( .A(n31059), .X(n31060) );
  inv_x1_sg U36831 ( .A(n34010), .X(n31061) );
  inv_x1_sg U36832 ( .A(n31061), .X(n31062) );
  inv_x1_sg U36833 ( .A(n31061), .X(n31063) );
  inv_x1_sg U36834 ( .A(n31062), .X(n31064) );
  inv_x1_sg U36835 ( .A(n29677), .X(n31065) );
  inv_x1_sg U36836 ( .A(n34015), .X(n31066) );
  inv_x1_sg U36837 ( .A(n31066), .X(n31067) );
  inv_x1_sg U36838 ( .A(n31066), .X(n31068) );
  inv_x1_sg U36839 ( .A(n31067), .X(n31069) );
  inv_x1_sg U36840 ( .A(n29678), .X(n31070) );
  inv_x1_sg U36841 ( .A(n34020), .X(n31071) );
  inv_x1_sg U36842 ( .A(n31071), .X(n31072) );
  inv_x1_sg U36843 ( .A(n31071), .X(n31073) );
  inv_x1_sg U36844 ( .A(n31073), .X(n31074) );
  inv_x1_sg U36845 ( .A(n31072), .X(n31075) );
  inv_x1_sg U36846 ( .A(n34027), .X(n31076) );
  inv_x1_sg U36847 ( .A(n31076), .X(n31077) );
  inv_x1_sg U36848 ( .A(n31076), .X(n31078) );
  inv_x1_sg U36849 ( .A(n31078), .X(n31079) );
  inv_x1_sg U36850 ( .A(n31077), .X(n31080) );
  inv_x1_sg U36851 ( .A(n34032), .X(n31081) );
  inv_x1_sg U36852 ( .A(n31081), .X(n31082) );
  inv_x1_sg U36853 ( .A(n31081), .X(n31083) );
  inv_x1_sg U36854 ( .A(n31083), .X(n31084) );
  inv_x1_sg U36855 ( .A(n31082), .X(n31085) );
  inv_x1_sg U36856 ( .A(n34037), .X(n31086) );
  inv_x1_sg U36857 ( .A(n31086), .X(n31087) );
  inv_x1_sg U36858 ( .A(n31086), .X(n31088) );
  inv_x1_sg U36859 ( .A(n31088), .X(n31089) );
  inv_x1_sg U36860 ( .A(n31087), .X(n31090) );
  inv_x1_sg U36861 ( .A(n31676), .X(n31091) );
  inv_x1_sg U36862 ( .A(n31091), .X(n31092) );
  inv_x1_sg U36863 ( .A(n35369), .X(n31093) );
  inv_x1_sg U36864 ( .A(n35386), .X(n31094) );
  inv_x1_sg U36865 ( .A(n35340), .X(n31095) );
  inv_x1_sg U36866 ( .A(n35324), .X(n31096) );
  inv_x1_sg U36867 ( .A(n35324), .X(n31097) );
  inv_x1_sg U36868 ( .A(n31610), .X(n31098) );
  inv_x1_sg U36869 ( .A(n31612), .X(n31099) );
  inv_x1_sg U36870 ( .A(n31611), .X(n31100) );
  inv_x1_sg U36871 ( .A(n31613), .X(n31101) );
  inv_x1_sg U36872 ( .A(n31615), .X(n31102) );
  inv_x1_sg U36873 ( .A(n31101), .X(n31103) );
  inv_x1_sg U36874 ( .A(n31616), .X(n31104) );
  inv_x1_sg U36875 ( .A(n29686), .X(n31105) );
  inv_x1_sg U36876 ( .A(n31104), .X(n31106) );
  inv_x1_sg U36877 ( .A(n35685), .X(n31107) );
  inv_x1_sg U36878 ( .A(n35415), .X(n31108) );
  inv_x1_sg U36879 ( .A(n35062), .X(n31109) );
  inv_x1_sg U36880 ( .A(n26590), .X(n31110) );
  inv_x1_sg U36881 ( .A(n31588), .X(n31111) );
  inv_x1_sg U36882 ( .A(n35035), .X(n31112) );
  inv_x1_sg U36883 ( .A(n31557), .X(n31113) );
  inv_x1_sg U36884 ( .A(n31113), .X(n31114) );
  inv_x1_sg U36885 ( .A(n31114), .X(n31115) );
  inv_x1_sg U36886 ( .A(n31114), .X(n31116) );
  inv_x1_sg U36887 ( .A(\filter_0/i_pointer[3] ), .X(n31117) );
  inv_x1_sg U36888 ( .A(n31117), .X(n31118) );
  inv_x1_sg U36889 ( .A(n35258), .X(n31119) );
  inv_x1_sg U36890 ( .A(\filter_0/i_pointer[0] ), .X(n31120) );
  inv_x1_sg U36891 ( .A(n31120), .X(n31121) );
  inv_x1_sg U36892 ( .A(\filter_0/w_pointer[3] ), .X(n31122) );
  inv_x1_sg U36893 ( .A(n31122), .X(n31123) );
  inv_x1_sg U36894 ( .A(n35256), .X(n31124) );
  inv_x1_sg U36895 ( .A(\shifter_0/reg_i_7[0] ), .X(n31125) );
  inv_x1_sg U36896 ( .A(n31125), .X(n31126) );
  inv_x1_sg U36897 ( .A(\shifter_0/reg_i_7[1] ), .X(n31127) );
  inv_x1_sg U36898 ( .A(n31127), .X(n31128) );
  inv_x1_sg U36899 ( .A(\shifter_0/reg_i_7[3] ), .X(n31129) );
  inv_x1_sg U36900 ( .A(n31129), .X(n31130) );
  inv_x1_sg U36901 ( .A(n35255), .X(n31131) );
  inv_x1_sg U36902 ( .A(\shifter_0/reg_i_7[5] ), .X(n31132) );
  inv_x1_sg U36903 ( .A(n31132), .X(n31133) );
  inv_x1_sg U36904 ( .A(\shifter_0/reg_i_7[6] ), .X(n31134) );
  inv_x1_sg U36905 ( .A(n31134), .X(n31135) );
  inv_x1_sg U36906 ( .A(\shifter_0/reg_i_7[7] ), .X(n31136) );
  inv_x1_sg U36907 ( .A(n31136), .X(n31137) );
  inv_x1_sg U36908 ( .A(\shifter_0/reg_i_7[8] ), .X(n31138) );
  inv_x1_sg U36909 ( .A(n31138), .X(n31139) );
  inv_x1_sg U36910 ( .A(\shifter_0/reg_i_7[9] ), .X(n31140) );
  inv_x1_sg U36911 ( .A(n31140), .X(n31141) );
  inv_x1_sg U36912 ( .A(\shifter_0/reg_i_7[10] ), .X(n31142) );
  inv_x1_sg U36913 ( .A(n31142), .X(n31143) );
  inv_x1_sg U36914 ( .A(\shifter_0/reg_i_7[11] ), .X(n31144) );
  inv_x1_sg U36915 ( .A(n31144), .X(n31145) );
  inv_x1_sg U36916 ( .A(\shifter_0/reg_i_7[12] ), .X(n31146) );
  inv_x1_sg U36917 ( .A(n31146), .X(n31147) );
  inv_x1_sg U36918 ( .A(\shifter_0/reg_i_7[13] ), .X(n31148) );
  inv_x1_sg U36919 ( .A(n31148), .X(n31149) );
  inv_x1_sg U36920 ( .A(\shifter_0/reg_i_7[14] ), .X(n31150) );
  inv_x1_sg U36921 ( .A(n31150), .X(n31151) );
  inv_x1_sg U36922 ( .A(\shifter_0/reg_i_7[15] ), .X(n31152) );
  inv_x1_sg U36923 ( .A(n31152), .X(n31153) );
  inv_x1_sg U36924 ( .A(\shifter_0/reg_i_7[16] ), .X(n31154) );
  inv_x1_sg U36925 ( .A(n31154), .X(n31155) );
  inv_x1_sg U36926 ( .A(\shifter_0/reg_i_7[19] ), .X(n31156) );
  inv_x1_sg U36927 ( .A(n31156), .X(n31157) );
  inv_x1_sg U36928 ( .A(n35254), .X(n31158) );
  inv_x1_sg U36929 ( .A(n35253), .X(n31159) );
  inv_x1_sg U36930 ( .A(\shifter_0/reg_w_7[0] ), .X(n31160) );
  inv_x1_sg U36931 ( .A(n31160), .X(n31161) );
  inv_x1_sg U36932 ( .A(\shifter_0/reg_w_7[1] ), .X(n31162) );
  inv_x1_sg U36933 ( .A(n31162), .X(n31163) );
  inv_x1_sg U36934 ( .A(\shifter_0/reg_w_7[2] ), .X(n31164) );
  inv_x1_sg U36935 ( .A(n31164), .X(n31165) );
  inv_x1_sg U36936 ( .A(\shifter_0/reg_w_7[3] ), .X(n31166) );
  inv_x1_sg U36937 ( .A(n31166), .X(n31167) );
  inv_x1_sg U36938 ( .A(\shifter_0/reg_w_7[4] ), .X(n31168) );
  inv_x1_sg U36939 ( .A(n31168), .X(n31169) );
  inv_x1_sg U36940 ( .A(\shifter_0/reg_w_7[5] ), .X(n31170) );
  inv_x1_sg U36941 ( .A(n31170), .X(n31171) );
  inv_x1_sg U36942 ( .A(\shifter_0/reg_w_7[6] ), .X(n31172) );
  inv_x1_sg U36943 ( .A(n31172), .X(n31173) );
  inv_x1_sg U36944 ( .A(\shifter_0/reg_w_7[7] ), .X(n31174) );
  inv_x1_sg U36945 ( .A(n31174), .X(n31175) );
  inv_x1_sg U36946 ( .A(\shifter_0/reg_w_7[8] ), .X(n31176) );
  inv_x1_sg U36947 ( .A(n31176), .X(n31177) );
  inv_x1_sg U36948 ( .A(\shifter_0/reg_w_7[9] ), .X(n31178) );
  inv_x1_sg U36949 ( .A(n31178), .X(n31179) );
  inv_x1_sg U36950 ( .A(\shifter_0/reg_w_7[10] ), .X(n31180) );
  inv_x1_sg U36951 ( .A(n31180), .X(n31181) );
  inv_x1_sg U36952 ( .A(\shifter_0/reg_w_7[11] ), .X(n31182) );
  inv_x1_sg U36953 ( .A(n31182), .X(n31183) );
  inv_x1_sg U36954 ( .A(\shifter_0/reg_w_7[12] ), .X(n31184) );
  inv_x1_sg U36955 ( .A(n31184), .X(n31185) );
  inv_x1_sg U36956 ( .A(\shifter_0/reg_w_7[13] ), .X(n31186) );
  inv_x1_sg U36957 ( .A(n31186), .X(n31187) );
  inv_x1_sg U36958 ( .A(\shifter_0/reg_w_7[14] ), .X(n31188) );
  inv_x1_sg U36959 ( .A(n31188), .X(n31189) );
  inv_x1_sg U36960 ( .A(\shifter_0/reg_w_7[15] ), .X(n31190) );
  inv_x1_sg U36961 ( .A(n31190), .X(n31191) );
  inv_x1_sg U36962 ( .A(\shifter_0/reg_w_7[16] ), .X(n31192) );
  inv_x1_sg U36963 ( .A(n31192), .X(n31193) );
  inv_x1_sg U36964 ( .A(\shifter_0/reg_w_7[17] ), .X(n31194) );
  inv_x1_sg U36965 ( .A(n31194), .X(n31195) );
  inv_x1_sg U36966 ( .A(\shifter_0/reg_w_7[18] ), .X(n31196) );
  inv_x1_sg U36967 ( .A(n31196), .X(n31197) );
  inv_x1_sg U36968 ( .A(\shifter_0/reg_w_7[19] ), .X(n31198) );
  inv_x1_sg U36969 ( .A(n31198), .X(n31199) );
  inv_x1_sg U36970 ( .A(n35252), .X(n31200) );
  nand_x8_sg U36971 ( .A(n26574), .B(n35527), .X(n35628) );
  inv_x1_sg U36972 ( .A(n26347), .X(n31202) );
  inv_x1_sg U36973 ( .A(n32002), .X(n31203) );
  inv_x1_sg U36974 ( .A(\filter_0/N12 ), .X(n31204) );
  inv_x1_sg U36975 ( .A(n35684), .X(n31205) );
  inv_x1_sg U36976 ( .A(n35381), .X(n31206) );
  inv_x1_sg U36977 ( .A(n35381), .X(n31207) );
  inv_x1_sg U36978 ( .A(n31109), .X(n31208) );
  inv_x1_sg U36979 ( .A(n31606), .X(n31209) );
  inv_x1_sg U36980 ( .A(n31607), .X(n31210) );
  inv_x1_sg U36981 ( .A(n35056), .X(n31211) );
  inv_x1_sg U36982 ( .A(n30604), .X(n31212) );
  inv_x1_sg U36983 ( .A(n35014), .X(n31213) );
  inv_x1_sg U36984 ( .A(n30564), .X(n31214) );
  inv_x1_sg U36985 ( .A(n30564), .X(n31215) );
  nor_x1_sg U36986 ( .A(n20893), .B(n19609), .X(n31216) );
  inv_x1_sg U36987 ( .A(n29671), .X(n31217) );
  inv_x1_sg U36988 ( .A(n30545), .X(n31218) );
  inv_x1_sg U36989 ( .A(n35248), .X(n31219) );
  inv_x1_sg U36990 ( .A(n31559), .X(n31220) );
  inv_x1_sg U36991 ( .A(n34990), .X(n31221) );
  inv_x1_sg U36992 ( .A(n34991), .X(n31222) );
  inv_x1_sg U36993 ( .A(n31113), .X(n31223) );
  inv_x1_sg U36994 ( .A(n31115), .X(n31224) );
  inv_x1_sg U36995 ( .A(n34972), .X(n31225) );
  inv_x1_sg U36996 ( .A(n31545), .X(n31226) );
  inv_x1_sg U36997 ( .A(n30607), .X(n31227) );
  inv_x1_sg U36998 ( .A(n34969), .X(n31228) );
  inv_x1_sg U36999 ( .A(n31228), .X(n31229) );
  inv_x1_sg U37000 ( .A(n31229), .X(n31230) );
  inv_x1_sg U37001 ( .A(n29679), .X(n31231) );
  inv_x1_sg U37002 ( .A(n31609), .X(n31232) );
  inv_x1_sg U37003 ( .A(n34963), .X(n31233) );
  inv_x1_sg U37004 ( .A(n34956), .X(n31234) );
  inv_x1_sg U37005 ( .A(n31234), .X(n31235) );
  inv_x1_sg U37006 ( .A(n34957), .X(n31236) );
  inv_x1_sg U37007 ( .A(n31607), .X(n31237) );
  inv_x1_sg U37008 ( .A(n35056), .X(n31238) );
  inv_x1_sg U37009 ( .A(n34910), .X(n31239) );
  inv_x1_sg U37010 ( .A(n31239), .X(n31240) );
  inv_x1_sg U37011 ( .A(n31239), .X(n31241) );
  inv_x1_sg U37012 ( .A(n29680), .X(n31242) );
  inv_x1_sg U37013 ( .A(n29680), .X(n31243) );
  inv_x1_sg U37014 ( .A(n34905), .X(n31244) );
  inv_x1_sg U37015 ( .A(n31244), .X(n31245) );
  inv_x1_sg U37016 ( .A(n31244), .X(n31246) );
  inv_x1_sg U37017 ( .A(n29681), .X(n31247) );
  inv_x1_sg U37018 ( .A(n31246), .X(n31248) );
  inv_x1_sg U37019 ( .A(n31253), .X(n31249) );
  inv_x1_sg U37020 ( .A(n34868), .X(n31250) );
  inv_x1_sg U37021 ( .A(n31253), .X(n31251) );
  inv_x1_sg U37022 ( .A(n30202), .X(n31252) );
  inv_x1_sg U37023 ( .A(n26350), .X(n31253) );
  inv_x1_sg U37024 ( .A(n34841), .X(n31254) );
  inv_x1_sg U37025 ( .A(n31254), .X(n31255) );
  inv_x1_sg U37026 ( .A(n31254), .X(n31256) );
  inv_x1_sg U37027 ( .A(n31255), .X(n31257) );
  inv_x1_sg U37028 ( .A(n31255), .X(n31258) );
  inv_x1_sg U37029 ( .A(n34836), .X(n31259) );
  inv_x1_sg U37030 ( .A(n31259), .X(n31260) );
  inv_x1_sg U37031 ( .A(n31259), .X(n31261) );
  inv_x1_sg U37032 ( .A(n31261), .X(n31262) );
  inv_x1_sg U37033 ( .A(n31260), .X(n31263) );
  inv_x1_sg U37034 ( .A(n29899), .X(n31264) );
  inv_x1_sg U37035 ( .A(n31259), .X(n31265) );
  inv_x1_sg U37036 ( .A(n31264), .X(n31266) );
  inv_x1_sg U37037 ( .A(n31264), .X(n31267) );
  inv_x1_sg U37038 ( .A(n34836), .X(n31268) );
  inv_x1_sg U37039 ( .A(n31268), .X(n31269) );
  inv_x1_sg U37040 ( .A(n31268), .X(n31270) );
  inv_x1_sg U37041 ( .A(n30380), .X(n31271) );
  inv_x1_sg U37042 ( .A(n30380), .X(n31272) );
  inv_x1_sg U37043 ( .A(n34822), .X(n31273) );
  inv_x1_sg U37044 ( .A(n31273), .X(n31274) );
  inv_x1_sg U37045 ( .A(n31273), .X(n31275) );
  inv_x1_sg U37046 ( .A(n31274), .X(n31276) );
  inv_x1_sg U37047 ( .A(n30377), .X(n31277) );
  inv_x1_sg U37048 ( .A(n34817), .X(n31278) );
  inv_x1_sg U37049 ( .A(n31278), .X(n31279) );
  inv_x1_sg U37050 ( .A(n31278), .X(n31280) );
  inv_x1_sg U37051 ( .A(n31280), .X(n31281) );
  inv_x1_sg U37052 ( .A(n31280), .X(n31282) );
  inv_x1_sg U37053 ( .A(n35060), .X(n31283) );
  inv_x1_sg U37054 ( .A(n34916), .X(n31284) );
  inv_x1_sg U37055 ( .A(n31284), .X(n31285) );
  inv_x1_sg U37056 ( .A(n31284), .X(n31286) );
  inv_x1_sg U37057 ( .A(n31959), .X(n31287) );
  inv_x1_sg U37058 ( .A(n31287), .X(n31288) );
  inv_x1_sg U37059 ( .A(n31287), .X(n31289) );
  inv_x1_sg U37060 ( .A(n31289), .X(n31290) );
  inv_x1_sg U37061 ( .A(n31289), .X(n31291) );
  inv_x1_sg U37062 ( .A(n35066), .X(n31292) );
  inv_x1_sg U37063 ( .A(n30165), .X(n31293) );
  inv_x1_sg U37064 ( .A(n31110), .X(n31294) );
  inv_x1_sg U37065 ( .A(n31110), .X(n31295) );
  inv_x1_sg U37066 ( .A(n31605), .X(n31296) );
  inv_x1_sg U37067 ( .A(n35071), .X(n31297) );
  inv_x1_sg U37068 ( .A(\shifter_0/pointer[3] ), .X(n31298) );
  inv_x1_sg U37069 ( .A(n31298), .X(n31299) );
  inv_x1_sg U37070 ( .A(n35263), .X(n31300) );
  inv_x1_sg U37071 ( .A(n35416), .X(n31301) );
  inv_x1_sg U37072 ( .A(n31301), .X(n31302) );
  inv_x1_sg U37073 ( .A(n34543), .X(n31303) );
  inv_x1_sg U37074 ( .A(n15053), .X(n31304) );
  inv_x1_sg U37075 ( .A(n34383), .X(n31305) );
  inv_x1_sg U37076 ( .A(n30365), .X(n31306) );
  inv_x1_sg U37077 ( .A(n35483), .X(n31307) );
  inv_x1_sg U37078 ( .A(n34378), .X(n31308) );
  inv_x1_sg U37079 ( .A(n30363), .X(n31309) );
  inv_x1_sg U37080 ( .A(n35458), .X(n31310) );
  inv_x1_sg U37081 ( .A(n34373), .X(n31311) );
  inv_x1_sg U37082 ( .A(n30361), .X(n31312) );
  inv_x1_sg U37083 ( .A(n11641), .X(n31313) );
  inv_x1_sg U37084 ( .A(n34368), .X(n31314) );
  inv_x1_sg U37085 ( .A(n30359), .X(n31315) );
  inv_x1_sg U37086 ( .A(n11536), .X(n31316) );
  inv_x1_sg U37087 ( .A(n34363), .X(n31317) );
  inv_x1_sg U37088 ( .A(n30357), .X(n31318) );
  inv_x1_sg U37089 ( .A(n11586), .X(n31319) );
  inv_x1_sg U37090 ( .A(n34358), .X(n31320) );
  inv_x1_sg U37091 ( .A(n30355), .X(n31321) );
  inv_x1_sg U37092 ( .A(n11562), .X(n31322) );
  inv_x1_sg U37093 ( .A(n34353), .X(n31323) );
  inv_x1_sg U37094 ( .A(n30353), .X(n31324) );
  inv_x1_sg U37095 ( .A(n35631), .X(n31325) );
  inv_x1_sg U37096 ( .A(n34348), .X(n31326) );
  inv_x1_sg U37097 ( .A(n30351), .X(n31327) );
  inv_x1_sg U37098 ( .A(n13368), .X(n31328) );
  inv_x1_sg U37099 ( .A(n34343), .X(n31329) );
  inv_x1_sg U37100 ( .A(n30349), .X(n31330) );
  inv_x1_sg U37101 ( .A(n15187), .X(n31331) );
  inv_x1_sg U37102 ( .A(n34338), .X(n31332) );
  inv_x1_sg U37103 ( .A(n30347), .X(n31333) );
  inv_x1_sg U37104 ( .A(n15047), .X(n31334) );
  inv_x1_sg U37105 ( .A(n34333), .X(n31335) );
  inv_x1_sg U37106 ( .A(n30345), .X(n31336) );
  inv_x1_sg U37107 ( .A(n35595), .X(n31337) );
  inv_x1_sg U37108 ( .A(n34328), .X(n31338) );
  inv_x1_sg U37109 ( .A(n30343), .X(n31339) );
  inv_x1_sg U37110 ( .A(n35596), .X(n31340) );
  inv_x1_sg U37111 ( .A(n34323), .X(n31341) );
  inv_x1_sg U37112 ( .A(n30341), .X(n31342) );
  inv_x1_sg U37113 ( .A(n35597), .X(n31343) );
  inv_x1_sg U37114 ( .A(n34318), .X(n31344) );
  inv_x1_sg U37115 ( .A(n30339), .X(n31345) );
  inv_x1_sg U37116 ( .A(n35598), .X(n31346) );
  inv_x1_sg U37117 ( .A(n34313), .X(n31347) );
  inv_x1_sg U37118 ( .A(n30337), .X(n31348) );
  inv_x1_sg U37119 ( .A(n35599), .X(n31349) );
  inv_x1_sg U37120 ( .A(n34308), .X(n31350) );
  inv_x1_sg U37121 ( .A(n30335), .X(n31351) );
  inv_x1_sg U37122 ( .A(n15046), .X(n31352) );
  inv_x1_sg U37123 ( .A(n34303), .X(n31353) );
  inv_x1_sg U37124 ( .A(n30333), .X(n31354) );
  inv_x1_sg U37125 ( .A(n15050), .X(n31355) );
  inv_x1_sg U37126 ( .A(n34298), .X(n31356) );
  inv_x1_sg U37127 ( .A(n30331), .X(n31357) );
  inv_x1_sg U37128 ( .A(n15179), .X(n31358) );
  inv_x1_sg U37129 ( .A(n34293), .X(n31359) );
  inv_x1_sg U37130 ( .A(n30329), .X(n31360) );
  inv_x1_sg U37131 ( .A(n15184), .X(n31361) );
  inv_x1_sg U37132 ( .A(n34288), .X(n31362) );
  inv_x1_sg U37133 ( .A(n30327), .X(n31363) );
  inv_x1_sg U37134 ( .A(n11535), .X(n31364) );
  inv_x1_sg U37135 ( .A(n34283), .X(n31365) );
  inv_x1_sg U37136 ( .A(n30325), .X(n31366) );
  inv_x1_sg U37137 ( .A(n11667), .X(n31367) );
  inv_x1_sg U37138 ( .A(n34278), .X(n31368) );
  inv_x1_sg U37139 ( .A(n30323), .X(n31369) );
  inv_x1_sg U37140 ( .A(n13367), .X(n31370) );
  inv_x1_sg U37141 ( .A(n34273), .X(n31371) );
  inv_x1_sg U37142 ( .A(n30321), .X(n31372) );
  inv_x1_sg U37143 ( .A(n13804), .X(n31373) );
  inv_x1_sg U37144 ( .A(n34268), .X(n31374) );
  inv_x1_sg U37145 ( .A(n30318), .X(n31375) );
  inv_x1_sg U37146 ( .A(n13805), .X(n31376) );
  inv_x1_sg U37147 ( .A(n34263), .X(n31377) );
  inv_x1_sg U37148 ( .A(n30315), .X(n31378) );
  inv_x1_sg U37149 ( .A(n13816), .X(n31379) );
  inv_x1_sg U37150 ( .A(n34258), .X(n31380) );
  inv_x1_sg U37151 ( .A(n30312), .X(n31381) );
  inv_x1_sg U37152 ( .A(n35650), .X(n31382) );
  inv_x1_sg U37153 ( .A(n34253), .X(n31383) );
  inv_x1_sg U37154 ( .A(n30309), .X(n31384) );
  inv_x1_sg U37155 ( .A(n35632), .X(n31385) );
  inv_x1_sg U37156 ( .A(n34248), .X(n31386) );
  inv_x1_sg U37157 ( .A(n30307), .X(n31387) );
  inv_x1_sg U37158 ( .A(n35630), .X(n31388) );
  inv_x1_sg U37159 ( .A(n34243), .X(n31389) );
  inv_x1_sg U37160 ( .A(n30305), .X(n31390) );
  inv_x1_sg U37161 ( .A(n35629), .X(n31391) );
  inv_x1_sg U37162 ( .A(n34238), .X(n31392) );
  inv_x1_sg U37163 ( .A(n30303), .X(n31393) );
  inv_x1_sg U37164 ( .A(n12533), .X(n31394) );
  inv_x1_sg U37165 ( .A(n34233), .X(n31395) );
  inv_x1_sg U37166 ( .A(n30301), .X(n31396) );
  inv_x1_sg U37167 ( .A(n35633), .X(n31397) );
  inv_x1_sg U37168 ( .A(n34228), .X(n31398) );
  inv_x1_sg U37169 ( .A(n30299), .X(n31399) );
  inv_x1_sg U37170 ( .A(n12531), .X(n31400) );
  inv_x1_sg U37171 ( .A(n34223), .X(n31401) );
  inv_x1_sg U37172 ( .A(n30296), .X(n31402) );
  inv_x1_sg U37173 ( .A(n13787), .X(n31403) );
  inv_x1_sg U37174 ( .A(n34218), .X(n31404) );
  inv_x1_sg U37175 ( .A(n30293), .X(n31405) );
  inv_x1_sg U37176 ( .A(n35645), .X(n31406) );
  inv_x1_sg U37177 ( .A(n34213), .X(n31407) );
  inv_x1_sg U37178 ( .A(n30291), .X(n31408) );
  inv_x1_sg U37179 ( .A(n35644), .X(n31409) );
  inv_x1_sg U37180 ( .A(n34208), .X(n31410) );
  inv_x1_sg U37181 ( .A(n30289), .X(n31411) );
  inv_x1_sg U37182 ( .A(n13808), .X(n31412) );
  inv_x1_sg U37183 ( .A(n34203), .X(n31413) );
  inv_x1_sg U37184 ( .A(n30286), .X(n31414) );
  inv_x1_sg U37185 ( .A(n15037), .X(n31415) );
  inv_x1_sg U37186 ( .A(n34198), .X(n31416) );
  inv_x1_sg U37187 ( .A(n30284), .X(n31417) );
  inv_x1_sg U37188 ( .A(n15038), .X(n31418) );
  inv_x1_sg U37189 ( .A(n34193), .X(n31419) );
  inv_x1_sg U37190 ( .A(n30282), .X(n31420) );
  inv_x1_sg U37191 ( .A(n15039), .X(n31421) );
  inv_x1_sg U37192 ( .A(n34188), .X(n31422) );
  inv_x1_sg U37193 ( .A(n30280), .X(n31423) );
  inv_x1_sg U37194 ( .A(n15170), .X(n31424) );
  inv_x1_sg U37195 ( .A(n34183), .X(n31425) );
  inv_x1_sg U37196 ( .A(n30278), .X(n31426) );
  inv_x1_sg U37197 ( .A(n15172), .X(n31427) );
  inv_x1_sg U37198 ( .A(n34178), .X(n31428) );
  inv_x1_sg U37199 ( .A(n30276), .X(n31429) );
  inv_x1_sg U37200 ( .A(n15049), .X(n31430) );
  inv_x1_sg U37201 ( .A(n34173), .X(n31431) );
  inv_x1_sg U37202 ( .A(n30274), .X(n31432) );
  inv_x1_sg U37203 ( .A(n15055), .X(n31433) );
  inv_x1_sg U37204 ( .A(n34168), .X(n31434) );
  inv_x1_sg U37205 ( .A(n30272), .X(n31435) );
  inv_x1_sg U37206 ( .A(n15182), .X(n31436) );
  inv_x1_sg U37207 ( .A(n34163), .X(n31437) );
  inv_x1_sg U37208 ( .A(n30270), .X(n31438) );
  inv_x1_sg U37209 ( .A(n15190), .X(n31439) );
  inv_x1_sg U37210 ( .A(n34158), .X(n31440) );
  inv_x1_sg U37211 ( .A(n30268), .X(n31441) );
  inv_x1_sg U37212 ( .A(n15044), .X(n31442) );
  inv_x1_sg U37213 ( .A(n34153), .X(n31443) );
  inv_x1_sg U37214 ( .A(n30266), .X(n31444) );
  inv_x1_sg U37215 ( .A(n15048), .X(n31445) );
  inv_x1_sg U37216 ( .A(n34148), .X(n31446) );
  inv_x1_sg U37217 ( .A(n30264), .X(n31447) );
  inv_x1_sg U37218 ( .A(n15177), .X(n31448) );
  inv_x1_sg U37219 ( .A(n34143), .X(n31449) );
  inv_x1_sg U37220 ( .A(n30262), .X(n31450) );
  inv_x1_sg U37221 ( .A(n15180), .X(n31451) );
  inv_x1_sg U37222 ( .A(n34138), .X(n31452) );
  inv_x1_sg U37223 ( .A(n30260), .X(n31453) );
  inv_x1_sg U37224 ( .A(n15181), .X(n31454) );
  inv_x1_sg U37225 ( .A(n34133), .X(n31455) );
  inv_x1_sg U37226 ( .A(n30258), .X(n31456) );
  inv_x1_sg U37227 ( .A(n15171), .X(n31457) );
  inv_x1_sg U37228 ( .A(n34128), .X(n31458) );
  inv_x1_sg U37229 ( .A(n31457), .X(n31459) );
  inv_x1_sg U37230 ( .A(n35461), .X(n31460) );
  inv_x1_sg U37231 ( .A(n11710), .X(n31461) );
  inv_x1_sg U37232 ( .A(n31460), .X(n31462) );
  inv_x1_sg U37233 ( .A(n35462), .X(n31463) );
  inv_x1_sg U37234 ( .A(n11791), .X(n31464) );
  inv_x1_sg U37235 ( .A(n31463), .X(n31465) );
  inv_x1_sg U37236 ( .A(n35464), .X(n31466) );
  inv_x1_sg U37237 ( .A(n11737), .X(n31467) );
  inv_x1_sg U37238 ( .A(n31466), .X(n31468) );
  inv_x1_sg U37239 ( .A(n35606), .X(n31469) );
  inv_x1_sg U37240 ( .A(n35600), .X(n31470) );
  inv_x1_sg U37241 ( .A(n31469), .X(n31471) );
  inv_x1_sg U37242 ( .A(n34107), .X(n31472) );
  inv_x1_sg U37243 ( .A(n34413), .X(n31473) );
  inv_x1_sg U37244 ( .A(n31472), .X(n31474) );
  inv_x1_sg U37245 ( .A(n31473), .X(n31475) );
  inv_x1_sg U37246 ( .A(n31474), .X(n31476) );
  inv_x1_sg U37247 ( .A(n34927), .X(n31477) );
  inv_x1_sg U37248 ( .A(n31477), .X(n31478) );
  inv_x1_sg U37249 ( .A(n31477), .X(n31479) );
  inv_x1_sg U37250 ( .A(n31478), .X(n31480) );
  inv_x1_sg U37251 ( .A(n29682), .X(n31481) );
  inv_x1_sg U37252 ( .A(n34100), .X(n31482) );
  inv_x1_sg U37253 ( .A(n34412), .X(n31483) );
  inv_x1_sg U37254 ( .A(n31482), .X(n31484) );
  inv_x1_sg U37255 ( .A(n31483), .X(n31485) );
  inv_x1_sg U37256 ( .A(n31484), .X(n31486) );
  inv_x1_sg U37257 ( .A(n29684), .X(n31487) );
  inv_x1_sg U37258 ( .A(n31107), .X(n31488) );
  inv_x1_sg U37259 ( .A(n35363), .X(n31489) );
  inv_x1_sg U37260 ( .A(n35349), .X(n31490) );
  inv_x1_sg U37261 ( .A(n35375), .X(n31491) );
  inv_x1_sg U37262 ( .A(n35319), .X(n31492) );
  inv_x1_sg U37263 ( .A(n13221), .X(n31493) );
  inv_x1_sg U37264 ( .A(n30038), .X(n31494) );
  inv_x1_sg U37265 ( .A(n34085), .X(n31495) );
  inv_x1_sg U37266 ( .A(n33982), .X(n31496) );
  inv_x1_sg U37267 ( .A(n31496), .X(n31497) );
  inv_x1_sg U37268 ( .A(n33977), .X(n31498) );
  inv_x1_sg U37269 ( .A(n31498), .X(n31499) );
  inv_x1_sg U37270 ( .A(n33976), .X(n31500) );
  inv_x1_sg U37271 ( .A(n31500), .X(n31501) );
  inv_x1_sg U37272 ( .A(n33972), .X(n31502) );
  inv_x1_sg U37273 ( .A(n31502), .X(n31503) );
  inv_x1_sg U37274 ( .A(n33971), .X(n31504) );
  inv_x1_sg U37275 ( .A(n31504), .X(n31505) );
  inv_x1_sg U37276 ( .A(n30913), .X(n31506) );
  inv_x1_sg U37277 ( .A(n35314), .X(n31507) );
  inv_x1_sg U37278 ( .A(n33951), .X(n31508) );
  inv_x1_sg U37279 ( .A(n31508), .X(n31509) );
  inv_x1_sg U37280 ( .A(n33950), .X(n31510) );
  inv_x1_sg U37281 ( .A(n31510), .X(n31511) );
  inv_x1_sg U37282 ( .A(n33946), .X(n31512) );
  inv_x1_sg U37283 ( .A(n31512), .X(n31513) );
  inv_x1_sg U37284 ( .A(n33945), .X(n31514) );
  inv_x1_sg U37285 ( .A(n31514), .X(n31515) );
  inv_x1_sg U37286 ( .A(n30922), .X(n31516) );
  inv_x1_sg U37287 ( .A(n30922), .X(n31517) );
  inv_x1_sg U37288 ( .A(n30924), .X(n31518) );
  inv_x1_sg U37289 ( .A(n30924), .X(n31519) );
  inv_x1_sg U37290 ( .A(n30926), .X(n31520) );
  inv_x1_sg U37291 ( .A(n30926), .X(n31521) );
  inv_x1_sg U37292 ( .A(n30928), .X(n31522) );
  inv_x1_sg U37293 ( .A(n30928), .X(n31523) );
  inv_x1_sg U37294 ( .A(n30930), .X(n31524) );
  inv_x1_sg U37295 ( .A(n30930), .X(n31525) );
  inv_x1_sg U37296 ( .A(n30932), .X(n31526) );
  inv_x1_sg U37297 ( .A(n30932), .X(n31527) );
  inv_x1_sg U37298 ( .A(n30934), .X(n31528) );
  inv_x1_sg U37299 ( .A(n30934), .X(n31529) );
  inv_x1_sg U37300 ( .A(n30936), .X(n31530) );
  inv_x1_sg U37301 ( .A(n30936), .X(n31531) );
  inv_x1_sg U37302 ( .A(n30938), .X(n31532) );
  inv_x1_sg U37303 ( .A(n30938), .X(n31533) );
  inv_x1_sg U37304 ( .A(n34970), .X(n31534) );
  inv_x1_sg U37305 ( .A(n31545), .X(n31535) );
  inv_x1_sg U37306 ( .A(n34973), .X(n31536) );
  inv_x1_sg U37307 ( .A(n31230), .X(n31537) );
  inv_x1_sg U37308 ( .A(n30607), .X(n31538) );
  inv_x1_sg U37309 ( .A(n34970), .X(n31539) );
  inv_x1_sg U37310 ( .A(n34973), .X(n31540) );
  inv_x1_sg U37311 ( .A(n30607), .X(n31541) );
  inv_x1_sg U37312 ( .A(n34972), .X(n31542) );
  inv_x1_sg U37313 ( .A(n31544), .X(n31543) );
  inv_x1_sg U37314 ( .A(n31229), .X(n31544) );
  inv_x1_sg U37315 ( .A(n29679), .X(n31545) );
  inv_x1_sg U37316 ( .A(n31544), .X(n31546) );
  inv_x1_sg U37317 ( .A(n34973), .X(n31547) );
  inv_x1_sg U37318 ( .A(n31205), .X(n31548) );
  inv_x1_sg U37319 ( .A(n31559), .X(n31549) );
  inv_x1_sg U37320 ( .A(n31558), .X(n31550) );
  inv_x1_sg U37321 ( .A(n31116), .X(n31551) );
  inv_x1_sg U37322 ( .A(n31556), .X(n31552) );
  inv_x1_sg U37323 ( .A(n31205), .X(n31553) );
  inv_x1_sg U37324 ( .A(n34991), .X(n31554) );
  inv_x1_sg U37325 ( .A(n31116), .X(n31555) );
  inv_x1_sg U37326 ( .A(n35684), .X(n31556) );
  inv_x1_sg U37327 ( .A(n31556), .X(n31557) );
  inv_x1_sg U37328 ( .A(n31557), .X(n31558) );
  inv_x1_sg U37329 ( .A(n34969), .X(n31559) );
  inv_x1_sg U37330 ( .A(n35248), .X(n31560) );
  inv_x1_sg U37331 ( .A(n31115), .X(n31561) );
  inv_x1_sg U37332 ( .A(n30601), .X(n31562) );
  inv_x1_sg U37333 ( .A(n31589), .X(n31563) );
  inv_x1_sg U37334 ( .A(n31575), .X(n31564) );
  inv_x1_sg U37335 ( .A(n31218), .X(n31565) );
  inv_x1_sg U37336 ( .A(n35011), .X(n31566) );
  inv_x1_sg U37337 ( .A(n30603), .X(n31567) );
  inv_x1_sg U37338 ( .A(n30601), .X(n31568) );
  inv_x1_sg U37339 ( .A(n31575), .X(n31569) );
  inv_x1_sg U37340 ( .A(n35034), .X(n31570) );
  inv_x1_sg U37341 ( .A(n30604), .X(n31571) );
  inv_x1_sg U37342 ( .A(n35033), .X(n31572) );
  inv_x1_sg U37343 ( .A(n35032), .X(n31573) );
  inv_x1_sg U37344 ( .A(n31216), .X(n31574) );
  inv_x1_sg U37345 ( .A(n35594), .X(n31575) );
  inv_x1_sg U37346 ( .A(n35013), .X(n31576) );
  inv_x1_sg U37347 ( .A(n35012), .X(n31577) );
  inv_x1_sg U37348 ( .A(n30601), .X(n31578) );
  inv_x1_sg U37349 ( .A(n31218), .X(n31579) );
  inv_x1_sg U37350 ( .A(n31588), .X(n31580) );
  inv_x1_sg U37351 ( .A(n31588), .X(n31581) );
  inv_x1_sg U37352 ( .A(n30239), .X(n31582) );
  inv_x1_sg U37353 ( .A(n35011), .X(n31583) );
  inv_x1_sg U37354 ( .A(n35014), .X(n31584) );
  inv_x1_sg U37355 ( .A(n30606), .X(n31585) );
  inv_x1_sg U37356 ( .A(n30606), .X(n31586) );
  inv_x1_sg U37357 ( .A(n31589), .X(n31587) );
  inv_x1_sg U37358 ( .A(n33065), .X(n31588) );
  inv_x1_sg U37359 ( .A(n29671), .X(n31589) );
  inv_x1_sg U37360 ( .A(n30603), .X(n31590) );
  inv_x1_sg U37361 ( .A(n30239), .X(n31591) );
  inv_x1_sg U37362 ( .A(\filter_0/i_pointer[1] ), .X(n31592) );
  inv_x1_sg U37363 ( .A(n31592), .X(n31593) );
  inv_x1_sg U37364 ( .A(n35268), .X(n31594) );
  inv_x1_sg U37365 ( .A(n31670), .X(n31595) );
  inv_x1_sg U37366 ( .A(\shifter_0/i_pointer[1] ), .X(n31596) );
  inv_x1_sg U37367 ( .A(n31596), .X(n31597) );
  inv_x1_sg U37368 ( .A(\shifter_0/pointer[1] ), .X(n31598) );
  inv_x1_sg U37369 ( .A(n31598), .X(n31599) );
  inv_x1_sg U37370 ( .A(n32222), .X(n31600) );
  inv_x1_sg U37371 ( .A(n19600), .X(n31601) );
  inv_x1_sg U37372 ( .A(n42409), .X(n31602) );
  inv_x1_sg U37373 ( .A(n31602), .X(n31603) );
  inv_x1_sg U37374 ( .A(n31602), .X(n31604) );
  inv_x1_sg U37375 ( .A(n26590), .X(n31605) );
  inv_x1_sg U37376 ( .A(n35062), .X(n31606) );
  inv_x1_sg U37377 ( .A(n35415), .X(n31607) );
  inv_x1_sg U37378 ( .A(n35247), .X(n31608) );
  inv_x1_sg U37379 ( .A(n35685), .X(n31609) );
  inv_x1_sg U37380 ( .A(n30121), .X(n31610) );
  inv_x1_sg U37381 ( .A(n31610), .X(n31611) );
  inv_x1_sg U37382 ( .A(n31610), .X(n31612) );
  inv_x1_sg U37383 ( .A(n35455), .X(n31613) );
  inv_x1_sg U37384 ( .A(n31613), .X(n31614) );
  inv_x1_sg U37385 ( .A(n31613), .X(n31615) );
  inv_x1_sg U37386 ( .A(n30118), .X(n31616) );
  inv_x1_sg U37387 ( .A(n31616), .X(n31617) );
  inv_x1_sg U37388 ( .A(n31616), .X(n31618) );
  inv_x1_sg U37389 ( .A(n34867), .X(n31619) );
  inv_x1_sg U37390 ( .A(n34867), .X(n31620) );
  inv_x1_sg U37391 ( .A(n30202), .X(n31621) );
  inv_x1_sg U37392 ( .A(n31620), .X(n31622) );
  inv_x1_sg U37393 ( .A(n31104), .X(n31623) );
  inv_x1_sg U37394 ( .A(n29686), .X(n31624) );
  inv_x1_sg U37395 ( .A(n31615), .X(n31625) );
  inv_x1_sg U37396 ( .A(n31101), .X(n31626) );
  inv_x1_sg U37397 ( .A(n31611), .X(n31627) );
  inv_x1_sg U37398 ( .A(n31098), .X(n31628) );
  inv_x1_sg U37399 ( .A(n33981), .X(n31629) );
  inv_x1_sg U37400 ( .A(n31629), .X(n31630) );
  inv_x1_sg U37401 ( .A(n31629), .X(n31631) );
  inv_x1_sg U37402 ( .A(n33980), .X(n31632) );
  inv_x1_sg U37403 ( .A(n31632), .X(n31633) );
  inv_x1_sg U37404 ( .A(n31632), .X(n31634) );
  inv_x1_sg U37405 ( .A(n33979), .X(n31635) );
  inv_x1_sg U37406 ( .A(n31635), .X(n31636) );
  inv_x1_sg U37407 ( .A(n31635), .X(n31637) );
  inv_x1_sg U37408 ( .A(n33975), .X(n31638) );
  inv_x1_sg U37409 ( .A(n31638), .X(n31639) );
  inv_x1_sg U37410 ( .A(n31638), .X(n31640) );
  inv_x1_sg U37411 ( .A(n33974), .X(n31641) );
  inv_x1_sg U37412 ( .A(n31641), .X(n31642) );
  inv_x1_sg U37413 ( .A(n31641), .X(n31643) );
  inv_x1_sg U37414 ( .A(n33970), .X(n31644) );
  inv_x1_sg U37415 ( .A(n31644), .X(n31645) );
  inv_x1_sg U37416 ( .A(n31644), .X(n31646) );
  inv_x1_sg U37417 ( .A(n30914), .X(n31647) );
  inv_x1_sg U37418 ( .A(n31647), .X(n31648) );
  inv_x1_sg U37419 ( .A(n31647), .X(n31649) );
  inv_x1_sg U37420 ( .A(n30911), .X(n31650) );
  inv_x1_sg U37421 ( .A(n33963), .X(n31651) );
  inv_x1_sg U37422 ( .A(n30912), .X(n31652) );
  inv_x1_sg U37423 ( .A(n33958), .X(n31653) );
  inv_x1_sg U37424 ( .A(\filter_0/N12 ), .X(n31654) );
  inv_x1_sg U37425 ( .A(n31654), .X(n31655) );
  inv_x1_sg U37426 ( .A(n31654), .X(n31656) );
  inv_x1_sg U37427 ( .A(n30584), .X(n31657) );
  inv_x1_sg U37428 ( .A(n30584), .X(n31658) );
  inv_x1_sg U37429 ( .A(n35271), .X(n31659) );
  inv_x1_sg U37430 ( .A(n15052), .X(n31660) );
  inv_x1_sg U37431 ( .A(n31660), .X(n31661) );
  inv_x1_sg U37432 ( .A(n31660), .X(n31662) );
  nand_x1_sg U37433 ( .A(n32169), .B(n32935), .X(n31663) );
  inv_x1_sg U37434 ( .A(n19588), .X(n31664) );
  inv_x1_sg U37435 ( .A(n31664), .X(n31665) );
  inv_x1_sg U37436 ( .A(n31664), .X(n31666) );
  inv_x1_sg U37437 ( .A(n35301), .X(n31667) );
  inv_x1_sg U37438 ( .A(n31667), .X(n31668) );
  inv_x1_sg U37439 ( .A(n31667), .X(n31669) );
  inv_x1_sg U37440 ( .A(n31667), .X(n31670) );
  inv_x1_sg U37441 ( .A(n30880), .X(n31671) );
  inv_x1_sg U37442 ( .A(n30880), .X(n31672) );
  inv_x1_sg U37443 ( .A(n30885), .X(n31673) );
  inv_x1_sg U37444 ( .A(n30885), .X(n31674) );
  inv_x1_sg U37445 ( .A(n30893), .X(n31675) );
  inv_x1_sg U37446 ( .A(n34044), .X(n31676) );
  inv_x1_sg U37447 ( .A(n31088), .X(n31677) );
  inv_x1_sg U37448 ( .A(n31087), .X(n31678) );
  inv_x1_sg U37449 ( .A(n31083), .X(n31679) );
  inv_x1_sg U37450 ( .A(n31082), .X(n31680) );
  inv_x1_sg U37451 ( .A(n31078), .X(n31681) );
  inv_x1_sg U37452 ( .A(n31077), .X(n31682) );
  inv_x1_sg U37453 ( .A(n31073), .X(n31683) );
  inv_x1_sg U37454 ( .A(n31072), .X(n31684) );
  inv_x1_sg U37455 ( .A(n31068), .X(n31685) );
  inv_x1_sg U37456 ( .A(n29678), .X(n31686) );
  inv_x1_sg U37457 ( .A(n31063), .X(n31687) );
  inv_x1_sg U37458 ( .A(n29677), .X(n31688) );
  inv_x1_sg U37459 ( .A(n34003), .X(n31689) );
  inv_x1_sg U37460 ( .A(n34003), .X(n31690) );
  inv_x1_sg U37461 ( .A(n33998), .X(n31691) );
  inv_x1_sg U37462 ( .A(n33998), .X(n31692) );
  inv_x1_sg U37463 ( .A(n33992), .X(n31693) );
  inv_x1_sg U37464 ( .A(n33988), .X(n31694) );
  inv_x1_sg U37465 ( .A(n33983), .X(n31695) );
  inv_x1_sg U37466 ( .A(n30910), .X(n31696) );
  inv_x1_sg U37467 ( .A(\shifter_0/i_pointer[2] ), .X(n31697) );
  inv_x1_sg U37468 ( .A(n31697), .X(n31698) );
  inv_x1_sg U37469 ( .A(n31697), .X(n31699) );
  inv_x1_sg U37470 ( .A(\shifter_0/w_pointer[2] ), .X(n31700) );
  inv_x1_sg U37471 ( .A(n31700), .X(n31701) );
  inv_x1_sg U37472 ( .A(n31700), .X(n31702) );
  inv_x1_sg U37473 ( .A(n32067), .X(n31703) );
  inv_x1_sg U37474 ( .A(n31703), .X(n31704) );
  inv_x1_sg U37475 ( .A(n31703), .X(n31705) );
  inv_x1_sg U37476 ( .A(n31703), .X(n31706) );
  inv_x1_sg U37477 ( .A(n35303), .X(n31707) );
  inv_x1_sg U37478 ( .A(n31707), .X(n31708) );
  inv_x1_sg U37479 ( .A(n31707), .X(n31709) );
  inv_x1_sg U37480 ( .A(n35300), .X(n31710) );
  inv_x1_sg U37481 ( .A(n31710), .X(n31711) );
  inv_x1_sg U37482 ( .A(n31710), .X(n31712) );
  inv_x1_sg U37483 ( .A(n31710), .X(n31713) );
  inv_x1_sg U37484 ( .A(n35299), .X(n31714) );
  inv_x1_sg U37485 ( .A(n31714), .X(n31715) );
  inv_x1_sg U37486 ( .A(n31714), .X(n31716) );
  inv_x1_sg U37487 ( .A(n31714), .X(n31717) );
  inv_x1_sg U37488 ( .A(n35296), .X(n31718) );
  inv_x1_sg U37489 ( .A(n31718), .X(n31719) );
  inv_x1_sg U37490 ( .A(n31718), .X(n31720) );
  inv_x1_sg U37491 ( .A(n31718), .X(n31721) );
  inv_x1_sg U37492 ( .A(n35293), .X(n31722) );
  inv_x1_sg U37493 ( .A(n31722), .X(n31723) );
  inv_x1_sg U37494 ( .A(n31722), .X(n31724) );
  inv_x1_sg U37495 ( .A(n31722), .X(n31725) );
  inv_x1_sg U37496 ( .A(n35292), .X(n31726) );
  inv_x1_sg U37497 ( .A(n31726), .X(n31727) );
  inv_x1_sg U37498 ( .A(n31726), .X(n31728) );
  inv_x1_sg U37499 ( .A(n31726), .X(n31729) );
  inv_x1_sg U37500 ( .A(n35291), .X(n31730) );
  inv_x1_sg U37501 ( .A(n31730), .X(n31731) );
  inv_x1_sg U37502 ( .A(n31730), .X(n31732) );
  inv_x1_sg U37503 ( .A(n31730), .X(n31733) );
  inv_x1_sg U37504 ( .A(n35289), .X(n31734) );
  inv_x1_sg U37505 ( .A(n31734), .X(n31735) );
  inv_x1_sg U37506 ( .A(n31734), .X(n31736) );
  inv_x1_sg U37507 ( .A(n31734), .X(n31737) );
  inv_x1_sg U37508 ( .A(n35287), .X(n31738) );
  inv_x1_sg U37509 ( .A(n31738), .X(n31739) );
  inv_x1_sg U37510 ( .A(n31738), .X(n31740) );
  inv_x1_sg U37511 ( .A(n31738), .X(n31741) );
  inv_x1_sg U37512 ( .A(n35283), .X(n31742) );
  inv_x1_sg U37513 ( .A(n31742), .X(n31743) );
  inv_x1_sg U37514 ( .A(n31742), .X(n31744) );
  inv_x1_sg U37515 ( .A(n31742), .X(n31745) );
  inv_x1_sg U37516 ( .A(n30631), .X(n31746) );
  inv_x1_sg U37517 ( .A(n30631), .X(n31747) );
  inv_x1_sg U37518 ( .A(n34868), .X(n31748) );
  inv_x1_sg U37519 ( .A(n31619), .X(n31749) );
  inv_x1_sg U37520 ( .A(n34407), .X(n31750) );
  inv_x1_sg U37521 ( .A(n30856), .X(n31751) );
  inv_x1_sg U37522 ( .A(n34402), .X(n31752) );
  inv_x1_sg U37523 ( .A(n31304), .X(n31753) );
  inv_x1_sg U37524 ( .A(n31304), .X(n31754) );
  inv_x1_sg U37525 ( .A(n31307), .X(n31755) );
  inv_x1_sg U37526 ( .A(n31307), .X(n31756) );
  inv_x1_sg U37527 ( .A(n31310), .X(n31757) );
  inv_x1_sg U37528 ( .A(n31310), .X(n31758) );
  inv_x1_sg U37529 ( .A(n31313), .X(n31759) );
  inv_x1_sg U37530 ( .A(n31313), .X(n31760) );
  inv_x1_sg U37531 ( .A(n31316), .X(n31761) );
  inv_x1_sg U37532 ( .A(n31316), .X(n31762) );
  inv_x1_sg U37533 ( .A(n31319), .X(n31763) );
  inv_x1_sg U37534 ( .A(n31319), .X(n31764) );
  inv_x1_sg U37535 ( .A(n31322), .X(n31765) );
  inv_x1_sg U37536 ( .A(n31322), .X(n31766) );
  inv_x1_sg U37537 ( .A(n31325), .X(n31767) );
  inv_x1_sg U37538 ( .A(n31325), .X(n31768) );
  inv_x1_sg U37539 ( .A(n31328), .X(n31769) );
  inv_x1_sg U37540 ( .A(n31328), .X(n31770) );
  inv_x1_sg U37541 ( .A(n31331), .X(n31771) );
  inv_x1_sg U37542 ( .A(n31331), .X(n31772) );
  inv_x1_sg U37543 ( .A(n31334), .X(n31773) );
  inv_x1_sg U37544 ( .A(n31334), .X(n31774) );
  inv_x1_sg U37545 ( .A(n31337), .X(n31775) );
  inv_x1_sg U37546 ( .A(n31337), .X(n31776) );
  inv_x1_sg U37547 ( .A(n31340), .X(n31777) );
  inv_x1_sg U37548 ( .A(n31340), .X(n31778) );
  inv_x1_sg U37549 ( .A(n31343), .X(n31779) );
  inv_x1_sg U37550 ( .A(n31343), .X(n31780) );
  inv_x1_sg U37551 ( .A(n31346), .X(n31781) );
  inv_x1_sg U37552 ( .A(n31346), .X(n31782) );
  inv_x1_sg U37553 ( .A(n31349), .X(n31783) );
  inv_x1_sg U37554 ( .A(n31349), .X(n31784) );
  inv_x1_sg U37555 ( .A(n31352), .X(n31785) );
  inv_x1_sg U37556 ( .A(n31352), .X(n31786) );
  inv_x1_sg U37557 ( .A(n31355), .X(n31787) );
  inv_x1_sg U37558 ( .A(n31355), .X(n31788) );
  inv_x1_sg U37559 ( .A(n31358), .X(n31789) );
  inv_x1_sg U37560 ( .A(n31358), .X(n31790) );
  inv_x1_sg U37561 ( .A(n31361), .X(n31791) );
  inv_x1_sg U37562 ( .A(n31361), .X(n31792) );
  inv_x1_sg U37563 ( .A(n31364), .X(n31793) );
  inv_x1_sg U37564 ( .A(n31364), .X(n31794) );
  inv_x1_sg U37565 ( .A(n31367), .X(n31795) );
  inv_x1_sg U37566 ( .A(n31367), .X(n31796) );
  inv_x1_sg U37567 ( .A(n31370), .X(n31797) );
  inv_x1_sg U37568 ( .A(n31370), .X(n31798) );
  inv_x1_sg U37569 ( .A(n31373), .X(n31799) );
  inv_x1_sg U37570 ( .A(n31376), .X(n31800) );
  inv_x1_sg U37571 ( .A(n31379), .X(n31801) );
  inv_x1_sg U37572 ( .A(n31382), .X(n31802) );
  inv_x1_sg U37573 ( .A(n31385), .X(n31803) );
  inv_x1_sg U37574 ( .A(n31385), .X(n31804) );
  inv_x1_sg U37575 ( .A(n31388), .X(n31805) );
  inv_x1_sg U37576 ( .A(n31388), .X(n31806) );
  inv_x1_sg U37577 ( .A(n31391), .X(n31807) );
  inv_x1_sg U37578 ( .A(n31391), .X(n31808) );
  inv_x1_sg U37579 ( .A(n31394), .X(n31809) );
  inv_x1_sg U37580 ( .A(n31394), .X(n31810) );
  inv_x1_sg U37581 ( .A(n31397), .X(n31811) );
  inv_x1_sg U37582 ( .A(n31397), .X(n31812) );
  inv_x1_sg U37583 ( .A(n31400), .X(n31813) );
  inv_x1_sg U37584 ( .A(n31403), .X(n31814) );
  inv_x1_sg U37585 ( .A(n31406), .X(n31815) );
  inv_x1_sg U37586 ( .A(n31406), .X(n31816) );
  inv_x1_sg U37587 ( .A(n31409), .X(n31817) );
  inv_x1_sg U37588 ( .A(n31409), .X(n31818) );
  inv_x1_sg U37589 ( .A(n31412), .X(n31819) );
  inv_x1_sg U37590 ( .A(n31415), .X(n31820) );
  inv_x1_sg U37591 ( .A(n31415), .X(n31821) );
  inv_x1_sg U37592 ( .A(n31418), .X(n31822) );
  inv_x1_sg U37593 ( .A(n31418), .X(n31823) );
  inv_x1_sg U37594 ( .A(n31421), .X(n31824) );
  inv_x1_sg U37595 ( .A(n31421), .X(n31825) );
  inv_x1_sg U37596 ( .A(n31424), .X(n31826) );
  inv_x1_sg U37597 ( .A(n31424), .X(n31827) );
  inv_x1_sg U37598 ( .A(n31427), .X(n31828) );
  inv_x1_sg U37599 ( .A(n31427), .X(n31829) );
  inv_x1_sg U37600 ( .A(n31430), .X(n31830) );
  inv_x1_sg U37601 ( .A(n31430), .X(n31831) );
  inv_x1_sg U37602 ( .A(n31433), .X(n31832) );
  inv_x1_sg U37603 ( .A(n31433), .X(n31833) );
  inv_x1_sg U37604 ( .A(n31436), .X(n31834) );
  inv_x1_sg U37605 ( .A(n31436), .X(n31835) );
  inv_x1_sg U37606 ( .A(n31439), .X(n31836) );
  inv_x1_sg U37607 ( .A(n31439), .X(n31837) );
  inv_x1_sg U37608 ( .A(n31442), .X(n31838) );
  inv_x1_sg U37609 ( .A(n31442), .X(n31839) );
  inv_x1_sg U37610 ( .A(n31445), .X(n31840) );
  inv_x1_sg U37611 ( .A(n31445), .X(n31841) );
  inv_x1_sg U37612 ( .A(n31448), .X(n31842) );
  inv_x1_sg U37613 ( .A(n31448), .X(n31843) );
  inv_x1_sg U37614 ( .A(n31451), .X(n31844) );
  inv_x1_sg U37615 ( .A(n31451), .X(n31845) );
  inv_x1_sg U37616 ( .A(n31454), .X(n31846) );
  inv_x1_sg U37617 ( .A(n31454), .X(n31847) );
  inv_x1_sg U37618 ( .A(n30059), .X(n31848) );
  inv_x1_sg U37619 ( .A(n30059), .X(n31849) );
  inv_x1_sg U37620 ( .A(n30056), .X(n31850) );
  inv_x1_sg U37621 ( .A(n30056), .X(n31851) );
  inv_x1_sg U37622 ( .A(n30053), .X(n31852) );
  inv_x1_sg U37623 ( .A(n30053), .X(n31853) );
  inv_x1_sg U37624 ( .A(n30050), .X(n31854) );
  inv_x1_sg U37625 ( .A(n30050), .X(n31855) );
  inv_x1_sg U37626 ( .A(n30047), .X(n31856) );
  inv_x1_sg U37627 ( .A(n30047), .X(n31857) );
  inv_x1_sg U37628 ( .A(n31474), .X(n31858) );
  inv_x1_sg U37629 ( .A(n31474), .X(n31859) );
  inv_x1_sg U37630 ( .A(n31484), .X(n31860) );
  inv_x1_sg U37631 ( .A(n31484), .X(n31861) );
  inv_x1_sg U37632 ( .A(n34093), .X(n31862) );
  inv_x1_sg U37633 ( .A(n34093), .X(n31863) );
  inv_x1_sg U37634 ( .A(n34090), .X(n31864) );
  inv_x1_sg U37635 ( .A(n34090), .X(n31865) );
  inv_x1_sg U37636 ( .A(n34085), .X(n31866) );
  inv_x1_sg U37637 ( .A(n30038), .X(n31867) );
  inv_x1_sg U37638 ( .A(n34079), .X(n31868) );
  inv_x1_sg U37639 ( .A(n34079), .X(n31869) );
  inv_x1_sg U37640 ( .A(n34075), .X(n31870) );
  inv_x1_sg U37641 ( .A(n34075), .X(n31871) );
  inv_x1_sg U37642 ( .A(n34071), .X(n31872) );
  inv_x1_sg U37643 ( .A(n34071), .X(n31873) );
  inv_x1_sg U37644 ( .A(\filter_0/N16 ), .X(n31874) );
  inv_x1_sg U37645 ( .A(n31874), .X(n31875) );
  inv_x1_sg U37646 ( .A(n31874), .X(n31876) );
  inv_x1_sg U37647 ( .A(\filter_0/w_pointer[1] ), .X(n31877) );
  inv_x1_sg U37648 ( .A(n31877), .X(n31878) );
  inv_x1_sg U37649 ( .A(n31877), .X(n31879) );
  inv_x1_sg U37650 ( .A(n31877), .X(n31880) );
  inv_x1_sg U37651 ( .A(\shifter_0/w_pointer[3] ), .X(n31881) );
  inv_x1_sg U37652 ( .A(n31881), .X(n31882) );
  inv_x1_sg U37653 ( .A(n31881), .X(n31883) );
  inv_x1_sg U37654 ( .A(n31881), .X(n31884) );
  nand_x2_sg U37655 ( .A(n29668), .B(n42410), .X(n31885) );
  nand_x4_sg U37656 ( .A(n29668), .B(n42410), .X(n31886) );
  nand_x8_sg U37657 ( .A(n29668), .B(n42410), .X(n26584) );
  inv_x1_sg U37658 ( .A(n35297), .X(n31887) );
  inv_x1_sg U37659 ( .A(n31887), .X(n31888) );
  inv_x1_sg U37660 ( .A(n31887), .X(n31889) );
  inv_x1_sg U37661 ( .A(n31887), .X(n31890) );
  inv_x1_sg U37662 ( .A(n35286), .X(n31891) );
  inv_x1_sg U37663 ( .A(n31891), .X(n31892) );
  inv_x1_sg U37664 ( .A(n31891), .X(n31893) );
  inv_x1_sg U37665 ( .A(n31891), .X(n31894) );
  inv_x1_sg U37666 ( .A(n35285), .X(n31895) );
  inv_x1_sg U37667 ( .A(n31895), .X(n31896) );
  inv_x1_sg U37668 ( .A(n31895), .X(n31897) );
  inv_x1_sg U37669 ( .A(n31895), .X(n31898) );
  inv_x1_sg U37670 ( .A(n35282), .X(n31899) );
  inv_x1_sg U37671 ( .A(n31899), .X(n31900) );
  inv_x1_sg U37672 ( .A(n31899), .X(n31901) );
  inv_x1_sg U37673 ( .A(n31899), .X(n31902) );
  inv_x1_sg U37674 ( .A(n32338), .X(n31903) );
  inv_x1_sg U37675 ( .A(n31903), .X(n31904) );
  inv_x1_sg U37676 ( .A(n31903), .X(n31905) );
  inv_x1_sg U37677 ( .A(n31903), .X(n31906) );
  inv_x1_sg U37678 ( .A(n32337), .X(n31907) );
  inv_x1_sg U37679 ( .A(n31907), .X(n31908) );
  inv_x1_sg U37680 ( .A(n31907), .X(n31909) );
  inv_x1_sg U37681 ( .A(n31907), .X(n31910) );
  inv_x1_sg U37682 ( .A(n31605), .X(n31911) );
  inv_x1_sg U37683 ( .A(n35071), .X(n31912) );
  inv_x1_sg U37684 ( .A(n26590), .X(n31913) );
  inv_x1_sg U37685 ( .A(n31913), .X(n31914) );
  inv_x1_sg U37686 ( .A(n31913), .X(n31915) );
  inv_x1_sg U37687 ( .A(n31913), .X(n31916) );
  inv_x1_sg U37688 ( .A(n31606), .X(n31917) );
  inv_x1_sg U37689 ( .A(n35066), .X(n31918) );
  inv_x1_sg U37690 ( .A(n31293), .X(n31919) );
  inv_x1_sg U37691 ( .A(n31919), .X(n31920) );
  inv_x1_sg U37692 ( .A(n31919), .X(n31921) );
  inv_x1_sg U37693 ( .A(n31919), .X(n31922) );
  inv_x1_sg U37694 ( .A(n34900), .X(n31923) );
  inv_x1_sg U37695 ( .A(n31923), .X(n31924) );
  inv_x1_sg U37696 ( .A(n31923), .X(n31925) );
  inv_x1_sg U37697 ( .A(n31923), .X(n31926) );
  inv_x1_sg U37698 ( .A(n30791), .X(n31927) );
  inv_x1_sg U37699 ( .A(n30791), .X(n31928) );
  inv_x1_sg U37700 ( .A(n30797), .X(n31929) );
  inv_x1_sg U37701 ( .A(n34497), .X(n31930) );
  inv_x1_sg U37702 ( .A(n30800), .X(n31931) );
  inv_x1_sg U37703 ( .A(n34492), .X(n31932) );
  inv_x1_sg U37704 ( .A(n30804), .X(n31933) );
  inv_x1_sg U37705 ( .A(n30804), .X(n31934) );
  inv_x1_sg U37706 ( .A(n34488), .X(n31935) );
  inv_x1_sg U37707 ( .A(n31935), .X(n31936) );
  inv_x1_sg U37708 ( .A(n31935), .X(n31937) );
  inv_x1_sg U37709 ( .A(n31935), .X(n31938) );
  inv_x1_sg U37710 ( .A(n30808), .X(n31939) );
  inv_x1_sg U37711 ( .A(n30808), .X(n31940) );
  inv_x1_sg U37712 ( .A(n34483), .X(n31941) );
  inv_x1_sg U37713 ( .A(n31941), .X(n31942) );
  inv_x1_sg U37714 ( .A(n31941), .X(n31943) );
  inv_x1_sg U37715 ( .A(n31941), .X(n31944) );
  inv_x1_sg U37716 ( .A(n30812), .X(n31945) );
  inv_x1_sg U37717 ( .A(n30812), .X(n31946) );
  inv_x1_sg U37718 ( .A(n34478), .X(n31947) );
  inv_x1_sg U37719 ( .A(n31947), .X(n31948) );
  inv_x1_sg U37720 ( .A(n31947), .X(n31949) );
  inv_x1_sg U37721 ( .A(n31947), .X(n31950) );
  inv_x1_sg U37722 ( .A(n30817), .X(n31951) );
  inv_x1_sg U37723 ( .A(n30817), .X(n31952) );
  inv_x1_sg U37724 ( .A(n34471), .X(n31953) );
  inv_x1_sg U37725 ( .A(n31953), .X(n31954) );
  inv_x1_sg U37726 ( .A(n31953), .X(n31955) );
  inv_x1_sg U37727 ( .A(n31953), .X(n31956) );
  inv_x1_sg U37728 ( .A(n30821), .X(n31957) );
  inv_x1_sg U37729 ( .A(n30821), .X(n31958) );
  inv_x1_sg U37730 ( .A(n34466), .X(n31959) );
  inv_x1_sg U37731 ( .A(n31959), .X(n31960) );
  inv_x1_sg U37732 ( .A(n31959), .X(n31961) );
  inv_x1_sg U37733 ( .A(n31959), .X(n31962) );
  inv_x1_sg U37734 ( .A(n30827), .X(n31963) );
  inv_x1_sg U37735 ( .A(n30827), .X(n31964) );
  inv_x1_sg U37736 ( .A(n34459), .X(n31965) );
  inv_x1_sg U37737 ( .A(n31965), .X(n31966) );
  inv_x1_sg U37738 ( .A(n31965), .X(n31967) );
  inv_x1_sg U37739 ( .A(n31965), .X(n31968) );
  inv_x1_sg U37740 ( .A(n30831), .X(n31969) );
  inv_x1_sg U37741 ( .A(n30831), .X(n31970) );
  inv_x1_sg U37742 ( .A(n34454), .X(n31971) );
  inv_x1_sg U37743 ( .A(n31971), .X(n31972) );
  inv_x1_sg U37744 ( .A(n31971), .X(n31973) );
  inv_x1_sg U37745 ( .A(n31971), .X(n31974) );
  inv_x1_sg U37746 ( .A(n34436), .X(n31975) );
  inv_x1_sg U37747 ( .A(n30841), .X(n31976) );
  inv_x1_sg U37748 ( .A(n34437), .X(n31977) );
  inv_x1_sg U37749 ( .A(n31977), .X(n31978) );
  inv_x1_sg U37750 ( .A(n31977), .X(n31979) );
  inv_x1_sg U37751 ( .A(n31977), .X(n31980) );
  inv_x1_sg U37752 ( .A(n30849), .X(n31981) );
  inv_x1_sg U37753 ( .A(n34416), .X(n31982) );
  inv_x1_sg U37754 ( .A(n30849), .X(n31983) );
  inv_x1_sg U37755 ( .A(n34416), .X(n31984) );
  inv_x1_sg U37756 ( .A(n30042), .X(n31985) );
  inv_x1_sg U37757 ( .A(n34107), .X(n31986) );
  inv_x1_sg U37758 ( .A(n34414), .X(n31987) );
  inv_x1_sg U37759 ( .A(n31987), .X(n31988) );
  inv_x1_sg U37760 ( .A(n31987), .X(n31989) );
  inv_x1_sg U37761 ( .A(n31987), .X(n31990) );
  inv_x1_sg U37762 ( .A(n34408), .X(n31991) );
  inv_x1_sg U37763 ( .A(n31991), .X(n31992) );
  inv_x1_sg U37764 ( .A(n31991), .X(n31993) );
  inv_x1_sg U37765 ( .A(n31991), .X(n31994) );
  inv_x1_sg U37766 ( .A(n34404), .X(n31995) );
  inv_x1_sg U37767 ( .A(n31995), .X(n31996) );
  inv_x1_sg U37768 ( .A(n31995), .X(n31997) );
  inv_x1_sg U37769 ( .A(n31995), .X(n31998) );
  inv_x1_sg U37770 ( .A(\filter_0/N15 ), .X(n31999) );
  inv_x1_sg U37771 ( .A(n31999), .X(n32000) );
  inv_x1_sg U37772 ( .A(n31999), .X(n32001) );
  inv_x1_sg U37773 ( .A(n31999), .X(n32002) );
  inv_x1_sg U37774 ( .A(\shifter_0/i_pointer[3] ), .X(n32003) );
  inv_x1_sg U37775 ( .A(n32003), .X(n32004) );
  inv_x1_sg U37776 ( .A(n32003), .X(n32005) );
  inv_x1_sg U37777 ( .A(n32003), .X(n32006) );
  inv_x1_sg U37778 ( .A(n35313), .X(n32009) );
  inv_x1_sg U37779 ( .A(n32009), .X(n32010) );
  inv_x1_sg U37780 ( .A(n32009), .X(n32011) );
  inv_x1_sg U37781 ( .A(n32009), .X(n32012) );
  inv_x1_sg U37782 ( .A(n35311), .X(n32013) );
  inv_x1_sg U37783 ( .A(n32013), .X(n32014) );
  inv_x1_sg U37784 ( .A(n32013), .X(n32015) );
  inv_x1_sg U37785 ( .A(n32013), .X(n32016) );
  inv_x1_sg U37786 ( .A(n35310), .X(n32017) );
  inv_x1_sg U37787 ( .A(n32017), .X(n32018) );
  inv_x1_sg U37788 ( .A(n32017), .X(n32019) );
  inv_x1_sg U37789 ( .A(n32017), .X(n32020) );
  inv_x1_sg U37790 ( .A(n30038), .X(n32021) );
  inv_x1_sg U37791 ( .A(n32021), .X(n32022) );
  inv_x1_sg U37792 ( .A(n32021), .X(n32023) );
  inv_x1_sg U37793 ( .A(n32021), .X(n32024) );
  inv_x1_sg U37794 ( .A(n35294), .X(n32025) );
  inv_x1_sg U37795 ( .A(n32025), .X(n32026) );
  inv_x1_sg U37796 ( .A(n32025), .X(n32027) );
  inv_x1_sg U37797 ( .A(n32025), .X(n32028) );
  inv_x1_sg U37798 ( .A(n35288), .X(n32029) );
  inv_x1_sg U37799 ( .A(n32029), .X(n32030) );
  inv_x1_sg U37800 ( .A(n32029), .X(n32031) );
  inv_x1_sg U37801 ( .A(n32029), .X(n32032) );
  inv_x1_sg U37802 ( .A(n35281), .X(n32033) );
  inv_x1_sg U37803 ( .A(n32033), .X(n32034) );
  inv_x1_sg U37804 ( .A(n32033), .X(n32035) );
  inv_x1_sg U37805 ( .A(n32033), .X(n32036) );
  inv_x1_sg U37806 ( .A(n35276), .X(n32037) );
  inv_x1_sg U37807 ( .A(n35276), .X(n32038) );
  inv_x1_sg U37808 ( .A(n35275), .X(n32039) );
  inv_x1_sg U37809 ( .A(n32039), .X(n32040) );
  inv_x1_sg U37810 ( .A(n32039), .X(n32041) );
  inv_x1_sg U37811 ( .A(n32039), .X(n32042) );
  inv_x1_sg U37812 ( .A(n35156), .X(n32043) );
  inv_x1_sg U37813 ( .A(n32043), .X(n32044) );
  inv_x1_sg U37814 ( .A(n32043), .X(n32045) );
  inv_x1_sg U37815 ( .A(n32043), .X(n32046) );
  inv_x1_sg U37816 ( .A(n35155), .X(n32047) );
  inv_x1_sg U37817 ( .A(n32047), .X(n32048) );
  inv_x1_sg U37818 ( .A(n32047), .X(n32049) );
  inv_x1_sg U37819 ( .A(n32047), .X(n32050) );
  inv_x1_sg U37820 ( .A(n35157), .X(n32051) );
  inv_x1_sg U37821 ( .A(n35157), .X(n32052) );
  inv_x1_sg U37822 ( .A(n31301), .X(n32053) );
  inv_x1_sg U37823 ( .A(n34543), .X(n32054) );
  inv_x1_sg U37824 ( .A(n31598), .X(n32055) );
  inv_x1_sg U37825 ( .A(n32055), .X(n32056) );
  inv_x1_sg U37826 ( .A(n32055), .X(n32057) );
  inv_x1_sg U37827 ( .A(n32055), .X(n32058) );
  inv_x1_sg U37828 ( .A(n29676), .X(n32059) );
  inv_x1_sg U37829 ( .A(n34538), .X(n32060) );
  inv_x1_sg U37830 ( .A(n31022), .X(n32061) );
  inv_x1_sg U37831 ( .A(n32061), .X(n32062) );
  inv_x1_sg U37832 ( .A(n32061), .X(n32063) );
  inv_x1_sg U37833 ( .A(n32061), .X(n32064) );
  inv_x1_sg U37834 ( .A(n34533), .X(n32065) );
  inv_x1_sg U37835 ( .A(n31018), .X(n32066) );
  inv_x1_sg U37836 ( .A(n34534), .X(n32067) );
  inv_x1_sg U37837 ( .A(n32067), .X(n32068) );
  inv_x1_sg U37838 ( .A(n32067), .X(n32069) );
  inv_x1_sg U37839 ( .A(n32067), .X(n32070) );
  inv_x1_sg U37840 ( .A(n31015), .X(n32071) );
  inv_x1_sg U37841 ( .A(n31015), .X(n32072) );
  inv_x1_sg U37842 ( .A(n30132), .X(n32073) );
  inv_x1_sg U37843 ( .A(n32073), .X(n32074) );
  inv_x1_sg U37844 ( .A(n32073), .X(n32075) );
  inv_x1_sg U37845 ( .A(n32073), .X(n32076) );
  inv_x1_sg U37846 ( .A(n31010), .X(n32077) );
  inv_x1_sg U37847 ( .A(n31009), .X(n32078) );
  inv_x1_sg U37848 ( .A(n34525), .X(n32079) );
  inv_x1_sg U37849 ( .A(n32079), .X(n32080) );
  inv_x1_sg U37850 ( .A(n32079), .X(n32081) );
  inv_x1_sg U37851 ( .A(n32079), .X(n32082) );
  inv_x1_sg U37852 ( .A(n31005), .X(n32083) );
  inv_x1_sg U37853 ( .A(n31004), .X(n32084) );
  inv_x1_sg U37854 ( .A(n34521), .X(n32085) );
  inv_x1_sg U37855 ( .A(n32085), .X(n32086) );
  inv_x1_sg U37856 ( .A(n32085), .X(n32087) );
  inv_x1_sg U37857 ( .A(n32085), .X(n32088) );
  inv_x1_sg U37858 ( .A(n34508), .X(n32089) );
  inv_x1_sg U37859 ( .A(n32089), .X(n32090) );
  inv_x1_sg U37860 ( .A(n32089), .X(n32091) );
  inv_x1_sg U37861 ( .A(n32089), .X(n32092) );
  inv_x1_sg U37862 ( .A(n34943), .X(n32093) );
  inv_x1_sg U37863 ( .A(n32093), .X(n32094) );
  inv_x1_sg U37864 ( .A(n32093), .X(n32095) );
  inv_x1_sg U37865 ( .A(n32093), .X(n32096) );
  inv_x1_sg U37866 ( .A(n30660), .X(n32097) );
  inv_x1_sg U37867 ( .A(n32097), .X(n32098) );
  inv_x1_sg U37868 ( .A(n32097), .X(n32099) );
  inv_x1_sg U37869 ( .A(n32097), .X(n32100) );
  inv_x1_sg U37870 ( .A(n30846), .X(n32101) );
  inv_x1_sg U37871 ( .A(n34426), .X(n32102) );
  inv_x1_sg U37872 ( .A(n32102), .X(n32103) );
  inv_x1_sg U37873 ( .A(n32103), .X(n32104) );
  inv_x1_sg U37874 ( .A(n32103), .X(n32105) );
  inv_x1_sg U37875 ( .A(n32103), .X(n32106) );
  inv_x1_sg U37876 ( .A(n30848), .X(n32107) );
  inv_x1_sg U37877 ( .A(n34421), .X(n32108) );
  inv_x1_sg U37878 ( .A(n34425), .X(n32109) );
  inv_x1_sg U37879 ( .A(n32109), .X(n32110) );
  inv_x1_sg U37880 ( .A(n32109), .X(n32111) );
  inv_x1_sg U37881 ( .A(n32109), .X(n32112) );
  inv_x1_sg U37882 ( .A(n15104), .X(n32113) );
  inv_x1_sg U37883 ( .A(n32113), .X(n32114) );
  inv_x1_sg U37884 ( .A(n32113), .X(n32115) );
  inv_x1_sg U37885 ( .A(n32113), .X(n32116) );
  inv_x1_sg U37886 ( .A(n15090), .X(n32117) );
  inv_x1_sg U37887 ( .A(n32117), .X(n32118) );
  inv_x1_sg U37888 ( .A(n32117), .X(n32119) );
  inv_x1_sg U37889 ( .A(n32117), .X(n32120) );
  inv_x1_sg U37890 ( .A(n15093), .X(n32121) );
  inv_x1_sg U37891 ( .A(n32121), .X(n32122) );
  inv_x1_sg U37892 ( .A(n32121), .X(n32123) );
  inv_x1_sg U37893 ( .A(n32121), .X(n32124) );
  inv_x1_sg U37894 ( .A(n15095), .X(n32125) );
  inv_x1_sg U37895 ( .A(n32125), .X(n32126) );
  inv_x1_sg U37896 ( .A(n32125), .X(n32127) );
  inv_x1_sg U37897 ( .A(n32125), .X(n32128) );
  inv_x1_sg U37898 ( .A(n15089), .X(n32129) );
  inv_x1_sg U37899 ( .A(n32129), .X(n32130) );
  inv_x1_sg U37900 ( .A(n32129), .X(n32131) );
  inv_x1_sg U37901 ( .A(n32129), .X(n32132) );
  inv_x1_sg U37902 ( .A(n15101), .X(n32133) );
  inv_x1_sg U37903 ( .A(n32133), .X(n32134) );
  inv_x1_sg U37904 ( .A(n32133), .X(n32135) );
  inv_x1_sg U37905 ( .A(n32133), .X(n32136) );
  inv_x1_sg U37906 ( .A(n34897), .X(n32137) );
  inv_x1_sg U37907 ( .A(n32137), .X(n32138) );
  inv_x1_sg U37908 ( .A(n32137), .X(n32139) );
  inv_x1_sg U37909 ( .A(n32137), .X(n32140) );
  inv_x1_sg U37910 ( .A(n32137), .X(n32141) );
  inv_x1_sg U37911 ( .A(n34595), .X(n32142) );
  inv_x1_sg U37912 ( .A(n32142), .X(n32143) );
  inv_x1_sg U37913 ( .A(n32142), .X(n32144) );
  inv_x1_sg U37914 ( .A(n32142), .X(n32145) );
  inv_x1_sg U37915 ( .A(n32142), .X(n32146) );
  inv_x1_sg U37916 ( .A(n34590), .X(n32147) );
  inv_x1_sg U37917 ( .A(n32147), .X(n32148) );
  inv_x1_sg U37918 ( .A(n32147), .X(n32149) );
  inv_x1_sg U37919 ( .A(n32147), .X(n32150) );
  inv_x1_sg U37920 ( .A(n32147), .X(n32151) );
  inv_x1_sg U37921 ( .A(n32349), .X(n32152) );
  inv_x1_sg U37922 ( .A(n32152), .X(n32153) );
  inv_x1_sg U37923 ( .A(n32152), .X(n32154) );
  inv_x1_sg U37924 ( .A(n32152), .X(n32155) );
  inv_x1_sg U37925 ( .A(n32152), .X(n32156) );
  inv_x1_sg U37926 ( .A(n34558), .X(n32157) );
  inv_x1_sg U37927 ( .A(n32157), .X(n32158) );
  inv_x1_sg U37928 ( .A(n32157), .X(n32159) );
  inv_x1_sg U37929 ( .A(n32157), .X(n32160) );
  inv_x1_sg U37930 ( .A(n32157), .X(n32161) );
  inv_x1_sg U37931 ( .A(n34557), .X(n32162) );
  inv_x1_sg U37932 ( .A(n32162), .X(n32163) );
  inv_x1_sg U37933 ( .A(n32162), .X(n32164) );
  inv_x1_sg U37934 ( .A(n32162), .X(n32165) );
  inv_x1_sg U37935 ( .A(n32162), .X(n32166) );
  inv_x1_sg U37936 ( .A(n31298), .X(n32167) );
  inv_x1_sg U37937 ( .A(n35263), .X(n32168) );
  inv_x1_sg U37938 ( .A(n34547), .X(n32169) );
  inv_x1_sg U37939 ( .A(n32398), .X(n32170) );
  inv_x1_sg U37940 ( .A(n30142), .X(n32171) );
  inv_x1_sg U37941 ( .A(n30143), .X(n32172) );
  inv_x1_sg U37942 ( .A(n34520), .X(n32173) );
  inv_x1_sg U37943 ( .A(n32173), .X(n32174) );
  inv_x1_sg U37944 ( .A(n32173), .X(n32175) );
  inv_x1_sg U37945 ( .A(n32173), .X(n32176) );
  inv_x1_sg U37946 ( .A(n30787), .X(n32177) );
  inv_x1_sg U37947 ( .A(n34512), .X(n32178) );
  inv_x1_sg U37948 ( .A(n30794), .X(n32179) );
  inv_x1_sg U37949 ( .A(n30794), .X(n32180) );
  inv_x1_sg U37950 ( .A(n34504), .X(n32181) );
  inv_x1_sg U37951 ( .A(n32181), .X(n32182) );
  inv_x1_sg U37952 ( .A(n32181), .X(n32183) );
  inv_x1_sg U37953 ( .A(n32181), .X(n32184) );
  inv_x1_sg U37954 ( .A(n32181), .X(n32185) );
  inv_x1_sg U37955 ( .A(n34446), .X(n32186) );
  inv_x1_sg U37956 ( .A(n34450), .X(n32187) );
  inv_x1_sg U37957 ( .A(n32187), .X(n32188) );
  inv_x1_sg U37958 ( .A(n32187), .X(n32189) );
  inv_x1_sg U37959 ( .A(n32187), .X(n32190) );
  inv_x1_sg U37960 ( .A(n32187), .X(n32191) );
  inv_x1_sg U37961 ( .A(n34441), .X(n32192) );
  inv_x1_sg U37962 ( .A(n34443), .X(n32193) );
  inv_x1_sg U37963 ( .A(n32193), .X(n32194) );
  inv_x1_sg U37964 ( .A(n32193), .X(n32195) );
  inv_x1_sg U37965 ( .A(n32193), .X(n32196) );
  inv_x1_sg U37966 ( .A(n32193), .X(n32197) );
  inv_x1_sg U37967 ( .A(n34431), .X(n32198) );
  inv_x1_sg U37968 ( .A(n34433), .X(n32199) );
  inv_x1_sg U37969 ( .A(n32199), .X(n32200) );
  inv_x1_sg U37970 ( .A(n32199), .X(n32201) );
  inv_x1_sg U37971 ( .A(n32199), .X(n32202) );
  inv_x1_sg U37972 ( .A(n32199), .X(n32203) );
  inv_x1_sg U37973 ( .A(n15105), .X(n32204) );
  inv_x1_sg U37974 ( .A(n32204), .X(n32205) );
  inv_x1_sg U37975 ( .A(n32204), .X(n32206) );
  inv_x1_sg U37976 ( .A(n32204), .X(n32207) );
  inv_x1_sg U37977 ( .A(n32204), .X(n32208) );
  inv_x1_sg U37978 ( .A(n28259), .X(n32209) );
  inv_x1_sg U37979 ( .A(n32209), .X(n32210) );
  inv_x1_sg U37980 ( .A(n32209), .X(n32211) );
  inv_x1_sg U37981 ( .A(n32209), .X(n32212) );
  inv_x1_sg U37982 ( .A(n32156), .X(n32213) );
  inv_x1_sg U37983 ( .A(n32213), .X(n32214) );
  inv_x1_sg U37984 ( .A(n32213), .X(n32215) );
  inv_x1_sg U37985 ( .A(n32213), .X(n32216) );
  inv_x1_sg U37986 ( .A(n32213), .X(n32217) );
  inv_x1_sg U37987 ( .A(n35307), .X(n32218) );
  inv_x1_sg U37988 ( .A(n32218), .X(n32219) );
  inv_x1_sg U37989 ( .A(n32218), .X(n32220) );
  inv_x1_sg U37990 ( .A(n32218), .X(n32221) );
  inv_x1_sg U37991 ( .A(n32218), .X(n32222) );
  inv_x1_sg U37992 ( .A(n35485), .X(n32223) );
  inv_x1_sg U37993 ( .A(n32008), .X(n32224) );
  inv_x1_sg U37994 ( .A(n34619), .X(n32225) );
  inv_x1_sg U37995 ( .A(n32225), .X(n32226) );
  inv_x1_sg U37996 ( .A(n32225), .X(n32227) );
  inv_x1_sg U37997 ( .A(n32225), .X(n32228) );
  inv_x1_sg U37998 ( .A(n32225), .X(n32229) );
  inv_x1_sg U37999 ( .A(n34618), .X(n32230) );
  inv_x1_sg U38000 ( .A(n32230), .X(n32231) );
  inv_x1_sg U38001 ( .A(n32230), .X(n32232) );
  inv_x1_sg U38002 ( .A(n32230), .X(n32233) );
  inv_x1_sg U38003 ( .A(n32230), .X(n32234) );
  inv_x1_sg U38004 ( .A(n34617), .X(n32235) );
  inv_x1_sg U38005 ( .A(n32235), .X(n32236) );
  inv_x1_sg U38006 ( .A(n32235), .X(n32237) );
  inv_x1_sg U38007 ( .A(n32235), .X(n32238) );
  inv_x1_sg U38008 ( .A(n32235), .X(n32239) );
  inv_x1_sg U38009 ( .A(n34614), .X(n32240) );
  inv_x1_sg U38010 ( .A(n32240), .X(n32241) );
  inv_x1_sg U38011 ( .A(n32240), .X(n32242) );
  inv_x1_sg U38012 ( .A(n32240), .X(n32243) );
  inv_x1_sg U38013 ( .A(n32240), .X(n32244) );
  inv_x1_sg U38014 ( .A(n34613), .X(n32245) );
  inv_x1_sg U38015 ( .A(n32245), .X(n32246) );
  inv_x1_sg U38016 ( .A(n32245), .X(n32247) );
  inv_x1_sg U38017 ( .A(n32245), .X(n32248) );
  inv_x1_sg U38018 ( .A(n32245), .X(n32249) );
  inv_x1_sg U38019 ( .A(n34612), .X(n32250) );
  inv_x1_sg U38020 ( .A(n32250), .X(n32251) );
  inv_x1_sg U38021 ( .A(n32250), .X(n32252) );
  inv_x1_sg U38022 ( .A(n32250), .X(n32253) );
  inv_x1_sg U38023 ( .A(n32250), .X(n32254) );
  inv_x1_sg U38024 ( .A(n30776), .X(n32255) );
  inv_x1_sg U38025 ( .A(n34605), .X(n32256) );
  inv_x1_sg U38026 ( .A(n30775), .X(n32257) );
  inv_x1_sg U38027 ( .A(n32257), .X(n32258) );
  inv_x1_sg U38028 ( .A(n32257), .X(n32259) );
  inv_x1_sg U38029 ( .A(n32257), .X(n32260) );
  inv_x1_sg U38030 ( .A(n32257), .X(n32261) );
  inv_x1_sg U38031 ( .A(n34606), .X(n32262) );
  inv_x1_sg U38032 ( .A(n32262), .X(n32263) );
  inv_x1_sg U38033 ( .A(n32262), .X(n32264) );
  inv_x1_sg U38034 ( .A(n32262), .X(n32265) );
  inv_x1_sg U38035 ( .A(n32262), .X(n32266) );
  inv_x1_sg U38036 ( .A(n30778), .X(n32267) );
  inv_x1_sg U38037 ( .A(n34600), .X(n32268) );
  inv_x1_sg U38038 ( .A(n34602), .X(n32269) );
  inv_x1_sg U38039 ( .A(n32269), .X(n32270) );
  inv_x1_sg U38040 ( .A(n32269), .X(n32271) );
  inv_x1_sg U38041 ( .A(n32269), .X(n32272) );
  inv_x1_sg U38042 ( .A(n32269), .X(n32273) );
  inv_x1_sg U38043 ( .A(n34601), .X(n32274) );
  inv_x1_sg U38044 ( .A(n32274), .X(n32275) );
  inv_x1_sg U38045 ( .A(n32274), .X(n32276) );
  inv_x1_sg U38046 ( .A(n32274), .X(n32277) );
  inv_x1_sg U38047 ( .A(n32274), .X(n32278) );
  inv_x1_sg U38048 ( .A(n34599), .X(n32279) );
  inv_x1_sg U38049 ( .A(n32279), .X(n32280) );
  inv_x1_sg U38050 ( .A(n32279), .X(n32281) );
  inv_x1_sg U38051 ( .A(n32279), .X(n32282) );
  inv_x1_sg U38052 ( .A(n32279), .X(n32283) );
  inv_x1_sg U38053 ( .A(n34598), .X(n32284) );
  inv_x1_sg U38054 ( .A(n32284), .X(n32285) );
  inv_x1_sg U38055 ( .A(n32284), .X(n32286) );
  inv_x1_sg U38056 ( .A(n32284), .X(n32287) );
  inv_x1_sg U38057 ( .A(n32284), .X(n32288) );
  inv_x1_sg U38058 ( .A(n34597), .X(n32289) );
  inv_x1_sg U38059 ( .A(n32289), .X(n32290) );
  inv_x1_sg U38060 ( .A(n32289), .X(n32291) );
  inv_x1_sg U38061 ( .A(n32289), .X(n32292) );
  inv_x1_sg U38062 ( .A(n32289), .X(n32293) );
  inv_x1_sg U38063 ( .A(n34594), .X(n32294) );
  inv_x1_sg U38064 ( .A(n32294), .X(n32295) );
  inv_x1_sg U38065 ( .A(n32294), .X(n32296) );
  inv_x1_sg U38066 ( .A(n32294), .X(n32297) );
  inv_x1_sg U38067 ( .A(n32294), .X(n32298) );
  inv_x1_sg U38068 ( .A(n34593), .X(n32299) );
  inv_x1_sg U38069 ( .A(n32299), .X(n32300) );
  inv_x1_sg U38070 ( .A(n32299), .X(n32301) );
  inv_x1_sg U38071 ( .A(n32299), .X(n32302) );
  inv_x1_sg U38072 ( .A(n32299), .X(n32303) );
  inv_x1_sg U38073 ( .A(n34592), .X(n32304) );
  inv_x1_sg U38074 ( .A(n32304), .X(n32305) );
  inv_x1_sg U38075 ( .A(n32304), .X(n32306) );
  inv_x1_sg U38076 ( .A(n32304), .X(n32307) );
  inv_x1_sg U38077 ( .A(n32304), .X(n32308) );
  inv_x1_sg U38078 ( .A(n34589), .X(n32309) );
  inv_x1_sg U38079 ( .A(n32309), .X(n32310) );
  inv_x1_sg U38080 ( .A(n32309), .X(n32311) );
  inv_x1_sg U38081 ( .A(n32309), .X(n32312) );
  inv_x1_sg U38082 ( .A(n32309), .X(n32313) );
  inv_x1_sg U38083 ( .A(n34588), .X(n32314) );
  inv_x1_sg U38084 ( .A(n32314), .X(n32315) );
  inv_x1_sg U38085 ( .A(n32314), .X(n32316) );
  inv_x1_sg U38086 ( .A(n32314), .X(n32317) );
  inv_x1_sg U38087 ( .A(n32314), .X(n32318) );
  inv_x1_sg U38088 ( .A(n32350), .X(n32319) );
  inv_x1_sg U38089 ( .A(n32319), .X(n32320) );
  inv_x1_sg U38090 ( .A(n32319), .X(n32321) );
  inv_x1_sg U38091 ( .A(n32319), .X(n32322) );
  inv_x1_sg U38092 ( .A(n32319), .X(n32323) );
  inv_x1_sg U38093 ( .A(n35157), .X(n32324) );
  inv_x1_sg U38094 ( .A(n32324), .X(n32325) );
  inv_x1_sg U38095 ( .A(n32324), .X(n32326) );
  inv_x1_sg U38096 ( .A(n32324), .X(n32327) );
  inv_x1_sg U38097 ( .A(n32324), .X(n32328) );
  inv_x1_sg U38098 ( .A(n34586), .X(n32329) );
  inv_x1_sg U38099 ( .A(n32329), .X(n32330) );
  inv_x1_sg U38100 ( .A(n32329), .X(n32331) );
  inv_x1_sg U38101 ( .A(n32329), .X(n32332) );
  inv_x1_sg U38102 ( .A(n32329), .X(n32333) );
  inv_x1_sg U38103 ( .A(n34585), .X(n32334) );
  inv_x1_sg U38104 ( .A(n32334), .X(n32335) );
  inv_x1_sg U38105 ( .A(n32334), .X(n32336) );
  inv_x1_sg U38106 ( .A(n32334), .X(n32337) );
  inv_x1_sg U38107 ( .A(n32334), .X(n32338) );
  inv_x1_sg U38108 ( .A(n34579), .X(n32339) );
  inv_x1_sg U38109 ( .A(n30779), .X(n32340) );
  inv_x1_sg U38110 ( .A(n34581), .X(n32341) );
  inv_x1_sg U38111 ( .A(n32341), .X(n32342) );
  inv_x1_sg U38112 ( .A(n32341), .X(n32343) );
  inv_x1_sg U38113 ( .A(n32341), .X(n32344) );
  inv_x1_sg U38114 ( .A(n32341), .X(n32345) );
  inv_x1_sg U38115 ( .A(n32327), .X(n32346) );
  inv_x1_sg U38116 ( .A(n32346), .X(n32347) );
  inv_x1_sg U38117 ( .A(n32346), .X(n32348) );
  inv_x1_sg U38118 ( .A(n32346), .X(n32349) );
  inv_x1_sg U38119 ( .A(n32346), .X(n32350) );
  inv_x1_sg U38120 ( .A(n34574), .X(n32351) );
  inv_x1_sg U38121 ( .A(n30780), .X(n32352) );
  inv_x1_sg U38122 ( .A(n34576), .X(n32353) );
  inv_x1_sg U38123 ( .A(n32353), .X(n32354) );
  inv_x1_sg U38124 ( .A(n32353), .X(n32355) );
  inv_x1_sg U38125 ( .A(n32353), .X(n32356) );
  inv_x1_sg U38126 ( .A(n32353), .X(n32357) );
  inv_x1_sg U38127 ( .A(n32141), .X(n32358) );
  inv_x1_sg U38128 ( .A(n32358), .X(n32359) );
  inv_x1_sg U38129 ( .A(n32358), .X(n32360) );
  inv_x1_sg U38130 ( .A(n32358), .X(n32361) );
  inv_x1_sg U38131 ( .A(n32358), .X(n32362) );
  inv_x1_sg U38132 ( .A(n34569), .X(n32363) );
  inv_x1_sg U38133 ( .A(n30781), .X(n32364) );
  inv_x1_sg U38134 ( .A(n32139), .X(n32365) );
  inv_x1_sg U38135 ( .A(n32365), .X(n32366) );
  inv_x1_sg U38136 ( .A(n32365), .X(n32367) );
  inv_x1_sg U38137 ( .A(n32365), .X(n32368) );
  inv_x1_sg U38138 ( .A(n32365), .X(n32369) );
  inv_x1_sg U38139 ( .A(n32332), .X(n32370) );
  inv_x1_sg U38140 ( .A(n32370), .X(n32371) );
  inv_x1_sg U38141 ( .A(n32370), .X(n32372) );
  inv_x1_sg U38142 ( .A(n32370), .X(n32373) );
  inv_x1_sg U38143 ( .A(n32370), .X(n32374) );
  inv_x1_sg U38144 ( .A(n34564), .X(n32375) );
  inv_x1_sg U38145 ( .A(n30783), .X(n32376) );
  inv_x1_sg U38146 ( .A(n34566), .X(n32377) );
  inv_x1_sg U38147 ( .A(n32377), .X(n32378) );
  inv_x1_sg U38148 ( .A(n32377), .X(n32379) );
  inv_x1_sg U38149 ( .A(n32377), .X(n32380) );
  inv_x1_sg U38150 ( .A(n32377), .X(n32381) );
  inv_x1_sg U38151 ( .A(n34565), .X(n32382) );
  inv_x1_sg U38152 ( .A(n32382), .X(n32383) );
  inv_x1_sg U38153 ( .A(n32382), .X(n32384) );
  inv_x1_sg U38154 ( .A(n32382), .X(n32385) );
  inv_x1_sg U38155 ( .A(n32382), .X(n32386) );
  inv_x1_sg U38156 ( .A(n30141), .X(n32387) );
  inv_x1_sg U38157 ( .A(n31300), .X(n32388) );
  inv_x1_sg U38158 ( .A(n32387), .X(n32389) );
  inv_x1_sg U38159 ( .A(n32389), .X(n32390) );
  inv_x1_sg U38160 ( .A(n32389), .X(n32391) );
  inv_x1_sg U38161 ( .A(n32389), .X(n32392) );
  inv_x1_sg U38162 ( .A(n32389), .X(n32393) );
  inv_x1_sg U38163 ( .A(n32393), .X(n32394) );
  inv_x1_sg U38164 ( .A(n32394), .X(n32395) );
  inv_x1_sg U38165 ( .A(n32394), .X(n32396) );
  inv_x1_sg U38166 ( .A(n32394), .X(n32397) );
  inv_x1_sg U38167 ( .A(n32394), .X(n32398) );
  inv_x1_sg U38168 ( .A(n34556), .X(n32399) );
  inv_x1_sg U38169 ( .A(n32399), .X(n32400) );
  inv_x1_sg U38170 ( .A(n32399), .X(n32401) );
  inv_x1_sg U38171 ( .A(n32399), .X(n32402) );
  inv_x1_sg U38172 ( .A(n32399), .X(n32403) );
  inv_x1_sg U38173 ( .A(n34555), .X(n32404) );
  inv_x1_sg U38174 ( .A(n32404), .X(n32405) );
  inv_x1_sg U38175 ( .A(n32404), .X(n32406) );
  inv_x1_sg U38176 ( .A(n32404), .X(n32407) );
  inv_x1_sg U38177 ( .A(n32404), .X(n32408) );
  inv_x1_sg U38178 ( .A(n34519), .X(n32409) );
  inv_x1_sg U38179 ( .A(n32409), .X(n32410) );
  inv_x1_sg U38180 ( .A(n32409), .X(n32411) );
  inv_x1_sg U38181 ( .A(n32409), .X(n32412) );
  inv_x1_sg U38182 ( .A(n34518), .X(n32413) );
  inv_x1_sg U38183 ( .A(n32413), .X(n32414) );
  inv_x1_sg U38184 ( .A(n32413), .X(n32415) );
  inv_x1_sg U38185 ( .A(n32413), .X(n32416) );
  inv_x1_sg U38186 ( .A(n32413), .X(n32417) );
  inv_x1_sg U38187 ( .A(n32178), .X(n32418) );
  inv_x1_sg U38188 ( .A(n32418), .X(n32419) );
  inv_x1_sg U38189 ( .A(n32418), .X(n32420) );
  inv_x1_sg U38190 ( .A(n32418), .X(n32421) );
  inv_x1_sg U38191 ( .A(n32418), .X(n32422) );
  inv_x1_sg U38192 ( .A(n35308), .X(n32423) );
  inv_x1_sg U38193 ( .A(n32423), .X(n32424) );
  inv_x1_sg U38194 ( .A(n32423), .X(n32425) );
  inv_x1_sg U38195 ( .A(n32423), .X(n32426) );
  inv_x1_sg U38196 ( .A(n32423), .X(n32427) );
  inv_x1_sg U38197 ( .A(n30731), .X(n32428) );
  inv_x1_sg U38198 ( .A(n34694), .X(n32429) );
  inv_x1_sg U38199 ( .A(n30734), .X(n32430) );
  inv_x1_sg U38200 ( .A(n30734), .X(n32431) );
  inv_x1_sg U38201 ( .A(n30737), .X(n32432) );
  inv_x1_sg U38202 ( .A(n34684), .X(n32433) );
  inv_x1_sg U38203 ( .A(n30740), .X(n32434) );
  inv_x1_sg U38204 ( .A(n30740), .X(n32435) );
  inv_x1_sg U38205 ( .A(n30743), .X(n32436) );
  inv_x1_sg U38206 ( .A(n30743), .X(n32437) );
  inv_x1_sg U38207 ( .A(n30746), .X(n32438) );
  inv_x1_sg U38208 ( .A(n30746), .X(n32439) );
  inv_x1_sg U38209 ( .A(n30750), .X(n32440) );
  inv_x1_sg U38210 ( .A(n34664), .X(n32441) );
  inv_x1_sg U38211 ( .A(n34661), .X(n32442) );
  inv_x1_sg U38212 ( .A(n34661), .X(n32443) );
  inv_x1_sg U38213 ( .A(n30753), .X(n32444) );
  inv_x1_sg U38214 ( .A(n34656), .X(n32445) );
  inv_x1_sg U38215 ( .A(n32445), .X(n32446) );
  inv_x1_sg U38216 ( .A(n32445), .X(n32447) );
  inv_x1_sg U38217 ( .A(n32445), .X(n32448) );
  inv_x1_sg U38218 ( .A(n32445), .X(n32449) );
  inv_x1_sg U38219 ( .A(n30756), .X(n32450) );
  inv_x1_sg U38220 ( .A(n34649), .X(n32451) );
  inv_x1_sg U38221 ( .A(n34651), .X(n32452) );
  inv_x1_sg U38222 ( .A(n32452), .X(n32453) );
  inv_x1_sg U38223 ( .A(n32452), .X(n32454) );
  inv_x1_sg U38224 ( .A(n32452), .X(n32455) );
  inv_x1_sg U38225 ( .A(n32452), .X(n32456) );
  inv_x1_sg U38226 ( .A(n30759), .X(n32457) );
  inv_x1_sg U38227 ( .A(n30759), .X(n32458) );
  inv_x1_sg U38228 ( .A(n34646), .X(n32459) );
  inv_x1_sg U38229 ( .A(n32459), .X(n32460) );
  inv_x1_sg U38230 ( .A(n32459), .X(n32461) );
  inv_x1_sg U38231 ( .A(n32459), .X(n32462) );
  inv_x1_sg U38232 ( .A(n32459), .X(n32463) );
  inv_x1_sg U38233 ( .A(n30763), .X(n32464) );
  inv_x1_sg U38234 ( .A(n30763), .X(n32465) );
  inv_x1_sg U38235 ( .A(n34641), .X(n32466) );
  inv_x1_sg U38236 ( .A(n32466), .X(n32467) );
  inv_x1_sg U38237 ( .A(n32466), .X(n32468) );
  inv_x1_sg U38238 ( .A(n32466), .X(n32469) );
  inv_x1_sg U38239 ( .A(n32466), .X(n32470) );
  inv_x1_sg U38240 ( .A(n30766), .X(n32471) );
  inv_x1_sg U38241 ( .A(n30766), .X(n32472) );
  inv_x1_sg U38242 ( .A(n34634), .X(n32473) );
  inv_x1_sg U38243 ( .A(n32473), .X(n32474) );
  inv_x1_sg U38244 ( .A(n32473), .X(n32475) );
  inv_x1_sg U38245 ( .A(n32473), .X(n32476) );
  inv_x1_sg U38246 ( .A(n32473), .X(n32477) );
  inv_x1_sg U38247 ( .A(n30769), .X(n32478) );
  inv_x1_sg U38248 ( .A(n30769), .X(n32479) );
  inv_x1_sg U38249 ( .A(n34629), .X(n32480) );
  inv_x1_sg U38250 ( .A(n32480), .X(n32481) );
  inv_x1_sg U38251 ( .A(n32480), .X(n32482) );
  inv_x1_sg U38252 ( .A(n32480), .X(n32483) );
  inv_x1_sg U38253 ( .A(n32480), .X(n32484) );
  inv_x1_sg U38254 ( .A(n30774), .X(n32485) );
  inv_x1_sg U38255 ( .A(n30774), .X(n32486) );
  inv_x1_sg U38256 ( .A(n34624), .X(n32487) );
  inv_x1_sg U38257 ( .A(n32487), .X(n32488) );
  inv_x1_sg U38258 ( .A(n32487), .X(n32489) );
  inv_x1_sg U38259 ( .A(n32487), .X(n32490) );
  inv_x1_sg U38260 ( .A(n32487), .X(n32491) );
  inv_x1_sg U38261 ( .A(n34616), .X(n32492) );
  inv_x1_sg U38262 ( .A(n32492), .X(n32493) );
  inv_x1_sg U38263 ( .A(n32492), .X(n32494) );
  inv_x1_sg U38264 ( .A(n32492), .X(n32495) );
  inv_x1_sg U38265 ( .A(n32492), .X(n32496) );
  inv_x1_sg U38266 ( .A(n34611), .X(n32497) );
  inv_x1_sg U38267 ( .A(n32497), .X(n32498) );
  inv_x1_sg U38268 ( .A(n32497), .X(n32499) );
  inv_x1_sg U38269 ( .A(n32497), .X(n32500) );
  inv_x1_sg U38270 ( .A(n32497), .X(n32501) );
  inv_x1_sg U38271 ( .A(n29669), .X(n32502) );
  inv_x1_sg U38272 ( .A(n32502), .X(n32503) );
  inv_x1_sg U38273 ( .A(n32502), .X(n32504) );
  inv_x1_sg U38274 ( .A(n32502), .X(n32505) );
  inv_x1_sg U38275 ( .A(n31664), .X(n32506) );
  inv_x1_sg U38276 ( .A(n32506), .X(n32507) );
  inv_x1_sg U38277 ( .A(n32506), .X(n32508) );
  inv_x1_sg U38278 ( .A(n32506), .X(n32509) );
  inv_x1_sg U38279 ( .A(n32506), .X(n32510) );
  inv_x1_sg U38280 ( .A(n35314), .X(n32511) );
  inv_x1_sg U38281 ( .A(n32511), .X(n32512) );
  inv_x1_sg U38282 ( .A(n32511), .X(n32513) );
  inv_x1_sg U38283 ( .A(n32511), .X(n32514) );
  inv_x1_sg U38284 ( .A(n32511), .X(n32515) );
  inv_x1_sg U38285 ( .A(n32061), .X(n32516) );
  inv_x1_sg U38286 ( .A(n32516), .X(n32517) );
  inv_x1_sg U38287 ( .A(n32516), .X(n32518) );
  inv_x1_sg U38288 ( .A(n32516), .X(n32519) );
  inv_x1_sg U38289 ( .A(n32516), .X(n32520) );
  inv_x1_sg U38290 ( .A(n30643), .X(n32521) );
  inv_x1_sg U38291 ( .A(n30643), .X(n32522) );
  inv_x1_sg U38292 ( .A(n34802), .X(n32523) );
  inv_x1_sg U38293 ( .A(n32523), .X(n32524) );
  inv_x1_sg U38294 ( .A(n32523), .X(n32525) );
  inv_x1_sg U38295 ( .A(n32523), .X(n32526) );
  inv_x1_sg U38296 ( .A(n32523), .X(n32527) );
  inv_x1_sg U38297 ( .A(n30646), .X(n32528) );
  inv_x1_sg U38298 ( .A(n34795), .X(n32529) );
  inv_x1_sg U38299 ( .A(n34797), .X(n32530) );
  inv_x1_sg U38300 ( .A(n32530), .X(n32531) );
  inv_x1_sg U38301 ( .A(n32530), .X(n32532) );
  inv_x1_sg U38302 ( .A(n32530), .X(n32533) );
  inv_x1_sg U38303 ( .A(n32530), .X(n32534) );
  inv_x1_sg U38304 ( .A(n30188), .X(n32535) );
  inv_x1_sg U38305 ( .A(n32535), .X(n32536) );
  inv_x1_sg U38306 ( .A(n32535), .X(n32537) );
  inv_x1_sg U38307 ( .A(n32535), .X(n32538) );
  inv_x1_sg U38308 ( .A(n32535), .X(n32539) );
  inv_x1_sg U38309 ( .A(n30650), .X(n32540) );
  inv_x1_sg U38310 ( .A(n30650), .X(n32541) );
  inv_x1_sg U38311 ( .A(n34792), .X(n32542) );
  inv_x1_sg U38312 ( .A(n32542), .X(n32543) );
  inv_x1_sg U38313 ( .A(n32542), .X(n32544) );
  inv_x1_sg U38314 ( .A(n32542), .X(n32545) );
  inv_x1_sg U38315 ( .A(n32542), .X(n32546) );
  inv_x1_sg U38316 ( .A(n34791), .X(n32547) );
  inv_x1_sg U38317 ( .A(n32547), .X(n32548) );
  inv_x1_sg U38318 ( .A(n32547), .X(n32549) );
  inv_x1_sg U38319 ( .A(n32547), .X(n32550) );
  inv_x1_sg U38320 ( .A(n32547), .X(n32551) );
  inv_x1_sg U38321 ( .A(n30654), .X(n32552) );
  inv_x1_sg U38322 ( .A(n30654), .X(n32553) );
  inv_x1_sg U38323 ( .A(n34787), .X(n32554) );
  inv_x1_sg U38324 ( .A(n32554), .X(n32555) );
  inv_x1_sg U38325 ( .A(n32554), .X(n32556) );
  inv_x1_sg U38326 ( .A(n32554), .X(n32557) );
  inv_x1_sg U38327 ( .A(n32554), .X(n32558) );
  inv_x1_sg U38328 ( .A(n34786), .X(n32559) );
  inv_x1_sg U38329 ( .A(n32559), .X(n32560) );
  inv_x1_sg U38330 ( .A(n32559), .X(n32561) );
  inv_x1_sg U38331 ( .A(n32559), .X(n32562) );
  inv_x1_sg U38332 ( .A(n32559), .X(n32563) );
  inv_x1_sg U38333 ( .A(n30658), .X(n32564) );
  inv_x1_sg U38334 ( .A(n30658), .X(n32565) );
  inv_x1_sg U38335 ( .A(n34782), .X(n32566) );
  inv_x1_sg U38336 ( .A(n32566), .X(n32567) );
  inv_x1_sg U38337 ( .A(n32566), .X(n32568) );
  inv_x1_sg U38338 ( .A(n32566), .X(n32569) );
  inv_x1_sg U38339 ( .A(n32566), .X(n32570) );
  inv_x1_sg U38340 ( .A(n34781), .X(n32571) );
  inv_x1_sg U38341 ( .A(n32571), .X(n32572) );
  inv_x1_sg U38342 ( .A(n32571), .X(n32573) );
  inv_x1_sg U38343 ( .A(n32571), .X(n32574) );
  inv_x1_sg U38344 ( .A(n32571), .X(n32575) );
  inv_x1_sg U38345 ( .A(n30662), .X(n32576) );
  inv_x1_sg U38346 ( .A(n30662), .X(n32577) );
  inv_x1_sg U38347 ( .A(n34776), .X(n32578) );
  inv_x1_sg U38348 ( .A(n32578), .X(n32579) );
  inv_x1_sg U38349 ( .A(n32578), .X(n32580) );
  inv_x1_sg U38350 ( .A(n32578), .X(n32581) );
  inv_x1_sg U38351 ( .A(n32578), .X(n32582) );
  inv_x1_sg U38352 ( .A(n34777), .X(n32583) );
  inv_x1_sg U38353 ( .A(n32583), .X(n32584) );
  inv_x1_sg U38354 ( .A(n32583), .X(n32585) );
  inv_x1_sg U38355 ( .A(n32583), .X(n32586) );
  inv_x1_sg U38356 ( .A(n32583), .X(n32587) );
  inv_x1_sg U38357 ( .A(n30666), .X(n32588) );
  inv_x1_sg U38358 ( .A(n30666), .X(n32589) );
  inv_x1_sg U38359 ( .A(n34771), .X(n32590) );
  inv_x1_sg U38360 ( .A(n32590), .X(n32591) );
  inv_x1_sg U38361 ( .A(n32590), .X(n32592) );
  inv_x1_sg U38362 ( .A(n32590), .X(n32593) );
  inv_x1_sg U38363 ( .A(n32590), .X(n32594) );
  inv_x1_sg U38364 ( .A(n34772), .X(n32595) );
  inv_x1_sg U38365 ( .A(n32595), .X(n32596) );
  inv_x1_sg U38366 ( .A(n32595), .X(n32597) );
  inv_x1_sg U38367 ( .A(n32595), .X(n32598) );
  inv_x1_sg U38368 ( .A(n32595), .X(n32599) );
  inv_x1_sg U38369 ( .A(n30670), .X(n32600) );
  inv_x1_sg U38370 ( .A(n30670), .X(n32601) );
  inv_x1_sg U38371 ( .A(n34766), .X(n32602) );
  inv_x1_sg U38372 ( .A(n32602), .X(n32603) );
  inv_x1_sg U38373 ( .A(n32602), .X(n32604) );
  inv_x1_sg U38374 ( .A(n32602), .X(n32605) );
  inv_x1_sg U38375 ( .A(n32602), .X(n32606) );
  inv_x1_sg U38376 ( .A(n34767), .X(n32607) );
  inv_x1_sg U38377 ( .A(n32607), .X(n32608) );
  inv_x1_sg U38378 ( .A(n32607), .X(n32609) );
  inv_x1_sg U38379 ( .A(n32607), .X(n32610) );
  inv_x1_sg U38380 ( .A(n32607), .X(n32611) );
  inv_x1_sg U38381 ( .A(n30675), .X(n32612) );
  inv_x1_sg U38382 ( .A(n30675), .X(n32613) );
  inv_x1_sg U38383 ( .A(n34762), .X(n32614) );
  inv_x1_sg U38384 ( .A(n32614), .X(n32615) );
  inv_x1_sg U38385 ( .A(n32614), .X(n32616) );
  inv_x1_sg U38386 ( .A(n32614), .X(n32617) );
  inv_x1_sg U38387 ( .A(n32614), .X(n32618) );
  inv_x1_sg U38388 ( .A(n34761), .X(n32619) );
  inv_x1_sg U38389 ( .A(n32619), .X(n32620) );
  inv_x1_sg U38390 ( .A(n32619), .X(n32621) );
  inv_x1_sg U38391 ( .A(n32619), .X(n32622) );
  inv_x1_sg U38392 ( .A(n32619), .X(n32623) );
  inv_x1_sg U38393 ( .A(n30679), .X(n32624) );
  inv_x1_sg U38394 ( .A(n30679), .X(n32625) );
  inv_x1_sg U38395 ( .A(n34757), .X(n32626) );
  inv_x1_sg U38396 ( .A(n32626), .X(n32627) );
  inv_x1_sg U38397 ( .A(n32626), .X(n32628) );
  inv_x1_sg U38398 ( .A(n32626), .X(n32629) );
  inv_x1_sg U38399 ( .A(n32626), .X(n32630) );
  inv_x1_sg U38400 ( .A(n34756), .X(n32631) );
  inv_x1_sg U38401 ( .A(n32631), .X(n32632) );
  inv_x1_sg U38402 ( .A(n32631), .X(n32633) );
  inv_x1_sg U38403 ( .A(n32631), .X(n32634) );
  inv_x1_sg U38404 ( .A(n32631), .X(n32635) );
  inv_x1_sg U38405 ( .A(n30683), .X(n32636) );
  inv_x1_sg U38406 ( .A(n30683), .X(n32637) );
  inv_x1_sg U38407 ( .A(n34752), .X(n32638) );
  inv_x1_sg U38408 ( .A(n32638), .X(n32639) );
  inv_x1_sg U38409 ( .A(n32638), .X(n32640) );
  inv_x1_sg U38410 ( .A(n32638), .X(n32641) );
  inv_x1_sg U38411 ( .A(n32638), .X(n32642) );
  inv_x1_sg U38412 ( .A(n34751), .X(n32643) );
  inv_x1_sg U38413 ( .A(n32643), .X(n32644) );
  inv_x1_sg U38414 ( .A(n32643), .X(n32645) );
  inv_x1_sg U38415 ( .A(n32643), .X(n32646) );
  inv_x1_sg U38416 ( .A(n32643), .X(n32647) );
  inv_x1_sg U38417 ( .A(n30687), .X(n32648) );
  inv_x1_sg U38418 ( .A(n30687), .X(n32649) );
  inv_x1_sg U38419 ( .A(n34747), .X(n32650) );
  inv_x1_sg U38420 ( .A(n32650), .X(n32651) );
  inv_x1_sg U38421 ( .A(n32650), .X(n32652) );
  inv_x1_sg U38422 ( .A(n32650), .X(n32653) );
  inv_x1_sg U38423 ( .A(n32650), .X(n32654) );
  inv_x1_sg U38424 ( .A(n34746), .X(n32655) );
  inv_x1_sg U38425 ( .A(n32655), .X(n32656) );
  inv_x1_sg U38426 ( .A(n32655), .X(n32657) );
  inv_x1_sg U38427 ( .A(n32655), .X(n32658) );
  inv_x1_sg U38428 ( .A(n32655), .X(n32659) );
  inv_x1_sg U38429 ( .A(n30691), .X(n32660) );
  inv_x1_sg U38430 ( .A(n30691), .X(n32661) );
  inv_x1_sg U38431 ( .A(n34742), .X(n32662) );
  inv_x1_sg U38432 ( .A(n32662), .X(n32663) );
  inv_x1_sg U38433 ( .A(n32662), .X(n32664) );
  inv_x1_sg U38434 ( .A(n32662), .X(n32665) );
  inv_x1_sg U38435 ( .A(n32662), .X(n32666) );
  inv_x1_sg U38436 ( .A(n34741), .X(n32667) );
  inv_x1_sg U38437 ( .A(n32667), .X(n32668) );
  inv_x1_sg U38438 ( .A(n32667), .X(n32669) );
  inv_x1_sg U38439 ( .A(n32667), .X(n32670) );
  inv_x1_sg U38440 ( .A(n32667), .X(n32671) );
  inv_x1_sg U38441 ( .A(n30695), .X(n32672) );
  inv_x1_sg U38442 ( .A(n30695), .X(n32673) );
  inv_x1_sg U38443 ( .A(n34737), .X(n32674) );
  inv_x1_sg U38444 ( .A(n32674), .X(n32675) );
  inv_x1_sg U38445 ( .A(n32674), .X(n32676) );
  inv_x1_sg U38446 ( .A(n32674), .X(n32677) );
  inv_x1_sg U38447 ( .A(n32674), .X(n32678) );
  inv_x1_sg U38448 ( .A(n34736), .X(n32679) );
  inv_x1_sg U38449 ( .A(n32679), .X(n32680) );
  inv_x1_sg U38450 ( .A(n32679), .X(n32681) );
  inv_x1_sg U38451 ( .A(n32679), .X(n32682) );
  inv_x1_sg U38452 ( .A(n32679), .X(n32683) );
  inv_x1_sg U38453 ( .A(n30699), .X(n32684) );
  inv_x1_sg U38454 ( .A(n30699), .X(n32685) );
  inv_x1_sg U38455 ( .A(n34732), .X(n32686) );
  inv_x1_sg U38456 ( .A(n32686), .X(n32687) );
  inv_x1_sg U38457 ( .A(n32686), .X(n32688) );
  inv_x1_sg U38458 ( .A(n32686), .X(n32689) );
  inv_x1_sg U38459 ( .A(n32686), .X(n32690) );
  inv_x1_sg U38460 ( .A(n34731), .X(n32691) );
  inv_x1_sg U38461 ( .A(n32691), .X(n32692) );
  inv_x1_sg U38462 ( .A(n32691), .X(n32693) );
  inv_x1_sg U38463 ( .A(n32691), .X(n32694) );
  inv_x1_sg U38464 ( .A(n32691), .X(n32695) );
  inv_x1_sg U38465 ( .A(n30703), .X(n32696) );
  inv_x1_sg U38466 ( .A(n29672), .X(n32697) );
  inv_x1_sg U38467 ( .A(n34727), .X(n32698) );
  inv_x1_sg U38468 ( .A(n32698), .X(n32699) );
  inv_x1_sg U38469 ( .A(n32698), .X(n32700) );
  inv_x1_sg U38470 ( .A(n32698), .X(n32701) );
  inv_x1_sg U38471 ( .A(n32698), .X(n32702) );
  inv_x1_sg U38472 ( .A(n34728), .X(n32703) );
  inv_x1_sg U38473 ( .A(n32703), .X(n32704) );
  inv_x1_sg U38474 ( .A(n32703), .X(n32705) );
  inv_x1_sg U38475 ( .A(n32703), .X(n32706) );
  inv_x1_sg U38476 ( .A(n32703), .X(n32707) );
  inv_x1_sg U38477 ( .A(n30710), .X(n32708) );
  inv_x1_sg U38478 ( .A(n30710), .X(n32709) );
  inv_x1_sg U38479 ( .A(n34722), .X(n32710) );
  inv_x1_sg U38480 ( .A(n32710), .X(n32711) );
  inv_x1_sg U38481 ( .A(n32710), .X(n32712) );
  inv_x1_sg U38482 ( .A(n32710), .X(n32713) );
  inv_x1_sg U38483 ( .A(n32710), .X(n32714) );
  inv_x1_sg U38484 ( .A(n34721), .X(n32715) );
  inv_x1_sg U38485 ( .A(n32715), .X(n32716) );
  inv_x1_sg U38486 ( .A(n32715), .X(n32717) );
  inv_x1_sg U38487 ( .A(n32715), .X(n32718) );
  inv_x1_sg U38488 ( .A(n32715), .X(n32719) );
  inv_x1_sg U38489 ( .A(n30714), .X(n32720) );
  inv_x1_sg U38490 ( .A(n30714), .X(n32721) );
  inv_x1_sg U38491 ( .A(n34717), .X(n32722) );
  inv_x1_sg U38492 ( .A(n32722), .X(n32723) );
  inv_x1_sg U38493 ( .A(n32722), .X(n32724) );
  inv_x1_sg U38494 ( .A(n32722), .X(n32725) );
  inv_x1_sg U38495 ( .A(n32722), .X(n32726) );
  inv_x1_sg U38496 ( .A(n34716), .X(n32727) );
  inv_x1_sg U38497 ( .A(n32727), .X(n32728) );
  inv_x1_sg U38498 ( .A(n32727), .X(n32729) );
  inv_x1_sg U38499 ( .A(n32727), .X(n32730) );
  inv_x1_sg U38500 ( .A(n32727), .X(n32731) );
  inv_x1_sg U38501 ( .A(n35340), .X(n32732) );
  inv_x1_sg U38502 ( .A(n35369), .X(n32733) );
  inv_x1_sg U38503 ( .A(n34710), .X(n32734) );
  inv_x1_sg U38504 ( .A(n32734), .X(n32735) );
  inv_x1_sg U38505 ( .A(n32734), .X(n32736) );
  inv_x1_sg U38506 ( .A(n32734), .X(n32737) );
  inv_x1_sg U38507 ( .A(n32734), .X(n32738) );
  inv_x1_sg U38508 ( .A(n34709), .X(n32739) );
  inv_x1_sg U38509 ( .A(n32739), .X(n32740) );
  inv_x1_sg U38510 ( .A(n32739), .X(n32741) );
  inv_x1_sg U38511 ( .A(n32739), .X(n32742) );
  inv_x1_sg U38512 ( .A(n32739), .X(n32743) );
  inv_x1_sg U38513 ( .A(n35178), .X(n32744) );
  inv_x1_sg U38514 ( .A(n35384), .X(n32745) );
  inv_x1_sg U38515 ( .A(n34706), .X(n32746) );
  inv_x1_sg U38516 ( .A(n32746), .X(n32747) );
  inv_x1_sg U38517 ( .A(n32746), .X(n32748) );
  inv_x1_sg U38518 ( .A(n32746), .X(n32749) );
  inv_x1_sg U38519 ( .A(n32746), .X(n32750) );
  inv_x1_sg U38520 ( .A(n34705), .X(n32751) );
  inv_x1_sg U38521 ( .A(n32751), .X(n32752) );
  inv_x1_sg U38522 ( .A(n32751), .X(n32753) );
  inv_x1_sg U38523 ( .A(n32751), .X(n32754) );
  inv_x1_sg U38524 ( .A(n32751), .X(n32755) );
  inv_x1_sg U38525 ( .A(n30728), .X(n32756) );
  inv_x1_sg U38526 ( .A(n30728), .X(n32757) );
  inv_x1_sg U38527 ( .A(n34701), .X(n32758) );
  inv_x1_sg U38528 ( .A(n32758), .X(n32759) );
  inv_x1_sg U38529 ( .A(n32758), .X(n32760) );
  inv_x1_sg U38530 ( .A(n32758), .X(n32761) );
  inv_x1_sg U38531 ( .A(n32758), .X(n32762) );
  inv_x1_sg U38532 ( .A(n34702), .X(n32763) );
  inv_x1_sg U38533 ( .A(n32763), .X(n32764) );
  inv_x1_sg U38534 ( .A(n32763), .X(n32765) );
  inv_x1_sg U38535 ( .A(n32763), .X(n32766) );
  inv_x1_sg U38536 ( .A(n32763), .X(n32767) );
  inv_x1_sg U38537 ( .A(n34696), .X(n32768) );
  inv_x1_sg U38538 ( .A(n32768), .X(n32769) );
  inv_x1_sg U38539 ( .A(n32768), .X(n32770) );
  inv_x1_sg U38540 ( .A(n32768), .X(n32771) );
  inv_x1_sg U38541 ( .A(n32768), .X(n32772) );
  inv_x1_sg U38542 ( .A(n34695), .X(n32773) );
  inv_x1_sg U38543 ( .A(n32773), .X(n32774) );
  inv_x1_sg U38544 ( .A(n32773), .X(n32775) );
  inv_x1_sg U38545 ( .A(n32773), .X(n32776) );
  inv_x1_sg U38546 ( .A(n32773), .X(n32777) );
  inv_x1_sg U38547 ( .A(n34691), .X(n32778) );
  inv_x1_sg U38548 ( .A(n32778), .X(n32779) );
  inv_x1_sg U38549 ( .A(n32778), .X(n32780) );
  inv_x1_sg U38550 ( .A(n32778), .X(n32781) );
  inv_x1_sg U38551 ( .A(n32778), .X(n32782) );
  inv_x1_sg U38552 ( .A(n34690), .X(n32783) );
  inv_x1_sg U38553 ( .A(n32783), .X(n32784) );
  inv_x1_sg U38554 ( .A(n32783), .X(n32785) );
  inv_x1_sg U38555 ( .A(n32783), .X(n32786) );
  inv_x1_sg U38556 ( .A(n32783), .X(n32787) );
  inv_x1_sg U38557 ( .A(n34686), .X(n32788) );
  inv_x1_sg U38558 ( .A(n32788), .X(n32789) );
  inv_x1_sg U38559 ( .A(n32788), .X(n32790) );
  inv_x1_sg U38560 ( .A(n32788), .X(n32791) );
  inv_x1_sg U38561 ( .A(n32788), .X(n32792) );
  inv_x1_sg U38562 ( .A(n34685), .X(n32793) );
  inv_x1_sg U38563 ( .A(n32793), .X(n32794) );
  inv_x1_sg U38564 ( .A(n32793), .X(n32795) );
  inv_x1_sg U38565 ( .A(n32793), .X(n32796) );
  inv_x1_sg U38566 ( .A(n32793), .X(n32797) );
  inv_x1_sg U38567 ( .A(n34680), .X(n32798) );
  inv_x1_sg U38568 ( .A(n32798), .X(n32799) );
  inv_x1_sg U38569 ( .A(n32798), .X(n32800) );
  inv_x1_sg U38570 ( .A(n32798), .X(n32801) );
  inv_x1_sg U38571 ( .A(n32798), .X(n32802) );
  inv_x1_sg U38572 ( .A(n34681), .X(n32803) );
  inv_x1_sg U38573 ( .A(n32803), .X(n32804) );
  inv_x1_sg U38574 ( .A(n32803), .X(n32805) );
  inv_x1_sg U38575 ( .A(n32803), .X(n32806) );
  inv_x1_sg U38576 ( .A(n32803), .X(n32807) );
  inv_x1_sg U38577 ( .A(n34676), .X(n32808) );
  inv_x1_sg U38578 ( .A(n32808), .X(n32809) );
  inv_x1_sg U38579 ( .A(n32808), .X(n32810) );
  inv_x1_sg U38580 ( .A(n32808), .X(n32811) );
  inv_x1_sg U38581 ( .A(n32808), .X(n32812) );
  inv_x1_sg U38582 ( .A(n34675), .X(n32813) );
  inv_x1_sg U38583 ( .A(n32813), .X(n32814) );
  inv_x1_sg U38584 ( .A(n32813), .X(n32815) );
  inv_x1_sg U38585 ( .A(n32813), .X(n32816) );
  inv_x1_sg U38586 ( .A(n32813), .X(n32817) );
  inv_x1_sg U38587 ( .A(n34670), .X(n32818) );
  inv_x1_sg U38588 ( .A(n32818), .X(n32819) );
  inv_x1_sg U38589 ( .A(n32818), .X(n32820) );
  inv_x1_sg U38590 ( .A(n32818), .X(n32821) );
  inv_x1_sg U38591 ( .A(n32818), .X(n32822) );
  inv_x1_sg U38592 ( .A(n34671), .X(n32823) );
  inv_x1_sg U38593 ( .A(n32823), .X(n32824) );
  inv_x1_sg U38594 ( .A(n32823), .X(n32825) );
  inv_x1_sg U38595 ( .A(n32823), .X(n32826) );
  inv_x1_sg U38596 ( .A(n32823), .X(n32827) );
  inv_x1_sg U38597 ( .A(n34665), .X(n32828) );
  inv_x1_sg U38598 ( .A(n32828), .X(n32829) );
  inv_x1_sg U38599 ( .A(n32828), .X(n32830) );
  inv_x1_sg U38600 ( .A(n32828), .X(n32831) );
  inv_x1_sg U38601 ( .A(n32828), .X(n32832) );
  inv_x1_sg U38602 ( .A(n34666), .X(n32833) );
  inv_x1_sg U38603 ( .A(n32833), .X(n32834) );
  inv_x1_sg U38604 ( .A(n32833), .X(n32835) );
  inv_x1_sg U38605 ( .A(n32833), .X(n32836) );
  inv_x1_sg U38606 ( .A(n32833), .X(n32837) );
  inv_x1_sg U38607 ( .A(n30752), .X(n32838) );
  inv_x1_sg U38608 ( .A(n32838), .X(n32839) );
  inv_x1_sg U38609 ( .A(n32838), .X(n32840) );
  inv_x1_sg U38610 ( .A(n32838), .X(n32841) );
  inv_x1_sg U38611 ( .A(n32838), .X(n32842) );
  inv_x1_sg U38612 ( .A(n30752), .X(n32843) );
  inv_x1_sg U38613 ( .A(n32843), .X(n32844) );
  inv_x1_sg U38614 ( .A(n32843), .X(n32845) );
  inv_x1_sg U38615 ( .A(n32843), .X(n32846) );
  inv_x1_sg U38616 ( .A(n32843), .X(n32847) );
  inv_x1_sg U38617 ( .A(n34655), .X(n32848) );
  inv_x1_sg U38618 ( .A(n32848), .X(n32849) );
  inv_x1_sg U38619 ( .A(n32848), .X(n32850) );
  inv_x1_sg U38620 ( .A(n32848), .X(n32851) );
  inv_x1_sg U38621 ( .A(n32848), .X(n32852) );
  inv_x1_sg U38622 ( .A(n34650), .X(n32853) );
  inv_x1_sg U38623 ( .A(n32853), .X(n32854) );
  inv_x1_sg U38624 ( .A(n32853), .X(n32855) );
  inv_x1_sg U38625 ( .A(n32853), .X(n32856) );
  inv_x1_sg U38626 ( .A(n32853), .X(n32857) );
  inv_x1_sg U38627 ( .A(n34645), .X(n32858) );
  inv_x1_sg U38628 ( .A(n32858), .X(n32859) );
  inv_x1_sg U38629 ( .A(n32858), .X(n32860) );
  inv_x1_sg U38630 ( .A(n32858), .X(n32861) );
  inv_x1_sg U38631 ( .A(n32858), .X(n32862) );
  inv_x1_sg U38632 ( .A(n34640), .X(n32863) );
  inv_x1_sg U38633 ( .A(n32863), .X(n32864) );
  inv_x1_sg U38634 ( .A(n32863), .X(n32865) );
  inv_x1_sg U38635 ( .A(n32863), .X(n32866) );
  inv_x1_sg U38636 ( .A(n32863), .X(n32867) );
  inv_x1_sg U38637 ( .A(n34633), .X(n32868) );
  inv_x1_sg U38638 ( .A(n32868), .X(n32869) );
  inv_x1_sg U38639 ( .A(n32868), .X(n32870) );
  inv_x1_sg U38640 ( .A(n32868), .X(n32871) );
  inv_x1_sg U38641 ( .A(n32868), .X(n32872) );
  inv_x1_sg U38642 ( .A(n34628), .X(n32873) );
  inv_x1_sg U38643 ( .A(n32873), .X(n32874) );
  inv_x1_sg U38644 ( .A(n32873), .X(n32875) );
  inv_x1_sg U38645 ( .A(n32873), .X(n32876) );
  inv_x1_sg U38646 ( .A(n32873), .X(n32877) );
  inv_x1_sg U38647 ( .A(n34623), .X(n32878) );
  inv_x1_sg U38648 ( .A(n32878), .X(n32879) );
  inv_x1_sg U38649 ( .A(n32878), .X(n32880) );
  inv_x1_sg U38650 ( .A(n32878), .X(n32881) );
  inv_x1_sg U38651 ( .A(n32878), .X(n32882) );
  inv_x1_sg U38652 ( .A(n26579), .X(n32883) );
  inv_x1_sg U38653 ( .A(n32883), .X(n32884) );
  inv_x1_sg U38654 ( .A(n32883), .X(n32885) );
  inv_x1_sg U38655 ( .A(n32883), .X(n32886) );
  inv_x1_sg U38656 ( .A(n32883), .X(n32887) );
  inv_x1_sg U38657 ( .A(n30199), .X(n32888) );
  inv_x1_sg U38658 ( .A(n35417), .X(n32889) );
  inv_x1_sg U38659 ( .A(n34856), .X(n32890) );
  inv_x1_sg U38660 ( .A(n32890), .X(n32891) );
  inv_x1_sg U38661 ( .A(n32890), .X(n32892) );
  inv_x1_sg U38662 ( .A(n32890), .X(n32893) );
  inv_x1_sg U38663 ( .A(n32890), .X(n32894) );
  inv_x1_sg U38664 ( .A(n34857), .X(n32895) );
  inv_x1_sg U38665 ( .A(n32895), .X(n32896) );
  inv_x1_sg U38666 ( .A(n32895), .X(n32897) );
  inv_x1_sg U38667 ( .A(n32895), .X(n32898) );
  inv_x1_sg U38668 ( .A(n32895), .X(n32899) );
  inv_x1_sg U38669 ( .A(n34801), .X(n32900) );
  inv_x1_sg U38670 ( .A(n32900), .X(n32901) );
  inv_x1_sg U38671 ( .A(n32900), .X(n32902) );
  inv_x1_sg U38672 ( .A(n32900), .X(n32903) );
  inv_x1_sg U38673 ( .A(n32900), .X(n32904) );
  inv_x1_sg U38674 ( .A(n12438), .X(n32905) );
  inv_x1_sg U38675 ( .A(n32905), .X(n32906) );
  inv_x1_sg U38676 ( .A(n32905), .X(n32907) );
  inv_x1_sg U38677 ( .A(n32905), .X(n32908) );
  inv_x1_sg U38678 ( .A(n32905), .X(n32909) );
  inv_x1_sg U38679 ( .A(n13104), .X(n32910) );
  inv_x1_sg U38680 ( .A(n32910), .X(n32911) );
  inv_x1_sg U38681 ( .A(n32910), .X(n32912) );
  inv_x1_sg U38682 ( .A(n32910), .X(n32913) );
  inv_x1_sg U38683 ( .A(n32910), .X(n32914) );
  inv_x1_sg U38684 ( .A(n35374), .X(n32915) );
  inv_x1_sg U38685 ( .A(n32915), .X(n32916) );
  inv_x1_sg U38686 ( .A(n32915), .X(n32917) );
  inv_x1_sg U38687 ( .A(n32915), .X(n32918) );
  inv_x1_sg U38688 ( .A(n32915), .X(n32919) );
  inv_x1_sg U38689 ( .A(n35315), .X(n32920) );
  inv_x1_sg U38690 ( .A(n32920), .X(n32921) );
  inv_x1_sg U38691 ( .A(n32920), .X(n32922) );
  inv_x1_sg U38692 ( .A(n32920), .X(n32923) );
  inv_x1_sg U38693 ( .A(n32920), .X(n32924) );
  inv_x1_sg U38694 ( .A(n30962), .X(n32925) );
  inv_x1_sg U38695 ( .A(n30635), .X(n32926) );
  inv_x1_sg U38696 ( .A(n34854), .X(n32927) );
  inv_x1_sg U38697 ( .A(n32927), .X(n32928) );
  inv_x1_sg U38698 ( .A(n32927), .X(n32929) );
  inv_x1_sg U38699 ( .A(n32927), .X(n32930) );
  inv_x1_sg U38700 ( .A(n32927), .X(n32931) );
  inv_x1_sg U38701 ( .A(\shifter_0/pointer[2] ), .X(n32932) );
  inv_x1_sg U38702 ( .A(\shifter_0/pointer[2] ), .X(n32933) );
  inv_x1_sg U38703 ( .A(\shifter_0/pointer[2] ), .X(n32934) );
  inv_x1_sg U38704 ( .A(n32932), .X(n32935) );
  inv_x1_sg U38705 ( .A(n32934), .X(n32936) );
  inv_x1_sg U38706 ( .A(n32933), .X(n32937) );
  inv_x1_sg U38707 ( .A(n32934), .X(n32938) );
  inv_x1_sg U38708 ( .A(n32932), .X(n32939) );
  inv_x1_sg U38709 ( .A(n32933), .X(n32940) );
  inv_x1_sg U38710 ( .A(n31255), .X(n32941) );
  inv_x1_sg U38711 ( .A(n31256), .X(n32942) );
  inv_x1_sg U38712 ( .A(n31261), .X(n32943) );
  inv_x1_sg U38713 ( .A(n31260), .X(n32944) );
  inv_x1_sg U38714 ( .A(n31265), .X(n32945) );
  inv_x1_sg U38715 ( .A(n31265), .X(n32946) );
  inv_x1_sg U38716 ( .A(n31270), .X(n32947) );
  inv_x1_sg U38717 ( .A(n31270), .X(n32948) );
  inv_x1_sg U38718 ( .A(n31275), .X(n32949) );
  inv_x1_sg U38719 ( .A(n31274), .X(n32950) );
  inv_x1_sg U38720 ( .A(n34823), .X(n32951) );
  inv_x1_sg U38721 ( .A(n32951), .X(n32952) );
  inv_x1_sg U38722 ( .A(n32951), .X(n32953) );
  inv_x1_sg U38723 ( .A(n32951), .X(n32954) );
  inv_x1_sg U38724 ( .A(n32951), .X(n32955) );
  inv_x1_sg U38725 ( .A(n30372), .X(n32956) );
  inv_x1_sg U38726 ( .A(n30372), .X(n32957) );
  inv_x1_sg U38727 ( .A(n34818), .X(n32958) );
  inv_x1_sg U38728 ( .A(n32958), .X(n32959) );
  inv_x1_sg U38729 ( .A(n32958), .X(n32960) );
  inv_x1_sg U38730 ( .A(n32958), .X(n32961) );
  inv_x1_sg U38731 ( .A(n32958), .X(n32962) );
  inv_x1_sg U38732 ( .A(n30369), .X(n32963) );
  inv_x1_sg U38733 ( .A(n30369), .X(n32964) );
  inv_x1_sg U38734 ( .A(n34814), .X(n32965) );
  inv_x1_sg U38735 ( .A(n32965), .X(n32966) );
  inv_x1_sg U38736 ( .A(n32965), .X(n32967) );
  inv_x1_sg U38737 ( .A(n32965), .X(n32968) );
  inv_x1_sg U38738 ( .A(n32965), .X(n32969) );
  inv_x1_sg U38739 ( .A(n30366), .X(n32970) );
  inv_x1_sg U38740 ( .A(n30366), .X(n32971) );
  inv_x1_sg U38741 ( .A(n34810), .X(n32972) );
  inv_x1_sg U38742 ( .A(n29795), .X(n32973) );
  inv_x1_sg U38743 ( .A(n32972), .X(n32974) );
  inv_x1_sg U38744 ( .A(n32972), .X(n32975) );
  inv_x1_sg U38745 ( .A(n29795), .X(n32976) );
  inv_x1_sg U38746 ( .A(n34809), .X(n32977) );
  inv_x1_sg U38747 ( .A(n29797), .X(n32978) );
  inv_x1_sg U38748 ( .A(n32977), .X(n32979) );
  inv_x1_sg U38749 ( .A(n32977), .X(n32980) );
  inv_x1_sg U38750 ( .A(n32977), .X(n32981) );
  inv_x1_sg U38751 ( .A(n41321), .X(n32982) );
  inv_x1_sg U38752 ( .A(n32982), .X(n32983) );
  inv_x1_sg U38753 ( .A(n32982), .X(n32984) );
  inv_x1_sg U38754 ( .A(n32982), .X(n32985) );
  inv_x1_sg U38755 ( .A(n32982), .X(n32986) );
  inv_x1_sg U38756 ( .A(n35408), .X(n32987) );
  inv_x1_sg U38757 ( .A(n32987), .X(n32988) );
  inv_x1_sg U38758 ( .A(n32987), .X(n32989) );
  inv_x1_sg U38759 ( .A(n32987), .X(n32990) );
  inv_x1_sg U38760 ( .A(n32987), .X(n32991) );
  inv_x1_sg U38761 ( .A(n35407), .X(n32992) );
  inv_x1_sg U38762 ( .A(n32992), .X(n32993) );
  inv_x1_sg U38763 ( .A(n32992), .X(n32994) );
  inv_x1_sg U38764 ( .A(n32992), .X(n32995) );
  inv_x1_sg U38765 ( .A(n32992), .X(n32996) );
  inv_x1_sg U38766 ( .A(n35406), .X(n32997) );
  inv_x1_sg U38767 ( .A(n32997), .X(n32998) );
  inv_x1_sg U38768 ( .A(n32997), .X(n32999) );
  inv_x1_sg U38769 ( .A(n32997), .X(n33000) );
  inv_x1_sg U38770 ( .A(n32997), .X(n33001) );
  inv_x1_sg U38771 ( .A(n35405), .X(n33002) );
  inv_x1_sg U38772 ( .A(n33002), .X(n33003) );
  inv_x1_sg U38773 ( .A(n33002), .X(n33004) );
  inv_x1_sg U38774 ( .A(n33002), .X(n33005) );
  inv_x1_sg U38775 ( .A(n33002), .X(n33006) );
  inv_x1_sg U38776 ( .A(n35246), .X(n33007) );
  inv_x1_sg U38777 ( .A(n33007), .X(n33008) );
  inv_x1_sg U38778 ( .A(n33007), .X(n33009) );
  inv_x1_sg U38779 ( .A(n33007), .X(n33010) );
  inv_x1_sg U38780 ( .A(n33007), .X(n33011) );
  inv_x1_sg U38781 ( .A(n35245), .X(n33012) );
  inv_x1_sg U38782 ( .A(n33012), .X(n33013) );
  inv_x1_sg U38783 ( .A(n33012), .X(n33014) );
  inv_x1_sg U38784 ( .A(n33012), .X(n33015) );
  inv_x1_sg U38785 ( .A(n33012), .X(n33016) );
  inv_x1_sg U38786 ( .A(n35244), .X(n33017) );
  inv_x1_sg U38787 ( .A(n33017), .X(n33018) );
  inv_x1_sg U38788 ( .A(n33017), .X(n33019) );
  inv_x1_sg U38789 ( .A(n33017), .X(n33020) );
  inv_x1_sg U38790 ( .A(n33017), .X(n33021) );
  inv_x1_sg U38791 ( .A(n35243), .X(n33022) );
  inv_x1_sg U38792 ( .A(n33022), .X(n33023) );
  inv_x1_sg U38793 ( .A(n33022), .X(n33024) );
  inv_x1_sg U38794 ( .A(n33022), .X(n33025) );
  inv_x1_sg U38795 ( .A(n33022), .X(n33026) );
  inv_x1_sg U38796 ( .A(n35242), .X(n33027) );
  inv_x1_sg U38797 ( .A(n33027), .X(n33028) );
  inv_x1_sg U38798 ( .A(n33027), .X(n33029) );
  inv_x1_sg U38799 ( .A(n33027), .X(n33030) );
  inv_x1_sg U38800 ( .A(n33027), .X(n33031) );
  inv_x1_sg U38801 ( .A(n35241), .X(n33032) );
  inv_x1_sg U38802 ( .A(n33032), .X(n33033) );
  inv_x1_sg U38803 ( .A(n33032), .X(n33034) );
  inv_x1_sg U38804 ( .A(n33032), .X(n33035) );
  inv_x1_sg U38805 ( .A(n33032), .X(n33036) );
  inv_x1_sg U38806 ( .A(n35409), .X(n33037) );
  inv_x1_sg U38807 ( .A(n33037), .X(n33038) );
  inv_x1_sg U38808 ( .A(n33037), .X(n33039) );
  inv_x1_sg U38809 ( .A(n33037), .X(n33040) );
  inv_x1_sg U38810 ( .A(n35031), .X(n33041) );
  inv_x1_sg U38811 ( .A(n30245), .X(n33042) );
  inv_x1_sg U38812 ( .A(n35047), .X(n33043) );
  inv_x1_sg U38813 ( .A(n33043), .X(n33044) );
  inv_x1_sg U38814 ( .A(n33043), .X(n33045) );
  inv_x1_sg U38815 ( .A(n33043), .X(n33046) );
  inv_x1_sg U38816 ( .A(n33043), .X(n33047) );
  inv_x1_sg U38817 ( .A(n31591), .X(n33048) );
  inv_x1_sg U38818 ( .A(n33048), .X(n33049) );
  inv_x1_sg U38819 ( .A(n33048), .X(n33050) );
  inv_x1_sg U38820 ( .A(n33048), .X(n33051) );
  inv_x1_sg U38821 ( .A(n33048), .X(n33052) );
  inv_x1_sg U38822 ( .A(n35031), .X(n33053) );
  inv_x1_sg U38823 ( .A(n30604), .X(n33054) );
  inv_x1_sg U38824 ( .A(n35044), .X(n33055) );
  inv_x1_sg U38825 ( .A(n29803), .X(n33056) );
  inv_x1_sg U38826 ( .A(n29803), .X(n33057) );
  inv_x1_sg U38827 ( .A(n33055), .X(n33058) );
  inv_x1_sg U38828 ( .A(n33055), .X(n33059) );
  inv_x1_sg U38829 ( .A(n30246), .X(n33060) );
  inv_x1_sg U38830 ( .A(n29806), .X(n33061) );
  inv_x1_sg U38831 ( .A(n29806), .X(n33062) );
  inv_x1_sg U38832 ( .A(n33060), .X(n33063) );
  inv_x1_sg U38833 ( .A(n33060), .X(n33064) );
  inv_x1_sg U38834 ( .A(n35013), .X(n33065) );
  inv_x1_sg U38835 ( .A(n31112), .X(n33066) );
  inv_x1_sg U38836 ( .A(n30605), .X(n33067) );
  inv_x1_sg U38837 ( .A(n29809), .X(n33068) );
  inv_x1_sg U38838 ( .A(n29809), .X(n33069) );
  inv_x1_sg U38839 ( .A(n33067), .X(n33070) );
  inv_x1_sg U38840 ( .A(n33067), .X(n33071) );
  inv_x1_sg U38841 ( .A(n31572), .X(n33072) );
  inv_x1_sg U38842 ( .A(n29812), .X(n33073) );
  inv_x1_sg U38843 ( .A(n29812), .X(n33074) );
  inv_x1_sg U38844 ( .A(n33072), .X(n33075) );
  inv_x1_sg U38845 ( .A(n33072), .X(n33076) );
  inv_x1_sg U38846 ( .A(n30601), .X(n33077) );
  inv_x1_sg U38847 ( .A(n30606), .X(n33078) );
  inv_x1_sg U38848 ( .A(n31111), .X(n33079) );
  inv_x1_sg U38849 ( .A(n29817), .X(n33080) );
  inv_x1_sg U38850 ( .A(n29817), .X(n33081) );
  inv_x1_sg U38851 ( .A(n33079), .X(n33082) );
  inv_x1_sg U38852 ( .A(n33079), .X(n33083) );
  inv_x1_sg U38853 ( .A(n35036), .X(n33084) );
  inv_x1_sg U38854 ( .A(n29820), .X(n33085) );
  inv_x1_sg U38855 ( .A(n33084), .X(n33086) );
  inv_x1_sg U38856 ( .A(n29820), .X(n33087) );
  inv_x1_sg U38857 ( .A(n33084), .X(n33088) );
  inv_x1_sg U38858 ( .A(n30239), .X(n33089) );
  inv_x1_sg U38859 ( .A(n35014), .X(n33090) );
  inv_x1_sg U38860 ( .A(n35027), .X(n33091) );
  inv_x1_sg U38861 ( .A(n33091), .X(n33092) );
  inv_x1_sg U38862 ( .A(n30242), .X(n33093) );
  inv_x1_sg U38863 ( .A(n33091), .X(n33094) );
  inv_x1_sg U38864 ( .A(n33091), .X(n33095) );
  inv_x1_sg U38865 ( .A(n30244), .X(n33096) );
  inv_x1_sg U38866 ( .A(n33096), .X(n33097) );
  inv_x1_sg U38867 ( .A(n29823), .X(n33098) );
  inv_x1_sg U38868 ( .A(n33096), .X(n33099) );
  inv_x1_sg U38869 ( .A(n29823), .X(n33100) );
  inv_x1_sg U38870 ( .A(n35013), .X(n33101) );
  inv_x1_sg U38871 ( .A(n31575), .X(n33102) );
  inv_x1_sg U38872 ( .A(n35024), .X(n33103) );
  inv_x1_sg U38873 ( .A(n33103), .X(n33104) );
  inv_x1_sg U38874 ( .A(n33103), .X(n33105) );
  inv_x1_sg U38875 ( .A(n33103), .X(n33106) );
  inv_x1_sg U38876 ( .A(n33103), .X(n33107) );
  inv_x1_sg U38877 ( .A(n30241), .X(n33108) );
  inv_x1_sg U38878 ( .A(n33108), .X(n33109) );
  inv_x1_sg U38879 ( .A(n33108), .X(n33110) );
  inv_x1_sg U38880 ( .A(n33108), .X(n33111) );
  inv_x1_sg U38881 ( .A(n29828), .X(n33112) );
  inv_x1_sg U38882 ( .A(n35011), .X(n33113) );
  inv_x1_sg U38883 ( .A(n31589), .X(n33114) );
  inv_x1_sg U38884 ( .A(n35019), .X(n33115) );
  inv_x1_sg U38885 ( .A(n33115), .X(n33116) );
  inv_x1_sg U38886 ( .A(n33115), .X(n33117) );
  inv_x1_sg U38887 ( .A(n33115), .X(n33118) );
  inv_x1_sg U38888 ( .A(n29832), .X(n33119) );
  inv_x1_sg U38889 ( .A(n31577), .X(n33120) );
  inv_x1_sg U38890 ( .A(n33120), .X(n33121) );
  inv_x1_sg U38891 ( .A(n33120), .X(n33122) );
  inv_x1_sg U38892 ( .A(n33120), .X(n33123) );
  inv_x1_sg U38893 ( .A(n33120), .X(n33124) );
  inv_x1_sg U38894 ( .A(n35034), .X(n33125) );
  inv_x1_sg U38895 ( .A(n31574), .X(n33126) );
  inv_x1_sg U38896 ( .A(n35021), .X(n33127) );
  inv_x1_sg U38897 ( .A(n29835), .X(n33128) );
  inv_x1_sg U38898 ( .A(n29835), .X(n33129) );
  inv_x1_sg U38899 ( .A(n33127), .X(n33130) );
  inv_x1_sg U38900 ( .A(n33127), .X(n33131) );
  inv_x1_sg U38901 ( .A(n34993), .X(n33132) );
  inv_x1_sg U38902 ( .A(n31558), .X(n33133) );
  inv_x1_sg U38903 ( .A(n35006), .X(n33134) );
  inv_x1_sg U38904 ( .A(n29838), .X(n33135) );
  inv_x1_sg U38905 ( .A(n33134), .X(n33136) );
  inv_x1_sg U38906 ( .A(n33134), .X(n33137) );
  inv_x1_sg U38907 ( .A(n33134), .X(n33138) );
  inv_x1_sg U38908 ( .A(n35007), .X(n33139) );
  inv_x1_sg U38909 ( .A(n29841), .X(n33140) );
  inv_x1_sg U38910 ( .A(n33139), .X(n33141) );
  inv_x1_sg U38911 ( .A(n33139), .X(n33142) );
  inv_x1_sg U38912 ( .A(n33139), .X(n33143) );
  inv_x1_sg U38913 ( .A(n34993), .X(n33144) );
  inv_x1_sg U38914 ( .A(n31559), .X(n33145) );
  inv_x1_sg U38915 ( .A(n35003), .X(n33146) );
  inv_x1_sg U38916 ( .A(n33146), .X(n33147) );
  inv_x1_sg U38917 ( .A(n30237), .X(n33148) );
  inv_x1_sg U38918 ( .A(n33146), .X(n33149) );
  inv_x1_sg U38919 ( .A(n33146), .X(n33150) );
  inv_x1_sg U38920 ( .A(n35002), .X(n33151) );
  inv_x1_sg U38921 ( .A(n30235), .X(n33152) );
  inv_x1_sg U38922 ( .A(n33151), .X(n33153) );
  inv_x1_sg U38923 ( .A(n30235), .X(n33154) );
  inv_x1_sg U38924 ( .A(n33151), .X(n33155) );
  inv_x1_sg U38925 ( .A(n31113), .X(n33156) );
  inv_x1_sg U38926 ( .A(n34990), .X(n33157) );
  inv_x1_sg U38927 ( .A(n34999), .X(n33158) );
  inv_x1_sg U38928 ( .A(n33158), .X(n33159) );
  inv_x1_sg U38929 ( .A(n33158), .X(n33160) );
  inv_x1_sg U38930 ( .A(n33158), .X(n33161) );
  inv_x1_sg U38931 ( .A(n30232), .X(n33162) );
  inv_x1_sg U38932 ( .A(n30232), .X(n33163) );
  inv_x1_sg U38933 ( .A(n29848), .X(n33164) );
  inv_x1_sg U38934 ( .A(n30232), .X(n33165) );
  inv_x1_sg U38935 ( .A(n29848), .X(n33166) );
  inv_x1_sg U38936 ( .A(n34992), .X(n33167) );
  inv_x1_sg U38937 ( .A(n35248), .X(n33168) );
  inv_x1_sg U38938 ( .A(n34995), .X(n33169) );
  inv_x1_sg U38939 ( .A(n33169), .X(n33170) );
  inv_x1_sg U38940 ( .A(n33169), .X(n33171) );
  inv_x1_sg U38941 ( .A(n33169), .X(n33172) );
  inv_x1_sg U38942 ( .A(n33169), .X(n33173) );
  inv_x1_sg U38943 ( .A(n34994), .X(n33174) );
  inv_x1_sg U38944 ( .A(n33174), .X(n33175) );
  inv_x1_sg U38945 ( .A(n33174), .X(n33176) );
  inv_x1_sg U38946 ( .A(n33174), .X(n33177) );
  inv_x1_sg U38947 ( .A(n30229), .X(n33178) );
  inv_x1_sg U38948 ( .A(n30607), .X(n33179) );
  inv_x1_sg U38949 ( .A(n30969), .X(n33180) );
  inv_x1_sg U38950 ( .A(n30228), .X(n33181) );
  inv_x1_sg U38951 ( .A(n29852), .X(n33182) );
  inv_x1_sg U38952 ( .A(n33181), .X(n33183) );
  inv_x1_sg U38953 ( .A(n29852), .X(n33184) );
  inv_x1_sg U38954 ( .A(n33181), .X(n33185) );
  inv_x1_sg U38955 ( .A(n34986), .X(n33186) );
  inv_x1_sg U38956 ( .A(n29855), .X(n33187) );
  inv_x1_sg U38957 ( .A(n33186), .X(n33188) );
  inv_x1_sg U38958 ( .A(n33186), .X(n33189) );
  inv_x1_sg U38959 ( .A(n33186), .X(n33190) );
  inv_x1_sg U38960 ( .A(n30217), .X(n33191) );
  inv_x1_sg U38961 ( .A(n30217), .X(n33192) );
  inv_x1_sg U38962 ( .A(n34983), .X(n33193) );
  inv_x1_sg U38963 ( .A(n30225), .X(n33194) );
  inv_x1_sg U38964 ( .A(n30225), .X(n33195) );
  inv_x1_sg U38965 ( .A(n33193), .X(n33196) );
  inv_x1_sg U38966 ( .A(n33193), .X(n33197) );
  inv_x1_sg U38967 ( .A(n34982), .X(n33198) );
  inv_x1_sg U38968 ( .A(n29859), .X(n33199) );
  inv_x1_sg U38969 ( .A(n33198), .X(n33200) );
  inv_x1_sg U38970 ( .A(n33198), .X(n33201) );
  inv_x1_sg U38971 ( .A(n33198), .X(n33202) );
  inv_x1_sg U38972 ( .A(n34970), .X(n33203) );
  inv_x1_sg U38973 ( .A(n30969), .X(n33204) );
  inv_x1_sg U38974 ( .A(n34979), .X(n33205) );
  inv_x1_sg U38975 ( .A(n33205), .X(n33206) );
  inv_x1_sg U38976 ( .A(n33205), .X(n33207) );
  inv_x1_sg U38977 ( .A(n29862), .X(n33208) );
  inv_x1_sg U38978 ( .A(n33205), .X(n33209) );
  inv_x1_sg U38979 ( .A(n34978), .X(n33210) );
  inv_x1_sg U38980 ( .A(n30221), .X(n33211) );
  inv_x1_sg U38981 ( .A(n30221), .X(n33212) );
  inv_x1_sg U38982 ( .A(n33210), .X(n33213) );
  inv_x1_sg U38983 ( .A(n33210), .X(n33214) );
  inv_x1_sg U38984 ( .A(n31231), .X(n33215) );
  inv_x1_sg U38985 ( .A(n34972), .X(n33216) );
  inv_x1_sg U38986 ( .A(n34975), .X(n33217) );
  inv_x1_sg U38987 ( .A(n29866), .X(n33218) );
  inv_x1_sg U38988 ( .A(n29866), .X(n33219) );
  inv_x1_sg U38989 ( .A(n33217), .X(n33220) );
  inv_x1_sg U38990 ( .A(n33217), .X(n33221) );
  inv_x1_sg U38991 ( .A(n34841), .X(n33222) );
  inv_x1_sg U38992 ( .A(n34831), .X(n33223) );
  inv_x1_sg U38993 ( .A(n34841), .X(n33224) );
  inv_x1_sg U38994 ( .A(n34841), .X(n33225) );
  inv_x1_sg U38995 ( .A(n34842), .X(n33226) );
  inv_x1_sg U38996 ( .A(n33226), .X(n33227) );
  inv_x1_sg U38997 ( .A(n33226), .X(n33228) );
  inv_x1_sg U38998 ( .A(n33226), .X(n33229) );
  inv_x1_sg U38999 ( .A(n33226), .X(n33230) );
  inv_x1_sg U39000 ( .A(n34838), .X(n33231) );
  inv_x1_sg U39001 ( .A(n33231), .X(n33232) );
  inv_x1_sg U39002 ( .A(n33231), .X(n33233) );
  inv_x1_sg U39003 ( .A(n33231), .X(n33234) );
  inv_x1_sg U39004 ( .A(n33231), .X(n33235) );
  inv_x1_sg U39005 ( .A(n34837), .X(n33236) );
  inv_x1_sg U39006 ( .A(n33236), .X(n33237) );
  inv_x1_sg U39007 ( .A(n33236), .X(n33238) );
  inv_x1_sg U39008 ( .A(n33236), .X(n33239) );
  inv_x1_sg U39009 ( .A(n33236), .X(n33240) );
  inv_x1_sg U39010 ( .A(n34833), .X(n33241) );
  inv_x1_sg U39011 ( .A(n29896), .X(n33242) );
  inv_x1_sg U39012 ( .A(n33241), .X(n33243) );
  inv_x1_sg U39013 ( .A(n33241), .X(n33244) );
  inv_x1_sg U39014 ( .A(n33241), .X(n33245) );
  inv_x1_sg U39015 ( .A(n29900), .X(n33246) );
  inv_x1_sg U39016 ( .A(n29870), .X(n33247) );
  inv_x1_sg U39017 ( .A(n29870), .X(n33248) );
  inv_x1_sg U39018 ( .A(n29896), .X(n33249) );
  inv_x1_sg U39019 ( .A(n29900), .X(n33250) );
  inv_x1_sg U39020 ( .A(n33241), .X(n33251) );
  inv_x1_sg U39021 ( .A(n31269), .X(n33252) );
  inv_x1_sg U39022 ( .A(n29900), .X(n33253) );
  inv_x1_sg U39023 ( .A(n34827), .X(n33254) );
  inv_x1_sg U39024 ( .A(n29902), .X(n33255) );
  inv_x1_sg U39025 ( .A(n29902), .X(n33256) );
  inv_x1_sg U39026 ( .A(n33254), .X(n33257) );
  inv_x1_sg U39027 ( .A(n33254), .X(n33258) );
  inv_x1_sg U39028 ( .A(n34824), .X(n33259) );
  inv_x1_sg U39029 ( .A(n29904), .X(n33260) );
  inv_x1_sg U39030 ( .A(n29904), .X(n33261) );
  inv_x1_sg U39031 ( .A(n33259), .X(n33262) );
  inv_x1_sg U39032 ( .A(n33259), .X(n33263) );
  inv_x1_sg U39033 ( .A(n34819), .X(n33264) );
  inv_x1_sg U39034 ( .A(n33264), .X(n33265) );
  inv_x1_sg U39035 ( .A(n33264), .X(n33266) );
  inv_x1_sg U39036 ( .A(n33264), .X(n33267) );
  inv_x1_sg U39037 ( .A(n33264), .X(n33268) );
  inv_x1_sg U39038 ( .A(n34813), .X(n33269) );
  inv_x1_sg U39039 ( .A(n33269), .X(n33270) );
  inv_x1_sg U39040 ( .A(n33269), .X(n33271) );
  inv_x1_sg U39041 ( .A(n33269), .X(n33272) );
  inv_x1_sg U39042 ( .A(n33269), .X(n33273) );
  inv_x1_sg U39043 ( .A(n35642), .X(n33274) );
  inv_x1_sg U39044 ( .A(n33274), .X(n33275) );
  inv_x1_sg U39045 ( .A(n29908), .X(n33276) );
  inv_x1_sg U39046 ( .A(n33274), .X(n33277) );
  inv_x1_sg U39047 ( .A(n29908), .X(n33278) );
  inv_x1_sg U39048 ( .A(n35648), .X(n33279) );
  inv_x1_sg U39049 ( .A(n33279), .X(n33280) );
  inv_x1_sg U39050 ( .A(n29910), .X(n33281) );
  inv_x1_sg U39051 ( .A(n33279), .X(n33282) );
  inv_x1_sg U39052 ( .A(n29910), .X(n33283) );
  inv_x1_sg U39053 ( .A(n12976), .X(n33284) );
  inv_x1_sg U39054 ( .A(n33284), .X(n33285) );
  inv_x1_sg U39055 ( .A(n29912), .X(n33286) );
  inv_x1_sg U39056 ( .A(n33284), .X(n33287) );
  inv_x1_sg U39057 ( .A(n29912), .X(n33288) );
  inv_x1_sg U39058 ( .A(n12353), .X(n33289) );
  inv_x1_sg U39059 ( .A(n33289), .X(n33290) );
  inv_x1_sg U39060 ( .A(n29914), .X(n33291) );
  inv_x1_sg U39061 ( .A(n33289), .X(n33292) );
  inv_x1_sg U39062 ( .A(n29914), .X(n33293) );
  inv_x1_sg U39063 ( .A(n35659), .X(n33294) );
  inv_x1_sg U39064 ( .A(n33294), .X(n33295) );
  inv_x1_sg U39065 ( .A(n33294), .X(n33296) );
  inv_x1_sg U39066 ( .A(n33294), .X(n33297) );
  inv_x1_sg U39067 ( .A(n33294), .X(n33298) );
  inv_x1_sg U39068 ( .A(n29492), .X(n33299) );
  inv_x1_sg U39069 ( .A(n33299), .X(n33300) );
  inv_x1_sg U39070 ( .A(n33299), .X(n33301) );
  inv_x1_sg U39071 ( .A(n33299), .X(n33302) );
  inv_x1_sg U39072 ( .A(n33299), .X(n33303) );
  inv_x1_sg U39073 ( .A(n28978), .X(n33304) );
  inv_x1_sg U39074 ( .A(n33304), .X(n33305) );
  inv_x1_sg U39075 ( .A(n33304), .X(n33306) );
  inv_x1_sg U39076 ( .A(n33304), .X(n33307) );
  inv_x1_sg U39077 ( .A(n33304), .X(n33308) );
  inv_x1_sg U39078 ( .A(n35662), .X(n33309) );
  inv_x1_sg U39079 ( .A(n33309), .X(n33310) );
  inv_x1_sg U39080 ( .A(n33309), .X(n33311) );
  inv_x1_sg U39081 ( .A(n33309), .X(n33312) );
  inv_x1_sg U39082 ( .A(n33309), .X(n33313) );
  inv_x1_sg U39083 ( .A(n35668), .X(n33314) );
  inv_x1_sg U39084 ( .A(n33314), .X(n33315) );
  inv_x1_sg U39085 ( .A(n33314), .X(n33316) );
  inv_x1_sg U39086 ( .A(n33314), .X(n33317) );
  inv_x1_sg U39087 ( .A(n33314), .X(n33318) );
  inv_x1_sg U39088 ( .A(n35670), .X(n33319) );
  inv_x1_sg U39089 ( .A(n33319), .X(n33320) );
  inv_x1_sg U39090 ( .A(n33319), .X(n33321) );
  inv_x1_sg U39091 ( .A(n33319), .X(n33322) );
  inv_x1_sg U39092 ( .A(n33319), .X(n33323) );
  inv_x1_sg U39093 ( .A(n35658), .X(n33324) );
  inv_x1_sg U39094 ( .A(n33324), .X(n33325) );
  inv_x1_sg U39095 ( .A(n33324), .X(n33326) );
  inv_x1_sg U39096 ( .A(n33324), .X(n33327) );
  inv_x1_sg U39097 ( .A(n33324), .X(n33328) );
  inv_x1_sg U39098 ( .A(n35660), .X(n33329) );
  inv_x1_sg U39099 ( .A(n33329), .X(n33330) );
  inv_x1_sg U39100 ( .A(n33329), .X(n33331) );
  inv_x1_sg U39101 ( .A(n33329), .X(n33332) );
  inv_x1_sg U39102 ( .A(n33329), .X(n33333) );
  inv_x1_sg U39103 ( .A(n35671), .X(n33334) );
  inv_x1_sg U39104 ( .A(n33334), .X(n33335) );
  inv_x1_sg U39105 ( .A(n33334), .X(n33336) );
  inv_x1_sg U39106 ( .A(n33334), .X(n33337) );
  inv_x1_sg U39107 ( .A(n33334), .X(n33338) );
  inv_x1_sg U39108 ( .A(n35674), .X(n33339) );
  inv_x1_sg U39109 ( .A(n33339), .X(n33340) );
  inv_x1_sg U39110 ( .A(n33339), .X(n33341) );
  inv_x1_sg U39111 ( .A(n33339), .X(n33342) );
  inv_x1_sg U39112 ( .A(n33339), .X(n33343) );
  inv_x1_sg U39113 ( .A(n28452), .X(n33344) );
  inv_x1_sg U39114 ( .A(n33344), .X(n33345) );
  inv_x1_sg U39115 ( .A(n33344), .X(n33346) );
  inv_x1_sg U39116 ( .A(n33344), .X(n33347) );
  inv_x1_sg U39117 ( .A(n33344), .X(n33348) );
  inv_x1_sg U39118 ( .A(n35681), .X(n33349) );
  inv_x1_sg U39119 ( .A(n33349), .X(n33350) );
  inv_x1_sg U39120 ( .A(n33349), .X(n33351) );
  inv_x1_sg U39121 ( .A(n33349), .X(n33352) );
  inv_x1_sg U39122 ( .A(n33349), .X(n33353) );
  inv_x1_sg U39123 ( .A(n35672), .X(n33354) );
  inv_x1_sg U39124 ( .A(n33354), .X(n33355) );
  inv_x1_sg U39125 ( .A(n33354), .X(n33356) );
  inv_x1_sg U39126 ( .A(n33354), .X(n33357) );
  inv_x1_sg U39127 ( .A(n33354), .X(n33358) );
  inv_x1_sg U39128 ( .A(n28621), .X(n33359) );
  inv_x1_sg U39129 ( .A(n33359), .X(n33360) );
  inv_x1_sg U39130 ( .A(n33359), .X(n33361) );
  inv_x1_sg U39131 ( .A(n33359), .X(n33362) );
  inv_x1_sg U39132 ( .A(n33359), .X(n33363) );
  inv_x1_sg U39133 ( .A(n35680), .X(n33364) );
  inv_x1_sg U39134 ( .A(n33364), .X(n33365) );
  inv_x1_sg U39135 ( .A(n33364), .X(n33366) );
  inv_x1_sg U39136 ( .A(n33364), .X(n33367) );
  inv_x1_sg U39137 ( .A(n33364), .X(n33368) );
  inv_x1_sg U39138 ( .A(n28705), .X(n33369) );
  inv_x1_sg U39139 ( .A(n33369), .X(n33370) );
  inv_x1_sg U39140 ( .A(n33369), .X(n33371) );
  inv_x1_sg U39141 ( .A(n33369), .X(n33372) );
  inv_x1_sg U39142 ( .A(n33369), .X(n33373) );
  inv_x1_sg U39143 ( .A(n35673), .X(n33374) );
  inv_x1_sg U39144 ( .A(n33374), .X(n33375) );
  inv_x1_sg U39145 ( .A(n33374), .X(n33376) );
  inv_x1_sg U39146 ( .A(n33374), .X(n33377) );
  inv_x1_sg U39147 ( .A(n33374), .X(n33378) );
  inv_x1_sg U39148 ( .A(n35675), .X(n33379) );
  inv_x1_sg U39149 ( .A(n33379), .X(n33380) );
  inv_x1_sg U39150 ( .A(n33379), .X(n33381) );
  inv_x1_sg U39151 ( .A(n33379), .X(n33382) );
  inv_x1_sg U39152 ( .A(n33379), .X(n33383) );
  inv_x1_sg U39153 ( .A(n35678), .X(n33384) );
  inv_x1_sg U39154 ( .A(n33384), .X(n33385) );
  inv_x1_sg U39155 ( .A(n33384), .X(n33386) );
  inv_x1_sg U39156 ( .A(n33384), .X(n33387) );
  inv_x1_sg U39157 ( .A(n33384), .X(n33388) );
  inv_x1_sg U39158 ( .A(n29623), .X(n33389) );
  inv_x1_sg U39159 ( .A(n33389), .X(n33390) );
  inv_x1_sg U39160 ( .A(n33389), .X(n33391) );
  inv_x1_sg U39161 ( .A(n33389), .X(n33392) );
  inv_x1_sg U39162 ( .A(n33389), .X(n33393) );
  inv_x1_sg U39163 ( .A(n35664), .X(n33394) );
  inv_x1_sg U39164 ( .A(n33394), .X(n33395) );
  inv_x1_sg U39165 ( .A(n33394), .X(n33396) );
  inv_x1_sg U39166 ( .A(n33394), .X(n33397) );
  inv_x1_sg U39167 ( .A(n33394), .X(n33398) );
  inv_x1_sg U39168 ( .A(n29447), .X(n33399) );
  inv_x1_sg U39169 ( .A(n33399), .X(n33400) );
  inv_x1_sg U39170 ( .A(n33399), .X(n33401) );
  inv_x1_sg U39171 ( .A(n33399), .X(n33402) );
  inv_x1_sg U39172 ( .A(n33399), .X(n33403) );
  inv_x1_sg U39173 ( .A(n35663), .X(n33404) );
  inv_x1_sg U39174 ( .A(n33404), .X(n33405) );
  inv_x1_sg U39175 ( .A(n33404), .X(n33406) );
  inv_x1_sg U39176 ( .A(n33404), .X(n33407) );
  inv_x1_sg U39177 ( .A(n33404), .X(n33408) );
  inv_x1_sg U39178 ( .A(n12134), .X(n33409) );
  inv_x1_sg U39179 ( .A(n33409), .X(n33410) );
  inv_x1_sg U39180 ( .A(n29962), .X(n33411) );
  inv_x1_sg U39181 ( .A(n33409), .X(n33412) );
  inv_x1_sg U39182 ( .A(n29962), .X(n33413) );
  inv_x1_sg U39183 ( .A(n11906), .X(n33414) );
  inv_x1_sg U39184 ( .A(n33414), .X(n33415) );
  inv_x1_sg U39185 ( .A(n29964), .X(n33416) );
  inv_x1_sg U39186 ( .A(n33414), .X(n33417) );
  inv_x1_sg U39187 ( .A(n29964), .X(n33418) );
  inv_x1_sg U39188 ( .A(n11895), .X(n33419) );
  inv_x1_sg U39189 ( .A(n33419), .X(n33420) );
  inv_x1_sg U39190 ( .A(n29966), .X(n33421) );
  inv_x1_sg U39191 ( .A(n33419), .X(n33422) );
  inv_x1_sg U39192 ( .A(n29966), .X(n33423) );
  inv_x1_sg U39193 ( .A(n35651), .X(n33424) );
  inv_x1_sg U39194 ( .A(n33424), .X(n33425) );
  inv_x1_sg U39195 ( .A(n29968), .X(n33426) );
  inv_x1_sg U39196 ( .A(n33424), .X(n33427) );
  inv_x1_sg U39197 ( .A(n29968), .X(n33428) );
  inv_x1_sg U39198 ( .A(n35676), .X(n33429) );
  inv_x1_sg U39199 ( .A(n33429), .X(n33430) );
  inv_x1_sg U39200 ( .A(n33429), .X(n33431) );
  inv_x1_sg U39201 ( .A(n33429), .X(n33432) );
  inv_x1_sg U39202 ( .A(n33429), .X(n33433) );
  inv_x1_sg U39203 ( .A(n35665), .X(n33434) );
  inv_x1_sg U39204 ( .A(n33434), .X(n33435) );
  inv_x1_sg U39205 ( .A(n33434), .X(n33436) );
  inv_x1_sg U39206 ( .A(n33434), .X(n33437) );
  inv_x1_sg U39207 ( .A(n33434), .X(n33438) );
  inv_x1_sg U39208 ( .A(n35661), .X(n33439) );
  inv_x1_sg U39209 ( .A(n33439), .X(n33440) );
  inv_x1_sg U39210 ( .A(n33439), .X(n33441) );
  inv_x1_sg U39211 ( .A(n33439), .X(n33442) );
  inv_x1_sg U39212 ( .A(n33439), .X(n33443) );
  inv_x1_sg U39213 ( .A(n35679), .X(n33444) );
  inv_x1_sg U39214 ( .A(n33444), .X(n33445) );
  inv_x1_sg U39215 ( .A(n33444), .X(n33446) );
  inv_x1_sg U39216 ( .A(n33444), .X(n33447) );
  inv_x1_sg U39217 ( .A(n33444), .X(n33448) );
  inv_x1_sg U39218 ( .A(n35669), .X(n33449) );
  inv_x1_sg U39219 ( .A(n33449), .X(n33450) );
  inv_x1_sg U39220 ( .A(n33449), .X(n33451) );
  inv_x1_sg U39221 ( .A(n33449), .X(n33452) );
  inv_x1_sg U39222 ( .A(n33449), .X(n33453) );
  inv_x1_sg U39223 ( .A(n35667), .X(n33454) );
  inv_x1_sg U39224 ( .A(n33454), .X(n33455) );
  inv_x1_sg U39225 ( .A(n33454), .X(n33456) );
  inv_x1_sg U39226 ( .A(n33454), .X(n33457) );
  inv_x1_sg U39227 ( .A(n33454), .X(n33458) );
  inv_x1_sg U39228 ( .A(n35666), .X(n33459) );
  inv_x1_sg U39229 ( .A(n33459), .X(n33460) );
  inv_x1_sg U39230 ( .A(n33459), .X(n33461) );
  inv_x1_sg U39231 ( .A(n33459), .X(n33462) );
  inv_x1_sg U39232 ( .A(n33459), .X(n33463) );
  inv_x1_sg U39233 ( .A(n29064), .X(n33464) );
  inv_x1_sg U39234 ( .A(n33464), .X(n33465) );
  inv_x1_sg U39235 ( .A(n33464), .X(n33466) );
  inv_x1_sg U39236 ( .A(n33464), .X(n33467) );
  inv_x1_sg U39237 ( .A(n33464), .X(n33468) );
  inv_x1_sg U39238 ( .A(n35677), .X(n33469) );
  inv_x1_sg U39239 ( .A(n33469), .X(n33470) );
  inv_x1_sg U39240 ( .A(n33469), .X(n33471) );
  inv_x1_sg U39241 ( .A(n33469), .X(n33472) );
  inv_x1_sg U39242 ( .A(n33469), .X(n33473) );
  nand_x1_sg U39243 ( .A(n29487), .B(n29018), .X(n33474) );
  inv_x1_sg U39244 ( .A(n33477), .X(n33475) );
  inv_x1_sg U39245 ( .A(n33477), .X(n33476) );
  inv_x1_sg U39246 ( .A(n33474), .X(n33477) );
  inv_x1_sg U39247 ( .A(n33474), .X(n33478) );
  inv_x1_sg U39248 ( .A(n33477), .X(n33479) );
  inv_x1_sg U39249 ( .A(n33478), .X(n33480) );
  inv_x1_sg U39250 ( .A(n33478), .X(n33481) );
  nand_x1_sg U39251 ( .A(n29487), .B(n29061), .X(n33482) );
  inv_x1_sg U39252 ( .A(n33485), .X(n33483) );
  inv_x1_sg U39253 ( .A(n33485), .X(n33484) );
  inv_x1_sg U39254 ( .A(n33482), .X(n33485) );
  inv_x1_sg U39255 ( .A(n33482), .X(n33486) );
  inv_x1_sg U39256 ( .A(n33485), .X(n33487) );
  inv_x1_sg U39257 ( .A(n33486), .X(n33488) );
  inv_x1_sg U39258 ( .A(n33486), .X(n33489) );
  nand_x1_sg U39259 ( .A(n29018), .B(n35562), .X(n33490) );
  inv_x1_sg U39260 ( .A(n33493), .X(n33491) );
  inv_x1_sg U39261 ( .A(n33493), .X(n33492) );
  inv_x1_sg U39262 ( .A(n33490), .X(n33493) );
  inv_x1_sg U39263 ( .A(n33490), .X(n33494) );
  inv_x1_sg U39264 ( .A(n33493), .X(n33495) );
  inv_x1_sg U39265 ( .A(n33494), .X(n33496) );
  inv_x1_sg U39266 ( .A(n33494), .X(n33497) );
  nand_x1_sg U39267 ( .A(n29018), .B(n29317), .X(n33498) );
  inv_x1_sg U39268 ( .A(n33501), .X(n33499) );
  inv_x1_sg U39269 ( .A(n33501), .X(n33500) );
  inv_x1_sg U39270 ( .A(n33498), .X(n33501) );
  inv_x1_sg U39271 ( .A(n33498), .X(n33502) );
  inv_x1_sg U39272 ( .A(n33501), .X(n33503) );
  inv_x1_sg U39273 ( .A(n33502), .X(n33504) );
  inv_x1_sg U39274 ( .A(n33502), .X(n33505) );
  nand_x1_sg U39275 ( .A(n29018), .B(n29148), .X(n33506) );
  inv_x1_sg U39276 ( .A(n33509), .X(n33507) );
  inv_x1_sg U39277 ( .A(n33509), .X(n33508) );
  inv_x1_sg U39278 ( .A(n33506), .X(n33509) );
  inv_x1_sg U39279 ( .A(n33506), .X(n33510) );
  inv_x1_sg U39280 ( .A(n33509), .X(n33511) );
  inv_x1_sg U39281 ( .A(n33510), .X(n33512) );
  inv_x1_sg U39282 ( .A(n33510), .X(n33513) );
  nand_x1_sg U39283 ( .A(n29061), .B(n35562), .X(n33514) );
  inv_x1_sg U39284 ( .A(n33517), .X(n33515) );
  inv_x1_sg U39285 ( .A(n33517), .X(n33516) );
  inv_x1_sg U39286 ( .A(n33514), .X(n33517) );
  inv_x1_sg U39287 ( .A(n33514), .X(n33518) );
  inv_x1_sg U39288 ( .A(n33517), .X(n33519) );
  inv_x1_sg U39289 ( .A(n33518), .X(n33520) );
  inv_x1_sg U39290 ( .A(n33518), .X(n33521) );
  inv_x1_sg U39291 ( .A(n14411), .X(n33522) );
  inv_x1_sg U39292 ( .A(n33522), .X(n33523) );
  inv_x1_sg U39293 ( .A(n33522), .X(n33524) );
  inv_x1_sg U39294 ( .A(n33522), .X(n33525) );
  nand_x1_sg U39295 ( .A(n28448), .B(n28788), .X(n33526) );
  inv_x1_sg U39296 ( .A(n33529), .X(n33527) );
  inv_x1_sg U39297 ( .A(n33529), .X(n33528) );
  inv_x1_sg U39298 ( .A(n33526), .X(n33529) );
  inv_x1_sg U39299 ( .A(n33526), .X(n33530) );
  inv_x1_sg U39300 ( .A(n33529), .X(n33531) );
  inv_x1_sg U39301 ( .A(n33530), .X(n33532) );
  inv_x1_sg U39302 ( .A(n33530), .X(n33533) );
  nand_x1_sg U39303 ( .A(n29147), .B(n29317), .X(n33534) );
  inv_x1_sg U39304 ( .A(n33537), .X(n33535) );
  inv_x1_sg U39305 ( .A(n33537), .X(n33536) );
  inv_x1_sg U39306 ( .A(n33534), .X(n33537) );
  inv_x1_sg U39307 ( .A(n33534), .X(n33538) );
  inv_x1_sg U39308 ( .A(n33537), .X(n33539) );
  inv_x1_sg U39309 ( .A(n33538), .X(n33540) );
  inv_x1_sg U39310 ( .A(n33538), .X(n33541) );
  nand_x1_sg U39311 ( .A(n28319), .B(n28618), .X(n33542) );
  inv_x1_sg U39312 ( .A(n33545), .X(n33543) );
  inv_x1_sg U39313 ( .A(n33545), .X(n33544) );
  inv_x1_sg U39314 ( .A(n33542), .X(n33545) );
  inv_x1_sg U39315 ( .A(n33542), .X(n33546) );
  inv_x1_sg U39316 ( .A(n33545), .X(n33547) );
  inv_x1_sg U39317 ( .A(n33546), .X(n33548) );
  inv_x1_sg U39318 ( .A(n33546), .X(n33549) );
  nand_x1_sg U39319 ( .A(n28319), .B(n28788), .X(n33550) );
  inv_x1_sg U39320 ( .A(n33553), .X(n33551) );
  inv_x1_sg U39321 ( .A(n33553), .X(n33552) );
  inv_x1_sg U39322 ( .A(n33550), .X(n33553) );
  inv_x1_sg U39323 ( .A(n33550), .X(n33554) );
  inv_x1_sg U39324 ( .A(n33553), .X(n33555) );
  inv_x1_sg U39325 ( .A(n33554), .X(n33556) );
  inv_x1_sg U39326 ( .A(n33554), .X(n33557) );
  nand_x1_sg U39327 ( .A(n28405), .B(n35511), .X(n33558) );
  inv_x1_sg U39328 ( .A(n33561), .X(n33559) );
  inv_x1_sg U39329 ( .A(n33561), .X(n33560) );
  inv_x1_sg U39330 ( .A(n33558), .X(n33561) );
  inv_x1_sg U39331 ( .A(n33558), .X(n33562) );
  inv_x1_sg U39332 ( .A(n33561), .X(n33563) );
  inv_x1_sg U39333 ( .A(n33562), .X(n33564) );
  inv_x1_sg U39334 ( .A(n33562), .X(n33565) );
  nand_x1_sg U39335 ( .A(n28405), .B(n28618), .X(n33566) );
  inv_x1_sg U39336 ( .A(n33569), .X(n33567) );
  inv_x1_sg U39337 ( .A(n33569), .X(n33568) );
  inv_x1_sg U39338 ( .A(n33566), .X(n33569) );
  inv_x1_sg U39339 ( .A(n33566), .X(n33570) );
  inv_x1_sg U39340 ( .A(n33569), .X(n33571) );
  inv_x1_sg U39341 ( .A(n33570), .X(n33572) );
  inv_x1_sg U39342 ( .A(n33570), .X(n33573) );
  nand_x1_sg U39343 ( .A(n28405), .B(n28788), .X(n33574) );
  inv_x1_sg U39344 ( .A(n33577), .X(n33575) );
  inv_x1_sg U39345 ( .A(n33577), .X(n33576) );
  inv_x1_sg U39346 ( .A(n33574), .X(n33577) );
  inv_x1_sg U39347 ( .A(n33574), .X(n33578) );
  inv_x1_sg U39348 ( .A(n33577), .X(n33579) );
  inv_x1_sg U39349 ( .A(n33578), .X(n33580) );
  inv_x1_sg U39350 ( .A(n33578), .X(n33581) );
  nand_x1_sg U39351 ( .A(n28448), .B(n35511), .X(n33582) );
  inv_x1_sg U39352 ( .A(n33585), .X(n33583) );
  inv_x1_sg U39353 ( .A(n33585), .X(n33584) );
  inv_x1_sg U39354 ( .A(n33582), .X(n33585) );
  inv_x1_sg U39355 ( .A(n33582), .X(n33586) );
  inv_x1_sg U39356 ( .A(n33585), .X(n33587) );
  inv_x1_sg U39357 ( .A(n33586), .X(n33588) );
  inv_x1_sg U39358 ( .A(n33586), .X(n33589) );
  nand_x1_sg U39359 ( .A(n29147), .B(n29148), .X(n33590) );
  inv_x1_sg U39360 ( .A(n33593), .X(n33591) );
  inv_x1_sg U39361 ( .A(n33593), .X(n33592) );
  inv_x1_sg U39362 ( .A(n33590), .X(n33593) );
  inv_x1_sg U39363 ( .A(n33590), .X(n33594) );
  inv_x1_sg U39364 ( .A(n33593), .X(n33595) );
  inv_x1_sg U39365 ( .A(n33594), .X(n33596) );
  inv_x1_sg U39366 ( .A(n33594), .X(n33597) );
  nand_x1_sg U39367 ( .A(n29487), .B(n29104), .X(n33598) );
  inv_x1_sg U39368 ( .A(n33601), .X(n33599) );
  inv_x1_sg U39369 ( .A(n33601), .X(n33600) );
  inv_x1_sg U39370 ( .A(n33598), .X(n33601) );
  inv_x1_sg U39371 ( .A(n33598), .X(n33602) );
  inv_x1_sg U39372 ( .A(n33601), .X(n33603) );
  inv_x1_sg U39373 ( .A(n33602), .X(n33604) );
  inv_x1_sg U39374 ( .A(n33602), .X(n33605) );
  nand_x1_sg U39375 ( .A(n29104), .B(n29148), .X(n33606) );
  inv_x1_sg U39376 ( .A(n33609), .X(n33607) );
  inv_x1_sg U39377 ( .A(n33609), .X(n33608) );
  inv_x1_sg U39378 ( .A(n33606), .X(n33609) );
  inv_x1_sg U39379 ( .A(n33606), .X(n33610) );
  inv_x1_sg U39380 ( .A(n33609), .X(n33611) );
  inv_x1_sg U39381 ( .A(n33610), .X(n33612) );
  inv_x1_sg U39382 ( .A(n33610), .X(n33613) );
  nand_x1_sg U39383 ( .A(n29104), .B(n35562), .X(n33614) );
  inv_x1_sg U39384 ( .A(n33617), .X(n33615) );
  inv_x1_sg U39385 ( .A(n33617), .X(n33616) );
  inv_x1_sg U39386 ( .A(n33614), .X(n33617) );
  inv_x1_sg U39387 ( .A(n33614), .X(n33618) );
  inv_x1_sg U39388 ( .A(n33617), .X(n33619) );
  inv_x1_sg U39389 ( .A(n33618), .X(n33620) );
  inv_x1_sg U39390 ( .A(n33618), .X(n33621) );
  nand_x1_sg U39391 ( .A(n29104), .B(n29317), .X(n33622) );
  inv_x1_sg U39392 ( .A(n33625), .X(n33623) );
  inv_x1_sg U39393 ( .A(n33625), .X(n33624) );
  inv_x1_sg U39394 ( .A(n33622), .X(n33625) );
  inv_x1_sg U39395 ( .A(n33622), .X(n33626) );
  inv_x1_sg U39396 ( .A(n33625), .X(n33627) );
  inv_x1_sg U39397 ( .A(n33626), .X(n33628) );
  inv_x1_sg U39398 ( .A(n33626), .X(n33629) );
  inv_x1_sg U39399 ( .A(n35635), .X(n33630) );
  inv_x1_sg U39400 ( .A(n33630), .X(n33631) );
  inv_x1_sg U39401 ( .A(n33630), .X(n33632) );
  inv_x1_sg U39402 ( .A(n33630), .X(n33633) );
  inv_x1_sg U39403 ( .A(n35621), .X(n33634) );
  inv_x1_sg U39404 ( .A(n33634), .X(n33635) );
  inv_x1_sg U39405 ( .A(n33634), .X(n33636) );
  inv_x1_sg U39406 ( .A(n33634), .X(n33637) );
  nand_x1_sg U39407 ( .A(n28362), .B(n35511), .X(n33638) );
  inv_x1_sg U39408 ( .A(n33641), .X(n33639) );
  inv_x1_sg U39409 ( .A(n33641), .X(n33640) );
  inv_x1_sg U39410 ( .A(n33638), .X(n33641) );
  inv_x1_sg U39411 ( .A(n33638), .X(n33642) );
  inv_x1_sg U39412 ( .A(n33641), .X(n33643) );
  inv_x1_sg U39413 ( .A(n33642), .X(n33644) );
  inv_x1_sg U39414 ( .A(n33642), .X(n33645) );
  nand_x1_sg U39415 ( .A(n28362), .B(n28618), .X(n33646) );
  inv_x1_sg U39416 ( .A(n33649), .X(n33647) );
  inv_x1_sg U39417 ( .A(n33649), .X(n33648) );
  inv_x1_sg U39418 ( .A(n33646), .X(n33649) );
  inv_x1_sg U39419 ( .A(n33646), .X(n33650) );
  inv_x1_sg U39420 ( .A(n33649), .X(n33651) );
  inv_x1_sg U39421 ( .A(n33650), .X(n33652) );
  inv_x1_sg U39422 ( .A(n33650), .X(n33653) );
  nand_x1_sg U39423 ( .A(n29061), .B(n29148), .X(n33654) );
  inv_x1_sg U39424 ( .A(n33657), .X(n33655) );
  inv_x1_sg U39425 ( .A(n33657), .X(n33656) );
  inv_x1_sg U39426 ( .A(n33654), .X(n33657) );
  inv_x1_sg U39427 ( .A(n33654), .X(n33658) );
  inv_x1_sg U39428 ( .A(n33657), .X(n33659) );
  inv_x1_sg U39429 ( .A(n33658), .X(n33660) );
  inv_x1_sg U39430 ( .A(n33658), .X(n33661) );
  nand_x1_sg U39431 ( .A(n28362), .B(n28788), .X(n33662) );
  inv_x1_sg U39432 ( .A(n33665), .X(n33663) );
  inv_x1_sg U39433 ( .A(n33665), .X(n33664) );
  inv_x1_sg U39434 ( .A(n33662), .X(n33665) );
  inv_x1_sg U39435 ( .A(n33662), .X(n33666) );
  inv_x1_sg U39436 ( .A(n33665), .X(n33667) );
  inv_x1_sg U39437 ( .A(n33666), .X(n33668) );
  inv_x1_sg U39438 ( .A(n33666), .X(n33669) );
  nand_x1_sg U39439 ( .A(n29061), .B(n29317), .X(n33670) );
  inv_x1_sg U39440 ( .A(n33673), .X(n33671) );
  inv_x1_sg U39441 ( .A(n33673), .X(n33672) );
  inv_x1_sg U39442 ( .A(n33670), .X(n33673) );
  inv_x1_sg U39443 ( .A(n33670), .X(n33674) );
  inv_x1_sg U39444 ( .A(n33673), .X(n33675) );
  inv_x1_sg U39445 ( .A(n33674), .X(n33676) );
  inv_x1_sg U39446 ( .A(n33674), .X(n33677) );
  nand_x1_sg U39447 ( .A(n28448), .B(n28618), .X(n33678) );
  inv_x1_sg U39448 ( .A(n33681), .X(n33679) );
  inv_x1_sg U39449 ( .A(n33681), .X(n33680) );
  inv_x1_sg U39450 ( .A(n33678), .X(n33681) );
  inv_x1_sg U39451 ( .A(n33678), .X(n33682) );
  inv_x1_sg U39452 ( .A(n33681), .X(n33683) );
  inv_x1_sg U39453 ( .A(n33682), .X(n33684) );
  inv_x1_sg U39454 ( .A(n33682), .X(n33685) );
  nand_x1_sg U39455 ( .A(n28319), .B(n35511), .X(n33686) );
  inv_x1_sg U39456 ( .A(n33689), .X(n33687) );
  inv_x1_sg U39457 ( .A(n33689), .X(n33688) );
  inv_x1_sg U39458 ( .A(n33686), .X(n33689) );
  inv_x1_sg U39459 ( .A(n33686), .X(n33690) );
  inv_x1_sg U39460 ( .A(n33689), .X(n33691) );
  inv_x1_sg U39461 ( .A(n33690), .X(n33692) );
  inv_x1_sg U39462 ( .A(n33690), .X(n33693) );
  nand_x1_sg U39463 ( .A(n29147), .B(n29487), .X(n33694) );
  inv_x1_sg U39464 ( .A(n33697), .X(n33695) );
  inv_x1_sg U39465 ( .A(n33697), .X(n33696) );
  inv_x1_sg U39466 ( .A(n33694), .X(n33697) );
  inv_x1_sg U39467 ( .A(n33694), .X(n33698) );
  inv_x1_sg U39468 ( .A(n33697), .X(n33699) );
  inv_x1_sg U39469 ( .A(n33698), .X(n33700) );
  inv_x1_sg U39470 ( .A(n33698), .X(n33701) );
  nand_x1_sg U39471 ( .A(n29147), .B(n35562), .X(n33702) );
  inv_x1_sg U39472 ( .A(n33705), .X(n33703) );
  inv_x1_sg U39473 ( .A(n33705), .X(n33704) );
  inv_x1_sg U39474 ( .A(n33702), .X(n33705) );
  inv_x1_sg U39475 ( .A(n33702), .X(n33706) );
  inv_x1_sg U39476 ( .A(n33705), .X(n33707) );
  inv_x1_sg U39477 ( .A(n33706), .X(n33708) );
  inv_x1_sg U39478 ( .A(n33706), .X(n33709) );
  inv_x1_sg U39479 ( .A(n35624), .X(n33710) );
  inv_x1_sg U39480 ( .A(n33710), .X(n33711) );
  inv_x1_sg U39481 ( .A(n33710), .X(n33712) );
  inv_x1_sg U39482 ( .A(n33710), .X(n33713) );
  inv_x1_sg U39483 ( .A(n33710), .X(n33714) );
  inv_x1_sg U39484 ( .A(n35622), .X(n33715) );
  inv_x1_sg U39485 ( .A(n33715), .X(n33716) );
  inv_x1_sg U39486 ( .A(n33715), .X(n33717) );
  inv_x1_sg U39487 ( .A(n33715), .X(n33718) );
  inv_x1_sg U39488 ( .A(n35638), .X(n33719) );
  inv_x1_sg U39489 ( .A(n33719), .X(n33720) );
  inv_x1_sg U39490 ( .A(n33719), .X(n33721) );
  inv_x1_sg U39491 ( .A(n33719), .X(n33722) );
  inv_x1_sg U39492 ( .A(n35636), .X(n33723) );
  inv_x1_sg U39493 ( .A(n33723), .X(n33724) );
  inv_x1_sg U39494 ( .A(n33723), .X(n33725) );
  inv_x1_sg U39495 ( .A(n33723), .X(n33726) );
  inv_x1_sg U39496 ( .A(n35623), .X(n33727) );
  inv_x1_sg U39497 ( .A(n33727), .X(n33728) );
  inv_x1_sg U39498 ( .A(n33727), .X(n33729) );
  inv_x1_sg U39499 ( .A(n33727), .X(n33730) );
  inv_x1_sg U39500 ( .A(n33727), .X(n33731) );
  inv_x1_sg U39501 ( .A(n35639), .X(n33732) );
  inv_x1_sg U39502 ( .A(n33732), .X(n33733) );
  inv_x1_sg U39503 ( .A(n33732), .X(n33734) );
  inv_x1_sg U39504 ( .A(n33732), .X(n33735) );
  inv_x1_sg U39505 ( .A(n35637), .X(n33736) );
  inv_x1_sg U39506 ( .A(n33736), .X(n33737) );
  inv_x1_sg U39507 ( .A(n33736), .X(n33738) );
  inv_x1_sg U39508 ( .A(n33736), .X(n33739) );
  inv_x1_sg U39509 ( .A(n35620), .X(n33740) );
  inv_x1_sg U39510 ( .A(n33740), .X(n33741) );
  inv_x1_sg U39511 ( .A(n33740), .X(n33742) );
  inv_x1_sg U39512 ( .A(n33740), .X(n33743) );
  inv_x1_sg U39513 ( .A(n35649), .X(n33744) );
  inv_x1_sg U39514 ( .A(n33744), .X(n33745) );
  inv_x1_sg U39515 ( .A(n33744), .X(n33746) );
  inv_x1_sg U39516 ( .A(n33744), .X(n33747) );
  inv_x1_sg U39517 ( .A(n33744), .X(n33748) );
  inv_x1_sg U39518 ( .A(n35652), .X(n33749) );
  inv_x1_sg U39519 ( .A(n33749), .X(n33750) );
  inv_x1_sg U39520 ( .A(n33749), .X(n33751) );
  inv_x1_sg U39521 ( .A(n33749), .X(n33752) );
  inv_x1_sg U39522 ( .A(n30008), .X(n33754) );
  inv_x1_sg U39523 ( .A(n30008), .X(n33755) );
  inv_x1_sg U39524 ( .A(n33753), .X(n33756) );
  inv_x1_sg U39525 ( .A(n33753), .X(n33757) );
  inv_x1_sg U39526 ( .A(n30011), .X(n33759) );
  inv_x1_sg U39527 ( .A(n30011), .X(n33760) );
  inv_x1_sg U39528 ( .A(n33758), .X(n33761) );
  inv_x1_sg U39529 ( .A(n33758), .X(n33762) );
  nand_x1_sg U39530 ( .A(n28405), .B(n28449), .X(n33763) );
  inv_x1_sg U39531 ( .A(n33766), .X(n33764) );
  inv_x1_sg U39532 ( .A(n33766), .X(n33765) );
  inv_x1_sg U39533 ( .A(n33763), .X(n33766) );
  inv_x1_sg U39534 ( .A(n33763), .X(n33767) );
  inv_x1_sg U39535 ( .A(n33766), .X(n33768) );
  inv_x1_sg U39536 ( .A(n33767), .X(n33769) );
  inv_x1_sg U39537 ( .A(n33767), .X(n33770) );
  nand_x1_sg U39538 ( .A(n28448), .B(n28449), .X(n33771) );
  inv_x1_sg U39539 ( .A(n33774), .X(n33772) );
  inv_x1_sg U39540 ( .A(n33774), .X(n33773) );
  inv_x1_sg U39541 ( .A(n33771), .X(n33774) );
  inv_x1_sg U39542 ( .A(n33771), .X(n33775) );
  inv_x1_sg U39543 ( .A(n33774), .X(n33776) );
  inv_x1_sg U39544 ( .A(n33775), .X(n33777) );
  inv_x1_sg U39545 ( .A(n33775), .X(n33778) );
  nand_x1_sg U39546 ( .A(n28362), .B(n28449), .X(n33779) );
  inv_x1_sg U39547 ( .A(n33782), .X(n33780) );
  inv_x1_sg U39548 ( .A(n33782), .X(n33781) );
  inv_x1_sg U39549 ( .A(n33779), .X(n33782) );
  inv_x1_sg U39550 ( .A(n33779), .X(n33783) );
  inv_x1_sg U39551 ( .A(n33782), .X(n33784) );
  inv_x1_sg U39552 ( .A(n33783), .X(n33785) );
  inv_x1_sg U39553 ( .A(n33783), .X(n33786) );
  nand_x1_sg U39554 ( .A(n28319), .B(n28449), .X(n33787) );
  inv_x1_sg U39555 ( .A(n33790), .X(n33788) );
  inv_x1_sg U39556 ( .A(n33790), .X(n33789) );
  inv_x1_sg U39557 ( .A(n33787), .X(n33790) );
  inv_x1_sg U39558 ( .A(n33787), .X(n33791) );
  inv_x1_sg U39559 ( .A(n33790), .X(n33792) );
  inv_x1_sg U39560 ( .A(n33791), .X(n33793) );
  inv_x1_sg U39561 ( .A(n33791), .X(n33794) );
  inv_x1_sg U39562 ( .A(n12842), .X(n33795) );
  inv_x1_sg U39563 ( .A(n33795), .X(n33796) );
  inv_x1_sg U39564 ( .A(n33795), .X(n33797) );
  inv_x1_sg U39565 ( .A(n33795), .X(n33798) );
  inv_x1_sg U39566 ( .A(n35410), .X(n33799) );
  inv_x1_sg U39567 ( .A(n33799), .X(n33800) );
  inv_x1_sg U39568 ( .A(n30984), .X(n33801) );
  inv_x1_sg U39569 ( .A(n33799), .X(n33802) );
  inv_x1_sg U39570 ( .A(n35261), .X(n33803) );
  inv_x1_sg U39571 ( .A(n30981), .X(n33804) );
  inv_x1_sg U39572 ( .A(n33803), .X(n33805) );
  inv_x1_sg U39573 ( .A(n30981), .X(n33806) );
  inv_x1_sg U39574 ( .A(n33803), .X(n33807) );
  inv_x1_sg U39575 ( .A(n35260), .X(n33808) );
  inv_x1_sg U39576 ( .A(n30978), .X(n33809) );
  inv_x1_sg U39577 ( .A(n33808), .X(n33810) );
  inv_x1_sg U39578 ( .A(n30978), .X(n33811) );
  inv_x1_sg U39579 ( .A(n33808), .X(n33812) );
  inv_x1_sg U39580 ( .A(n35259), .X(n33813) );
  inv_x1_sg U39581 ( .A(n30975), .X(n33814) );
  inv_x1_sg U39582 ( .A(n33813), .X(n33815) );
  inv_x1_sg U39583 ( .A(n30975), .X(n33816) );
  inv_x1_sg U39584 ( .A(n33813), .X(n33817) );
  inv_x1_sg U39585 ( .A(n35594), .X(n33818) );
  inv_x1_sg U39586 ( .A(n33818), .X(n33819) );
  inv_x1_sg U39587 ( .A(n33818), .X(n33820) );
  inv_x1_sg U39588 ( .A(n30972), .X(n33821) );
  inv_x1_sg U39589 ( .A(n33818), .X(n33822) );
  inv_x1_sg U39590 ( .A(n34974), .X(n33823) );
  inv_x1_sg U39591 ( .A(n33823), .X(n33824) );
  inv_x1_sg U39592 ( .A(n33823), .X(n33825) );
  inv_x1_sg U39593 ( .A(n33823), .X(n33826) );
  inv_x1_sg U39594 ( .A(n33823), .X(n33827) );
  inv_x1_sg U39595 ( .A(n34805), .X(n33828) );
  inv_x1_sg U39596 ( .A(n34805), .X(n33829) );
  inv_x1_sg U39597 ( .A(n33829), .X(n33830) );
  inv_x1_sg U39598 ( .A(n30966), .X(n33831) );
  inv_x1_sg U39599 ( .A(n30966), .X(n33832) );
  inv_x1_sg U39600 ( .A(n30966), .X(n33833) );
  inv_x1_sg U39601 ( .A(n33830), .X(n33834) );
  inv_x1_sg U39602 ( .A(n30965), .X(n33835) );
  inv_x1_sg U39603 ( .A(n30962), .X(n33836) );
  inv_x1_sg U39604 ( .A(n30962), .X(n33837) );
  inv_x1_sg U39605 ( .A(n33835), .X(n33838) );
  inv_x1_sg U39606 ( .A(n33835), .X(n33839) );
  inv_x1_sg U39607 ( .A(n31108), .X(n33840) );
  inv_x1_sg U39608 ( .A(n31108), .X(n33841) );
  inv_x1_sg U39609 ( .A(n30634), .X(n33842) );
  inv_x1_sg U39610 ( .A(n30634), .X(n33843) );
  inv_x1_sg U39611 ( .A(n34865), .X(n33844) );
  inv_x1_sg U39612 ( .A(n30959), .X(n33845) );
  inv_x1_sg U39613 ( .A(n30959), .X(n33846) );
  inv_x1_sg U39614 ( .A(n30959), .X(n33847) );
  inv_x1_sg U39615 ( .A(n33844), .X(n33848) );
  inv_x1_sg U39616 ( .A(n30201), .X(n33849) );
  inv_x1_sg U39617 ( .A(n30955), .X(n33850) );
  inv_x1_sg U39618 ( .A(n30955), .X(n33851) );
  inv_x1_sg U39619 ( .A(n30955), .X(n33852) );
  inv_x1_sg U39620 ( .A(n33849), .X(n33853) );
  inv_x1_sg U39621 ( .A(n34863), .X(n33854) );
  inv_x1_sg U39622 ( .A(n30951), .X(n33855) );
  inv_x1_sg U39623 ( .A(n30951), .X(n33856) );
  inv_x1_sg U39624 ( .A(n30951), .X(n33857) );
  inv_x1_sg U39625 ( .A(n33854), .X(n33858) );
  inv_x1_sg U39626 ( .A(n35646), .X(n33859) );
  inv_x1_sg U39627 ( .A(n30948), .X(n33860) );
  inv_x1_sg U39628 ( .A(n33859), .X(n33861) );
  inv_x1_sg U39629 ( .A(n30948), .X(n33862) );
  inv_x1_sg U39630 ( .A(n33859), .X(n33863) );
  inv_x1_sg U39631 ( .A(n35640), .X(n33864) );
  inv_x1_sg U39632 ( .A(n30945), .X(n33865) );
  inv_x1_sg U39633 ( .A(n33864), .X(n33866) );
  inv_x1_sg U39634 ( .A(n30945), .X(n33867) );
  inv_x1_sg U39635 ( .A(n33864), .X(n33868) );
  inv_x1_sg U39636 ( .A(n35641), .X(n33869) );
  inv_x1_sg U39637 ( .A(n30942), .X(n33870) );
  inv_x1_sg U39638 ( .A(n33869), .X(n33871) );
  inv_x1_sg U39639 ( .A(n30942), .X(n33872) );
  inv_x1_sg U39640 ( .A(n33869), .X(n33873) );
  inv_x1_sg U39641 ( .A(n35647), .X(n33874) );
  inv_x1_sg U39642 ( .A(n30939), .X(n33875) );
  inv_x1_sg U39643 ( .A(n33874), .X(n33876) );
  inv_x1_sg U39644 ( .A(n30939), .X(n33877) );
  inv_x1_sg U39645 ( .A(n33874), .X(n33878) );
  nor_x1_sg U39646 ( .A(n31202), .B(n31201), .X(n33879) );
  inv_x1_sg U39647 ( .A(n33880), .X(n33881) );
  inv_x1_sg U39648 ( .A(n33880), .X(n33882) );
  inv_x1_sg U39649 ( .A(n33883), .X(n33884) );
  inv_x1_sg U39650 ( .A(n33883), .X(n33885) );
  inv_x1_sg U39651 ( .A(n33886), .X(n33887) );
  inv_x1_sg U39652 ( .A(n33886), .X(n33888) );
  inv_x1_sg U39653 ( .A(n30626), .X(n33889) );
  inv_x1_sg U39654 ( .A(n30626), .X(n33890) );
  inv_x1_sg U39655 ( .A(n34888), .X(n33891) );
  inv_x1_sg U39656 ( .A(n33891), .X(n33892) );
  inv_x1_sg U39657 ( .A(n30938), .X(n33893) );
  inv_x1_sg U39658 ( .A(n33891), .X(n33894) );
  inv_x1_sg U39659 ( .A(n33891), .X(n33895) );
  inv_x1_sg U39660 ( .A(n30628), .X(n33896) );
  inv_x1_sg U39661 ( .A(n30628), .X(n33897) );
  inv_x1_sg U39662 ( .A(n34884), .X(n33898) );
  inv_x1_sg U39663 ( .A(n33898), .X(n33899) );
  inv_x1_sg U39664 ( .A(n30936), .X(n33900) );
  inv_x1_sg U39665 ( .A(n33898), .X(n33901) );
  inv_x1_sg U39666 ( .A(n33898), .X(n33902) );
  inv_x1_sg U39667 ( .A(n30630), .X(n33903) );
  inv_x1_sg U39668 ( .A(n30630), .X(n33904) );
  inv_x1_sg U39669 ( .A(n34878), .X(n33905) );
  inv_x1_sg U39670 ( .A(n33905), .X(n33906) );
  inv_x1_sg U39671 ( .A(n30934), .X(n33907) );
  inv_x1_sg U39672 ( .A(n33905), .X(n33908) );
  inv_x1_sg U39673 ( .A(n33905), .X(n33909) );
  inv_x1_sg U39674 ( .A(n34879), .X(n33910) );
  inv_x1_sg U39675 ( .A(n33910), .X(n33911) );
  inv_x1_sg U39676 ( .A(n30932), .X(n33912) );
  inv_x1_sg U39677 ( .A(n33910), .X(n33913) );
  inv_x1_sg U39678 ( .A(n33910), .X(n33914) );
  inv_x1_sg U39679 ( .A(n30618), .X(n33915) );
  inv_x1_sg U39680 ( .A(n30600), .X(n33916) );
  inv_x1_sg U39681 ( .A(n34889), .X(n33917) );
  inv_x1_sg U39682 ( .A(n33917), .X(n33918) );
  inv_x1_sg U39683 ( .A(n33917), .X(n33919) );
  inv_x1_sg U39684 ( .A(n30930), .X(n33920) );
  inv_x1_sg U39685 ( .A(n33917), .X(n33921) );
  inv_x1_sg U39686 ( .A(n30625), .X(n33922) );
  inv_x1_sg U39687 ( .A(n33922), .X(n33923) );
  inv_x1_sg U39688 ( .A(n33922), .X(n33924) );
  inv_x1_sg U39689 ( .A(n30928), .X(n33925) );
  inv_x1_sg U39690 ( .A(n33922), .X(n33926) );
  inv_x1_sg U39691 ( .A(n34883), .X(n33927) );
  inv_x1_sg U39692 ( .A(n33927), .X(n33928) );
  inv_x1_sg U39693 ( .A(n33927), .X(n33929) );
  inv_x1_sg U39694 ( .A(n30926), .X(n33930) );
  inv_x1_sg U39695 ( .A(n33927), .X(n33931) );
  inv_x1_sg U39696 ( .A(n34885), .X(n33932) );
  inv_x1_sg U39697 ( .A(n33932), .X(n33933) );
  inv_x1_sg U39698 ( .A(n33932), .X(n33934) );
  inv_x1_sg U39699 ( .A(n30924), .X(n33935) );
  inv_x1_sg U39700 ( .A(n33932), .X(n33936) );
  inv_x1_sg U39701 ( .A(n34880), .X(n33937) );
  inv_x1_sg U39702 ( .A(n33937), .X(n33938) );
  inv_x1_sg U39703 ( .A(n33937), .X(n33939) );
  inv_x1_sg U39704 ( .A(n33937), .X(n33940) );
  inv_x1_sg U39705 ( .A(n30922), .X(n33941) );
  inv_x1_sg U39706 ( .A(n30637), .X(n33942) );
  inv_x1_sg U39707 ( .A(n30637), .X(n33943) );
  inv_x1_sg U39708 ( .A(n34851), .X(n33944) );
  inv_x1_sg U39709 ( .A(n33944), .X(n33945) );
  inv_x1_sg U39710 ( .A(n33944), .X(n33946) );
  inv_x1_sg U39711 ( .A(n33944), .X(n33947) );
  inv_x1_sg U39712 ( .A(n33944), .X(n33948) );
  inv_x1_sg U39713 ( .A(n34850), .X(n33949) );
  inv_x1_sg U39714 ( .A(n33949), .X(n33950) );
  inv_x1_sg U39715 ( .A(n33949), .X(n33951) );
  inv_x1_sg U39716 ( .A(n33949), .X(n33952) );
  inv_x1_sg U39717 ( .A(n33949), .X(n33953) );
  inv_x1_sg U39718 ( .A(n30913), .X(n33954) );
  inv_x1_sg U39719 ( .A(n35314), .X(n33955) );
  inv_x1_sg U39720 ( .A(n30913), .X(n33956) );
  inv_x1_sg U39721 ( .A(n30913), .X(n33957) );
  inv_x1_sg U39722 ( .A(n35274), .X(n33958) );
  inv_x1_sg U39723 ( .A(n33958), .X(n33959) );
  inv_x1_sg U39724 ( .A(n30912), .X(n33960) );
  inv_x1_sg U39725 ( .A(n33958), .X(n33961) );
  inv_x1_sg U39726 ( .A(n33958), .X(n33962) );
  inv_x1_sg U39727 ( .A(n26587), .X(n33963) );
  inv_x1_sg U39728 ( .A(n30911), .X(n33964) );
  inv_x1_sg U39729 ( .A(n30911), .X(n33965) );
  inv_x1_sg U39730 ( .A(n33963), .X(n33966) );
  inv_x1_sg U39731 ( .A(n34892), .X(n33967) );
  inv_x1_sg U39732 ( .A(n30624), .X(n33968) );
  inv_x1_sg U39733 ( .A(n34894), .X(n33969) );
  inv_x1_sg U39734 ( .A(n33969), .X(n33970) );
  inv_x1_sg U39735 ( .A(n33969), .X(n33971) );
  inv_x1_sg U39736 ( .A(n33969), .X(n33972) );
  inv_x1_sg U39737 ( .A(n34893), .X(n33973) );
  inv_x1_sg U39738 ( .A(n33973), .X(n33974) );
  inv_x1_sg U39739 ( .A(n33973), .X(n33975) );
  inv_x1_sg U39740 ( .A(n33973), .X(n33976) );
  inv_x1_sg U39741 ( .A(n33973), .X(n33977) );
  inv_x1_sg U39742 ( .A(n34895), .X(n33978) );
  inv_x1_sg U39743 ( .A(n33978), .X(n33979) );
  inv_x1_sg U39744 ( .A(n33978), .X(n33980) );
  inv_x1_sg U39745 ( .A(n33978), .X(n33981) );
  inv_x1_sg U39746 ( .A(n33978), .X(n33982) );
  inv_x1_sg U39747 ( .A(n19590), .X(n33983) );
  inv_x1_sg U39748 ( .A(n33983), .X(n33984) );
  inv_x1_sg U39749 ( .A(n33983), .X(n33985) );
  inv_x1_sg U39750 ( .A(n30910), .X(n33986) );
  inv_x1_sg U39751 ( .A(n30910), .X(n33987) );
  inv_x1_sg U39752 ( .A(n35414), .X(n33988) );
  inv_x1_sg U39753 ( .A(n31047), .X(n33989) );
  inv_x1_sg U39754 ( .A(n33988), .X(n33990) );
  inv_x1_sg U39755 ( .A(n31047), .X(n33991) );
  inv_x1_sg U39756 ( .A(n35413), .X(n33992) );
  inv_x1_sg U39757 ( .A(n31050), .X(n33993) );
  inv_x1_sg U39758 ( .A(n33992), .X(n33994) );
  inv_x1_sg U39759 ( .A(n31050), .X(n33995) );
  inv_x1_sg U39760 ( .A(n35387), .X(n33996) );
  inv_x1_sg U39761 ( .A(n35364), .X(n33997) );
  inv_x1_sg U39762 ( .A(n35090), .X(n33998) );
  inv_x1_sg U39763 ( .A(n30907), .X(n33999) );
  inv_x1_sg U39764 ( .A(n33998), .X(n34000) );
  inv_x1_sg U39765 ( .A(n30907), .X(n34001) );
  inv_x1_sg U39766 ( .A(n33998), .X(n34002) );
  inv_x1_sg U39767 ( .A(n34660), .X(n34003) );
  inv_x1_sg U39768 ( .A(n30900), .X(n34004) );
  inv_x1_sg U39769 ( .A(n30900), .X(n34005) );
  inv_x1_sg U39770 ( .A(n34003), .X(n34006) );
  inv_x1_sg U39771 ( .A(n34003), .X(n34007) );
  inv_x1_sg U39772 ( .A(n31241), .X(n34008) );
  inv_x1_sg U39773 ( .A(n31241), .X(n34009) );
  inv_x1_sg U39774 ( .A(n34913), .X(n34010) );
  inv_x1_sg U39775 ( .A(n31062), .X(n34011) );
  inv_x1_sg U39776 ( .A(n31063), .X(n34012) );
  inv_x1_sg U39777 ( .A(n31063), .X(n34013) );
  inv_x1_sg U39778 ( .A(n31062), .X(n34014) );
  inv_x1_sg U39779 ( .A(n34912), .X(n34015) );
  inv_x1_sg U39780 ( .A(n31067), .X(n34016) );
  inv_x1_sg U39781 ( .A(n31068), .X(n34017) );
  inv_x1_sg U39782 ( .A(n31068), .X(n34018) );
  inv_x1_sg U39783 ( .A(n31067), .X(n34019) );
  inv_x1_sg U39784 ( .A(n34911), .X(n34020) );
  inv_x1_sg U39785 ( .A(n31073), .X(n34021) );
  inv_x1_sg U39786 ( .A(n31072), .X(n34022) );
  inv_x1_sg U39787 ( .A(n31073), .X(n34023) );
  inv_x1_sg U39788 ( .A(n31072), .X(n34024) );
  inv_x1_sg U39789 ( .A(n31246), .X(n34025) );
  inv_x1_sg U39790 ( .A(n31245), .X(n34026) );
  inv_x1_sg U39791 ( .A(n34908), .X(n34027) );
  inv_x1_sg U39792 ( .A(n31078), .X(n34028) );
  inv_x1_sg U39793 ( .A(n31077), .X(n34029) );
  inv_x1_sg U39794 ( .A(n31078), .X(n34030) );
  inv_x1_sg U39795 ( .A(n31077), .X(n34031) );
  inv_x1_sg U39796 ( .A(n34907), .X(n34032) );
  inv_x1_sg U39797 ( .A(n31083), .X(n34033) );
  inv_x1_sg U39798 ( .A(n31082), .X(n34034) );
  inv_x1_sg U39799 ( .A(n31083), .X(n34035) );
  inv_x1_sg U39800 ( .A(n31082), .X(n34036) );
  inv_x1_sg U39801 ( .A(n34906), .X(n34037) );
  inv_x1_sg U39802 ( .A(n31088), .X(n34038) );
  inv_x1_sg U39803 ( .A(n31087), .X(n34039) );
  inv_x1_sg U39804 ( .A(n31088), .X(n34040) );
  inv_x1_sg U39805 ( .A(n31087), .X(n34041) );
  inv_x1_sg U39806 ( .A(n35319), .X(n34042) );
  inv_x1_sg U39807 ( .A(n35375), .X(n34043) );
  inv_x1_sg U39808 ( .A(n30180), .X(n34044) );
  inv_x1_sg U39809 ( .A(n30893), .X(n34045) );
  inv_x1_sg U39810 ( .A(n34044), .X(n34046) );
  inv_x1_sg U39811 ( .A(n34044), .X(n34047) );
  inv_x1_sg U39812 ( .A(n34044), .X(n34048) );
  inv_x1_sg U39813 ( .A(n34659), .X(n34049) );
  inv_x1_sg U39814 ( .A(n34049), .X(n34050) );
  inv_x1_sg U39815 ( .A(n34049), .X(n34051) );
  inv_x1_sg U39816 ( .A(n34049), .X(n34052) );
  inv_x1_sg U39817 ( .A(n34049), .X(n34053) );
  inv_x1_sg U39818 ( .A(n30587), .X(n34054) );
  inv_x1_sg U39819 ( .A(n34054), .X(n34055) );
  inv_x1_sg U39820 ( .A(n34054), .X(n34056) );
  inv_x1_sg U39821 ( .A(n34054), .X(n34057) );
  inv_x1_sg U39822 ( .A(n34054), .X(n34058) );
  inv_x1_sg U39823 ( .A(n28318), .X(n34059) );
  inv_x1_sg U39824 ( .A(n28318), .X(n34060) );
  inv_x1_sg U39825 ( .A(n28318), .X(n34061) );
  inv_x1_sg U39826 ( .A(n34059), .X(n34062) );
  inv_x1_sg U39827 ( .A(n34059), .X(n34063) );
  inv_x1_sg U39828 ( .A(n34060), .X(n34064) );
  inv_x1_sg U39829 ( .A(n34060), .X(n34065) );
  inv_x1_sg U39830 ( .A(n34060), .X(n34066) );
  inv_x1_sg U39831 ( .A(n34060), .X(n34067) );
  inv_x1_sg U39832 ( .A(n34061), .X(n34068) );
  inv_x1_sg U39833 ( .A(n34061), .X(n34069) );
  inv_x1_sg U39834 ( .A(n34061), .X(n34070) );
  inv_x1_sg U39835 ( .A(n34655), .X(n34071) );
  inv_x1_sg U39836 ( .A(n30723), .X(n34072) );
  inv_x1_sg U39837 ( .A(n34071), .X(n34073) );
  inv_x1_sg U39838 ( .A(n34071), .X(n34074) );
  inv_x1_sg U39839 ( .A(n31095), .X(n34075) );
  inv_x1_sg U39840 ( .A(n34075), .X(n34076) );
  inv_x1_sg U39841 ( .A(n30719), .X(n34077) );
  inv_x1_sg U39842 ( .A(n34075), .X(n34078) );
  inv_x1_sg U39843 ( .A(n35084), .X(n34079) );
  inv_x1_sg U39844 ( .A(n34079), .X(n34080) );
  inv_x1_sg U39845 ( .A(n30704), .X(n34081) );
  inv_x1_sg U39846 ( .A(n34079), .X(n34082) );
  inv_x1_sg U39847 ( .A(n35178), .X(n34083) );
  inv_x1_sg U39848 ( .A(n35385), .X(n34084) );
  inv_x1_sg U39849 ( .A(n13221), .X(n34085) );
  inv_x1_sg U39850 ( .A(n34085), .X(n34086) );
  inv_x1_sg U39851 ( .A(n34085), .X(n34087) );
  inv_x1_sg U39852 ( .A(n31493), .X(n34088) );
  inv_x1_sg U39853 ( .A(n31493), .X(n34089) );
  inv_x1_sg U39854 ( .A(n35089), .X(n34090) );
  inv_x1_sg U39855 ( .A(n34090), .X(n34091) );
  inv_x1_sg U39856 ( .A(n34090), .X(n34092) );
  inv_x1_sg U39857 ( .A(n35085), .X(n34093) );
  inv_x1_sg U39858 ( .A(n30860), .X(n34094) );
  inv_x1_sg U39859 ( .A(n30860), .X(n34095) );
  inv_x1_sg U39860 ( .A(n34093), .X(n34096) );
  inv_x1_sg U39861 ( .A(n34093), .X(n34097) );
  inv_x1_sg U39862 ( .A(n34963), .X(n34098) );
  inv_x1_sg U39863 ( .A(n34963), .X(n34099) );
  inv_x1_sg U39864 ( .A(n34725), .X(n34100) );
  inv_x1_sg U39865 ( .A(n31483), .X(n34101) );
  inv_x1_sg U39866 ( .A(n30042), .X(n34102) );
  inv_x1_sg U39867 ( .A(n31234), .X(n34103) );
  inv_x1_sg U39868 ( .A(n31483), .X(n34104) );
  inv_x1_sg U39869 ( .A(n31479), .X(n34105) );
  inv_x1_sg U39870 ( .A(n31478), .X(n34106) );
  inv_x1_sg U39871 ( .A(n31233), .X(n34107) );
  inv_x1_sg U39872 ( .A(n30182), .X(n34108) );
  inv_x1_sg U39873 ( .A(n29672), .X(n34109) );
  inv_x1_sg U39874 ( .A(n31473), .X(n34110) );
  inv_x1_sg U39875 ( .A(n31473), .X(n34111) );
  inv_x1_sg U39876 ( .A(n35600), .X(n34112) );
  inv_x1_sg U39877 ( .A(n31469), .X(n34113) );
  inv_x1_sg U39878 ( .A(n31469), .X(n34114) );
  inv_x1_sg U39879 ( .A(n30047), .X(n34115) );
  inv_x1_sg U39880 ( .A(n11737), .X(n34116) );
  inv_x1_sg U39881 ( .A(n31466), .X(n34117) );
  inv_x1_sg U39882 ( .A(n31466), .X(n34118) );
  inv_x1_sg U39883 ( .A(n30050), .X(n34119) );
  inv_x1_sg U39884 ( .A(n11791), .X(n34120) );
  inv_x1_sg U39885 ( .A(n31463), .X(n34121) );
  inv_x1_sg U39886 ( .A(n31463), .X(n34122) );
  inv_x1_sg U39887 ( .A(n30053), .X(n34123) );
  inv_x1_sg U39888 ( .A(n11710), .X(n34124) );
  inv_x1_sg U39889 ( .A(n31460), .X(n34125) );
  inv_x1_sg U39890 ( .A(n31460), .X(n34126) );
  inv_x1_sg U39891 ( .A(n30056), .X(n34127) );
  inv_x1_sg U39892 ( .A(n15171), .X(n34128) );
  inv_x1_sg U39893 ( .A(n34128), .X(n34129) );
  inv_x1_sg U39894 ( .A(n31457), .X(n34130) );
  inv_x1_sg U39895 ( .A(n31457), .X(n34131) );
  inv_x1_sg U39896 ( .A(n34128), .X(n34132) );
  inv_x1_sg U39897 ( .A(n15181), .X(n34133) );
  inv_x1_sg U39898 ( .A(n34133), .X(n34134) );
  inv_x1_sg U39899 ( .A(n30258), .X(n34135) );
  inv_x1_sg U39900 ( .A(n30258), .X(n34136) );
  inv_x1_sg U39901 ( .A(n34133), .X(n34137) );
  inv_x1_sg U39902 ( .A(n15180), .X(n34138) );
  inv_x1_sg U39903 ( .A(n34138), .X(n34139) );
  inv_x1_sg U39904 ( .A(n30260), .X(n34140) );
  inv_x1_sg U39905 ( .A(n30260), .X(n34141) );
  inv_x1_sg U39906 ( .A(n34138), .X(n34142) );
  inv_x1_sg U39907 ( .A(n15177), .X(n34143) );
  inv_x1_sg U39908 ( .A(n34143), .X(n34144) );
  inv_x1_sg U39909 ( .A(n30262), .X(n34145) );
  inv_x1_sg U39910 ( .A(n30262), .X(n34146) );
  inv_x1_sg U39911 ( .A(n34143), .X(n34147) );
  inv_x1_sg U39912 ( .A(n15048), .X(n34148) );
  inv_x1_sg U39913 ( .A(n34148), .X(n34149) );
  inv_x1_sg U39914 ( .A(n30264), .X(n34150) );
  inv_x1_sg U39915 ( .A(n30264), .X(n34151) );
  inv_x1_sg U39916 ( .A(n34148), .X(n34152) );
  inv_x1_sg U39917 ( .A(n15044), .X(n34153) );
  inv_x1_sg U39918 ( .A(n34153), .X(n34154) );
  inv_x1_sg U39919 ( .A(n30266), .X(n34155) );
  inv_x1_sg U39920 ( .A(n30266), .X(n34156) );
  inv_x1_sg U39921 ( .A(n34153), .X(n34157) );
  inv_x1_sg U39922 ( .A(n15190), .X(n34158) );
  inv_x1_sg U39923 ( .A(n34158), .X(n34159) );
  inv_x1_sg U39924 ( .A(n30268), .X(n34160) );
  inv_x1_sg U39925 ( .A(n30268), .X(n34161) );
  inv_x1_sg U39926 ( .A(n34158), .X(n34162) );
  inv_x1_sg U39927 ( .A(n15182), .X(n34163) );
  inv_x1_sg U39928 ( .A(n34163), .X(n34164) );
  inv_x1_sg U39929 ( .A(n30270), .X(n34165) );
  inv_x1_sg U39930 ( .A(n30270), .X(n34166) );
  inv_x1_sg U39931 ( .A(n34163), .X(n34167) );
  inv_x1_sg U39932 ( .A(n15055), .X(n34168) );
  inv_x1_sg U39933 ( .A(n34168), .X(n34169) );
  inv_x1_sg U39934 ( .A(n30272), .X(n34170) );
  inv_x1_sg U39935 ( .A(n30272), .X(n34171) );
  inv_x1_sg U39936 ( .A(n34168), .X(n34172) );
  inv_x1_sg U39937 ( .A(n15049), .X(n34173) );
  inv_x1_sg U39938 ( .A(n34173), .X(n34174) );
  inv_x1_sg U39939 ( .A(n30274), .X(n34175) );
  inv_x1_sg U39940 ( .A(n30274), .X(n34176) );
  inv_x1_sg U39941 ( .A(n34173), .X(n34177) );
  inv_x1_sg U39942 ( .A(n15172), .X(n34178) );
  inv_x1_sg U39943 ( .A(n34178), .X(n34179) );
  inv_x1_sg U39944 ( .A(n30276), .X(n34180) );
  inv_x1_sg U39945 ( .A(n30276), .X(n34181) );
  inv_x1_sg U39946 ( .A(n34178), .X(n34182) );
  inv_x1_sg U39947 ( .A(n15170), .X(n34183) );
  inv_x1_sg U39948 ( .A(n34183), .X(n34184) );
  inv_x1_sg U39949 ( .A(n30278), .X(n34185) );
  inv_x1_sg U39950 ( .A(n30278), .X(n34186) );
  inv_x1_sg U39951 ( .A(n34183), .X(n34187) );
  inv_x1_sg U39952 ( .A(n15039), .X(n34188) );
  inv_x1_sg U39953 ( .A(n34188), .X(n34189) );
  inv_x1_sg U39954 ( .A(n30280), .X(n34190) );
  inv_x1_sg U39955 ( .A(n30280), .X(n34191) );
  inv_x1_sg U39956 ( .A(n34188), .X(n34192) );
  inv_x1_sg U39957 ( .A(n15038), .X(n34193) );
  inv_x1_sg U39958 ( .A(n34193), .X(n34194) );
  inv_x1_sg U39959 ( .A(n30282), .X(n34195) );
  inv_x1_sg U39960 ( .A(n30282), .X(n34196) );
  inv_x1_sg U39961 ( .A(n34193), .X(n34197) );
  inv_x1_sg U39962 ( .A(n15037), .X(n34198) );
  inv_x1_sg U39963 ( .A(n34198), .X(n34199) );
  inv_x1_sg U39964 ( .A(n30284), .X(n34200) );
  inv_x1_sg U39965 ( .A(n30284), .X(n34201) );
  inv_x1_sg U39966 ( .A(n34198), .X(n34202) );
  inv_x1_sg U39967 ( .A(n13808), .X(n34203) );
  inv_x1_sg U39968 ( .A(n34203), .X(n34204) );
  inv_x1_sg U39969 ( .A(n30286), .X(n34205) );
  inv_x1_sg U39970 ( .A(n30286), .X(n34206) );
  inv_x1_sg U39971 ( .A(n34203), .X(n34207) );
  inv_x1_sg U39972 ( .A(n35644), .X(n34208) );
  inv_x1_sg U39973 ( .A(n34208), .X(n34209) );
  inv_x1_sg U39974 ( .A(n30289), .X(n34210) );
  inv_x1_sg U39975 ( .A(n30289), .X(n34211) );
  inv_x1_sg U39976 ( .A(n34208), .X(n34212) );
  inv_x1_sg U39977 ( .A(n35645), .X(n34213) );
  inv_x1_sg U39978 ( .A(n34213), .X(n34214) );
  inv_x1_sg U39979 ( .A(n30291), .X(n34215) );
  inv_x1_sg U39980 ( .A(n30291), .X(n34216) );
  inv_x1_sg U39981 ( .A(n34213), .X(n34217) );
  inv_x1_sg U39982 ( .A(n13787), .X(n34218) );
  inv_x1_sg U39983 ( .A(n34218), .X(n34219) );
  inv_x1_sg U39984 ( .A(n30293), .X(n34220) );
  inv_x1_sg U39985 ( .A(n30293), .X(n34221) );
  inv_x1_sg U39986 ( .A(n34218), .X(n34222) );
  inv_x1_sg U39987 ( .A(n12531), .X(n34223) );
  inv_x1_sg U39988 ( .A(n34223), .X(n34224) );
  inv_x1_sg U39989 ( .A(n30296), .X(n34225) );
  inv_x1_sg U39990 ( .A(n30296), .X(n34226) );
  inv_x1_sg U39991 ( .A(n34223), .X(n34227) );
  inv_x1_sg U39992 ( .A(n35633), .X(n34228) );
  inv_x1_sg U39993 ( .A(n34228), .X(n34229) );
  inv_x1_sg U39994 ( .A(n30299), .X(n34230) );
  inv_x1_sg U39995 ( .A(n30299), .X(n34231) );
  inv_x1_sg U39996 ( .A(n34228), .X(n34232) );
  inv_x1_sg U39997 ( .A(n12533), .X(n34233) );
  inv_x1_sg U39998 ( .A(n34233), .X(n34234) );
  inv_x1_sg U39999 ( .A(n30301), .X(n34235) );
  inv_x1_sg U40000 ( .A(n30301), .X(n34236) );
  inv_x1_sg U40001 ( .A(n34233), .X(n34237) );
  inv_x1_sg U40002 ( .A(n35629), .X(n34238) );
  inv_x1_sg U40003 ( .A(n34238), .X(n34239) );
  inv_x1_sg U40004 ( .A(n30303), .X(n34240) );
  inv_x1_sg U40005 ( .A(n30303), .X(n34241) );
  inv_x1_sg U40006 ( .A(n34238), .X(n34242) );
  inv_x1_sg U40007 ( .A(n35630), .X(n34243) );
  inv_x1_sg U40008 ( .A(n34243), .X(n34244) );
  inv_x1_sg U40009 ( .A(n30305), .X(n34245) );
  inv_x1_sg U40010 ( .A(n30305), .X(n34246) );
  inv_x1_sg U40011 ( .A(n34243), .X(n34247) );
  inv_x1_sg U40012 ( .A(n35632), .X(n34248) );
  inv_x1_sg U40013 ( .A(n34248), .X(n34249) );
  inv_x1_sg U40014 ( .A(n30307), .X(n34250) );
  inv_x1_sg U40015 ( .A(n30307), .X(n34251) );
  inv_x1_sg U40016 ( .A(n34248), .X(n34252) );
  inv_x1_sg U40017 ( .A(n35650), .X(n34253) );
  inv_x1_sg U40018 ( .A(n34253), .X(n34254) );
  inv_x1_sg U40019 ( .A(n30309), .X(n34255) );
  inv_x1_sg U40020 ( .A(n30309), .X(n34256) );
  inv_x1_sg U40021 ( .A(n34253), .X(n34257) );
  inv_x1_sg U40022 ( .A(n13816), .X(n34258) );
  inv_x1_sg U40023 ( .A(n34258), .X(n34259) );
  inv_x1_sg U40024 ( .A(n30312), .X(n34260) );
  inv_x1_sg U40025 ( .A(n30312), .X(n34261) );
  inv_x1_sg U40026 ( .A(n34258), .X(n34262) );
  inv_x1_sg U40027 ( .A(n13805), .X(n34263) );
  inv_x1_sg U40028 ( .A(n34263), .X(n34264) );
  inv_x1_sg U40029 ( .A(n30315), .X(n34265) );
  inv_x1_sg U40030 ( .A(n30315), .X(n34266) );
  inv_x1_sg U40031 ( .A(n34263), .X(n34267) );
  inv_x1_sg U40032 ( .A(n13804), .X(n34268) );
  inv_x1_sg U40033 ( .A(n34268), .X(n34269) );
  inv_x1_sg U40034 ( .A(n30318), .X(n34270) );
  inv_x1_sg U40035 ( .A(n30318), .X(n34271) );
  inv_x1_sg U40036 ( .A(n34268), .X(n34272) );
  inv_x1_sg U40037 ( .A(n13367), .X(n34273) );
  inv_x1_sg U40038 ( .A(n34273), .X(n34274) );
  inv_x1_sg U40039 ( .A(n30321), .X(n34275) );
  inv_x1_sg U40040 ( .A(n30321), .X(n34276) );
  inv_x1_sg U40041 ( .A(n34273), .X(n34277) );
  inv_x1_sg U40042 ( .A(n11667), .X(n34278) );
  inv_x1_sg U40043 ( .A(n34278), .X(n34279) );
  inv_x1_sg U40044 ( .A(n30323), .X(n34280) );
  inv_x1_sg U40045 ( .A(n30323), .X(n34281) );
  inv_x1_sg U40046 ( .A(n34278), .X(n34282) );
  inv_x1_sg U40047 ( .A(n11535), .X(n34283) );
  inv_x1_sg U40048 ( .A(n34283), .X(n34284) );
  inv_x1_sg U40049 ( .A(n30325), .X(n34285) );
  inv_x1_sg U40050 ( .A(n30325), .X(n34286) );
  inv_x1_sg U40051 ( .A(n34283), .X(n34287) );
  inv_x1_sg U40052 ( .A(n15184), .X(n34288) );
  inv_x1_sg U40053 ( .A(n34288), .X(n34289) );
  inv_x1_sg U40054 ( .A(n30327), .X(n34290) );
  inv_x1_sg U40055 ( .A(n30327), .X(n34291) );
  inv_x1_sg U40056 ( .A(n34288), .X(n34292) );
  inv_x1_sg U40057 ( .A(n15179), .X(n34293) );
  inv_x1_sg U40058 ( .A(n34293), .X(n34294) );
  inv_x1_sg U40059 ( .A(n30329), .X(n34295) );
  inv_x1_sg U40060 ( .A(n30329), .X(n34296) );
  inv_x1_sg U40061 ( .A(n34293), .X(n34297) );
  inv_x1_sg U40062 ( .A(n15050), .X(n34298) );
  inv_x1_sg U40063 ( .A(n34298), .X(n34299) );
  inv_x1_sg U40064 ( .A(n30331), .X(n34300) );
  inv_x1_sg U40065 ( .A(n30331), .X(n34301) );
  inv_x1_sg U40066 ( .A(n34298), .X(n34302) );
  inv_x1_sg U40067 ( .A(n15046), .X(n34303) );
  inv_x1_sg U40068 ( .A(n34303), .X(n34304) );
  inv_x1_sg U40069 ( .A(n30333), .X(n34305) );
  inv_x1_sg U40070 ( .A(n30333), .X(n34306) );
  inv_x1_sg U40071 ( .A(n34303), .X(n34307) );
  inv_x1_sg U40072 ( .A(n35599), .X(n34308) );
  inv_x1_sg U40073 ( .A(n34308), .X(n34309) );
  inv_x1_sg U40074 ( .A(n30335), .X(n34310) );
  inv_x1_sg U40075 ( .A(n30335), .X(n34311) );
  inv_x1_sg U40076 ( .A(n34308), .X(n34312) );
  inv_x1_sg U40077 ( .A(n35598), .X(n34313) );
  inv_x1_sg U40078 ( .A(n34313), .X(n34314) );
  inv_x1_sg U40079 ( .A(n30337), .X(n34315) );
  inv_x1_sg U40080 ( .A(n30337), .X(n34316) );
  inv_x1_sg U40081 ( .A(n34313), .X(n34317) );
  inv_x1_sg U40082 ( .A(n35597), .X(n34318) );
  inv_x1_sg U40083 ( .A(n34318), .X(n34319) );
  inv_x1_sg U40084 ( .A(n30339), .X(n34320) );
  inv_x1_sg U40085 ( .A(n30339), .X(n34321) );
  inv_x1_sg U40086 ( .A(n34318), .X(n34322) );
  inv_x1_sg U40087 ( .A(n35596), .X(n34323) );
  inv_x1_sg U40088 ( .A(n34323), .X(n34324) );
  inv_x1_sg U40089 ( .A(n30341), .X(n34325) );
  inv_x1_sg U40090 ( .A(n30341), .X(n34326) );
  inv_x1_sg U40091 ( .A(n34323), .X(n34327) );
  inv_x1_sg U40092 ( .A(n35595), .X(n34328) );
  inv_x1_sg U40093 ( .A(n34328), .X(n34329) );
  inv_x1_sg U40094 ( .A(n30343), .X(n34330) );
  inv_x1_sg U40095 ( .A(n30343), .X(n34331) );
  inv_x1_sg U40096 ( .A(n34328), .X(n34332) );
  inv_x1_sg U40097 ( .A(n15047), .X(n34333) );
  inv_x1_sg U40098 ( .A(n34333), .X(n34334) );
  inv_x1_sg U40099 ( .A(n30345), .X(n34335) );
  inv_x1_sg U40100 ( .A(n30345), .X(n34336) );
  inv_x1_sg U40101 ( .A(n34333), .X(n34337) );
  inv_x1_sg U40102 ( .A(n15187), .X(n34338) );
  inv_x1_sg U40103 ( .A(n34338), .X(n34339) );
  inv_x1_sg U40104 ( .A(n30347), .X(n34340) );
  inv_x1_sg U40105 ( .A(n30347), .X(n34341) );
  inv_x1_sg U40106 ( .A(n34338), .X(n34342) );
  inv_x1_sg U40107 ( .A(n13368), .X(n34343) );
  inv_x1_sg U40108 ( .A(n34343), .X(n34344) );
  inv_x1_sg U40109 ( .A(n30349), .X(n34345) );
  inv_x1_sg U40110 ( .A(n30349), .X(n34346) );
  inv_x1_sg U40111 ( .A(n34343), .X(n34347) );
  inv_x1_sg U40112 ( .A(n35631), .X(n34348) );
  inv_x1_sg U40113 ( .A(n34348), .X(n34349) );
  inv_x1_sg U40114 ( .A(n30351), .X(n34350) );
  inv_x1_sg U40115 ( .A(n30351), .X(n34351) );
  inv_x1_sg U40116 ( .A(n34348), .X(n34352) );
  inv_x1_sg U40117 ( .A(n11562), .X(n34353) );
  inv_x1_sg U40118 ( .A(n34353), .X(n34354) );
  inv_x1_sg U40119 ( .A(n30353), .X(n34355) );
  inv_x1_sg U40120 ( .A(n30353), .X(n34356) );
  inv_x1_sg U40121 ( .A(n34353), .X(n34357) );
  inv_x1_sg U40122 ( .A(n11586), .X(n34358) );
  inv_x1_sg U40123 ( .A(n34358), .X(n34359) );
  inv_x1_sg U40124 ( .A(n30355), .X(n34360) );
  inv_x1_sg U40125 ( .A(n30355), .X(n34361) );
  inv_x1_sg U40126 ( .A(n34358), .X(n34362) );
  inv_x1_sg U40127 ( .A(n11536), .X(n34363) );
  inv_x1_sg U40128 ( .A(n34363), .X(n34364) );
  inv_x1_sg U40129 ( .A(n30357), .X(n34365) );
  inv_x1_sg U40130 ( .A(n30357), .X(n34366) );
  inv_x1_sg U40131 ( .A(n34363), .X(n34367) );
  inv_x1_sg U40132 ( .A(n11641), .X(n34368) );
  inv_x1_sg U40133 ( .A(n34368), .X(n34369) );
  inv_x1_sg U40134 ( .A(n30359), .X(n34370) );
  inv_x1_sg U40135 ( .A(n30359), .X(n34371) );
  inv_x1_sg U40136 ( .A(n34368), .X(n34372) );
  inv_x1_sg U40137 ( .A(n35458), .X(n34373) );
  inv_x1_sg U40138 ( .A(n34373), .X(n34374) );
  inv_x1_sg U40139 ( .A(n30361), .X(n34375) );
  inv_x1_sg U40140 ( .A(n30361), .X(n34376) );
  inv_x1_sg U40141 ( .A(n34373), .X(n34377) );
  inv_x1_sg U40142 ( .A(n35483), .X(n34378) );
  inv_x1_sg U40143 ( .A(n34378), .X(n34379) );
  inv_x1_sg U40144 ( .A(n30363), .X(n34380) );
  inv_x1_sg U40145 ( .A(n30363), .X(n34381) );
  inv_x1_sg U40146 ( .A(n34378), .X(n34382) );
  inv_x1_sg U40147 ( .A(n15053), .X(n34383) );
  inv_x1_sg U40148 ( .A(n34383), .X(n34384) );
  inv_x1_sg U40149 ( .A(n30365), .X(n34385) );
  inv_x1_sg U40150 ( .A(n30365), .X(n34386) );
  inv_x1_sg U40151 ( .A(n34383), .X(n34387) );
  nor_x1_sg U40152 ( .A(n35454), .B(n35459), .X(n34388) );
  nor_x1_sg U40153 ( .A(n35454), .B(n35628), .X(n34389) );
  inv_x1_sg U40154 ( .A(n34388), .X(n34390) );
  inv_x1_sg U40155 ( .A(n34390), .X(n34391) );
  inv_x1_sg U40156 ( .A(n34390), .X(n34392) );
  inv_x1_sg U40157 ( .A(n34390), .X(n34393) );
  inv_x1_sg U40158 ( .A(n34390), .X(n34394) );
  inv_x1_sg U40159 ( .A(n34389), .X(n34395) );
  inv_x1_sg U40160 ( .A(n33880), .X(n34396) );
  inv_x1_sg U40161 ( .A(n34395), .X(n34397) );
  inv_x1_sg U40162 ( .A(n34395), .X(n34398) );
  inv_x1_sg U40163 ( .A(n34395), .X(n34399) );
  inv_x1_sg U40164 ( .A(n33886), .X(n34400) );
  inv_x1_sg U40165 ( .A(n33883), .X(n34401) );
  inv_x1_sg U40166 ( .A(n12717), .X(n34402) );
  inv_x1_sg U40167 ( .A(n30858), .X(n34403) );
  inv_x1_sg U40168 ( .A(n34402), .X(n34404) );
  inv_x1_sg U40169 ( .A(n30858), .X(n34405) );
  inv_x1_sg U40170 ( .A(n34402), .X(n34406) );
  inv_x1_sg U40171 ( .A(n19591), .X(n34407) );
  inv_x1_sg U40172 ( .A(n34407), .X(n34408) );
  inv_x1_sg U40173 ( .A(n30856), .X(n34409) );
  inv_x1_sg U40174 ( .A(n34407), .X(n34410) );
  inv_x1_sg U40175 ( .A(n30856), .X(n34411) );
  inv_x1_sg U40176 ( .A(n34100), .X(n34412) );
  inv_x1_sg U40177 ( .A(n30181), .X(n34413) );
  inv_x1_sg U40178 ( .A(n34100), .X(n34414) );
  inv_x1_sg U40179 ( .A(n34107), .X(n34415) );
  inv_x1_sg U40180 ( .A(n35634), .X(n34416) );
  inv_x1_sg U40181 ( .A(n30852), .X(n34417) );
  inv_x1_sg U40182 ( .A(n30849), .X(n34418) );
  inv_x1_sg U40183 ( .A(n30852), .X(n34419) );
  inv_x1_sg U40184 ( .A(n34416), .X(n34420) );
  inv_x1_sg U40185 ( .A(n11611), .X(n34421) );
  inv_x1_sg U40186 ( .A(n30848), .X(n34422) );
  inv_x1_sg U40187 ( .A(n34421), .X(n34423) );
  inv_x1_sg U40188 ( .A(n30848), .X(n34424) );
  inv_x1_sg U40189 ( .A(n34421), .X(n34425) );
  inv_x1_sg U40190 ( .A(n13619), .X(n34426) );
  inv_x1_sg U40191 ( .A(n30846), .X(n34427) );
  inv_x1_sg U40192 ( .A(n34426), .X(n34428) );
  inv_x1_sg U40193 ( .A(n30846), .X(n34429) );
  inv_x1_sg U40194 ( .A(n34426), .X(n34430) );
  inv_x1_sg U40195 ( .A(n35657), .X(n34431) );
  inv_x1_sg U40196 ( .A(n34431), .X(n34432) );
  inv_x1_sg U40197 ( .A(n30842), .X(n34433) );
  inv_x1_sg U40198 ( .A(n34431), .X(n34434) );
  inv_x1_sg U40199 ( .A(n30842), .X(n34435) );
  inv_x1_sg U40200 ( .A(n19582), .X(n34436) );
  inv_x1_sg U40201 ( .A(n34436), .X(n34437) );
  inv_x1_sg U40202 ( .A(n30841), .X(n34438) );
  inv_x1_sg U40203 ( .A(n34436), .X(n34439) );
  inv_x1_sg U40204 ( .A(n30841), .X(n34440) );
  inv_x1_sg U40205 ( .A(n11561), .X(n34441) );
  inv_x1_sg U40206 ( .A(n34441), .X(n34442) );
  inv_x1_sg U40207 ( .A(n30836), .X(n34443) );
  inv_x1_sg U40208 ( .A(n34441), .X(n34444) );
  inv_x1_sg U40209 ( .A(n30836), .X(n34445) );
  inv_x1_sg U40210 ( .A(n35653), .X(n34446) );
  inv_x1_sg U40211 ( .A(n34446), .X(n34447) );
  inv_x1_sg U40212 ( .A(n30833), .X(n34448) );
  inv_x1_sg U40213 ( .A(n34446), .X(n34449) );
  inv_x1_sg U40214 ( .A(n30833), .X(n34450) );
  inv_x1_sg U40215 ( .A(n31098), .X(n34451) );
  inv_x1_sg U40216 ( .A(n31611), .X(n34452) );
  inv_x1_sg U40217 ( .A(n34934), .X(n34453) );
  inv_x1_sg U40218 ( .A(n34453), .X(n34454) );
  inv_x1_sg U40219 ( .A(n30831), .X(n34455) );
  inv_x1_sg U40220 ( .A(n29902), .X(n34456) );
  inv_x1_sg U40221 ( .A(n34453), .X(n34457) );
  inv_x1_sg U40222 ( .A(n34932), .X(n34458) );
  inv_x1_sg U40223 ( .A(n34458), .X(n34459) );
  inv_x1_sg U40224 ( .A(n30827), .X(n34460) );
  inv_x1_sg U40225 ( .A(n30118), .X(n34461) );
  inv_x1_sg U40226 ( .A(n34458), .X(n34462) );
  inv_x1_sg U40227 ( .A(n31615), .X(n34463) );
  inv_x1_sg U40228 ( .A(n31614), .X(n34464) );
  inv_x1_sg U40229 ( .A(n34923), .X(n34465) );
  inv_x1_sg U40230 ( .A(n34465), .X(n34466) );
  inv_x1_sg U40231 ( .A(n30821), .X(n34467) );
  inv_x1_sg U40232 ( .A(n30119), .X(n34468) );
  inv_x1_sg U40233 ( .A(n34465), .X(n34469) );
  inv_x1_sg U40234 ( .A(n34924), .X(n34470) );
  inv_x1_sg U40235 ( .A(n34470), .X(n34471) );
  inv_x1_sg U40236 ( .A(n30817), .X(n34472) );
  inv_x1_sg U40237 ( .A(n34470), .X(n34473) );
  inv_x1_sg U40238 ( .A(n34470), .X(n34474) );
  inv_x1_sg U40239 ( .A(n29686), .X(n34475) );
  inv_x1_sg U40240 ( .A(n31618), .X(n34476) );
  inv_x1_sg U40241 ( .A(n34921), .X(n34477) );
  inv_x1_sg U40242 ( .A(n34477), .X(n34478) );
  inv_x1_sg U40243 ( .A(n30812), .X(n34479) );
  inv_x1_sg U40244 ( .A(n30120), .X(n34480) );
  inv_x1_sg U40245 ( .A(n34477), .X(n34481) );
  inv_x1_sg U40246 ( .A(n34920), .X(n34482) );
  inv_x1_sg U40247 ( .A(n34482), .X(n34483) );
  inv_x1_sg U40248 ( .A(n30121), .X(n34484) );
  inv_x1_sg U40249 ( .A(n30808), .X(n34485) );
  inv_x1_sg U40250 ( .A(n34482), .X(n34486) );
  inv_x1_sg U40251 ( .A(n34919), .X(n34487) );
  inv_x1_sg U40252 ( .A(n34487), .X(n34488) );
  inv_x1_sg U40253 ( .A(n30804), .X(n34489) );
  inv_x1_sg U40254 ( .A(n30122), .X(n34490) );
  inv_x1_sg U40255 ( .A(n34487), .X(n34491) );
  inv_x1_sg U40256 ( .A(n34955), .X(n34492) );
  inv_x1_sg U40257 ( .A(n34492), .X(n34493) );
  inv_x1_sg U40258 ( .A(n30800), .X(n34494) );
  inv_x1_sg U40259 ( .A(n34492), .X(n34495) );
  inv_x1_sg U40260 ( .A(n30800), .X(n34496) );
  inv_x1_sg U40261 ( .A(n34949), .X(n34497) );
  inv_x1_sg U40262 ( .A(n34497), .X(n34498) );
  inv_x1_sg U40263 ( .A(n30797), .X(n34499) );
  inv_x1_sg U40264 ( .A(n34497), .X(n34500) );
  inv_x1_sg U40265 ( .A(n30797), .X(n34501) );
  inv_x1_sg U40266 ( .A(n34933), .X(n34502) );
  inv_x1_sg U40267 ( .A(n34502), .X(n34503) );
  inv_x1_sg U40268 ( .A(n34502), .X(n34504) );
  inv_x1_sg U40269 ( .A(n30126), .X(n34505) );
  inv_x1_sg U40270 ( .A(n30794), .X(n34506) );
  inv_x1_sg U40271 ( .A(n34925), .X(n34507) );
  inv_x1_sg U40272 ( .A(n34507), .X(n34508) );
  inv_x1_sg U40273 ( .A(n30791), .X(n34509) );
  inv_x1_sg U40274 ( .A(n30128), .X(n34510) );
  inv_x1_sg U40275 ( .A(n34507), .X(n34511) );
  inv_x1_sg U40276 ( .A(n11716), .X(n34512) );
  inv_x1_sg U40277 ( .A(n30787), .X(n34513) );
  inv_x1_sg U40278 ( .A(n34512), .X(n34514) );
  inv_x1_sg U40279 ( .A(n30787), .X(n34515) );
  inv_x1_sg U40280 ( .A(n34512), .X(n34516) );
  inv_x1_sg U40281 ( .A(n35655), .X(n34517) );
  inv_x1_sg U40282 ( .A(n34517), .X(n34518) );
  inv_x1_sg U40283 ( .A(n34517), .X(n34519) );
  inv_x1_sg U40284 ( .A(n34517), .X(n34520) );
  inv_x1_sg U40285 ( .A(n29682), .X(n34521) );
  inv_x1_sg U40286 ( .A(n31005), .X(n34522) );
  inv_x1_sg U40287 ( .A(n31005), .X(n34523) );
  inv_x1_sg U40288 ( .A(n31004), .X(n34524) );
  inv_x1_sg U40289 ( .A(n31009), .X(n34525) );
  inv_x1_sg U40290 ( .A(n31010), .X(n34526) );
  inv_x1_sg U40291 ( .A(n31010), .X(n34527) );
  inv_x1_sg U40292 ( .A(n31009), .X(n34528) );
  inv_x1_sg U40293 ( .A(n31014), .X(n34529) );
  inv_x1_sg U40294 ( .A(n31014), .X(n34530) );
  inv_x1_sg U40295 ( .A(n31015), .X(n34531) );
  inv_x1_sg U40296 ( .A(n31014), .X(n34532) );
  inv_x1_sg U40297 ( .A(n13224), .X(n34533) );
  inv_x1_sg U40298 ( .A(n34533), .X(n34534) );
  inv_x1_sg U40299 ( .A(n31018), .X(n34535) );
  inv_x1_sg U40300 ( .A(n34533), .X(n34536) );
  inv_x1_sg U40301 ( .A(n31018), .X(n34537) );
  inv_x1_sg U40302 ( .A(n19589), .X(n34538) );
  inv_x1_sg U40303 ( .A(n34538), .X(n34539) );
  inv_x1_sg U40304 ( .A(n34538), .X(n34540) );
  inv_x1_sg U40305 ( .A(n29676), .X(n34541) );
  inv_x1_sg U40306 ( .A(n29676), .X(n34542) );
  inv_x1_sg U40307 ( .A(n35416), .X(n34543) );
  inv_x1_sg U40308 ( .A(n31301), .X(n34544) );
  inv_x1_sg U40309 ( .A(n31301), .X(n34545) );
  inv_x1_sg U40310 ( .A(n34543), .X(n34546) );
  inv_x1_sg U40311 ( .A(\shifter_0/pointer[3] ), .X(n34547) );
  inv_x1_sg U40312 ( .A(n34547), .X(n34548) );
  inv_x1_sg U40313 ( .A(n31298), .X(n34549) );
  inv_x1_sg U40314 ( .A(n30142), .X(n34550) );
  inv_x1_sg U40315 ( .A(n35263), .X(n34551) );
  inv_x1_sg U40316 ( .A(n32051), .X(n34552) );
  inv_x1_sg U40317 ( .A(n35076), .X(n34553) );
  inv_x1_sg U40318 ( .A(n30754), .X(n34554) );
  inv_x1_sg U40319 ( .A(n34554), .X(n34555) );
  inv_x1_sg U40320 ( .A(n34554), .X(n34556) );
  inv_x1_sg U40321 ( .A(n34554), .X(n34557) );
  inv_x1_sg U40322 ( .A(n34554), .X(n34558) );
  inv_x1_sg U40323 ( .A(n32392), .X(n34559) );
  inv_x1_sg U40324 ( .A(n34559), .X(n34560) );
  inv_x1_sg U40325 ( .A(n34551), .X(n34561) );
  inv_x1_sg U40326 ( .A(n31300), .X(n34562) );
  inv_x1_sg U40327 ( .A(n32168), .X(n34563) );
  inv_x1_sg U40328 ( .A(n30596), .X(n34564) );
  inv_x1_sg U40329 ( .A(n34564), .X(n34565) );
  inv_x1_sg U40330 ( .A(n34564), .X(n34566) );
  inv_x1_sg U40331 ( .A(n30783), .X(n34567) );
  inv_x1_sg U40332 ( .A(n30783), .X(n34568) );
  inv_x1_sg U40333 ( .A(n35079), .X(n34569) );
  inv_x1_sg U40334 ( .A(n34569), .X(n34570) );
  inv_x1_sg U40335 ( .A(n34569), .X(n34571) );
  inv_x1_sg U40336 ( .A(n30781), .X(n34572) );
  inv_x1_sg U40337 ( .A(n30781), .X(n34573) );
  inv_x1_sg U40338 ( .A(n35078), .X(n34574) );
  inv_x1_sg U40339 ( .A(n34574), .X(n34575) );
  inv_x1_sg U40340 ( .A(n34574), .X(n34576) );
  inv_x1_sg U40341 ( .A(n30780), .X(n34577) );
  inv_x1_sg U40342 ( .A(n30780), .X(n34578) );
  inv_x1_sg U40343 ( .A(n35077), .X(n34579) );
  inv_x1_sg U40344 ( .A(n34579), .X(n34580) );
  inv_x1_sg U40345 ( .A(n34579), .X(n34581) );
  inv_x1_sg U40346 ( .A(n30779), .X(n34582) );
  inv_x1_sg U40347 ( .A(n30779), .X(n34583) );
  inv_x1_sg U40348 ( .A(n34552), .X(n34584) );
  inv_x1_sg U40349 ( .A(n34584), .X(n34585) );
  inv_x1_sg U40350 ( .A(n34584), .X(n34586) );
  inv_x1_sg U40351 ( .A(n30213), .X(n34587) );
  inv_x1_sg U40352 ( .A(n34587), .X(n34588) );
  inv_x1_sg U40353 ( .A(n34587), .X(n34589) );
  inv_x1_sg U40354 ( .A(n34587), .X(n34590) );
  inv_x1_sg U40355 ( .A(n30597), .X(n34591) );
  inv_x1_sg U40356 ( .A(n34591), .X(n34592) );
  inv_x1_sg U40357 ( .A(n34591), .X(n34593) );
  inv_x1_sg U40358 ( .A(n34591), .X(n34594) );
  inv_x1_sg U40359 ( .A(n34591), .X(n34595) );
  inv_x1_sg U40360 ( .A(n30208), .X(n34596) );
  inv_x1_sg U40361 ( .A(n34596), .X(n34597) );
  inv_x1_sg U40362 ( .A(n34596), .X(n34598) );
  inv_x1_sg U40363 ( .A(n34596), .X(n34599) );
  inv_x1_sg U40364 ( .A(n35466), .X(n34600) );
  inv_x1_sg U40365 ( .A(n34600), .X(n34601) );
  inv_x1_sg U40366 ( .A(n34600), .X(n34602) );
  inv_x1_sg U40367 ( .A(n29675), .X(n34603) );
  inv_x1_sg U40368 ( .A(n30778), .X(n34604) );
  inv_x1_sg U40369 ( .A(n30256), .X(n34605) );
  inv_x1_sg U40370 ( .A(n34605), .X(n34606) );
  inv_x1_sg U40371 ( .A(n34605), .X(n34607) );
  inv_x1_sg U40372 ( .A(n30776), .X(n34608) );
  inv_x1_sg U40373 ( .A(n30776), .X(n34609) );
  inv_x1_sg U40374 ( .A(n34902), .X(n34610) );
  inv_x1_sg U40375 ( .A(n34610), .X(n34611) );
  inv_x1_sg U40376 ( .A(n34610), .X(n34612) );
  inv_x1_sg U40377 ( .A(n34610), .X(n34613) );
  inv_x1_sg U40378 ( .A(n34610), .X(n34614) );
  inv_x1_sg U40379 ( .A(n34901), .X(n34615) );
  inv_x1_sg U40380 ( .A(n34615), .X(n34616) );
  inv_x1_sg U40381 ( .A(n34615), .X(n34617) );
  inv_x1_sg U40382 ( .A(n34615), .X(n34618) );
  inv_x1_sg U40383 ( .A(n34615), .X(n34619) );
  inv_x1_sg U40384 ( .A(n31605), .X(n34620) );
  inv_x1_sg U40385 ( .A(n35071), .X(n34621) );
  inv_x1_sg U40386 ( .A(n30250), .X(n34622) );
  inv_x1_sg U40387 ( .A(n34622), .X(n34623) );
  inv_x1_sg U40388 ( .A(n34622), .X(n34624) );
  inv_x1_sg U40389 ( .A(n30771), .X(n34625) );
  inv_x1_sg U40390 ( .A(n34622), .X(n34626) );
  inv_x1_sg U40391 ( .A(n31914), .X(n34627) );
  inv_x1_sg U40392 ( .A(n34627), .X(n34628) );
  inv_x1_sg U40393 ( .A(n34627), .X(n34629) );
  inv_x1_sg U40394 ( .A(n30163), .X(n34630) );
  inv_x1_sg U40395 ( .A(n30769), .X(n34631) );
  inv_x1_sg U40396 ( .A(n30251), .X(n34632) );
  inv_x1_sg U40397 ( .A(n29673), .X(n34633) );
  inv_x1_sg U40398 ( .A(n34632), .X(n34634) );
  inv_x1_sg U40399 ( .A(n34632), .X(n34635) );
  inv_x1_sg U40400 ( .A(n30766), .X(n34636) );
  inv_x1_sg U40401 ( .A(n31606), .X(n34637) );
  inv_x1_sg U40402 ( .A(n31109), .X(n34638) );
  inv_x1_sg U40403 ( .A(n30248), .X(n34639) );
  inv_x1_sg U40404 ( .A(n34639), .X(n34640) );
  inv_x1_sg U40405 ( .A(n34639), .X(n34641) );
  inv_x1_sg U40406 ( .A(n30760), .X(n34642) );
  inv_x1_sg U40407 ( .A(n34639), .X(n34643) );
  inv_x1_sg U40408 ( .A(n31920), .X(n34644) );
  inv_x1_sg U40409 ( .A(n34644), .X(n34645) );
  inv_x1_sg U40410 ( .A(n34644), .X(n34646) );
  inv_x1_sg U40411 ( .A(n34644), .X(n34647) );
  inv_x1_sg U40412 ( .A(n30759), .X(n34648) );
  inv_x1_sg U40413 ( .A(n34941), .X(n34649) );
  inv_x1_sg U40414 ( .A(n34649), .X(n34650) );
  inv_x1_sg U40415 ( .A(n30756), .X(n34651) );
  inv_x1_sg U40416 ( .A(n30756), .X(n34652) );
  inv_x1_sg U40417 ( .A(n34649), .X(n34653) );
  inv_x1_sg U40418 ( .A(n35683), .X(n34654) );
  inv_x1_sg U40419 ( .A(n30753), .X(n34655) );
  inv_x1_sg U40420 ( .A(n34654), .X(n34656) );
  inv_x1_sg U40421 ( .A(n34654), .X(n34657) );
  inv_x1_sg U40422 ( .A(n30753), .X(n34658) );
  inv_x1_sg U40423 ( .A(n35394), .X(n34659) );
  inv_x1_sg U40424 ( .A(n35238), .X(n34660) );
  inv_x1_sg U40425 ( .A(n35091), .X(n34661) );
  inv_x1_sg U40426 ( .A(n34661), .X(n34662) );
  inv_x1_sg U40427 ( .A(n34661), .X(n34663) );
  inv_x1_sg U40428 ( .A(n35092), .X(n34664) );
  inv_x1_sg U40429 ( .A(n34664), .X(n34665) );
  inv_x1_sg U40430 ( .A(n34664), .X(n34666) );
  inv_x1_sg U40431 ( .A(n30750), .X(n34667) );
  inv_x1_sg U40432 ( .A(n30750), .X(n34668) );
  inv_x1_sg U40433 ( .A(n35068), .X(n34669) );
  inv_x1_sg U40434 ( .A(n34669), .X(n34670) );
  inv_x1_sg U40435 ( .A(n30167), .X(n34671) );
  inv_x1_sg U40436 ( .A(n34669), .X(n34672) );
  inv_x1_sg U40437 ( .A(n30746), .X(n34673) );
  inv_x1_sg U40438 ( .A(n35064), .X(n34674) );
  inv_x1_sg U40439 ( .A(n30743), .X(n34675) );
  inv_x1_sg U40440 ( .A(n34674), .X(n34676) );
  inv_x1_sg U40441 ( .A(n34674), .X(n34677) );
  inv_x1_sg U40442 ( .A(n34674), .X(n34678) );
  inv_x1_sg U40443 ( .A(n35061), .X(n34679) );
  inv_x1_sg U40444 ( .A(n30740), .X(n34680) );
  inv_x1_sg U40445 ( .A(n34679), .X(n34681) );
  inv_x1_sg U40446 ( .A(n34679), .X(n34682) );
  inv_x1_sg U40447 ( .A(n34679), .X(n34683) );
  inv_x1_sg U40448 ( .A(n35065), .X(n34684) );
  inv_x1_sg U40449 ( .A(n30737), .X(n34685) );
  inv_x1_sg U40450 ( .A(n34684), .X(n34686) );
  inv_x1_sg U40451 ( .A(n34684), .X(n34687) );
  inv_x1_sg U40452 ( .A(n30737), .X(n34688) );
  inv_x1_sg U40453 ( .A(n35064), .X(n34689) );
  inv_x1_sg U40454 ( .A(n34689), .X(n34690) );
  inv_x1_sg U40455 ( .A(n30734), .X(n34691) );
  inv_x1_sg U40456 ( .A(n34689), .X(n34692) );
  inv_x1_sg U40457 ( .A(n34689), .X(n34693) );
  inv_x1_sg U40458 ( .A(n34942), .X(n34694) );
  inv_x1_sg U40459 ( .A(n34694), .X(n34695) );
  inv_x1_sg U40460 ( .A(n30731), .X(n34696) );
  inv_x1_sg U40461 ( .A(n30731), .X(n34697) );
  inv_x1_sg U40462 ( .A(n34694), .X(n34698) );
  inv_x1_sg U40463 ( .A(n35166), .X(n34699) );
  inv_x1_sg U40464 ( .A(n35088), .X(n34700) );
  inv_x1_sg U40465 ( .A(n34700), .X(n34701) );
  inv_x1_sg U40466 ( .A(n34700), .X(n34702) );
  inv_x1_sg U40467 ( .A(n34700), .X(n34703) );
  inv_x1_sg U40468 ( .A(n30728), .X(n34704) );
  inv_x1_sg U40469 ( .A(n35364), .X(n34705) );
  inv_x1_sg U40470 ( .A(n35385), .X(n34706) );
  inv_x1_sg U40471 ( .A(n35387), .X(n34707) );
  inv_x1_sg U40472 ( .A(n35166), .X(n34708) );
  inv_x1_sg U40473 ( .A(n35343), .X(n34709) );
  inv_x1_sg U40474 ( .A(n35383), .X(n34710) );
  inv_x1_sg U40475 ( .A(n35393), .X(n34711) );
  inv_x1_sg U40476 ( .A(n35386), .X(n34712) );
  inv_x1_sg U40477 ( .A(n35378), .X(n34713) );
  inv_x1_sg U40478 ( .A(n35349), .X(n34714) );
  inv_x1_sg U40479 ( .A(n35081), .X(n34715) );
  inv_x1_sg U40480 ( .A(n34715), .X(n34716) );
  inv_x1_sg U40481 ( .A(n34715), .X(n34717) );
  inv_x1_sg U40482 ( .A(n34715), .X(n34718) );
  inv_x1_sg U40483 ( .A(n34715), .X(n34719) );
  inv_x1_sg U40484 ( .A(n35082), .X(n34720) );
  inv_x1_sg U40485 ( .A(n34720), .X(n34721) );
  inv_x1_sg U40486 ( .A(n34720), .X(n34722) );
  inv_x1_sg U40487 ( .A(n34720), .X(n34723) );
  inv_x1_sg U40488 ( .A(n34720), .X(n34724) );
  inv_x1_sg U40489 ( .A(n31609), .X(n34725) );
  inv_x1_sg U40490 ( .A(n34967), .X(n34726) );
  inv_x1_sg U40491 ( .A(n34726), .X(n34727) );
  inv_x1_sg U40492 ( .A(n34726), .X(n34728) );
  inv_x1_sg U40493 ( .A(n34726), .X(n34729) );
  inv_x1_sg U40494 ( .A(n34726), .X(n34730) );
  inv_x1_sg U40495 ( .A(n30703), .X(n34731) );
  inv_x1_sg U40496 ( .A(n30700), .X(n34732) );
  inv_x1_sg U40497 ( .A(n30700), .X(n34733) );
  inv_x1_sg U40498 ( .A(n30699), .X(n34734) );
  inv_x1_sg U40499 ( .A(n34965), .X(n34735) );
  inv_x1_sg U40500 ( .A(n34735), .X(n34736) );
  inv_x1_sg U40501 ( .A(n34735), .X(n34737) );
  inv_x1_sg U40502 ( .A(n30695), .X(n34738) );
  inv_x1_sg U40503 ( .A(n30181), .X(n34739) );
  inv_x1_sg U40504 ( .A(n34959), .X(n34740) );
  inv_x1_sg U40505 ( .A(n34740), .X(n34741) );
  inv_x1_sg U40506 ( .A(n30182), .X(n34742) );
  inv_x1_sg U40507 ( .A(n34740), .X(n34743) );
  inv_x1_sg U40508 ( .A(n30691), .X(n34744) );
  inv_x1_sg U40509 ( .A(n34961), .X(n34745) );
  inv_x1_sg U40510 ( .A(n34745), .X(n34746) );
  inv_x1_sg U40511 ( .A(n34745), .X(n34747) );
  inv_x1_sg U40512 ( .A(n30687), .X(n34748) );
  inv_x1_sg U40513 ( .A(n34745), .X(n34749) );
  inv_x1_sg U40514 ( .A(n34960), .X(n34750) );
  inv_x1_sg U40515 ( .A(n34750), .X(n34751) );
  inv_x1_sg U40516 ( .A(n34750), .X(n34752) );
  inv_x1_sg U40517 ( .A(n30683), .X(n34753) );
  inv_x1_sg U40518 ( .A(n34750), .X(n34754) );
  inv_x1_sg U40519 ( .A(n34954), .X(n34755) );
  inv_x1_sg U40520 ( .A(n30184), .X(n34756) );
  inv_x1_sg U40521 ( .A(n34755), .X(n34757) );
  inv_x1_sg U40522 ( .A(n30679), .X(n34758) );
  inv_x1_sg U40523 ( .A(n30184), .X(n34759) );
  inv_x1_sg U40524 ( .A(n34953), .X(n34760) );
  inv_x1_sg U40525 ( .A(n34760), .X(n34761) );
  inv_x1_sg U40526 ( .A(n34760), .X(n34762) );
  inv_x1_sg U40527 ( .A(n30672), .X(n34763) );
  inv_x1_sg U40528 ( .A(n30672), .X(n34764) );
  inv_x1_sg U40529 ( .A(n30214), .X(n34765) );
  inv_x1_sg U40530 ( .A(n34765), .X(n34766) );
  inv_x1_sg U40531 ( .A(n34765), .X(n34767) );
  inv_x1_sg U40532 ( .A(n30670), .X(n34768) );
  inv_x1_sg U40533 ( .A(n34765), .X(n34769) );
  inv_x1_sg U40534 ( .A(n34951), .X(n34770) );
  inv_x1_sg U40535 ( .A(n34770), .X(n34771) );
  inv_x1_sg U40536 ( .A(n34770), .X(n34772) );
  inv_x1_sg U40537 ( .A(n30666), .X(n34773) );
  inv_x1_sg U40538 ( .A(n34770), .X(n34774) );
  inv_x1_sg U40539 ( .A(n30664), .X(n34775) );
  inv_x1_sg U40540 ( .A(n34775), .X(n34776) );
  inv_x1_sg U40541 ( .A(n34775), .X(n34777) );
  inv_x1_sg U40542 ( .A(n30662), .X(n34778) );
  inv_x1_sg U40543 ( .A(n34775), .X(n34779) );
  inv_x1_sg U40544 ( .A(n34945), .X(n34780) );
  inv_x1_sg U40545 ( .A(n34780), .X(n34781) );
  inv_x1_sg U40546 ( .A(n34780), .X(n34782) );
  inv_x1_sg U40547 ( .A(n30658), .X(n34783) );
  inv_x1_sg U40548 ( .A(n34780), .X(n34784) );
  inv_x1_sg U40549 ( .A(n34948), .X(n34785) );
  inv_x1_sg U40550 ( .A(n34785), .X(n34786) );
  inv_x1_sg U40551 ( .A(n34785), .X(n34787) );
  inv_x1_sg U40552 ( .A(n30654), .X(n34788) );
  inv_x1_sg U40553 ( .A(n34785), .X(n34789) );
  inv_x1_sg U40554 ( .A(n34947), .X(n34790) );
  inv_x1_sg U40555 ( .A(n34790), .X(n34791) );
  inv_x1_sg U40556 ( .A(n34790), .X(n34792) );
  inv_x1_sg U40557 ( .A(n30650), .X(n34793) );
  inv_x1_sg U40558 ( .A(n34790), .X(n34794) );
  inv_x1_sg U40559 ( .A(n26219), .X(n34795) );
  inv_x1_sg U40560 ( .A(n30646), .X(n34796) );
  inv_x1_sg U40561 ( .A(n34795), .X(n34797) );
  inv_x1_sg U40562 ( .A(n30646), .X(n34798) );
  inv_x1_sg U40563 ( .A(n34795), .X(n34799) );
  inv_x1_sg U40564 ( .A(n34958), .X(n34800) );
  inv_x1_sg U40565 ( .A(n30189), .X(n34801) );
  inv_x1_sg U40566 ( .A(n34800), .X(n34802) );
  inv_x1_sg U40567 ( .A(n34800), .X(n34803) );
  inv_x1_sg U40568 ( .A(n30643), .X(n34804) );
  inv_x1_sg U40569 ( .A(n34861), .X(n34805) );
  inv_x1_sg U40570 ( .A(n34805), .X(n34806) );
  inv_x1_sg U40571 ( .A(n30639), .X(n34807) );
  inv_x1_sg U40572 ( .A(n30639), .X(n34808) );
  inv_x1_sg U40573 ( .A(n31283), .X(n34809) );
  inv_x1_sg U40574 ( .A(n31288), .X(n34810) );
  inv_x1_sg U40575 ( .A(n31289), .X(n34811) );
  inv_x1_sg U40576 ( .A(n31289), .X(n34812) );
  inv_x1_sg U40577 ( .A(n31279), .X(n34813) );
  inv_x1_sg U40578 ( .A(n31283), .X(n34814) );
  inv_x1_sg U40579 ( .A(n31284), .X(n34815) );
  inv_x1_sg U40580 ( .A(n31284), .X(n34816) );
  inv_x1_sg U40581 ( .A(n35058), .X(n34817) );
  inv_x1_sg U40582 ( .A(n30374), .X(n34818) );
  inv_x1_sg U40583 ( .A(n31279), .X(n34819) );
  inv_x1_sg U40584 ( .A(n31280), .X(n34820) );
  inv_x1_sg U40585 ( .A(n31280), .X(n34821) );
  inv_x1_sg U40586 ( .A(n34915), .X(n34822) );
  inv_x1_sg U40587 ( .A(n31275), .X(n34823) );
  inv_x1_sg U40588 ( .A(n31274), .X(n34824) );
  inv_x1_sg U40589 ( .A(n30377), .X(n34825) );
  inv_x1_sg U40590 ( .A(n31275), .X(n34826) );
  inv_x1_sg U40591 ( .A(n31270), .X(n34827) );
  inv_x1_sg U40592 ( .A(n31269), .X(n34828) );
  inv_x1_sg U40593 ( .A(n31269), .X(n34829) );
  inv_x1_sg U40594 ( .A(n31269), .X(n34830) );
  inv_x1_sg U40595 ( .A(n35053), .X(n34831) );
  inv_x1_sg U40596 ( .A(n29686), .X(n34832) );
  inv_x1_sg U40597 ( .A(n34836), .X(n34833) );
  inv_x1_sg U40598 ( .A(n31265), .X(n34834) );
  inv_x1_sg U40599 ( .A(n31264), .X(n34835) );
  inv_x1_sg U40600 ( .A(n34918), .X(n34836) );
  inv_x1_sg U40601 ( .A(n30600), .X(n34837) );
  inv_x1_sg U40602 ( .A(n30600), .X(n34838) );
  inv_x1_sg U40603 ( .A(n31261), .X(n34839) );
  inv_x1_sg U40604 ( .A(n31260), .X(n34840) );
  inv_x1_sg U40605 ( .A(n34917), .X(n34841) );
  inv_x1_sg U40606 ( .A(n30618), .X(n34842) );
  inv_x1_sg U40607 ( .A(n34831), .X(n34843) );
  inv_x1_sg U40608 ( .A(n31256), .X(n34844) );
  inv_x1_sg U40609 ( .A(n31256), .X(n34845) );
  inv_x1_sg U40610 ( .A(n32052), .X(n34846) );
  inv_x1_sg U40611 ( .A(n32052), .X(n34847) );
  inv_x1_sg U40612 ( .A(n32347), .X(n34848) );
  inv_x1_sg U40613 ( .A(n34848), .X(n34849) );
  inv_x1_sg U40614 ( .A(n34848), .X(n34850) );
  inv_x1_sg U40615 ( .A(n34848), .X(n34851) );
  inv_x1_sg U40616 ( .A(n30637), .X(n34852) );
  inv_x1_sg U40617 ( .A(\shifter_0/pointer[0] ), .X(n34853) );
  inv_x1_sg U40618 ( .A(n34853), .X(n34854) );
  inv_x1_sg U40619 ( .A(n35417), .X(n34855) );
  inv_x1_sg U40620 ( .A(n34853), .X(n34856) );
  inv_x1_sg U40621 ( .A(n35417), .X(n34857) );
  inv_x1_sg U40622 ( .A(n34853), .X(n34858) );
  inv_x1_sg U40623 ( .A(\shifter_0/pointer[0] ), .X(n34859) );
  inv_x1_sg U40624 ( .A(n34855), .X(n34860) );
  inv_x1_sg U40625 ( .A(n30635), .X(n34861) );
  inv_x1_sg U40626 ( .A(n26352), .X(n34862) );
  inv_x1_sg U40627 ( .A(n34862), .X(n34863) );
  inv_x1_sg U40628 ( .A(n30634), .X(n34864) );
  inv_x1_sg U40629 ( .A(n34862), .X(n34865) );
  inv_x1_sg U40630 ( .A(n34862), .X(n34866) );
  nor_x1_sg U40631 ( .A(n35459), .B(n26206), .X(n34867) );
  inv_x1_sg U40632 ( .A(n34867), .X(n34868) );
  inv_x1_sg U40633 ( .A(n31619), .X(n34869) );
  inv_x1_sg U40634 ( .A(n30202), .X(n34870) );
  inv_x1_sg U40635 ( .A(n34868), .X(n34871) );
  inv_x1_sg U40636 ( .A(n30631), .X(n34872) );
  inv_x1_sg U40637 ( .A(n31620), .X(n34873) );
  inv_x1_sg U40638 ( .A(n31253), .X(n34874) );
  inv_x1_sg U40639 ( .A(n31253), .X(n34875) );
  inv_x1_sg U40640 ( .A(n31619), .X(n34876) );
  inv_x1_sg U40641 ( .A(n34904), .X(n34877) );
  inv_x1_sg U40642 ( .A(n34877), .X(n34878) );
  inv_x1_sg U40643 ( .A(n34877), .X(n34879) );
  inv_x1_sg U40644 ( .A(n34877), .X(n34880) );
  inv_x1_sg U40645 ( .A(n30630), .X(n34881) );
  inv_x1_sg U40646 ( .A(n35412), .X(n34882) );
  inv_x1_sg U40647 ( .A(n34882), .X(n34883) );
  inv_x1_sg U40648 ( .A(n34882), .X(n34884) );
  inv_x1_sg U40649 ( .A(n34882), .X(n34885) );
  inv_x1_sg U40650 ( .A(n30628), .X(n34886) );
  inv_x1_sg U40651 ( .A(n34903), .X(n34887) );
  inv_x1_sg U40652 ( .A(n34887), .X(n34888) );
  inv_x1_sg U40653 ( .A(n34887), .X(n34889) );
  inv_x1_sg U40654 ( .A(n34887), .X(n34890) );
  inv_x1_sg U40655 ( .A(n30626), .X(n34891) );
  inv_x1_sg U40656 ( .A(n34939), .X(n34892) );
  inv_x1_sg U40657 ( .A(n34892), .X(n34893) );
  inv_x1_sg U40658 ( .A(n30624), .X(n34894) );
  inv_x1_sg U40659 ( .A(n34892), .X(n34895) );
  inv_x1_sg U40660 ( .A(n30624), .X(n34896) );
  inv_x1_sg U40661 ( .A(n32051), .X(n34897) );
  inv_x1_sg U40662 ( .A(n35076), .X(n34898) );
  inv_x1_sg U40663 ( .A(n32359), .X(n34899) );
  inv_x1_sg U40664 ( .A(n34899), .X(n34900) );
  inv_x1_sg U40665 ( .A(n34899), .X(n34901) );
  inv_x1_sg U40666 ( .A(n34899), .X(n34902) );
  inv_x1_sg U40667 ( .A(n35485), .X(n34903) );
  inv_x1_sg U40668 ( .A(n32008), .X(n34904) );
  inv_x1_sg U40669 ( .A(n32275), .X(n34905) );
  inv_x1_sg U40670 ( .A(n31245), .X(n34906) );
  inv_x1_sg U40671 ( .A(n30778), .X(n34907) );
  inv_x1_sg U40672 ( .A(n31246), .X(n34908) );
  inv_x1_sg U40673 ( .A(n31245), .X(n34909) );
  inv_x1_sg U40674 ( .A(n32263), .X(n34910) );
  inv_x1_sg U40675 ( .A(n31240), .X(n34911) );
  inv_x1_sg U40676 ( .A(n30630), .X(n34912) );
  inv_x1_sg U40677 ( .A(n29680), .X(n34913) );
  inv_x1_sg U40678 ( .A(n29680), .X(n34914) );
  inv_x1_sg U40679 ( .A(n31108), .X(n34915) );
  inv_x1_sg U40680 ( .A(n31607), .X(n34916) );
  inv_x1_sg U40681 ( .A(n31608), .X(n34917) );
  inv_x1_sg U40682 ( .A(n35051), .X(n34918) );
  inv_x1_sg U40683 ( .A(n31104), .X(n34919) );
  inv_x1_sg U40684 ( .A(n31618), .X(n34920) );
  inv_x1_sg U40685 ( .A(n31617), .X(n34921) );
  inv_x1_sg U40686 ( .A(n31618), .X(n34922) );
  inv_x1_sg U40687 ( .A(n31101), .X(n34923) );
  inv_x1_sg U40688 ( .A(n29685), .X(n34924) );
  inv_x1_sg U40689 ( .A(n31614), .X(n34925) );
  inv_x1_sg U40690 ( .A(n31614), .X(n34926) );
  inv_x1_sg U40691 ( .A(n30822), .X(n34927) );
  inv_x1_sg U40692 ( .A(n31479), .X(n34928) );
  inv_x1_sg U40693 ( .A(n29682), .X(n34929) );
  inv_x1_sg U40694 ( .A(n31478), .X(n34930) );
  inv_x1_sg U40695 ( .A(n31478), .X(n34931) );
  inv_x1_sg U40696 ( .A(n31098), .X(n34932) );
  inv_x1_sg U40697 ( .A(n31611), .X(n34933) );
  inv_x1_sg U40698 ( .A(n31612), .X(n34934) );
  inv_x1_sg U40699 ( .A(n31612), .X(n34935) );
  inv_x1_sg U40700 ( .A(n32052), .X(n34936) );
  inv_x1_sg U40701 ( .A(n32051), .X(n34937) );
  inv_x1_sg U40702 ( .A(n34849), .X(n34938) );
  inv_x1_sg U40703 ( .A(n34938), .X(n34939) );
  inv_x1_sg U40704 ( .A(n34938), .X(n34940) );
  inv_x1_sg U40705 ( .A(n34938), .X(n34941) );
  inv_x1_sg U40706 ( .A(n34938), .X(n34942) );
  nor_x1_sg U40707 ( .A(n31604), .B(n33824), .X(n34943) );
  inv_x1_sg U40708 ( .A(n34943), .X(n34944) );
  inv_x1_sg U40709 ( .A(n30609), .X(n34945) );
  inv_x1_sg U40710 ( .A(n34944), .X(n34946) );
  inv_x1_sg U40711 ( .A(n34944), .X(n34947) );
  inv_x1_sg U40712 ( .A(n30609), .X(n34948) );
  inv_x1_sg U40713 ( .A(n34944), .X(n34949) );
  inv_x1_sg U40714 ( .A(n18763), .X(n34950) );
  inv_x1_sg U40715 ( .A(n34950), .X(n34951) );
  inv_x1_sg U40716 ( .A(n34950), .X(n34952) );
  inv_x1_sg U40717 ( .A(n30609), .X(n34953) );
  inv_x1_sg U40718 ( .A(n34950), .X(n34954) );
  inv_x1_sg U40719 ( .A(n34950), .X(n34955) );
  nor_x1_sg U40720 ( .A(n31603), .B(n33820), .X(n34956) );
  inv_x1_sg U40721 ( .A(n34956), .X(n34957) );
  inv_x1_sg U40722 ( .A(n34957), .X(n34958) );
  inv_x1_sg U40723 ( .A(n31234), .X(n34959) );
  inv_x1_sg U40724 ( .A(n31234), .X(n34960) );
  inv_x1_sg U40725 ( .A(n34957), .X(n34961) );
  inv_x1_sg U40726 ( .A(n34957), .X(n34962) );
  inv_x1_sg U40727 ( .A(n35685), .X(n34963) );
  inv_x1_sg U40728 ( .A(n31609), .X(n34964) );
  inv_x1_sg U40729 ( .A(n31107), .X(n34965) );
  inv_x1_sg U40730 ( .A(n31107), .X(n34966) );
  inv_x1_sg U40731 ( .A(n29684), .X(n34967) );
  inv_x1_sg U40732 ( .A(n29684), .X(n34968) );
  nor_x1_sg U40733 ( .A(n42537), .B(n31603), .X(n34969) );
  inv_x1_sg U40734 ( .A(n34969), .X(n34970) );
  inv_x1_sg U40735 ( .A(n31229), .X(n34971) );
  inv_x1_sg U40736 ( .A(n29679), .X(n34972) );
  inv_x1_sg U40737 ( .A(n31229), .X(n34973) );
  inv_x1_sg U40738 ( .A(n34970), .X(n34974) );
  inv_x1_sg U40739 ( .A(n31544), .X(n34975) );
  inv_x1_sg U40740 ( .A(n31544), .X(n34976) );
  inv_x1_sg U40741 ( .A(n31230), .X(n34977) );
  inv_x1_sg U40742 ( .A(n34973), .X(n34978) );
  inv_x1_sg U40743 ( .A(n31231), .X(n34979) );
  inv_x1_sg U40744 ( .A(n34971), .X(n34980) );
  inv_x1_sg U40745 ( .A(n31231), .X(n34981) );
  inv_x1_sg U40746 ( .A(n31230), .X(n34982) );
  inv_x1_sg U40747 ( .A(n31545), .X(n34983) );
  inv_x1_sg U40748 ( .A(n34971), .X(n34984) );
  inv_x1_sg U40749 ( .A(n34971), .X(n34985) );
  inv_x1_sg U40750 ( .A(n30217), .X(n34986) );
  inv_x1_sg U40751 ( .A(n30217), .X(n34987) );
  inv_x1_sg U40752 ( .A(n34972), .X(n34988) );
  inv_x1_sg U40753 ( .A(n31545), .X(n34989) );
  inv_x1_sg U40754 ( .A(n31114), .X(n34990) );
  inv_x1_sg U40755 ( .A(n31557), .X(n34991) );
  inv_x1_sg U40756 ( .A(n34969), .X(n34992) );
  inv_x1_sg U40757 ( .A(n31557), .X(n34993) );
  inv_x1_sg U40758 ( .A(n31205), .X(n34994) );
  inv_x1_sg U40759 ( .A(n31558), .X(n34995) );
  inv_x1_sg U40760 ( .A(n31115), .X(n34996) );
  inv_x1_sg U40761 ( .A(n31116), .X(n34997) );
  inv_x1_sg U40762 ( .A(n34993), .X(n34998) );
  inv_x1_sg U40763 ( .A(n31559), .X(n34999) );
  inv_x1_sg U40764 ( .A(n31116), .X(n35000) );
  inv_x1_sg U40765 ( .A(n34992), .X(n35001) );
  inv_x1_sg U40766 ( .A(n34990), .X(n35002) );
  inv_x1_sg U40767 ( .A(n34991), .X(n35003) );
  inv_x1_sg U40768 ( .A(n31558), .X(n35004) );
  inv_x1_sg U40769 ( .A(n34992), .X(n35005) );
  inv_x1_sg U40770 ( .A(n31115), .X(n35006) );
  inv_x1_sg U40771 ( .A(n31556), .X(n35007) );
  inv_x1_sg U40772 ( .A(n31556), .X(n35008) );
  inv_x1_sg U40773 ( .A(n34990), .X(n35009) );
  nor_x1_sg U40774 ( .A(n20893), .B(n19609), .X(n35010) );
  inv_x1_sg U40775 ( .A(n35010), .X(n35011) );
  inv_x1_sg U40776 ( .A(n31216), .X(n35012) );
  inv_x1_sg U40777 ( .A(n35594), .X(n35013) );
  inv_x1_sg U40778 ( .A(n30602), .X(n35014) );
  inv_x1_sg U40779 ( .A(n35011), .X(n35015) );
  inv_x1_sg U40780 ( .A(n35034), .X(n35016) );
  inv_x1_sg U40781 ( .A(n31574), .X(n35017) );
  inv_x1_sg U40782 ( .A(n30245), .X(n35018) );
  inv_x1_sg U40783 ( .A(n31217), .X(n35019) );
  inv_x1_sg U40784 ( .A(n35013), .X(n35020) );
  inv_x1_sg U40785 ( .A(n30239), .X(n35021) );
  inv_x1_sg U40786 ( .A(n35012), .X(n35022) );
  inv_x1_sg U40787 ( .A(n31218), .X(n35023) );
  inv_x1_sg U40788 ( .A(n30544), .X(n35024) );
  inv_x1_sg U40789 ( .A(n31218), .X(n35025) );
  inv_x1_sg U40790 ( .A(n31589), .X(n35026) );
  inv_x1_sg U40791 ( .A(n35014), .X(n35027) );
  inv_x1_sg U40792 ( .A(n31217), .X(n35028) );
  inv_x1_sg U40793 ( .A(n31217), .X(n35029) );
  inv_x1_sg U40794 ( .A(n31574), .X(n35030) );
  inv_x1_sg U40795 ( .A(n29683), .X(n35031) );
  inv_x1_sg U40796 ( .A(n35010), .X(n35032) );
  inv_x1_sg U40797 ( .A(n35010), .X(n35033) );
  inv_x1_sg U40798 ( .A(n31216), .X(n35034) );
  inv_x1_sg U40799 ( .A(n31588), .X(n35035) );
  inv_x1_sg U40800 ( .A(n35465), .X(n35036) );
  inv_x1_sg U40801 ( .A(n31112), .X(n35037) );
  inv_x1_sg U40802 ( .A(n30564), .X(n35038) );
  inv_x1_sg U40803 ( .A(n30544), .X(n35039) );
  inv_x1_sg U40804 ( .A(n35031), .X(n35040) );
  inv_x1_sg U40805 ( .A(n35032), .X(n35041) );
  inv_x1_sg U40806 ( .A(n35032), .X(n35042) );
  inv_x1_sg U40807 ( .A(n35032), .X(n35043) );
  inv_x1_sg U40808 ( .A(n35033), .X(n35044) );
  inv_x1_sg U40809 ( .A(n35465), .X(n35045) );
  inv_x1_sg U40810 ( .A(n35012), .X(n35046) );
  inv_x1_sg U40811 ( .A(n30603), .X(n35047) );
  inv_x1_sg U40812 ( .A(n31575), .X(n35048) );
  inv_x1_sg U40813 ( .A(n35465), .X(n35049) );
  inv_x1_sg U40814 ( .A(n30544), .X(n35050) );
  inv_x1_sg U40815 ( .A(n35247), .X(n35051) );
  inv_x1_sg U40816 ( .A(n35051), .X(n35052) );
  inv_x1_sg U40817 ( .A(n31608), .X(n35053) );
  inv_x1_sg U40818 ( .A(n31608), .X(n35054) );
  inv_x1_sg U40819 ( .A(n35051), .X(n35055) );
  inv_x1_sg U40820 ( .A(n35415), .X(n35056) );
  inv_x1_sg U40821 ( .A(n35056), .X(n35057) );
  inv_x1_sg U40822 ( .A(n35056), .X(n35058) );
  inv_x1_sg U40823 ( .A(n31607), .X(n35059) );
  inv_x1_sg U40824 ( .A(n31108), .X(n35060) );
  nor_x1_sg U40825 ( .A(n31885), .B(n35159), .X(n35061) );
  nor_x1_sg U40826 ( .A(n26584), .B(n35411), .X(n35062) );
  inv_x1_sg U40827 ( .A(n35061), .X(n35063) );
  inv_x1_sg U40828 ( .A(n35063), .X(n35064) );
  inv_x1_sg U40829 ( .A(n35063), .X(n35065) );
  inv_x1_sg U40830 ( .A(n35062), .X(n35066) );
  inv_x1_sg U40831 ( .A(n35066), .X(n35067) );
  inv_x1_sg U40832 ( .A(n31109), .X(n35068) );
  inv_x1_sg U40833 ( .A(n31606), .X(n35069) );
  inv_x1_sg U40834 ( .A(n35066), .X(n35070) );
  inv_x1_sg U40835 ( .A(n26590), .X(n35071) );
  inv_x1_sg U40836 ( .A(n35071), .X(n35072) );
  inv_x1_sg U40837 ( .A(n31110), .X(n35073) );
  inv_x1_sg U40838 ( .A(n31605), .X(n35074) );
  inv_x1_sg U40839 ( .A(n31110), .X(n35075) );
  inv_x1_sg U40840 ( .A(n35157), .X(n35076) );
  inv_x1_sg U40841 ( .A(n30781), .X(n35077) );
  inv_x1_sg U40842 ( .A(n35076), .X(n35078) );
  inv_x1_sg U40843 ( .A(n32052), .X(n35079) );
  inv_x1_sg U40844 ( .A(n35076), .X(n35080) );
  inv_x1_sg U40845 ( .A(n35188), .X(n35081) );
  inv_x1_sg U40846 ( .A(n35174), .X(n35082) );
  inv_x1_sg U40847 ( .A(n35180), .X(n35083) );
  inv_x1_sg U40848 ( .A(n35170), .X(n35084) );
  inv_x1_sg U40849 ( .A(n35365), .X(n35085) );
  inv_x1_sg U40850 ( .A(n35384), .X(n35086) );
  inv_x1_sg U40851 ( .A(n35174), .X(n35087) );
  inv_x1_sg U40852 ( .A(n35188), .X(n35088) );
  inv_x1_sg U40853 ( .A(n35226), .X(n35089) );
  inv_x1_sg U40854 ( .A(n35316), .X(n35090) );
  inv_x1_sg U40855 ( .A(n35180), .X(n35091) );
  inv_x1_sg U40856 ( .A(n35170), .X(n35092) );
  inv_x1_sg U40857 ( .A(n35360), .X(n35093) );
  inv_x1_sg U40858 ( .A(n35363), .X(n35094) );
  nand_x2_sg U40859 ( .A(n13359), .B(n13222), .X(n13358) );
  nand_x1_sg U40860 ( .A(n14508), .B(n13715), .X(n35095) );
  inv_x1_sg U40861 ( .A(n19606), .X(n42409) );
  inv_x1_sg U40862 ( .A(n33755), .X(n35409) );
  nor_x1_sg U40863 ( .A(n31599), .B(n31706), .X(n13619) );
  inv_x16_sg U40864 ( .A(reset), .X(n35527) );
  nor_x1_sg U40865 ( .A(n33779), .B(n34067), .X(n35677) );
  nor_x1_sg U40866 ( .A(n33614), .B(n34067), .X(n29064) );
  nand_x4_sg U40867 ( .A(n26575), .B(mask_output_filter_input_taken), .X(
        n26574) );
  nand_x16_sg U40868 ( .A(n26574), .B(n35528), .X(n35459) );
  nor_x1_sg U40869 ( .A(n31601), .B(n32220), .X(n35655) );
  nor_x1_sg U40870 ( .A(n31601), .B(n32518), .X(n35653) );
  nor_x1_sg U40871 ( .A(n32221), .B(n31663), .X(n11561) );
  inv_x1_sg U40872 ( .A(n15204), .X(n35096) );
  inv_x1_sg U40873 ( .A(n15068), .X(n35097) );
  inv_x1_sg U40874 ( .A(n12116), .X(n35098) );
  inv_x1_sg U40875 ( .A(n11635), .X(n35099) );
  inv_x1_sg U40876 ( .A(n19580), .X(n35100) );
  inv_x1_sg U40877 ( .A(n19579), .X(n35101) );
  inv_x1_sg U40878 ( .A(n13222), .X(n35102) );
  inv_x1_sg U40879 ( .A(n15045), .X(n35103) );
  inv_x1_sg U40880 ( .A(n15178), .X(n35104) );
  inv_x1_sg U40881 ( .A(n11609), .X(n35105) );
  inv_x1_sg U40882 ( .A(n11639), .X(n35106) );
  inv_x1_sg U40883 ( .A(\shifter_0/reg_w_15[19] ), .X(n35107) );
  inv_x1_sg U40884 ( .A(\shifter_0/reg_w_15[18] ), .X(n35108) );
  inv_x1_sg U40885 ( .A(\shifter_0/reg_w_15[15] ), .X(n35109) );
  inv_x1_sg U40886 ( .A(\shifter_0/reg_w_15[14] ), .X(n35110) );
  inv_x1_sg U40887 ( .A(\shifter_0/reg_w_15[13] ), .X(n35111) );
  inv_x1_sg U40888 ( .A(\shifter_0/reg_w_15[10] ), .X(n35112) );
  inv_x1_sg U40889 ( .A(\shifter_0/reg_w_15[7] ), .X(n35113) );
  inv_x1_sg U40890 ( .A(\shifter_0/reg_w_15[4] ), .X(n35114) );
  inv_x1_sg U40891 ( .A(\shifter_0/reg_w_15[1] ), .X(n35115) );
  inv_x1_sg U40892 ( .A(\shifter_0/reg_w_15[0] ), .X(n35116) );
  inv_x1_sg U40893 ( .A(\shifter_0/reg_w_3[19] ), .X(n35117) );
  inv_x1_sg U40894 ( .A(\shifter_0/reg_w_3[16] ), .X(n35118) );
  inv_x1_sg U40895 ( .A(\shifter_0/reg_w_3[15] ), .X(n35119) );
  inv_x1_sg U40896 ( .A(\shifter_0/reg_w_3[14] ), .X(n35120) );
  inv_x1_sg U40897 ( .A(\shifter_0/reg_w_3[11] ), .X(n35121) );
  inv_x1_sg U40898 ( .A(\shifter_0/reg_w_3[10] ), .X(n35122) );
  inv_x1_sg U40899 ( .A(\shifter_0/reg_w_3[7] ), .X(n35123) );
  inv_x1_sg U40900 ( .A(\shifter_0/reg_w_3[6] ), .X(n35124) );
  inv_x1_sg U40901 ( .A(\shifter_0/reg_w_3[5] ), .X(n35125) );
  inv_x1_sg U40902 ( .A(\shifter_0/reg_w_3[2] ), .X(n35126) );
  inv_x1_sg U40903 ( .A(\shifter_0/reg_w_3[1] ), .X(n35127) );
  inv_x1_sg U40904 ( .A(\shifter_0/reg_w_3[0] ), .X(n35128) );
  inv_x1_sg U40905 ( .A(\shifter_0/reg_i_15[19] ), .X(n35129) );
  inv_x1_sg U40906 ( .A(\shifter_0/reg_i_15[17] ), .X(n35130) );
  inv_x1_sg U40907 ( .A(\shifter_0/reg_i_15[15] ), .X(n35131) );
  inv_x1_sg U40908 ( .A(\shifter_0/reg_i_15[14] ), .X(n35132) );
  inv_x1_sg U40909 ( .A(\shifter_0/reg_i_15[13] ), .X(n35133) );
  inv_x1_sg U40910 ( .A(\shifter_0/reg_i_15[10] ), .X(n35134) );
  inv_x1_sg U40911 ( .A(\shifter_0/reg_i_15[7] ), .X(n35135) );
  inv_x1_sg U40912 ( .A(\shifter_0/reg_i_15[2] ), .X(n35136) );
  inv_x1_sg U40913 ( .A(\shifter_0/reg_i_15[1] ), .X(n35137) );
  inv_x1_sg U40914 ( .A(\shifter_0/reg_i_15[0] ), .X(n35138) );
  inv_x1_sg U40915 ( .A(\shifter_0/reg_i_7[18] ), .X(n35139) );
  inv_x1_sg U40916 ( .A(\shifter_0/reg_i_7[17] ), .X(n35140) );
  inv_x1_sg U40917 ( .A(\shifter_0/reg_i_7[2] ), .X(n35141) );
  inv_x1_sg U40918 ( .A(\shifter_0/reg_i_3[19] ), .X(n35142) );
  inv_x1_sg U40919 ( .A(\shifter_0/reg_i_3[16] ), .X(n35143) );
  inv_x1_sg U40920 ( .A(\shifter_0/reg_i_3[15] ), .X(n35144) );
  inv_x1_sg U40921 ( .A(\shifter_0/reg_i_3[14] ), .X(n35145) );
  inv_x1_sg U40922 ( .A(\shifter_0/reg_i_3[11] ), .X(n35146) );
  inv_x1_sg U40923 ( .A(\shifter_0/reg_i_3[10] ), .X(n35147) );
  inv_x1_sg U40924 ( .A(\shifter_0/reg_i_3[7] ), .X(n35148) );
  inv_x1_sg U40925 ( .A(\shifter_0/reg_i_3[6] ), .X(n35149) );
  inv_x1_sg U40926 ( .A(\shifter_0/reg_i_3[5] ), .X(n35150) );
  inv_x1_sg U40927 ( .A(\shifter_0/reg_i_3[2] ), .X(n35151) );
  inv_x1_sg U40928 ( .A(\shifter_0/reg_i_3[1] ), .X(n35152) );
  inv_x1_sg U40929 ( .A(\shifter_0/reg_i_3[0] ), .X(n35153) );
  inv_x1_sg U40930 ( .A(\filter_0/N13 ), .X(n35154) );
  inv_x1_sg U40931 ( .A(n35309), .X(n35155) );
  inv_x1_sg U40932 ( .A(n35312), .X(n35156) );
  inv_x1_sg U40933 ( .A(n26194), .X(n35157) );
  inv_x1_sg U40934 ( .A(\shifter_0/pointer[2] ), .X(n35158) );
  inv_x1_sg U40935 ( .A(n32007), .X(n35159) );
  inv_x1_sg U40936 ( .A(n35322), .X(n35160) );
  inv_x1_sg U40937 ( .A(n35322), .X(n35161) );
  inv_x1_sg U40938 ( .A(n35323), .X(n35162) );
  inv_x1_sg U40939 ( .A(n35323), .X(n35163) );
  inv_x1_sg U40940 ( .A(n35324), .X(n35164) );
  inv_x1_sg U40941 ( .A(n35324), .X(n35165) );
  inv_x1_sg U40942 ( .A(n30751), .X(n35166) );
  inv_x1_sg U40943 ( .A(n35166), .X(n35167) );
  inv_x1_sg U40944 ( .A(n32852), .X(n35168) );
  inv_x1_sg U40945 ( .A(n35168), .X(n35169) );
  inv_x1_sg U40946 ( .A(n32444), .X(n35170) );
  inv_x1_sg U40947 ( .A(n35170), .X(n35171) );
  inv_x1_sg U40948 ( .A(n32850), .X(n35172) );
  inv_x1_sg U40949 ( .A(n35172), .X(n35173) );
  inv_x1_sg U40950 ( .A(n35683), .X(n35174) );
  inv_x1_sg U40951 ( .A(n35174), .X(n35175) );
  inv_x1_sg U40952 ( .A(n32448), .X(n35176) );
  inv_x1_sg U40953 ( .A(n35176), .X(n35177) );
  inv_x1_sg U40954 ( .A(n34655), .X(n35178) );
  inv_x1_sg U40955 ( .A(n35178), .X(n35179) );
  inv_x1_sg U40956 ( .A(n34657), .X(n35180) );
  inv_x1_sg U40957 ( .A(n35180), .X(n35181) );
  inv_x1_sg U40958 ( .A(n35363), .X(n35182) );
  inv_x1_sg U40959 ( .A(n35363), .X(n35183) );
  inv_x1_sg U40960 ( .A(n35364), .X(n35184) );
  inv_x1_sg U40961 ( .A(n35364), .X(n35185) );
  inv_x1_sg U40962 ( .A(n35365), .X(n35186) );
  inv_x1_sg U40963 ( .A(n35365), .X(n35187) );
  inv_x1_sg U40964 ( .A(n30177), .X(n35188) );
  inv_x1_sg U40965 ( .A(n35188), .X(n35189) );
  inv_x1_sg U40966 ( .A(n32446), .X(n35190) );
  inv_x1_sg U40967 ( .A(n35190), .X(n35191) );
  inv_x1_sg U40968 ( .A(n32447), .X(n35192) );
  inv_x1_sg U40969 ( .A(n35192), .X(n35193) );
  inv_x1_sg U40970 ( .A(n35372), .X(n35194) );
  inv_x1_sg U40971 ( .A(n35372), .X(n35195) );
  inv_x1_sg U40972 ( .A(n32851), .X(n35196) );
  inv_x1_sg U40973 ( .A(n35196), .X(n35197) );
  inv_x1_sg U40974 ( .A(n35373), .X(n35198) );
  inv_x1_sg U40975 ( .A(n35373), .X(n35199) );
  inv_x1_sg U40976 ( .A(n35381), .X(n35200) );
  inv_x1_sg U40977 ( .A(n35381), .X(n35201) );
  inv_x1_sg U40978 ( .A(n35382), .X(n35202) );
  inv_x1_sg U40979 ( .A(n35382), .X(n35203) );
  inv_x1_sg U40980 ( .A(n35383), .X(n35204) );
  inv_x1_sg U40981 ( .A(n35383), .X(n35205) );
  inv_x1_sg U40982 ( .A(n35384), .X(n35206) );
  inv_x1_sg U40983 ( .A(n35384), .X(n35207) );
  inv_x1_sg U40984 ( .A(n35385), .X(n35208) );
  inv_x1_sg U40985 ( .A(n35385), .X(n35209) );
  inv_x1_sg U40986 ( .A(n35386), .X(n35210) );
  inv_x1_sg U40987 ( .A(n35386), .X(n35211) );
  inv_x1_sg U40988 ( .A(n35387), .X(n35212) );
  inv_x1_sg U40989 ( .A(n35387), .X(n35213) );
  inv_x1_sg U40990 ( .A(n35388), .X(n35214) );
  inv_x1_sg U40991 ( .A(n35388), .X(n35215) );
  inv_x1_sg U40992 ( .A(n35389), .X(n35216) );
  inv_x1_sg U40993 ( .A(n35389), .X(n35217) );
  inv_x1_sg U40994 ( .A(n35390), .X(n35218) );
  inv_x1_sg U40995 ( .A(n35390), .X(n35219) );
  inv_x1_sg U40996 ( .A(n35391), .X(n35220) );
  inv_x1_sg U40997 ( .A(n35391), .X(n35221) );
  inv_x1_sg U40998 ( .A(n35392), .X(n35222) );
  inv_x1_sg U40999 ( .A(n35392), .X(n35223) );
  inv_x1_sg U41000 ( .A(n35393), .X(n35224) );
  inv_x1_sg U41001 ( .A(n35393), .X(n35225) );
  inv_x1_sg U41002 ( .A(n34658), .X(n35226) );
  inv_x1_sg U41003 ( .A(n35226), .X(n35227) );
  inv_x1_sg U41004 ( .A(n35226), .X(n35228) );
  inv_x1_sg U41005 ( .A(n35400), .X(n35229) );
  inv_x1_sg U41006 ( .A(n35400), .X(n35230) );
  inv_x1_sg U41007 ( .A(n35401), .X(n35231) );
  inv_x1_sg U41008 ( .A(n35401), .X(n35232) );
  inv_x1_sg U41009 ( .A(n35401), .X(n35233) );
  inv_x1_sg U41010 ( .A(n35401), .X(n35234) );
  inv_x1_sg U41011 ( .A(n32448), .X(n35235) );
  inv_x1_sg U41012 ( .A(n35235), .X(n35236) );
  inv_x1_sg U41013 ( .A(n35235), .X(n35237) );
  inv_x1_sg U41014 ( .A(n34657), .X(n35238) );
  inv_x1_sg U41015 ( .A(n35238), .X(n35239) );
  inv_x1_sg U41016 ( .A(n35238), .X(n35240) );
  inv_x1_sg U41017 ( .A(n33726), .X(n35241) );
  inv_x1_sg U41018 ( .A(n33722), .X(n35242) );
  inv_x1_sg U41019 ( .A(n33735), .X(n35243) );
  inv_x1_sg U41020 ( .A(n33743), .X(n35244) );
  inv_x1_sg U41021 ( .A(n33739), .X(n35245) );
  inv_x1_sg U41022 ( .A(n33750), .X(n35246) );
  inv_x1_sg U41023 ( .A(n23629), .X(n35247) );
  inv_x1_sg U41024 ( .A(n35684), .X(n35248) );
  inv_x1_sg U41025 ( .A(n29620), .X(n35249) );
  inv_x1_sg U41026 ( .A(n28921), .X(n35250) );
  inv_x1_sg U41027 ( .A(shifter_state[0]), .X(n35251) );
  inv_x1_sg U41028 ( .A(n13098), .X(n35252) );
  inv_x1_sg U41029 ( .A(\shifter_0/reg_i_15[18] ), .X(n35253) );
  inv_x1_sg U41030 ( .A(\shifter_0/reg_i_15[4] ), .X(n35254) );
  inv_x1_sg U41031 ( .A(\shifter_0/reg_i_7[4] ), .X(n35255) );
  inv_x1_sg U41032 ( .A(\filter_0/w_pointer[2] ), .X(n35256) );
  inv_x1_sg U41033 ( .A(\filter_0/i_pointer[0] ), .X(n35257) );
  inv_x1_sg U41034 ( .A(\filter_0/i_pointer[2] ), .X(n35258) );
  inv_x1_sg U41035 ( .A(n33711), .X(n35259) );
  inv_x1_sg U41036 ( .A(n33745), .X(n35260) );
  inv_x1_sg U41037 ( .A(n33728), .X(n35261) );
  inv_x1_sg U41038 ( .A(n34440), .X(n35262) );
  inv_x1_sg U41039 ( .A(\shifter_0/pointer[3] ), .X(n35263) );
  inv_x1_sg U41040 ( .A(n35485), .X(n35264) );
  inv_x1_sg U41041 ( .A(n32008), .X(n35265) );
  inv_x1_sg U41042 ( .A(n21303), .X(n35266) );
  inv_x1_sg U41043 ( .A(\shifter_0/i_pointer[1] ), .X(n35267) );
  inv_x1_sg U41044 ( .A(\filter_0/N14 ), .X(n35268) );
  inv_x1_sg U41045 ( .A(\filter_0/i_pointer[1] ), .X(n35269) );
  inv_x1_sg U41046 ( .A(n28318), .X(n35270) );
  inv_x1_sg U41047 ( .A(\shifter_0/w_pointer[1] ), .X(n35271) );
  inv_x1_sg U41048 ( .A(n31657), .X(n35272) );
  inv_x1_sg U41049 ( .A(n31655), .X(n35273) );
  inv_x1_sg U41050 ( .A(n30020), .X(n35274) );
  inv_x1_sg U41051 ( .A(n35312), .X(n35275) );
  inv_x1_sg U41052 ( .A(n32290), .X(n35276) );
  inv_x1_sg U41053 ( .A(n35276), .X(n35277) );
  inv_x1_sg U41054 ( .A(n19600), .X(n35278) );
  inv_x1_sg U41055 ( .A(\shifter_0/w_pointer[2] ), .X(n35279) );
  inv_x1_sg U41056 ( .A(\shifter_0/i_pointer[2] ), .X(n35280) );
  inv_x1_sg U41057 ( .A(n35309), .X(n35281) );
  inv_x1_sg U41058 ( .A(n35298), .X(n35282) );
  inv_x1_sg U41059 ( .A(n35295), .X(n35283) );
  inv_x1_sg U41060 ( .A(n32854), .X(n35284) );
  inv_x1_sg U41061 ( .A(n35284), .X(n35285) );
  inv_x1_sg U41062 ( .A(n35284), .X(n35286) );
  inv_x1_sg U41063 ( .A(n35298), .X(n35287) );
  inv_x1_sg U41064 ( .A(n35276), .X(n35288) );
  inv_x1_sg U41065 ( .A(n35295), .X(n35289) );
  inv_x1_sg U41066 ( .A(n32320), .X(n35290) );
  inv_x1_sg U41067 ( .A(n35290), .X(n35291) );
  inv_x1_sg U41068 ( .A(n35290), .X(n35292) );
  inv_x1_sg U41069 ( .A(n35290), .X(n35293) );
  inv_x1_sg U41070 ( .A(n35284), .X(n35294) );
  inv_x1_sg U41071 ( .A(n32774), .X(n35295) );
  inv_x1_sg U41072 ( .A(n35295), .X(n35296) );
  inv_x1_sg U41073 ( .A(n35295), .X(n35297) );
  inv_x1_sg U41074 ( .A(n32335), .X(n35298) );
  inv_x1_sg U41075 ( .A(n35298), .X(n35299) );
  inv_x1_sg U41076 ( .A(n35298), .X(n35300) );
  inv_x1_sg U41077 ( .A(\shifter_0/i_pointer[0] ), .X(n35301) );
  inv_x1_sg U41078 ( .A(n31882), .X(n35302) );
  nand_x2_sg U41079 ( .A(n11764), .B(n11765), .X(n35600) );
  inv_x1_sg U41080 ( .A(\shifter_0/w_pointer[0] ), .X(n35303) );
  inv_x1_sg U41081 ( .A(n32004), .X(n35304) );
  inv_x1_sg U41082 ( .A(n31879), .X(n35305) );
  inv_x1_sg U41083 ( .A(n32000), .X(n35306) );
  inv_x1_sg U41084 ( .A(n20968), .X(n35307) );
  inv_x1_sg U41085 ( .A(n31886), .X(n35308) );
  inv_x1_sg U41086 ( .A(n32383), .X(n35309) );
  inv_x1_sg U41087 ( .A(n35309), .X(n35310) );
  inv_x1_sg U41088 ( .A(n35309), .X(n35311) );
  inv_x1_sg U41089 ( .A(n31924), .X(n35312) );
  inv_x1_sg U41090 ( .A(n35312), .X(n35313) );
  inv_x1_sg U41091 ( .A(n33956), .X(n35314) );
  inv_x1_sg U41092 ( .A(n32906), .X(n35315) );
  inv_x1_sg U41093 ( .A(n29759), .X(n35316) );
  inv_x1_sg U41094 ( .A(n35316), .X(n35317) );
  inv_x1_sg U41095 ( .A(n35316), .X(n35318) );
  inv_x1_sg U41096 ( .A(n34658), .X(n35319) );
  inv_x1_sg U41097 ( .A(n35319), .X(n35320) );
  inv_x1_sg U41098 ( .A(n35319), .X(n35321) );
  inv_x1_sg U41099 ( .A(n32447), .X(n35322) );
  inv_x1_sg U41100 ( .A(n32851), .X(n35323) );
  inv_x1_sg U41101 ( .A(n34655), .X(n35324) );
  inv_x1_sg U41102 ( .A(n32447), .X(n35325) );
  inv_x1_sg U41103 ( .A(n35325), .X(n35326) );
  inv_x1_sg U41104 ( .A(n35325), .X(n35327) );
  inv_x1_sg U41105 ( .A(n32852), .X(n35328) );
  inv_x1_sg U41106 ( .A(n35328), .X(n35329) );
  inv_x1_sg U41107 ( .A(n35328), .X(n35330) );
  inv_x1_sg U41108 ( .A(n29759), .X(n35331) );
  inv_x1_sg U41109 ( .A(n35331), .X(n35332) );
  inv_x1_sg U41110 ( .A(n35331), .X(n35333) );
  inv_x1_sg U41111 ( .A(n32851), .X(n35334) );
  inv_x1_sg U41112 ( .A(n35334), .X(n35335) );
  inv_x1_sg U41113 ( .A(n35334), .X(n35336) );
  inv_x1_sg U41114 ( .A(n32448), .X(n35337) );
  inv_x1_sg U41115 ( .A(n35337), .X(n35338) );
  inv_x1_sg U41116 ( .A(n35337), .X(n35339) );
  inv_x1_sg U41117 ( .A(n30752), .X(n35340) );
  inv_x1_sg U41118 ( .A(n35340), .X(n35341) );
  inv_x1_sg U41119 ( .A(n35340), .X(n35342) );
  inv_x1_sg U41120 ( .A(n34656), .X(n35343) );
  inv_x1_sg U41121 ( .A(n35343), .X(n35344) );
  inv_x1_sg U41122 ( .A(n35343), .X(n35345) );
  inv_x1_sg U41123 ( .A(n32850), .X(n35346) );
  inv_x1_sg U41124 ( .A(n35346), .X(n35347) );
  inv_x1_sg U41125 ( .A(n35346), .X(n35348) );
  inv_x1_sg U41126 ( .A(n29760), .X(n35349) );
  inv_x1_sg U41127 ( .A(n35349), .X(n35350) );
  inv_x1_sg U41128 ( .A(n35349), .X(n35351) );
  inv_x1_sg U41129 ( .A(n32849), .X(n35352) );
  inv_x1_sg U41130 ( .A(n35352), .X(n35353) );
  inv_x1_sg U41131 ( .A(n32849), .X(n35354) );
  inv_x1_sg U41132 ( .A(n35354), .X(n35355) );
  inv_x1_sg U41133 ( .A(n35354), .X(n35356) );
  inv_x1_sg U41134 ( .A(n32447), .X(n35357) );
  inv_x1_sg U41135 ( .A(n35357), .X(n35358) );
  inv_x1_sg U41136 ( .A(n35357), .X(n35359) );
  inv_x1_sg U41137 ( .A(n34658), .X(n35360) );
  inv_x1_sg U41138 ( .A(n35360), .X(n35361) );
  inv_x1_sg U41139 ( .A(n35360), .X(n35362) );
  inv_x1_sg U41140 ( .A(n34657), .X(n35363) );
  inv_x1_sg U41141 ( .A(n29759), .X(n35364) );
  inv_x1_sg U41142 ( .A(n32444), .X(n35365) );
  inv_x1_sg U41143 ( .A(n32850), .X(n35366) );
  inv_x1_sg U41144 ( .A(n35366), .X(n35367) );
  inv_x1_sg U41145 ( .A(n35366), .X(n35368) );
  inv_x1_sg U41146 ( .A(n30717), .X(n35369) );
  inv_x1_sg U41147 ( .A(n35369), .X(n35370) );
  inv_x1_sg U41148 ( .A(n35369), .X(n35371) );
  inv_x1_sg U41149 ( .A(n32851), .X(n35372) );
  inv_x1_sg U41150 ( .A(n32448), .X(n35373) );
  inv_x1_sg U41151 ( .A(n32911), .X(n35374) );
  inv_x1_sg U41152 ( .A(n29760), .X(n35375) );
  inv_x1_sg U41153 ( .A(n35375), .X(n35376) );
  inv_x1_sg U41154 ( .A(n35375), .X(n35377) );
  inv_x1_sg U41155 ( .A(n30594), .X(n35378) );
  inv_x1_sg U41156 ( .A(n35378), .X(n35379) );
  inv_x1_sg U41157 ( .A(n35378), .X(n35380) );
  inv_x1_sg U41158 ( .A(n30752), .X(n35381) );
  inv_x1_sg U41159 ( .A(n32850), .X(n35382) );
  inv_x1_sg U41160 ( .A(n34656), .X(n35383) );
  inv_x1_sg U41161 ( .A(n29759), .X(n35384) );
  inv_x1_sg U41162 ( .A(n32444), .X(n35385) );
  inv_x1_sg U41163 ( .A(n30751), .X(n35386) );
  inv_x1_sg U41164 ( .A(n34658), .X(n35387) );
  inv_x1_sg U41165 ( .A(n32852), .X(n35388) );
  inv_x1_sg U41166 ( .A(n32449), .X(n35389) );
  inv_x1_sg U41167 ( .A(n32446), .X(n35390) );
  inv_x1_sg U41168 ( .A(n32849), .X(n35391) );
  inv_x1_sg U41169 ( .A(n32852), .X(n35392) );
  inv_x1_sg U41170 ( .A(n34656), .X(n35393) );
  inv_x1_sg U41171 ( .A(n34657), .X(n35394) );
  inv_x1_sg U41172 ( .A(n35394), .X(n35395) );
  inv_x1_sg U41173 ( .A(n35394), .X(n35396) );
  inv_x1_sg U41174 ( .A(n32446), .X(n35397) );
  inv_x1_sg U41175 ( .A(n35397), .X(n35398) );
  inv_x1_sg U41176 ( .A(n35397), .X(n35399) );
  inv_x1_sg U41177 ( .A(n32449), .X(n35400) );
  inv_x1_sg U41178 ( .A(n32446), .X(n35401) );
  inv_x1_sg U41179 ( .A(n32449), .X(n35402) );
  inv_x1_sg U41180 ( .A(n35402), .X(n35403) );
  inv_x1_sg U41181 ( .A(n35402), .X(n35404) );
  inv_x1_sg U41182 ( .A(n33525), .X(n35405) );
  inv_x1_sg U41183 ( .A(n33637), .X(n35406) );
  inv_x1_sg U41184 ( .A(n33718), .X(n35407) );
  inv_x1_sg U41185 ( .A(n33798), .X(n35408) );
  inv_x1_sg U41186 ( .A(n33760), .X(n35410) );
  inv_x1_sg U41187 ( .A(n35485), .X(n35411) );
  inv_x1_sg U41188 ( .A(n32007), .X(n35412) );
  inv_x1_sg U41189 ( .A(n14496), .X(n35413) );
  inv_x1_sg U41190 ( .A(n14497), .X(n35414) );
  inv_x1_sg U41191 ( .A(n35455), .X(n35415) );
  inv_x1_sg U41192 ( .A(\shifter_0/pointer[1] ), .X(n35416) );
  inv_x1_sg U41193 ( .A(\shifter_0/pointer[0] ), .X(n35417) );
  nand_x1_sg U41194 ( .A(n32425), .B(n35103), .X(n28449) );
  inv_x16_sg U41195 ( .A(reset), .X(n35528) );
  nor_x1_sg U41196 ( .A(n21014), .B(n21015), .X(n21013) );
  nor_x1_sg U41197 ( .A(n13837), .B(n13838), .X(n13836) );
  nor_x1_sg U41198 ( .A(n13800), .B(n13801), .X(n13799) );
  nor_x1_sg U41199 ( .A(n13899), .B(n13900), .X(n13898) );
  nor_x1_sg U41200 ( .A(n13868), .B(n13869), .X(n13867) );
  nor_x1_sg U41201 ( .A(n13961), .B(n13962), .X(n13960) );
  nor_x1_sg U41202 ( .A(n13930), .B(n13931), .X(n13929) );
  nor_x1_sg U41203 ( .A(n14023), .B(n14024), .X(n14022) );
  nor_x1_sg U41204 ( .A(n13992), .B(n13993), .X(n13991) );
  nor_x1_sg U41205 ( .A(n14085), .B(n14086), .X(n14084) );
  nor_x1_sg U41206 ( .A(n14054), .B(n14055), .X(n14053) );
  nor_x1_sg U41207 ( .A(n14147), .B(n14148), .X(n14146) );
  nor_x1_sg U41208 ( .A(n14116), .B(n14117), .X(n14115) );
  nor_x1_sg U41209 ( .A(n14209), .B(n14210), .X(n14208) );
  nor_x1_sg U41210 ( .A(n14178), .B(n14179), .X(n14177) );
  nor_x1_sg U41211 ( .A(n14271), .B(n14272), .X(n14270) );
  nor_x1_sg U41212 ( .A(n14240), .B(n14241), .X(n14239) );
  nor_x1_sg U41213 ( .A(n14333), .B(n14334), .X(n14332) );
  nor_x1_sg U41214 ( .A(n14302), .B(n14303), .X(n14301) );
  nor_x1_sg U41215 ( .A(n14395), .B(n14396), .X(n14394) );
  nor_x1_sg U41216 ( .A(n14364), .B(n14365), .X(n14363) );
  nor_x1_sg U41217 ( .A(n14458), .B(n14459), .X(n14457) );
  nor_x1_sg U41218 ( .A(n14427), .B(n14428), .X(n14426) );
  nor_x1_sg U41219 ( .A(n14584), .B(n14585), .X(n14583) );
  nor_x1_sg U41220 ( .A(n14522), .B(n14523), .X(n14521) );
  nor_x1_sg U41221 ( .A(n14646), .B(n14647), .X(n14645) );
  nor_x1_sg U41222 ( .A(n14615), .B(n14616), .X(n14614) );
  nor_x1_sg U41223 ( .A(n14708), .B(n14709), .X(n14707) );
  nor_x1_sg U41224 ( .A(n14677), .B(n14678), .X(n14676) );
  nor_x1_sg U41225 ( .A(n14770), .B(n14771), .X(n14769) );
  nor_x1_sg U41226 ( .A(n14739), .B(n14740), .X(n14738) );
  nor_x1_sg U41227 ( .A(n14832), .B(n14833), .X(n14831) );
  nor_x1_sg U41228 ( .A(n14801), .B(n14802), .X(n14800) );
  nor_x1_sg U41229 ( .A(n14894), .B(n14895), .X(n14893) );
  nor_x1_sg U41230 ( .A(n14863), .B(n14864), .X(n14862) );
  nor_x1_sg U41231 ( .A(n15018), .B(n15019), .X(n15017) );
  nor_x1_sg U41232 ( .A(n14925), .B(n14926), .X(n14924) );
  nand_x2_sg U41233 ( .A(n11766), .B(n31659), .X(n11765) );
  nor_x1_sg U41234 ( .A(n20985), .B(n20986), .X(n20915) );
  nor_x1_sg U41235 ( .A(n20973), .B(n20974), .X(n20928) );
  nor_x1_sg U41236 ( .A(n20962), .B(n20963), .X(n20932) );
  nor_x1_sg U41237 ( .A(n20993), .B(n20994), .X(n20921) );
  nor_x1_sg U41238 ( .A(n21566), .B(n21567), .X(n21360) );
  nor_x1_sg U41239 ( .A(n21472), .B(n21473), .X(n21356) );
  nor_x1_sg U41240 ( .A(n21379), .B(n21380), .X(n21355) );
  nor_x1_sg U41241 ( .A(n21659), .B(n21660), .X(n21359) );
  nor_x1_sg U41242 ( .A(n33506), .B(n34067), .X(n35666) );
  nor_x1_sg U41243 ( .A(n33590), .B(n34065), .X(n35667) );
  nor_x1_sg U41244 ( .A(n33582), .B(n34068), .X(n35669) );
  nand_x4_sg U41245 ( .A(n21305), .B(n21306), .X(n21304) );
  nand_x1_sg U41246 ( .A(n30522), .B(n35510), .X(n15053) );
  nand_x4_sg U41247 ( .A(n15034), .B(n30527), .X(n35483) );
  nand_x4_sg U41248 ( .A(n21744), .B(n19606), .X(n21303) );
  nand_x4_sg U41249 ( .A(n15355), .B(n31594), .X(n15101) );
  nand_x1_sg U41250 ( .A(n13218), .B(n13219), .X(n13104) );
  nand_x1_sg U41251 ( .A(n12522), .B(n12523), .X(n12438) );
  nand_x4_sg U41252 ( .A(n11634), .B(n30534), .X(n35458) );
  nand_x4_sg U41253 ( .A(n15356), .B(\filter_0/N14 ), .X(n29669) );
  nand_x4_sg U41254 ( .A(n13606), .B(n13607), .X(n35638) );
  nand_x4_sg U41255 ( .A(n11662), .B(n11663), .X(n11641) );
  nand_x1_sg U41256 ( .A(n35582), .B(n15215), .X(n15204) );
  nand_x4_sg U41257 ( .A(n11557), .B(n11558), .X(n11536) );
  nand_x4_sg U41258 ( .A(n11607), .B(n11608), .X(n11586) );
  nand_x4_sg U41259 ( .A(n11583), .B(n11584), .X(n11562) );
  nand_x1_sg U41260 ( .A(n11792), .B(n11793), .X(n11791) );
  nand_x1_sg U41261 ( .A(n11738), .B(n11739), .X(n11737) );
  nand_x1_sg U41262 ( .A(n11711), .B(n11712), .X(n11710) );
  nand_x1_sg U41263 ( .A(n12832), .B(n35507), .X(n35622) );
  nand_x1_sg U41264 ( .A(n20894), .B(n35551), .X(n19609) );
  nand_x1_sg U41265 ( .A(n32424), .B(n29576), .X(n29018) );
  nand_x1_sg U41266 ( .A(n32427), .B(n28966), .X(n28448) );
  nand_x1_sg U41267 ( .A(n35582), .B(n15079), .X(n15068) );
  nand_x1_sg U41268 ( .A(n32426), .B(n29532), .X(n29061) );
  nor_x1_sg U41269 ( .A(n32508), .B(n32939), .X(n19591) );
  nand_x1_sg U41270 ( .A(n32425), .B(n29488), .X(n29104) );
  nand_x1_sg U41271 ( .A(n32424), .B(n28877), .X(n28319) );
  inv_x1_sg U41272 ( .A(n15051), .X(n42402) );
  inv_x1_sg U41273 ( .A(n15185), .X(n35530) );
  nand_x2_sg U41274 ( .A(n15186), .B(n31661), .X(n15185) );
  inv_x1_sg U41275 ( .A(n15191), .X(n35553) );
  nand_x2_sg U41276 ( .A(n15192), .B(n31661), .X(n15191) );
  inv_x1_sg U41277 ( .A(n32007), .X(n35466) );
  inv_x1_sg U41278 ( .A(n35628), .X(n35418) );
  nor_x1_sg U41279 ( .A(n21093), .B(n21094), .X(n21092) );
  nor_x1_sg U41280 ( .A(n21070), .B(n21071), .X(n21069) );
  nor_x1_sg U41281 ( .A(n21052), .B(n21053), .X(n21051) );
  nor_x1_sg U41282 ( .A(n21032), .B(n21033), .X(n21031) );
  nor_x1_sg U41283 ( .A(n21170), .B(n21171), .X(n21169) );
  nor_x1_sg U41284 ( .A(n21149), .B(n21150), .X(n21148) );
  nor_x1_sg U41285 ( .A(n21131), .B(n21132), .X(n21130) );
  nor_x1_sg U41286 ( .A(n21111), .B(n21112), .X(n21110) );
  nor_x1_sg U41287 ( .A(n21249), .B(n21250), .X(n21248) );
  nor_x1_sg U41288 ( .A(n21231), .B(n21232), .X(n21230) );
  nor_x1_sg U41289 ( .A(n21209), .B(n21210), .X(n21208) );
  nor_x1_sg U41290 ( .A(n21191), .B(n21192), .X(n21190) );
  nor_x1_sg U41291 ( .A(n21316), .B(n21317), .X(n21305) );
  nor_x1_sg U41292 ( .A(n21307), .B(n21308), .X(n21306) );
  nor_x1_sg U41293 ( .A(n21287), .B(n21288), .X(n21286) );
  nor_x1_sg U41294 ( .A(n21269), .B(n21270), .X(n21268) );
  nor_x1_sg U41295 ( .A(n21453), .B(n21454), .X(n21452) );
  nor_x1_sg U41296 ( .A(n21435), .B(n21436), .X(n21434) );
  nor_x1_sg U41297 ( .A(n21415), .B(n21416), .X(n21414) );
  nor_x1_sg U41298 ( .A(n21397), .B(n21398), .X(n21396) );
  nor_x1_sg U41299 ( .A(n21545), .B(n21546), .X(n21544) );
  nor_x1_sg U41300 ( .A(n21527), .B(n21528), .X(n21526) );
  nor_x1_sg U41301 ( .A(n21507), .B(n21508), .X(n21506) );
  nor_x1_sg U41302 ( .A(n21489), .B(n21490), .X(n21488) );
  nor_x1_sg U41303 ( .A(n21640), .B(n21641), .X(n21639) );
  nor_x1_sg U41304 ( .A(n21622), .B(n21623), .X(n21621) );
  nor_x1_sg U41305 ( .A(n21602), .B(n21603), .X(n21601) );
  nor_x1_sg U41306 ( .A(n21584), .B(n21585), .X(n21583) );
  nor_x1_sg U41307 ( .A(n21736), .B(n21737), .X(n21725) );
  nor_x1_sg U41308 ( .A(n21709), .B(n21710), .X(n21708) );
  nor_x1_sg U41309 ( .A(n21691), .B(n21692), .X(n21690) );
  nor_x1_sg U41310 ( .A(n21670), .B(n21671), .X(n21669) );
  nor_x1_sg U41311 ( .A(n14988), .B(n14989), .X(n14987) );
  nor_x1_sg U41312 ( .A(n14957), .B(n14958), .X(n14956) );
  nor_x1_sg U41313 ( .A(n14554), .B(n14555), .X(n14553) );
  nor_x1_sg U41314 ( .A(n14490), .B(n14491), .X(n14489) );
  inv_x1_sg U41315 ( .A(n12611), .X(n35419) );
  nand_x4_sg U41316 ( .A(n23632), .B(input_ready), .X(n23631) );
  nand_x1_sg U41317 ( .A(n12958), .B(n12959), .X(n35420) );
  nand_x1_sg U41318 ( .A(n12934), .B(n12935), .X(n35421) );
  nand_x1_sg U41319 ( .A(n12940), .B(n12941), .X(n35422) );
  nand_x1_sg U41320 ( .A(n12946), .B(n12947), .X(n35423) );
  nand_x1_sg U41321 ( .A(n12952), .B(n12953), .X(n35424) );
  nand_x1_sg U41322 ( .A(n12910), .B(n12911), .X(n35425) );
  nand_x1_sg U41323 ( .A(n12916), .B(n12917), .X(n35426) );
  nand_x1_sg U41324 ( .A(n12922), .B(n12923), .X(n35427) );
  nand_x1_sg U41325 ( .A(n12928), .B(n12929), .X(n35428) );
  nand_x1_sg U41326 ( .A(n12886), .B(n12887), .X(n35429) );
  nand_x1_sg U41327 ( .A(n12892), .B(n12893), .X(n35430) );
  nand_x1_sg U41328 ( .A(n12898), .B(n12899), .X(n35431) );
  nand_x1_sg U41329 ( .A(n12904), .B(n12905), .X(n35432) );
  nand_x1_sg U41330 ( .A(n12856), .B(n12857), .X(n35433) );
  nand_x1_sg U41331 ( .A(n12868), .B(n12869), .X(n35434) );
  nand_x1_sg U41332 ( .A(n12874), .B(n12875), .X(n35435) );
  nand_x1_sg U41333 ( .A(n12880), .B(n12881), .X(n35436) );
  nand_x1_sg U41334 ( .A(n12822), .B(n12823), .X(n35437) );
  nand_x1_sg U41335 ( .A(n12828), .B(n12829), .X(n35438) );
  nand_x1_sg U41336 ( .A(n12844), .B(n12845), .X(n35439) );
  nand_x1_sg U41337 ( .A(n12850), .B(n12851), .X(n35440) );
  nand_x1_sg U41338 ( .A(n12792), .B(n12793), .X(n35441) );
  nand_x1_sg U41339 ( .A(n12804), .B(n12805), .X(n35442) );
  nand_x1_sg U41340 ( .A(n12810), .B(n12811), .X(n35443) );
  nand_x1_sg U41341 ( .A(n12816), .B(n12817), .X(n35444) );
  nand_x1_sg U41342 ( .A(n12762), .B(n12763), .X(n35445) );
  nand_x1_sg U41343 ( .A(n12768), .B(n12769), .X(n35446) );
  nand_x1_sg U41344 ( .A(n12774), .B(n12775), .X(n35447) );
  nand_x1_sg U41345 ( .A(n12780), .B(n12781), .X(n35448) );
  nand_x1_sg U41346 ( .A(n12713), .B(n12714), .X(n35449) );
  nand_x1_sg U41347 ( .A(n12726), .B(n12727), .X(n35450) );
  nand_x1_sg U41348 ( .A(n12744), .B(n12745), .X(n35451) );
  nand_x1_sg U41349 ( .A(n12750), .B(n12751), .X(n35452) );
  nand_x1_sg U41350 ( .A(n14546), .B(n14547), .X(n35453) );
  inv_x1_sg U41351 ( .A(n26347), .X(n35454) );
  inv_x1_sg U41352 ( .A(n32108), .X(n35456) );
  inv_x1_sg U41353 ( .A(state[1]), .X(n35457) );
  inv_x1_sg U41354 ( .A(n32503), .X(n35460) );
  inv_x1_sg U41355 ( .A(n11710), .X(n35461) );
  inv_x1_sg U41356 ( .A(n11791), .X(n35462) );
  inv_x1_sg U41357 ( .A(n19594), .X(n35463) );
  inv_x1_sg U41358 ( .A(n11737), .X(n35464) );
  inv_x1_sg U41359 ( .A(n35048), .X(n35465) );
  nand_x1_sg U41360 ( .A(n14973), .B(n41520), .X(n35467) );
  nand_x1_sg U41361 ( .A(n14787), .B(n13750), .X(n35468) );
  nand_x1_sg U41362 ( .A(n14942), .B(n41521), .X(n35469) );
  nand_x1_sg U41363 ( .A(n14694), .B(n13738), .X(n35470) );
  nand_x1_sg U41364 ( .A(n14539), .B(n41522), .X(n35471) );
  nand_x1_sg U41365 ( .A(n14319), .B(n13686), .X(n35472) );
  nand_x1_sg U41366 ( .A(n14071), .B(n13654), .X(n35473) );
  nand_x1_sg U41367 ( .A(n13568), .B(n41326), .X(n35474) );
  nand_x1_sg U41368 ( .A(n13562), .B(n41327), .X(n35475) );
  nand_x1_sg U41369 ( .A(n13556), .B(n41328), .X(n35476) );
  nand_x1_sg U41370 ( .A(n13550), .B(n41329), .X(n35477) );
  nand_x1_sg U41371 ( .A(n13532), .B(n41332), .X(n35478) );
  nand_x1_sg U41372 ( .A(n13526), .B(n41333), .X(n35479) );
  nand_x1_sg U41373 ( .A(n13520), .B(n41334), .X(n35480) );
  nand_x1_sg U41374 ( .A(n13492), .B(n41337), .X(n35481) );
  nand_x1_sg U41375 ( .A(n13461), .B(n41350), .X(n35482) );
  nand_x2_sg U41376 ( .A(n21351), .B(n21352), .X(n35484) );
  nand_x1_sg U41377 ( .A(n13538), .B(n41331), .X(n35486) );
  nand_x1_sg U41378 ( .A(n13479), .B(n41338), .X(n35487) );
  nand_x1_sg U41379 ( .A(n13473), .B(n41342), .X(n35488) );
  nand_x1_sg U41380 ( .A(n13467), .B(n41346), .X(n35489) );
  nand_x1_sg U41381 ( .A(n13455), .B(n41354), .X(n35490) );
  nand_x1_sg U41382 ( .A(n13449), .B(n41358), .X(n35491) );
  nand_x1_sg U41383 ( .A(n13443), .B(n41362), .X(n35492) );
  nand_x1_sg U41384 ( .A(n13437), .B(n41366), .X(n35493) );
  nand_x1_sg U41385 ( .A(n13431), .B(n41370), .X(n35494) );
  nand_x1_sg U41386 ( .A(n14818), .B(n13754), .X(n35495) );
  nand_x1_sg U41387 ( .A(n14663), .B(n13734), .X(n35496) );
  nand_x1_sg U41388 ( .A(n14350), .B(n13690), .X(n35497) );
  nand_x1_sg U41389 ( .A(n14195), .B(n13670), .X(n35498) );
  nand_x1_sg U41390 ( .A(n14164), .B(n13666), .X(n35499) );
  nand_x1_sg U41391 ( .A(n14040), .B(n13650), .X(n35500) );
  nand_x1_sg U41392 ( .A(n13916), .B(n13634), .X(n35501) );
  nand_x1_sg U41393 ( .A(n13885), .B(n13630), .X(n35502) );
  inv_x1_sg U41394 ( .A(n15183), .X(n35504) );
  nand_x1_sg U41395 ( .A(n21481), .B(n32063), .X(n21478) );
  nand_x1_sg U41396 ( .A(n32425), .B(n28833), .X(n28362) );
  nand_x1_sg U41397 ( .A(n32427), .B(n28789), .X(n28405) );
  nand_x1_sg U41398 ( .A(n12834), .B(n12835), .X(n35507) );
  inv_x1_sg U41399 ( .A(n15284), .X(n35508) );
  inv_x1_sg U41400 ( .A(n15054), .X(n35510) );
  nand_x1_sg U41401 ( .A(n35529), .B(n35510), .X(n35631) );
  nand_x1_sg U41402 ( .A(n32426), .B(n29665), .X(n29147) );
  inv_x1_sg U41403 ( .A(n28964), .X(n35511) );
  nand_x1_sg U41404 ( .A(n34537), .B(n32926), .X(n13368) );
  inv_x1_sg U41405 ( .A(n15188), .X(n35515) );
  nand_x1_sg U41406 ( .A(n30520), .B(n35515), .X(n15187) );
  nand_x2_sg U41407 ( .A(n15189), .B(n31662), .X(n15188) );
  inv_x1_sg U41408 ( .A(n15056), .X(n35516) );
  nand_x1_sg U41409 ( .A(n15004), .B(n13776), .X(n35517) );
  nand_x1_sg U41410 ( .A(n14756), .B(n13746), .X(n35518) );
  nand_x1_sg U41411 ( .A(n14725), .B(n13742), .X(n35519) );
  nand_x1_sg U41412 ( .A(n14444), .B(n13708), .X(n35520) );
  nand_x1_sg U41413 ( .A(n14381), .B(n13694), .X(n35521) );
  nand_x1_sg U41414 ( .A(n14133), .B(n13662), .X(n35522) );
  nand_x1_sg U41415 ( .A(n13785), .B(n13617), .X(n35523) );
  nand_x1_sg U41416 ( .A(n13425), .B(n41374), .X(n35524) );
  nand_x1_sg U41417 ( .A(n13419), .B(n41378), .X(n35525) );
  nand_x1_sg U41418 ( .A(n13413), .B(n41382), .X(n35526) );
  nor_x1_sg U41419 ( .A(n33558), .B(n34064), .X(n35679) );
  nor_x1_sg U41420 ( .A(n33498), .B(n34064), .X(n35661) );
  nor_x1_sg U41421 ( .A(n33654), .B(n34069), .X(n35665) );
  inv_x16_sg U41422 ( .A(reset), .X(n42410) );
  inv_x1_sg U41423 ( .A(n28745), .X(n35529) );
  nand_x1_sg U41424 ( .A(n14911), .B(n13766), .X(n35531) );
  nand_x1_sg U41425 ( .A(n14880), .B(n13762), .X(n35532) );
  nand_x1_sg U41426 ( .A(n14849), .B(n13758), .X(n35533) );
  nand_x1_sg U41427 ( .A(n14632), .B(n13730), .X(n35534) );
  nand_x1_sg U41428 ( .A(n14601), .B(n13726), .X(n35535) );
  nand_x1_sg U41429 ( .A(n14570), .B(n13722), .X(n35536) );
  nand_x1_sg U41430 ( .A(n14413), .B(n13704), .X(n35537) );
  nand_x1_sg U41431 ( .A(n14288), .B(n13682), .X(n35538) );
  nand_x1_sg U41432 ( .A(n14257), .B(n13678), .X(n35539) );
  nand_x1_sg U41433 ( .A(n14226), .B(n13674), .X(n35540) );
  nand_x1_sg U41434 ( .A(n14102), .B(n13658), .X(n35541) );
  nand_x1_sg U41435 ( .A(n14009), .B(n13646), .X(n35542) );
  nand_x1_sg U41436 ( .A(n13978), .B(n13642), .X(n35543) );
  nand_x1_sg U41437 ( .A(n13947), .B(n13638), .X(n35544) );
  nand_x1_sg U41438 ( .A(n13854), .B(n13626), .X(n35545) );
  nand_x1_sg U41439 ( .A(n13823), .B(n13622), .X(n35546) );
  nand_x1_sg U41440 ( .A(n13407), .B(n41386), .X(n35547) );
  nand_x1_sg U41441 ( .A(n13377), .B(n41406), .X(n35548) );
  nand_x1_sg U41442 ( .A(n13363), .B(n41414), .X(n35549) );
  nand_x1_sg U41443 ( .A(n14475), .B(n41523), .X(n35550) );
  inv_x1_sg U41444 ( .A(shifter_state[1]), .X(n35551) );
  inv_x1_sg U41445 ( .A(n29444), .X(n35552) );
  nand_x1_sg U41446 ( .A(n13401), .B(n41390), .X(n35554) );
  nand_x1_sg U41447 ( .A(n13395), .B(n41394), .X(n35555) );
  nand_x1_sg U41448 ( .A(n13389), .B(n41398), .X(n35556) );
  nand_x1_sg U41449 ( .A(n13371), .B(n41410), .X(n35557) );
  nand_x1_sg U41450 ( .A(n13509), .B(n41335), .X(n35558) );
  nand_x1_sg U41451 ( .A(n13383), .B(n41402), .X(n35559) );
  inv_x1_sg U41452 ( .A(n29663), .X(n35562) );
  inv_x1_sg U41453 ( .A(n12840), .X(n35563) );
  nand_x1_sg U41454 ( .A(n30524), .B(n35510), .X(n15047) );
  nand_x1_sg U41455 ( .A(n15201), .B(n31878), .X(n35564) );
  nand_x1_sg U41456 ( .A(n15065), .B(n31593), .X(n35565) );
  inv_x1_sg U41457 ( .A(o_mask[0]), .X(n35566) );
  inv_x1_sg U41458 ( .A(o_mask[3]), .X(n35567) );
  inv_x1_sg U41459 ( .A(o_mask[4]), .X(n35568) );
  inv_x1_sg U41460 ( .A(o_mask[6]), .X(n35569) );
  inv_x1_sg U41461 ( .A(o_mask[7]), .X(n35570) );
  inv_x1_sg U41462 ( .A(o_mask[8]), .X(n35571) );
  inv_x1_sg U41463 ( .A(o_mask[9]), .X(n35572) );
  inv_x1_sg U41464 ( .A(o_mask[12]), .X(n35573) );
  inv_x1_sg U41465 ( .A(o_mask[15]), .X(n35574) );
  inv_x1_sg U41466 ( .A(o_mask[18]), .X(n35575) );
  inv_x1_sg U41467 ( .A(o_mask[19]), .X(n35576) );
  inv_x1_sg U41468 ( .A(o_mask[20]), .X(n35577) );
  inv_x1_sg U41469 ( .A(o_mask[23]), .X(n35578) );
  inv_x1_sg U41470 ( .A(o_mask[25]), .X(n35579) );
  inv_x1_sg U41471 ( .A(o_mask[28]), .X(n35580) );
  inv_x1_sg U41472 ( .A(o_mask[31]), .X(n35581) );
  inv_x1_sg U41473 ( .A(n29667), .X(n35582) );
  nor_x1_sg U41474 ( .A(n20893), .B(n19609), .X(n35594) );
  nand_x1_sg U41475 ( .A(n35552), .B(n35515), .X(n35595) );
  nand_x1_sg U41476 ( .A(n35552), .B(n35530), .X(n35596) );
  nand_x1_sg U41477 ( .A(n35249), .B(n35504), .X(n35597) );
  nand_x1_sg U41478 ( .A(n35529), .B(n35508), .X(n35598) );
  nand_x1_sg U41479 ( .A(n35250), .B(n35508), .X(n35599) );
  nand_x2_sg U41480 ( .A(n21196), .B(n21197), .X(n21191) );
  nand_x2_sg U41481 ( .A(n21193), .B(n21194), .X(n21192) );
  nand_x1_sg U41482 ( .A(n21204), .B(n21205), .X(n21199) );
  nand_x1_sg U41483 ( .A(n21282), .B(n21283), .X(n21277) );
  nand_x2_sg U41484 ( .A(n21274), .B(n21275), .X(n21269) );
  nand_x2_sg U41485 ( .A(n21236), .B(n21237), .X(n21231) );
  nand_x2_sg U41486 ( .A(n21233), .B(n21234), .X(n21232) );
  nand_x1_sg U41487 ( .A(n21244), .B(n21245), .X(n21239) );
  nand_x1_sg U41488 ( .A(n21106), .B(n21107), .X(n21101) );
  nand_x2_sg U41489 ( .A(n21098), .B(n21099), .X(n21093) );
  nand_x1_sg U41490 ( .A(n21124), .B(n21125), .X(n21119) );
  nand_x2_sg U41491 ( .A(n21116), .B(n21117), .X(n21111) );
  nand_x1_sg U41492 ( .A(n21162), .B(n21163), .X(n21157) );
  nand_x2_sg U41493 ( .A(n21154), .B(n21155), .X(n21149) );
  nand_x1_sg U41494 ( .A(n21027), .B(n21028), .X(n21022) );
  nand_x2_sg U41495 ( .A(n21019), .B(n21020), .X(n21014) );
  nand_x1_sg U41496 ( .A(n21045), .B(n21046), .X(n21040) );
  nand_x2_sg U41497 ( .A(n21037), .B(n21038), .X(n21032) );
  nand_x1_sg U41498 ( .A(n21083), .B(n21084), .X(n21078) );
  nand_x2_sg U41499 ( .A(n21075), .B(n21076), .X(n21070) );
  nand_x1_sg U41500 ( .A(n21704), .B(n42634), .X(n21699) );
  inv_x1_sg U41501 ( .A(n21705), .X(n42634) );
  nand_x2_sg U41502 ( .A(n21693), .B(n21694), .X(n21692) );
  nand_x2_sg U41503 ( .A(n21589), .B(n21590), .X(n21584) );
  nand_x2_sg U41504 ( .A(n21586), .B(n21587), .X(n21585) );
  nand_x1_sg U41505 ( .A(n21594), .B(n21595), .X(n21593) );
  nand_x2_sg U41506 ( .A(n21607), .B(n21608), .X(n21602) );
  nand_x2_sg U41507 ( .A(n21604), .B(n21605), .X(n21603) );
  nand_x1_sg U41508 ( .A(n21612), .B(n21613), .X(n21611) );
  nand_x1_sg U41509 ( .A(n21653), .B(n42616), .X(n21648) );
  inv_x1_sg U41510 ( .A(n21654), .X(n42616) );
  nand_x2_sg U41511 ( .A(n21642), .B(n21643), .X(n21641) );
  nand_x2_sg U41512 ( .A(n21494), .B(n21495), .X(n21489) );
  nand_x2_sg U41513 ( .A(n21491), .B(n21492), .X(n21490) );
  nand_x1_sg U41514 ( .A(n21502), .B(n21503), .X(n21497) );
  nand_x2_sg U41515 ( .A(n21512), .B(n21513), .X(n21507) );
  nand_x2_sg U41516 ( .A(n21509), .B(n21510), .X(n21508) );
  nand_x1_sg U41517 ( .A(n21520), .B(n21521), .X(n21515) );
  nand_x1_sg U41518 ( .A(n21558), .B(n21559), .X(n21553) );
  nand_x2_sg U41519 ( .A(n21550), .B(n21551), .X(n21545) );
  nand_x2_sg U41520 ( .A(n21402), .B(n21403), .X(n21397) );
  nand_x2_sg U41521 ( .A(n21399), .B(n21400), .X(n21398) );
  nand_x1_sg U41522 ( .A(n21410), .B(n21411), .X(n21405) );
  nand_x2_sg U41523 ( .A(n21420), .B(n21421), .X(n21415) );
  nand_x2_sg U41524 ( .A(n21417), .B(n21418), .X(n21416) );
  nand_x1_sg U41525 ( .A(n21428), .B(n21429), .X(n21423) );
  nand_x1_sg U41526 ( .A(n21466), .B(n21467), .X(n21461) );
  nand_x2_sg U41527 ( .A(n21458), .B(n21459), .X(n21453) );
  nand_x2_sg U41528 ( .A(n15332), .B(n15333), .X(n15331) );
  nand_x1_sg U41529 ( .A(n15344), .B(n42388), .X(n15339) );
  inv_x1_sg U41530 ( .A(n15349), .X(n42395) );
  nand_x2_sg U41531 ( .A(n15350), .B(n15351), .X(n15349) );
  nand_x1_sg U41532 ( .A(n15328), .B(n42370), .X(n15324) );
  inv_x1_sg U41533 ( .A(n15298), .X(n42379) );
  nand_x2_sg U41534 ( .A(n21175), .B(n21176), .X(n21170) );
  nand_x2_sg U41535 ( .A(n21172), .B(n21173), .X(n21171) );
  nand_x1_sg U41536 ( .A(n21183), .B(n21184), .X(n21178) );
  nand_x2_sg U41537 ( .A(n21214), .B(n21215), .X(n21209) );
  nand_x2_sg U41538 ( .A(n21211), .B(n21212), .X(n21210) );
  nand_x1_sg U41539 ( .A(n21222), .B(n21223), .X(n21217) );
  nor_x1_sg U41540 ( .A(n21199), .B(n21200), .X(n21189) );
  nand_x1_sg U41541 ( .A(n21300), .B(n21301), .X(n21295) );
  nand_x2_sg U41542 ( .A(n21292), .B(n21293), .X(n21287) );
  nand_x2_sg U41543 ( .A(n21254), .B(n21255), .X(n21249) );
  nand_x2_sg U41544 ( .A(n21251), .B(n21252), .X(n21250) );
  nand_x1_sg U41545 ( .A(n21262), .B(n21263), .X(n21257) );
  nor_x1_sg U41546 ( .A(n21277), .B(n21278), .X(n21267) );
  nand_x2_sg U41547 ( .A(n21271), .B(n21272), .X(n21270) );
  nor_x1_sg U41548 ( .A(n21239), .B(n21240), .X(n21229) );
  nand_x1_sg U41549 ( .A(n21065), .B(n21066), .X(n21060) );
  nand_x2_sg U41550 ( .A(n21057), .B(n21058), .X(n21052) );
  nand_x1_sg U41551 ( .A(n21144), .B(n21145), .X(n21139) );
  nand_x2_sg U41552 ( .A(n21136), .B(n21137), .X(n21131) );
  nor_x1_sg U41553 ( .A(n21101), .B(n21102), .X(n21091) );
  nand_x2_sg U41554 ( .A(n21095), .B(n21096), .X(n21094) );
  nor_x1_sg U41555 ( .A(n21119), .B(n21120), .X(n21109) );
  nand_x2_sg U41556 ( .A(n21113), .B(n21114), .X(n21112) );
  nor_x1_sg U41557 ( .A(n21157), .B(n21158), .X(n21147) );
  nand_x2_sg U41558 ( .A(n21151), .B(n21152), .X(n21150) );
  nor_x1_sg U41559 ( .A(n21022), .B(n21023), .X(n21012) );
  nand_x2_sg U41560 ( .A(n21016), .B(n21017), .X(n21015) );
  nor_x1_sg U41561 ( .A(n21040), .B(n21041), .X(n21030) );
  nand_x2_sg U41562 ( .A(n21034), .B(n21035), .X(n21033) );
  nor_x1_sg U41563 ( .A(n21078), .B(n21079), .X(n21068) );
  nand_x2_sg U41564 ( .A(n21072), .B(n21073), .X(n21071) );
  nand_x1_sg U41565 ( .A(n21683), .B(n42641), .X(n21678) );
  inv_x1_sg U41566 ( .A(n21684), .X(n42641) );
  nand_x2_sg U41567 ( .A(n21672), .B(n21673), .X(n21671) );
  nand_x1_sg U41568 ( .A(n21722), .B(n42648), .X(n21717) );
  inv_x1_sg U41569 ( .A(n21723), .X(n42648) );
  nand_x2_sg U41570 ( .A(n21711), .B(n21712), .X(n21710) );
  nor_x1_sg U41571 ( .A(n21699), .B(n21700), .X(n21689) );
  nand_x2_sg U41572 ( .A(n21696), .B(n21697), .X(n21691) );
  nand_x1_sg U41573 ( .A(n21635), .B(n42627), .X(n21630) );
  inv_x1_sg U41574 ( .A(n21636), .X(n42627) );
  nand_x2_sg U41575 ( .A(n21624), .B(n21625), .X(n21623) );
  nor_x1_sg U41576 ( .A(n21592), .B(n21593), .X(n21582) );
  nor_x1_sg U41577 ( .A(n21610), .B(n21611), .X(n21600) );
  nor_x1_sg U41578 ( .A(n21648), .B(n21649), .X(n21638) );
  nand_x2_sg U41579 ( .A(n21645), .B(n21646), .X(n21640) );
  nand_x2_sg U41580 ( .A(n21529), .B(n42604), .X(n21528) );
  inv_x1_sg U41581 ( .A(n21530), .X(n42604) );
  nand_x2_sg U41582 ( .A(n21532), .B(n21533), .X(n21527) );
  nand_x1_sg U41583 ( .A(n21537), .B(n21538), .X(n21536) );
  nor_x1_sg U41584 ( .A(n21497), .B(n21498), .X(n21487) );
  nor_x1_sg U41585 ( .A(n21515), .B(n21516), .X(n21505) );
  nor_x1_sg U41586 ( .A(n21553), .B(n21554), .X(n21543) );
  nand_x2_sg U41587 ( .A(n21547), .B(n21548), .X(n21546) );
  nand_x2_sg U41588 ( .A(n21440), .B(n21441), .X(n21435) );
  nand_x2_sg U41589 ( .A(n21437), .B(n21438), .X(n21436) );
  nand_x1_sg U41590 ( .A(n21448), .B(n21449), .X(n21443) );
  nor_x1_sg U41591 ( .A(n21405), .B(n21406), .X(n21395) );
  nor_x1_sg U41592 ( .A(n21423), .B(n21424), .X(n21413) );
  nor_x1_sg U41593 ( .A(n21461), .B(n21462), .X(n21451) );
  nand_x2_sg U41594 ( .A(n21455), .B(n21456), .X(n21454) );
  nand_x1_sg U41595 ( .A(n12612), .B(n12613), .X(n12611) );
  inv_x1_sg U41596 ( .A(n12704), .X(n41705) );
  nand_x2_sg U41597 ( .A(n15321), .B(n15322), .X(n15320) );
  nand_x2_sg U41598 ( .A(n42381), .B(n15323), .X(n15322) );
  nand_x2_sg U41599 ( .A(n42395), .B(n15338), .X(n15321) );
  inv_x1_sg U41600 ( .A(n15331), .X(n42381) );
  nand_x2_sg U41601 ( .A(n15288), .B(n15289), .X(n15287) );
  nand_x2_sg U41602 ( .A(n42394), .B(n15305), .X(n15288) );
  nand_x2_sg U41603 ( .A(n42379), .B(n15290), .X(n15289) );
  inv_x1_sg U41604 ( .A(n15314), .X(n42394) );
  nand_x1_sg U41605 ( .A(n15271), .B(n15272), .X(n15270) );
  nand_x2_sg U41606 ( .A(n15256), .B(n15257), .X(n15255) );
  nor_x1_sg U41607 ( .A(n21178), .B(n21179), .X(n21168) );
  nor_x1_sg U41608 ( .A(n21217), .B(n21218), .X(n21207) );
  nor_x1_sg U41609 ( .A(n21295), .B(n21296), .X(n21285) );
  nand_x2_sg U41610 ( .A(n21289), .B(n21290), .X(n21288) );
  nor_x1_sg U41611 ( .A(n21257), .B(n21258), .X(n21247) );
  nor_x1_sg U41612 ( .A(n21060), .B(n21061), .X(n21050) );
  nand_x2_sg U41613 ( .A(n21054), .B(n21055), .X(n21053) );
  nor_x1_sg U41614 ( .A(n21139), .B(n21140), .X(n21129) );
  nand_x2_sg U41615 ( .A(n21133), .B(n21134), .X(n21132) );
  nor_x1_sg U41616 ( .A(n21678), .B(n21679), .X(n21668) );
  nand_x2_sg U41617 ( .A(n21675), .B(n21676), .X(n21670) );
  nor_x1_sg U41618 ( .A(n21717), .B(n21718), .X(n21707) );
  nand_x2_sg U41619 ( .A(n21714), .B(n21715), .X(n21709) );
  nor_x1_sg U41620 ( .A(n21630), .B(n21631), .X(n21620) );
  nand_x2_sg U41621 ( .A(n21627), .B(n21628), .X(n21622) );
  nor_x1_sg U41622 ( .A(n21535), .B(n21536), .X(n21525) );
  nor_x1_sg U41623 ( .A(n21443), .B(n21444), .X(n21433) );
  inv_x1_sg U41624 ( .A(n34513), .X(n35656) );
  nand_x1_sg U41625 ( .A(n13802), .B(n13803), .X(n13801) );
  nand_x1_sg U41626 ( .A(n13839), .B(n13840), .X(n13838) );
  nand_x1_sg U41627 ( .A(n13870), .B(n13871), .X(n13869) );
  nand_x1_sg U41628 ( .A(n13901), .B(n13902), .X(n13900) );
  nand_x1_sg U41629 ( .A(n13932), .B(n13933), .X(n13931) );
  nand_x1_sg U41630 ( .A(n13963), .B(n13964), .X(n13962) );
  nand_x1_sg U41631 ( .A(n13994), .B(n13995), .X(n13993) );
  nand_x1_sg U41632 ( .A(n14025), .B(n14026), .X(n14024) );
  nand_x1_sg U41633 ( .A(n14056), .B(n14057), .X(n14055) );
  nand_x1_sg U41634 ( .A(n14087), .B(n14088), .X(n14086) );
  nand_x1_sg U41635 ( .A(n14118), .B(n14119), .X(n14117) );
  nand_x1_sg U41636 ( .A(n14149), .B(n14150), .X(n14148) );
  nand_x1_sg U41637 ( .A(n14180), .B(n14181), .X(n14179) );
  nand_x1_sg U41638 ( .A(n14211), .B(n14212), .X(n14210) );
  nand_x1_sg U41639 ( .A(n14242), .B(n14243), .X(n14241) );
  nand_x1_sg U41640 ( .A(n14273), .B(n14274), .X(n14272) );
  nand_x1_sg U41641 ( .A(n14304), .B(n14305), .X(n14303) );
  nand_x1_sg U41642 ( .A(n14335), .B(n14336), .X(n14334) );
  nand_x1_sg U41643 ( .A(n14366), .B(n14367), .X(n14365) );
  nand_x1_sg U41644 ( .A(n14397), .B(n14398), .X(n14396) );
  nand_x1_sg U41645 ( .A(n14429), .B(n14430), .X(n14428) );
  nand_x1_sg U41646 ( .A(n14460), .B(n14461), .X(n14459) );
  nand_x1_sg U41647 ( .A(n14524), .B(n14525), .X(n14523) );
  nand_x1_sg U41648 ( .A(n14586), .B(n14587), .X(n14585) );
  nand_x1_sg U41649 ( .A(n14617), .B(n14618), .X(n14616) );
  nand_x1_sg U41650 ( .A(n14648), .B(n14649), .X(n14647) );
  nand_x1_sg U41651 ( .A(n14679), .B(n14680), .X(n14678) );
  nand_x1_sg U41652 ( .A(n14710), .B(n14711), .X(n14709) );
  nand_x1_sg U41653 ( .A(n14741), .B(n14742), .X(n14740) );
  nand_x1_sg U41654 ( .A(n14772), .B(n14773), .X(n14771) );
  nand_x1_sg U41655 ( .A(n14803), .B(n14804), .X(n14802) );
  nand_x1_sg U41656 ( .A(n14834), .B(n14835), .X(n14833) );
  nand_x1_sg U41657 ( .A(n14865), .B(n14866), .X(n14864) );
  nand_x1_sg U41658 ( .A(n14896), .B(n14897), .X(n14895) );
  nand_x1_sg U41659 ( .A(n14927), .B(n14928), .X(n14926) );
  nand_x1_sg U41660 ( .A(n15020), .B(n15021), .X(n15019) );
  nand_x1_sg U41661 ( .A(n15045), .B(n42402), .X(n15046) );
  nand_x1_sg U41662 ( .A(n28965), .B(n42402), .X(n15050) );
  nand_x1_sg U41663 ( .A(n15142), .B(n15143), .X(n15141) );
  nand_x2_sg U41664 ( .A(n15127), .B(n15128), .X(n15126) );
  nand_x1_sg U41665 ( .A(n15091), .B(n42367), .X(n15085) );
  nand_x1_sg U41666 ( .A(n15178), .B(n35530), .X(n15179) );
  nand_x1_sg U41667 ( .A(n29664), .B(n35530), .X(n15184) );
  nand_x1_sg U41668 ( .A(n15225), .B(n42368), .X(n15221) );
  inv_x1_sg U41669 ( .A(n15228), .X(n42378) );
  nand_x2_sg U41670 ( .A(n15229), .B(n15230), .X(n15228) );
  nor_x1_sg U41671 ( .A(n15269), .B(n15270), .X(n15252) );
  nand_x2_sg U41672 ( .A(n15262), .B(n15263), .X(n15254) );
  nor_x1_sg U41673 ( .A(n15236), .B(n15237), .X(n15235) );
  inv_x1_sg U41674 ( .A(n20919), .X(n42542) );
  nand_x1_sg U41675 ( .A(n20989), .B(n20990), .X(n20985) );
  nand_x2_sg U41676 ( .A(n21225), .B(n21226), .X(n20919) );
  nand_x1_sg U41677 ( .A(n20999), .B(n21000), .X(n20993) );
  nand_x1_sg U41678 ( .A(n20969), .B(n20970), .X(n20962) );
  nand_x2_sg U41679 ( .A(n21087), .B(n21088), .X(n21086) );
  nand_x1_sg U41680 ( .A(n20979), .B(n20980), .X(n20973) );
  nand_x2_sg U41681 ( .A(n21008), .B(n21009), .X(n21007) );
  nand_x2_sg U41682 ( .A(n21318), .B(n21319), .X(n21317) );
  nand_x2_sg U41683 ( .A(n21321), .B(n21322), .X(n21316) );
  nand_x2_sg U41684 ( .A(n21312), .B(n21313), .X(n21307) );
  nand_x1_sg U41685 ( .A(n21663), .B(n21664), .X(n21659) );
  nand_x2_sg U41686 ( .A(n21578), .B(n21579), .X(n21577) );
  nand_x1_sg U41687 ( .A(n21572), .B(n21573), .X(n21566) );
  nand_x2_sg U41688 ( .A(n21483), .B(n21484), .X(n21482) );
  nand_x1_sg U41689 ( .A(n21478), .B(n21479), .X(n21472) );
  nand_x2_sg U41690 ( .A(n21391), .B(n21392), .X(n21390) );
  nand_x1_sg U41691 ( .A(n21385), .B(n21386), .X(n21379) );
  nand_x2_sg U41692 ( .A(n21738), .B(n21739), .X(n21737) );
  nand_x2_sg U41693 ( .A(n21741), .B(n21742), .X(n21736) );
  nand_x1_sg U41694 ( .A(n21729), .B(n21730), .X(n21728) );
  nand_x1_sg U41695 ( .A(n34447), .B(n11891), .X(n11888) );
  nand_x1_sg U41696 ( .A(n13806), .B(n13807), .X(n13800) );
  nand_x1_sg U41697 ( .A(n13841), .B(n13842), .X(n13837) );
  nand_x1_sg U41698 ( .A(n13872), .B(n13873), .X(n13868) );
  nor_x1_sg U41699 ( .A(n13907), .B(n13908), .X(n13897) );
  nand_x1_sg U41700 ( .A(n13903), .B(n13904), .X(n13899) );
  nor_x1_sg U41701 ( .A(n13938), .B(n13939), .X(n13928) );
  nand_x1_sg U41702 ( .A(n13934), .B(n13935), .X(n13930) );
  nand_x1_sg U41703 ( .A(n13965), .B(n13966), .X(n13961) );
  nand_x1_sg U41704 ( .A(n13996), .B(n13997), .X(n13992) );
  nand_x1_sg U41705 ( .A(n14027), .B(n14028), .X(n14023) );
  nand_x1_sg U41706 ( .A(n14058), .B(n14059), .X(n14054) );
  nand_x1_sg U41707 ( .A(n14089), .B(n14090), .X(n14085) );
  nand_x1_sg U41708 ( .A(n14120), .B(n14121), .X(n14116) );
  nand_x1_sg U41709 ( .A(n14151), .B(n14152), .X(n14147) );
  nand_x1_sg U41710 ( .A(n14182), .B(n14183), .X(n14178) );
  nand_x1_sg U41711 ( .A(n14213), .B(n14214), .X(n14209) );
  nand_x1_sg U41712 ( .A(n14244), .B(n14245), .X(n14240) );
  nand_x1_sg U41713 ( .A(n14275), .B(n14276), .X(n14271) );
  nand_x1_sg U41714 ( .A(n14306), .B(n14307), .X(n14302) );
  nor_x1_sg U41715 ( .A(n14341), .B(n14342), .X(n14331) );
  nand_x1_sg U41716 ( .A(n14337), .B(n14338), .X(n14333) );
  nor_x1_sg U41717 ( .A(n14372), .B(n14373), .X(n14362) );
  nand_x1_sg U41718 ( .A(n14368), .B(n14369), .X(n14364) );
  nand_x1_sg U41719 ( .A(n14399), .B(n14400), .X(n14395) );
  nand_x1_sg U41720 ( .A(n14431), .B(n14432), .X(n14427) );
  nand_x1_sg U41721 ( .A(n14462), .B(n14463), .X(n14458) );
  nand_x1_sg U41722 ( .A(n14500), .B(n14501), .X(n14499) );
  nand_x1_sg U41723 ( .A(n14494), .B(n14495), .X(n14490) );
  nand_x1_sg U41724 ( .A(n14526), .B(n14527), .X(n14522) );
  nand_x1_sg U41725 ( .A(n14562), .B(n14563), .X(n14561) );
  nand_x1_sg U41726 ( .A(n14558), .B(n14559), .X(n14554) );
  nand_x1_sg U41727 ( .A(n14588), .B(n14589), .X(n14584) );
  nand_x1_sg U41728 ( .A(n14619), .B(n14620), .X(n14615) );
  nand_x1_sg U41729 ( .A(n14650), .B(n14651), .X(n14646) );
  nor_x1_sg U41730 ( .A(n14685), .B(n14686), .X(n14675) );
  nand_x1_sg U41731 ( .A(n14681), .B(n14682), .X(n14677) );
  nor_x1_sg U41732 ( .A(n14716), .B(n14717), .X(n14706) );
  nand_x1_sg U41733 ( .A(n14712), .B(n14713), .X(n14708) );
  nand_x1_sg U41734 ( .A(n14743), .B(n14744), .X(n14739) );
  nand_x1_sg U41735 ( .A(n14774), .B(n14775), .X(n14770) );
  nor_x1_sg U41736 ( .A(n14809), .B(n14810), .X(n14799) );
  nand_x1_sg U41737 ( .A(n14805), .B(n14806), .X(n14801) );
  nor_x1_sg U41738 ( .A(n14840), .B(n14841), .X(n14830) );
  nand_x1_sg U41739 ( .A(n14836), .B(n14837), .X(n14832) );
  nand_x1_sg U41740 ( .A(n14867), .B(n14868), .X(n14863) );
  nand_x1_sg U41741 ( .A(n14898), .B(n14899), .X(n14894) );
  nor_x1_sg U41742 ( .A(n14933), .B(n14934), .X(n14923) );
  nand_x1_sg U41743 ( .A(n14929), .B(n14930), .X(n14925) );
  nand_x1_sg U41744 ( .A(n14965), .B(n14966), .X(n14964) );
  nand_x1_sg U41745 ( .A(n14961), .B(n14962), .X(n14957) );
  nand_x1_sg U41746 ( .A(n14996), .B(n14997), .X(n14995) );
  nand_x1_sg U41747 ( .A(n14992), .B(n14993), .X(n14988) );
  nand_x1_sg U41748 ( .A(n15022), .B(n15023), .X(n15018) );
  nand_x1_sg U41749 ( .A(n13291), .B(n35252), .X(n13287) );
  nand_x4_sg U41750 ( .A(n13609), .B(n13610), .X(n13606) );
  inv_x1_sg U41751 ( .A(n13786), .X(n35627) );
  inv_x1_sg U41752 ( .A(n13824), .X(n35626) );
  inv_x1_sg U41753 ( .A(n13855), .X(n35625) );
  inv_x1_sg U41754 ( .A(n13886), .X(n41288) );
  inv_x1_sg U41755 ( .A(n13917), .X(n41289) );
  inv_x1_sg U41756 ( .A(n13948), .X(n41290) );
  inv_x1_sg U41757 ( .A(n13979), .X(n41291) );
  inv_x1_sg U41758 ( .A(n14010), .X(n41292) );
  inv_x1_sg U41759 ( .A(n14041), .X(n41293) );
  inv_x1_sg U41760 ( .A(n14072), .X(n41294) );
  inv_x1_sg U41761 ( .A(n14103), .X(n41295) );
  inv_x1_sg U41762 ( .A(n14134), .X(n41296) );
  inv_x1_sg U41763 ( .A(n14165), .X(n41297) );
  inv_x1_sg U41764 ( .A(n14196), .X(n41298) );
  inv_x1_sg U41765 ( .A(n14227), .X(n41299) );
  inv_x1_sg U41766 ( .A(n14258), .X(n41300) );
  inv_x1_sg U41767 ( .A(n14289), .X(n41301) );
  inv_x1_sg U41768 ( .A(n14320), .X(n41302) );
  inv_x1_sg U41769 ( .A(n14351), .X(n41303) );
  inv_x1_sg U41770 ( .A(n14382), .X(n41304) );
  inv_x1_sg U41771 ( .A(n14414), .X(n41305) );
  inv_x1_sg U41772 ( .A(n14445), .X(n41306) );
  inv_x1_sg U41773 ( .A(n14476), .X(n41523) );
  inv_x1_sg U41774 ( .A(n14509), .X(n41307) );
  inv_x1_sg U41775 ( .A(n14540), .X(n41522) );
  inv_x1_sg U41776 ( .A(n14571), .X(n41308) );
  inv_x1_sg U41777 ( .A(n14602), .X(n41309) );
  inv_x1_sg U41778 ( .A(n14633), .X(n41310) );
  inv_x1_sg U41779 ( .A(n14664), .X(n41311) );
  inv_x1_sg U41780 ( .A(n14695), .X(n41312) );
  inv_x1_sg U41781 ( .A(n14726), .X(n41313) );
  inv_x1_sg U41782 ( .A(n14757), .X(n41314) );
  inv_x1_sg U41783 ( .A(n14788), .X(n41315) );
  inv_x1_sg U41784 ( .A(n14819), .X(n41316) );
  inv_x1_sg U41785 ( .A(n14850), .X(n41317) );
  inv_x1_sg U41786 ( .A(n14881), .X(n41318) );
  inv_x1_sg U41787 ( .A(n14912), .X(n41319) );
  inv_x1_sg U41788 ( .A(n14943), .X(n41521) );
  inv_x1_sg U41789 ( .A(n14974), .X(n41520) );
  inv_x1_sg U41790 ( .A(n15005), .X(n41320) );
  nor_x1_sg U41791 ( .A(n15140), .B(n15141), .X(n15123) );
  nand_x2_sg U41792 ( .A(n15133), .B(n15134), .X(n15125) );
  nor_x1_sg U41793 ( .A(n15107), .B(n15108), .X(n15106) );
  nand_x1_sg U41794 ( .A(n42377), .B(n15084), .X(n15083) );
  inv_x1_sg U41795 ( .A(n15096), .X(n42377) );
  nand_x2_sg U41796 ( .A(n15097), .B(n15098), .X(n15096) );
  nand_x1_sg U41797 ( .A(n15216), .B(n15217), .X(n15215) );
  nand_x1_sg U41798 ( .A(n15218), .B(n15219), .X(n15217) );
  nand_x1_sg U41799 ( .A(n42378), .B(n15220), .X(n15219) );
  nand_x2_sg U41800 ( .A(n20958), .B(n20959), .X(n20938) );
  nand_x2_sg U41801 ( .A(n21309), .B(n21310), .X(n21308) );
  nor_x1_sg U41802 ( .A(n21727), .B(n21728), .X(n21726) );
  nand_x1_sg U41803 ( .A(n11903), .B(n11904), .X(n11537) );
  nand_x1_sg U41804 ( .A(n11915), .B(n11916), .X(n11538) );
  nand_x1_sg U41805 ( .A(n11926), .B(n11927), .X(n11539) );
  nand_x1_sg U41806 ( .A(n11937), .B(n11938), .X(n11540) );
  nand_x1_sg U41807 ( .A(n11948), .B(n11949), .X(n11541) );
  nand_x1_sg U41808 ( .A(n11959), .B(n11960), .X(n11542) );
  nand_x1_sg U41809 ( .A(n11970), .B(n11971), .X(n11543) );
  nand_x1_sg U41810 ( .A(n11981), .B(n11982), .X(n11544) );
  nand_x1_sg U41811 ( .A(n11992), .B(n11993), .X(n11545) );
  nand_x1_sg U41812 ( .A(n12003), .B(n12004), .X(n11546) );
  nand_x1_sg U41813 ( .A(n12014), .B(n12015), .X(n11547) );
  nand_x1_sg U41814 ( .A(n12025), .B(n12026), .X(n11548) );
  nand_x1_sg U41815 ( .A(n12036), .B(n12037), .X(n11549) );
  nand_x1_sg U41816 ( .A(n12047), .B(n12048), .X(n11550) );
  nand_x1_sg U41817 ( .A(n12058), .B(n12059), .X(n11551) );
  nand_x1_sg U41818 ( .A(n12069), .B(n12070), .X(n11552) );
  nand_x1_sg U41819 ( .A(n12080), .B(n12081), .X(n11553) );
  nand_x1_sg U41820 ( .A(n12091), .B(n12092), .X(n11554) );
  nand_x1_sg U41821 ( .A(n12102), .B(n12103), .X(n11555) );
  nand_x1_sg U41822 ( .A(n12113), .B(n12114), .X(n11556) );
  nand_x1_sg U41823 ( .A(n12131), .B(n12132), .X(n11563) );
  nand_x1_sg U41824 ( .A(n12143), .B(n12144), .X(n11564) );
  nand_x1_sg U41825 ( .A(n12154), .B(n12155), .X(n11565) );
  nand_x1_sg U41826 ( .A(n12165), .B(n12166), .X(n11566) );
  nand_x1_sg U41827 ( .A(n12176), .B(n12177), .X(n11567) );
  nand_x1_sg U41828 ( .A(n12187), .B(n12188), .X(n11568) );
  nand_x1_sg U41829 ( .A(n12198), .B(n12199), .X(n11569) );
  nand_x1_sg U41830 ( .A(n12209), .B(n12210), .X(n11570) );
  nand_x1_sg U41831 ( .A(n12220), .B(n12221), .X(n11571) );
  nand_x1_sg U41832 ( .A(n12231), .B(n12232), .X(n11572) );
  nand_x1_sg U41833 ( .A(n12242), .B(n12243), .X(n11573) );
  nand_x1_sg U41834 ( .A(n12253), .B(n12254), .X(n11574) );
  nand_x1_sg U41835 ( .A(n12264), .B(n12265), .X(n11575) );
  nand_x1_sg U41836 ( .A(n12275), .B(n12276), .X(n11576) );
  nand_x1_sg U41837 ( .A(n12286), .B(n12287), .X(n11577) );
  nand_x1_sg U41838 ( .A(n12297), .B(n12298), .X(n11578) );
  nand_x1_sg U41839 ( .A(n12308), .B(n12309), .X(n11579) );
  nand_x1_sg U41840 ( .A(n12319), .B(n12320), .X(n11580) );
  nand_x1_sg U41841 ( .A(n12330), .B(n12331), .X(n11581) );
  nand_x1_sg U41842 ( .A(n12341), .B(n12342), .X(n11582) );
  nand_x1_sg U41843 ( .A(n41143), .B(n11902), .X(n11587) );
  nand_x1_sg U41844 ( .A(n41144), .B(n11914), .X(n11588) );
  nand_x1_sg U41845 ( .A(n41145), .B(n11925), .X(n11589) );
  nand_x1_sg U41846 ( .A(n41146), .B(n11936), .X(n11590) );
  nand_x1_sg U41847 ( .A(n41147), .B(n11947), .X(n11591) );
  nand_x1_sg U41848 ( .A(n41148), .B(n11958), .X(n11592) );
  nand_x1_sg U41849 ( .A(n41149), .B(n11969), .X(n11593) );
  nand_x1_sg U41850 ( .A(n41150), .B(n11980), .X(n11594) );
  nand_x1_sg U41851 ( .A(n41151), .B(n11991), .X(n11595) );
  nand_x1_sg U41852 ( .A(n41152), .B(n12002), .X(n11596) );
  nand_x1_sg U41853 ( .A(n41153), .B(n12013), .X(n11597) );
  nand_x1_sg U41854 ( .A(n41154), .B(n12024), .X(n11598) );
  nand_x1_sg U41855 ( .A(n41155), .B(n12035), .X(n11599) );
  nand_x1_sg U41856 ( .A(n41156), .B(n12046), .X(n11600) );
  nand_x1_sg U41857 ( .A(n41157), .B(n12057), .X(n11601) );
  nand_x1_sg U41858 ( .A(n41158), .B(n12068), .X(n11602) );
  nand_x1_sg U41859 ( .A(n41159), .B(n12079), .X(n11603) );
  nand_x1_sg U41860 ( .A(n41160), .B(n12090), .X(n11604) );
  nand_x1_sg U41861 ( .A(n41161), .B(n12101), .X(n11605) );
  nand_x1_sg U41862 ( .A(n41162), .B(n12112), .X(n11606) );
  nand_x1_sg U41863 ( .A(n41163), .B(n12130), .X(n11614) );
  nand_x1_sg U41864 ( .A(n41164), .B(n12142), .X(n11615) );
  nand_x1_sg U41865 ( .A(n41165), .B(n12153), .X(n11616) );
  nand_x1_sg U41866 ( .A(n41166), .B(n12164), .X(n11617) );
  nand_x1_sg U41867 ( .A(n41167), .B(n12175), .X(n11618) );
  nand_x1_sg U41868 ( .A(n41168), .B(n12186), .X(n11619) );
  nand_x1_sg U41869 ( .A(n41169), .B(n12197), .X(n11620) );
  nand_x1_sg U41870 ( .A(n41170), .B(n12208), .X(n11621) );
  nand_x1_sg U41871 ( .A(n41171), .B(n12219), .X(n11622) );
  nand_x1_sg U41872 ( .A(n41172), .B(n12230), .X(n11623) );
  nand_x1_sg U41873 ( .A(n41173), .B(n12241), .X(n11624) );
  nand_x1_sg U41874 ( .A(n41174), .B(n12252), .X(n11625) );
  nand_x1_sg U41875 ( .A(n41175), .B(n12263), .X(n11626) );
  nand_x1_sg U41876 ( .A(n41176), .B(n12274), .X(n11627) );
  nand_x1_sg U41877 ( .A(n41177), .B(n12285), .X(n11628) );
  nand_x1_sg U41878 ( .A(n41178), .B(n12296), .X(n11629) );
  nand_x1_sg U41879 ( .A(n41179), .B(n12307), .X(n11630) );
  nand_x1_sg U41880 ( .A(n41180), .B(n12318), .X(n11631) );
  nand_x1_sg U41881 ( .A(n41181), .B(n12329), .X(n11632) );
  nand_x1_sg U41882 ( .A(n41182), .B(n12340), .X(n11633) );
  nand_x1_sg U41883 ( .A(n41184), .B(n11901), .X(n11642) );
  nand_x1_sg U41884 ( .A(n41185), .B(n11913), .X(n11643) );
  nand_x1_sg U41885 ( .A(n41186), .B(n11924), .X(n11644) );
  nand_x1_sg U41886 ( .A(n41187), .B(n11935), .X(n11645) );
  nand_x1_sg U41887 ( .A(n41188), .B(n11946), .X(n11646) );
  nand_x1_sg U41888 ( .A(n41189), .B(n11957), .X(n11647) );
  nand_x1_sg U41889 ( .A(n41190), .B(n11968), .X(n11648) );
  nand_x1_sg U41890 ( .A(n41191), .B(n11979), .X(n11649) );
  nand_x1_sg U41891 ( .A(n41192), .B(n11990), .X(n11650) );
  nand_x1_sg U41892 ( .A(n41193), .B(n12001), .X(n11651) );
  nand_x1_sg U41893 ( .A(n41194), .B(n12012), .X(n11652) );
  nand_x1_sg U41894 ( .A(n41195), .B(n12023), .X(n11653) );
  nand_x1_sg U41895 ( .A(n41196), .B(n12034), .X(n11654) );
  nand_x1_sg U41896 ( .A(n41197), .B(n12045), .X(n11655) );
  nand_x1_sg U41897 ( .A(n41198), .B(n12056), .X(n11656) );
  nand_x1_sg U41898 ( .A(n41199), .B(n12067), .X(n11657) );
  nand_x1_sg U41899 ( .A(n41200), .B(n12078), .X(n11658) );
  nand_x1_sg U41900 ( .A(n41201), .B(n12089), .X(n11659) );
  nand_x1_sg U41901 ( .A(n41202), .B(n12100), .X(n11660) );
  nand_x1_sg U41902 ( .A(n41203), .B(n12111), .X(n11661) );
  nand_x1_sg U41903 ( .A(n41204), .B(n12129), .X(n11668) );
  nand_x1_sg U41904 ( .A(n41205), .B(n12141), .X(n11669) );
  nand_x1_sg U41905 ( .A(n41206), .B(n12152), .X(n11670) );
  nand_x1_sg U41906 ( .A(n41207), .B(n12163), .X(n11671) );
  nand_x1_sg U41907 ( .A(n41208), .B(n12174), .X(n11672) );
  nand_x1_sg U41908 ( .A(n41209), .B(n12185), .X(n11673) );
  nand_x1_sg U41909 ( .A(n41210), .B(n12196), .X(n11674) );
  nand_x1_sg U41910 ( .A(n41211), .B(n12207), .X(n11675) );
  nand_x1_sg U41911 ( .A(n41212), .B(n12218), .X(n11676) );
  nand_x1_sg U41912 ( .A(n41213), .B(n12229), .X(n11677) );
  nand_x1_sg U41913 ( .A(n41214), .B(n12240), .X(n11678) );
  nand_x1_sg U41914 ( .A(n41215), .B(n12251), .X(n11679) );
  nand_x1_sg U41915 ( .A(n41216), .B(n12262), .X(n11680) );
  nand_x1_sg U41916 ( .A(n41217), .B(n12273), .X(n11681) );
  nand_x1_sg U41917 ( .A(n41218), .B(n12284), .X(n11682) );
  nand_x1_sg U41918 ( .A(n41219), .B(n12295), .X(n11683) );
  nand_x1_sg U41919 ( .A(n41220), .B(n12306), .X(n11684) );
  nand_x1_sg U41920 ( .A(n41221), .B(n12317), .X(n11685) );
  nand_x1_sg U41921 ( .A(n41222), .B(n12328), .X(n11686) );
  nand_x1_sg U41922 ( .A(n41223), .B(n12339), .X(n11687) );
  nand_x1_sg U41923 ( .A(n41224), .B(n11900), .X(n11690) );
  nand_x1_sg U41924 ( .A(n41225), .B(n11912), .X(n11691) );
  nand_x1_sg U41925 ( .A(n41226), .B(n11923), .X(n11692) );
  nand_x1_sg U41926 ( .A(n41227), .B(n11934), .X(n11693) );
  nand_x1_sg U41927 ( .A(n41228), .B(n11945), .X(n11694) );
  nand_x1_sg U41928 ( .A(n41229), .B(n11956), .X(n11695) );
  nand_x1_sg U41929 ( .A(n41230), .B(n11967), .X(n11696) );
  nand_x1_sg U41930 ( .A(n41231), .B(n11978), .X(n11697) );
  nand_x1_sg U41931 ( .A(n41232), .B(n11989), .X(n11698) );
  nand_x1_sg U41932 ( .A(n41233), .B(n12000), .X(n11699) );
  nand_x1_sg U41933 ( .A(n41234), .B(n12011), .X(n11700) );
  nand_x1_sg U41934 ( .A(n41235), .B(n12022), .X(n11701) );
  nand_x1_sg U41935 ( .A(n41236), .B(n12033), .X(n11702) );
  nand_x1_sg U41936 ( .A(n41237), .B(n12044), .X(n11703) );
  nand_x1_sg U41937 ( .A(n41238), .B(n12055), .X(n11704) );
  nand_x1_sg U41938 ( .A(n41239), .B(n12066), .X(n11705) );
  nand_x1_sg U41939 ( .A(n41240), .B(n12077), .X(n11706) );
  nand_x1_sg U41940 ( .A(n41241), .B(n12088), .X(n11707) );
  nand_x1_sg U41941 ( .A(n41242), .B(n12099), .X(n11708) );
  nand_x1_sg U41942 ( .A(n41243), .B(n12110), .X(n11709) );
  nand_x1_sg U41943 ( .A(n41244), .B(n12128), .X(n11717) );
  nand_x1_sg U41944 ( .A(n41245), .B(n12140), .X(n11718) );
  nand_x1_sg U41945 ( .A(n41246), .B(n12151), .X(n11719) );
  nand_x1_sg U41946 ( .A(n41247), .B(n12162), .X(n11720) );
  nand_x1_sg U41947 ( .A(n41248), .B(n12173), .X(n11721) );
  nand_x1_sg U41948 ( .A(n41249), .B(n12184), .X(n11722) );
  nand_x1_sg U41949 ( .A(n41250), .B(n12195), .X(n11723) );
  nand_x1_sg U41950 ( .A(n41251), .B(n12206), .X(n11724) );
  nand_x1_sg U41951 ( .A(n41252), .B(n12217), .X(n11725) );
  nand_x1_sg U41952 ( .A(n41253), .B(n12228), .X(n11726) );
  nand_x1_sg U41953 ( .A(n41254), .B(n12239), .X(n11727) );
  nand_x1_sg U41954 ( .A(n41255), .B(n12250), .X(n11728) );
  nand_x1_sg U41955 ( .A(n41256), .B(n12261), .X(n11729) );
  nand_x1_sg U41956 ( .A(n41257), .B(n12272), .X(n11730) );
  nand_x1_sg U41957 ( .A(n41258), .B(n12283), .X(n11731) );
  nand_x1_sg U41958 ( .A(n41259), .B(n12294), .X(n11732) );
  nand_x1_sg U41959 ( .A(n41260), .B(n12305), .X(n11733) );
  nand_x1_sg U41960 ( .A(n41261), .B(n12316), .X(n11734) );
  nand_x1_sg U41961 ( .A(n41262), .B(n12327), .X(n11735) );
  nand_x1_sg U41962 ( .A(n41263), .B(n12338), .X(n11736) );
  nand_x1_sg U41963 ( .A(n41419), .B(n11899), .X(n11743) );
  nand_x1_sg U41964 ( .A(n41420), .B(n11911), .X(n11744) );
  nand_x1_sg U41965 ( .A(n41421), .B(n11922), .X(n11745) );
  nand_x1_sg U41966 ( .A(n41422), .B(n11933), .X(n11746) );
  nand_x1_sg U41967 ( .A(n41423), .B(n11944), .X(n11747) );
  nand_x1_sg U41968 ( .A(n41424), .B(n11955), .X(n11748) );
  nand_x1_sg U41969 ( .A(n41425), .B(n11966), .X(n11749) );
  nand_x1_sg U41970 ( .A(n41426), .B(n11977), .X(n11750) );
  nand_x1_sg U41971 ( .A(n41427), .B(n11988), .X(n11751) );
  nand_x1_sg U41972 ( .A(n41428), .B(n11999), .X(n11752) );
  nand_x1_sg U41973 ( .A(n41429), .B(n12010), .X(n11753) );
  nand_x1_sg U41974 ( .A(n41430), .B(n12021), .X(n11754) );
  nand_x1_sg U41975 ( .A(n41431), .B(n12032), .X(n11755) );
  nand_x1_sg U41976 ( .A(n41432), .B(n12043), .X(n11756) );
  nand_x1_sg U41977 ( .A(n41433), .B(n12054), .X(n11757) );
  nand_x1_sg U41978 ( .A(n41434), .B(n12065), .X(n11758) );
  nand_x1_sg U41979 ( .A(n41435), .B(n12076), .X(n11759) );
  nand_x1_sg U41980 ( .A(n41436), .B(n12087), .X(n11760) );
  nand_x1_sg U41981 ( .A(n41437), .B(n12098), .X(n11761) );
  nand_x1_sg U41982 ( .A(n41438), .B(n12109), .X(n11762) );
  nand_x1_sg U41983 ( .A(n41439), .B(n12127), .X(n11771) );
  nand_x1_sg U41984 ( .A(n41440), .B(n12139), .X(n11772) );
  nand_x1_sg U41985 ( .A(n41441), .B(n12150), .X(n11773) );
  nand_x1_sg U41986 ( .A(n41442), .B(n12161), .X(n11774) );
  nand_x1_sg U41987 ( .A(n41443), .B(n12172), .X(n11775) );
  nand_x1_sg U41988 ( .A(n41444), .B(n12183), .X(n11776) );
  nand_x1_sg U41989 ( .A(n41445), .B(n12194), .X(n11777) );
  nand_x1_sg U41990 ( .A(n41446), .B(n12205), .X(n11778) );
  nand_x1_sg U41991 ( .A(n41447), .B(n12216), .X(n11779) );
  nand_x1_sg U41992 ( .A(n41448), .B(n12227), .X(n11780) );
  nand_x1_sg U41993 ( .A(n41449), .B(n12238), .X(n11781) );
  nand_x1_sg U41994 ( .A(n41450), .B(n12249), .X(n11782) );
  nand_x1_sg U41995 ( .A(n41451), .B(n12260), .X(n11783) );
  nand_x1_sg U41996 ( .A(n41452), .B(n12271), .X(n11784) );
  nand_x1_sg U41997 ( .A(n41453), .B(n12282), .X(n11785) );
  nand_x1_sg U41998 ( .A(n41454), .B(n12293), .X(n11786) );
  nand_x1_sg U41999 ( .A(n41455), .B(n12304), .X(n11787) );
  nand_x1_sg U42000 ( .A(n41456), .B(n12315), .X(n11788) );
  nand_x1_sg U42001 ( .A(n41457), .B(n12326), .X(n11789) );
  nand_x1_sg U42002 ( .A(n41458), .B(n12337), .X(n11790) );
  nand_x2_sg U42003 ( .A(n12529), .B(n12530), .X(n12528) );
  nand_x2_sg U42004 ( .A(n12535), .B(n12536), .X(n12534) );
  nand_x2_sg U42005 ( .A(n12539), .B(n12540), .X(n12538) );
  nand_x2_sg U42006 ( .A(n12543), .B(n12544), .X(n12542) );
  nand_x2_sg U42007 ( .A(n12547), .B(n12548), .X(n12546) );
  nand_x2_sg U42008 ( .A(n12551), .B(n12552), .X(n12550) );
  nand_x2_sg U42009 ( .A(n12555), .B(n12556), .X(n12554) );
  nand_x2_sg U42010 ( .A(n12559), .B(n12560), .X(n12558) );
  nand_x2_sg U42011 ( .A(n12563), .B(n12564), .X(n12562) );
  nand_x2_sg U42012 ( .A(n12567), .B(n12568), .X(n12566) );
  nand_x2_sg U42013 ( .A(n12571), .B(n12572), .X(n12570) );
  nand_x2_sg U42014 ( .A(n12575), .B(n12576), .X(n12574) );
  nand_x2_sg U42015 ( .A(n12579), .B(n12580), .X(n12578) );
  nand_x2_sg U42016 ( .A(n12583), .B(n12584), .X(n12582) );
  nand_x2_sg U42017 ( .A(n12587), .B(n12588), .X(n12586) );
  nand_x2_sg U42018 ( .A(n12591), .B(n12592), .X(n12590) );
  nand_x2_sg U42019 ( .A(n12595), .B(n12596), .X(n12594) );
  nand_x2_sg U42020 ( .A(n12599), .B(n12600), .X(n12598) );
  nand_x2_sg U42021 ( .A(n12603), .B(n12604), .X(n12602) );
  nand_x2_sg U42022 ( .A(n12607), .B(n12608), .X(n12606) );
  nand_x2_sg U42023 ( .A(n12620), .B(n12621), .X(n12619) );
  nand_x2_sg U42024 ( .A(n12624), .B(n12625), .X(n12623) );
  nand_x2_sg U42025 ( .A(n12628), .B(n12629), .X(n12627) );
  nand_x2_sg U42026 ( .A(n12633), .B(n12634), .X(n12632) );
  nand_x2_sg U42027 ( .A(n12637), .B(n12638), .X(n12636) );
  nand_x2_sg U42028 ( .A(n12642), .B(n12643), .X(n12641) );
  nand_x2_sg U42029 ( .A(n12646), .B(n12647), .X(n12645) );
  nand_x2_sg U42030 ( .A(n12650), .B(n12651), .X(n12649) );
  nand_x2_sg U42031 ( .A(n12654), .B(n12655), .X(n12653) );
  nand_x2_sg U42032 ( .A(n12658), .B(n12659), .X(n12657) );
  nand_x2_sg U42033 ( .A(n12662), .B(n12663), .X(n12661) );
  nand_x2_sg U42034 ( .A(n12666), .B(n12667), .X(n12665) );
  nand_x2_sg U42035 ( .A(n12670), .B(n12671), .X(n12669) );
  nand_x2_sg U42036 ( .A(n12674), .B(n12675), .X(n12673) );
  nand_x2_sg U42037 ( .A(n12678), .B(n12679), .X(n12677) );
  nand_x2_sg U42038 ( .A(n12682), .B(n12683), .X(n12681) );
  nand_x2_sg U42039 ( .A(n12686), .B(n12687), .X(n12685) );
  nand_x2_sg U42040 ( .A(n12690), .B(n12691), .X(n12689) );
  nand_x2_sg U42041 ( .A(n12695), .B(n12696), .X(n12694) );
  nand_x2_sg U42042 ( .A(n12700), .B(n12701), .X(n12699) );
  nand_x1_sg U42043 ( .A(n12720), .B(n12721), .X(n12719) );
  nand_x4_sg U42044 ( .A(n12732), .B(n12733), .X(n12731) );
  nand_x1_sg U42045 ( .A(n12738), .B(n12739), .X(n12737) );
  nand_x1_sg U42046 ( .A(n12756), .B(n12757), .X(n12755) );
  nand_x1_sg U42047 ( .A(n12786), .B(n12787), .X(n12785) );
  nand_x1_sg U42048 ( .A(n12798), .B(n12799), .X(n12797) );
  nand_x4_sg U42049 ( .A(n12862), .B(n12863), .X(n12861) );
  nand_x4_sg U42050 ( .A(n13792), .B(n13793), .X(n12972) );
  nand_x4_sg U42051 ( .A(n13829), .B(n13830), .X(n12980) );
  nand_x4_sg U42052 ( .A(n13860), .B(n13861), .X(n12986) );
  nand_x4_sg U42053 ( .A(n13891), .B(n13892), .X(n12992) );
  nand_x4_sg U42054 ( .A(n13922), .B(n13923), .X(n12998) );
  nand_x4_sg U42055 ( .A(n13953), .B(n13954), .X(n13004) );
  nand_x4_sg U42056 ( .A(n13984), .B(n13985), .X(n13010) );
  nand_x4_sg U42057 ( .A(n14015), .B(n14016), .X(n13016) );
  nand_x4_sg U42058 ( .A(n14046), .B(n14047), .X(n13022) );
  nand_x4_sg U42059 ( .A(n14077), .B(n14078), .X(n13028) );
  nand_x4_sg U42060 ( .A(n14108), .B(n14109), .X(n13034) );
  nand_x4_sg U42061 ( .A(n14139), .B(n14140), .X(n13040) );
  nand_x4_sg U42062 ( .A(n14170), .B(n14171), .X(n13046) );
  nand_x4_sg U42063 ( .A(n14201), .B(n14202), .X(n13052) );
  nand_x4_sg U42064 ( .A(n14232), .B(n14233), .X(n13058) );
  nand_x4_sg U42065 ( .A(n14263), .B(n14264), .X(n13064) );
  nand_x4_sg U42066 ( .A(n14294), .B(n14295), .X(n13070) );
  nand_x4_sg U42067 ( .A(n14325), .B(n14326), .X(n13076) );
  nand_x4_sg U42068 ( .A(n14356), .B(n14357), .X(n13082) );
  nand_x4_sg U42069 ( .A(n14387), .B(n14388), .X(n13088) );
  nand_x4_sg U42070 ( .A(n14419), .B(n14420), .X(n13103) );
  nand_x4_sg U42071 ( .A(n14450), .B(n14451), .X(n13111) );
  nor_x1_sg U42072 ( .A(n14498), .B(n14499), .X(n14488) );
  nand_x1_sg U42073 ( .A(n14492), .B(n14493), .X(n14491) );
  nand_x1_sg U42074 ( .A(n14482), .B(n14483), .X(n13117) );
  inv_x1_sg U42075 ( .A(n14484), .X(n41120) );
  nand_x4_sg U42076 ( .A(n14514), .B(n14515), .X(n13122) );
  nor_x1_sg U42077 ( .A(n14560), .B(n14561), .X(n14552) );
  nand_x1_sg U42078 ( .A(n14556), .B(n14557), .X(n14555) );
  nand_x4_sg U42079 ( .A(n14576), .B(n14577), .X(n13133) );
  nand_x4_sg U42080 ( .A(n14607), .B(n14608), .X(n13139) );
  nand_x4_sg U42081 ( .A(n14638), .B(n14639), .X(n13145) );
  nand_x4_sg U42082 ( .A(n14669), .B(n14670), .X(n13151) );
  nand_x4_sg U42083 ( .A(n14700), .B(n14701), .X(n13157) );
  nand_x4_sg U42084 ( .A(n14731), .B(n14732), .X(n13163) );
  nand_x4_sg U42085 ( .A(n14762), .B(n14763), .X(n13169) );
  nand_x4_sg U42086 ( .A(n14793), .B(n14794), .X(n13175) );
  nand_x4_sg U42087 ( .A(n14824), .B(n14825), .X(n13181) );
  nand_x4_sg U42088 ( .A(n14855), .B(n14856), .X(n13187) );
  nand_x4_sg U42089 ( .A(n14886), .B(n14887), .X(n13193) );
  nand_x4_sg U42090 ( .A(n14917), .B(n14918), .X(n13199) );
  nor_x1_sg U42091 ( .A(n14963), .B(n14964), .X(n14955) );
  nand_x1_sg U42092 ( .A(n14959), .B(n14960), .X(n14958) );
  nand_x1_sg U42093 ( .A(n14949), .B(n14950), .X(n13205) );
  nor_x1_sg U42094 ( .A(n14994), .B(n14995), .X(n14986) );
  nand_x1_sg U42095 ( .A(n14990), .B(n14991), .X(n14989) );
  nand_x1_sg U42096 ( .A(n14980), .B(n14981), .X(n13210) );
  nand_x4_sg U42097 ( .A(n15010), .B(n15011), .X(n13215) );
  nand_x1_sg U42098 ( .A(n41414), .B(n13229), .X(n13228) );
  nand_x1_sg U42099 ( .A(n41410), .B(n13232), .X(n13231) );
  nand_x1_sg U42100 ( .A(n41406), .B(n13235), .X(n13234) );
  nand_x1_sg U42101 ( .A(n41402), .B(n13238), .X(n13237) );
  nand_x1_sg U42102 ( .A(n41398), .B(n13241), .X(n13240) );
  nand_x1_sg U42103 ( .A(n41394), .B(n13244), .X(n13243) );
  nand_x1_sg U42104 ( .A(n41390), .B(n13247), .X(n13246) );
  nand_x1_sg U42105 ( .A(n41386), .B(n13250), .X(n13249) );
  nand_x1_sg U42106 ( .A(n41382), .B(n13253), .X(n13252) );
  nand_x1_sg U42107 ( .A(n41378), .B(n13256), .X(n13255) );
  nand_x1_sg U42108 ( .A(n41374), .B(n13259), .X(n13258) );
  nand_x1_sg U42109 ( .A(n41370), .B(n13262), .X(n13261) );
  nand_x1_sg U42110 ( .A(n41366), .B(n13265), .X(n13264) );
  nand_x1_sg U42111 ( .A(n41362), .B(n13268), .X(n13267) );
  nand_x1_sg U42112 ( .A(n41358), .B(n13271), .X(n13270) );
  nand_x1_sg U42113 ( .A(n41354), .B(n13274), .X(n13273) );
  nand_x1_sg U42114 ( .A(n41350), .B(n13277), .X(n13276) );
  nand_x1_sg U42115 ( .A(n41346), .B(n13280), .X(n13279) );
  nand_x1_sg U42116 ( .A(n41342), .B(n13283), .X(n13282) );
  nand_x1_sg U42117 ( .A(n41338), .B(n13286), .X(n13285) );
  nand_x1_sg U42118 ( .A(n41337), .B(n13295), .X(n13294) );
  nand_x1_sg U42119 ( .A(n41336), .B(n13298), .X(n13297) );
  nand_x1_sg U42120 ( .A(n41335), .B(n13305), .X(n13304) );
  nand_x1_sg U42121 ( .A(n41334), .B(n13312), .X(n13311) );
  nand_x1_sg U42122 ( .A(n41333), .B(n13315), .X(n13314) );
  nand_x1_sg U42123 ( .A(n41332), .B(n13318), .X(n13317) );
  nand_x1_sg U42124 ( .A(n41331), .B(n13321), .X(n13320) );
  nand_x1_sg U42125 ( .A(n41330), .B(n13324), .X(n13323) );
  nand_x1_sg U42126 ( .A(n41329), .B(n13327), .X(n13326) );
  nand_x1_sg U42127 ( .A(n41328), .B(n13330), .X(n13329) );
  nand_x1_sg U42128 ( .A(n41327), .B(n13333), .X(n13332) );
  nand_x1_sg U42129 ( .A(n41326), .B(n13336), .X(n13335) );
  nand_x1_sg U42130 ( .A(n41325), .B(n13339), .X(n13338) );
  nand_x1_sg U42131 ( .A(n41324), .B(n13342), .X(n13341) );
  nand_x1_sg U42132 ( .A(n41323), .B(n13345), .X(n13344) );
  nand_x1_sg U42133 ( .A(n41322), .B(n13356), .X(n13355) );
  nand_x1_sg U42134 ( .A(n13363), .B(n41414), .X(n13362) );
  nand_x1_sg U42135 ( .A(n13371), .B(n41410), .X(n13370) );
  nand_x1_sg U42136 ( .A(n13377), .B(n41406), .X(n13376) );
  nand_x1_sg U42137 ( .A(n13383), .B(n41402), .X(n13382) );
  nand_x1_sg U42138 ( .A(n13389), .B(n41398), .X(n13388) );
  nand_x1_sg U42139 ( .A(n13395), .B(n41394), .X(n13394) );
  nand_x1_sg U42140 ( .A(n13401), .B(n41390), .X(n13400) );
  nand_x1_sg U42141 ( .A(n13407), .B(n41386), .X(n13406) );
  nand_x1_sg U42142 ( .A(n13413), .B(n41382), .X(n13412) );
  nand_x1_sg U42143 ( .A(n13419), .B(n41378), .X(n13418) );
  nand_x1_sg U42144 ( .A(n13425), .B(n41374), .X(n13424) );
  nand_x1_sg U42145 ( .A(n13431), .B(n41370), .X(n13430) );
  nand_x1_sg U42146 ( .A(n13437), .B(n41366), .X(n13436) );
  nand_x1_sg U42147 ( .A(n13443), .B(n41362), .X(n13442) );
  nand_x1_sg U42148 ( .A(n13449), .B(n41358), .X(n13448) );
  nand_x1_sg U42149 ( .A(n13455), .B(n41354), .X(n13454) );
  nand_x1_sg U42150 ( .A(n13461), .B(n41350), .X(n13460) );
  nand_x1_sg U42151 ( .A(n13467), .B(n41346), .X(n13466) );
  nand_x1_sg U42152 ( .A(n13473), .B(n41342), .X(n13472) );
  nand_x1_sg U42153 ( .A(n13479), .B(n41338), .X(n13478) );
  nand_x1_sg U42154 ( .A(n13492), .B(n41337), .X(n13491) );
  nand_x1_sg U42155 ( .A(n13498), .B(n41336), .X(n13497) );
  nand_x1_sg U42156 ( .A(n13509), .B(n41335), .X(n13508) );
  nand_x1_sg U42157 ( .A(n13520), .B(n41334), .X(n13519) );
  nand_x1_sg U42158 ( .A(n13526), .B(n41333), .X(n13525) );
  nand_x1_sg U42159 ( .A(n13532), .B(n41332), .X(n13531) );
  nand_x1_sg U42160 ( .A(n13538), .B(n41331), .X(n13537) );
  nand_x1_sg U42161 ( .A(n13544), .B(n41330), .X(n13543) );
  nand_x1_sg U42162 ( .A(n13550), .B(n41329), .X(n13549) );
  nand_x1_sg U42163 ( .A(n13556), .B(n41328), .X(n13555) );
  nand_x1_sg U42164 ( .A(n13562), .B(n41327), .X(n13561) );
  nand_x1_sg U42165 ( .A(n13568), .B(n41326), .X(n13567) );
  nand_x1_sg U42166 ( .A(n13574), .B(n41325), .X(n13573) );
  nand_x1_sg U42167 ( .A(n13580), .B(n41324), .X(n13579) );
  nand_x1_sg U42168 ( .A(n13586), .B(n41323), .X(n13585) );
  nand_x1_sg U42169 ( .A(n13602), .B(n41322), .X(n13601) );
  nand_x1_sg U42170 ( .A(n13617), .B(n13618), .X(n13616) );
  nand_x1_sg U42171 ( .A(n13622), .B(n13623), .X(n13621) );
  nand_x1_sg U42172 ( .A(n13626), .B(n13627), .X(n13625) );
  nand_x1_sg U42173 ( .A(n13630), .B(n13631), .X(n13629) );
  nand_x1_sg U42174 ( .A(n13634), .B(n13635), .X(n13633) );
  nand_x1_sg U42175 ( .A(n13638), .B(n13639), .X(n13637) );
  nand_x1_sg U42176 ( .A(n13642), .B(n13643), .X(n13641) );
  nand_x1_sg U42177 ( .A(n13646), .B(n13647), .X(n13645) );
  nand_x1_sg U42178 ( .A(n13650), .B(n13651), .X(n13649) );
  nand_x1_sg U42179 ( .A(n13654), .B(n13655), .X(n13653) );
  nand_x1_sg U42180 ( .A(n13658), .B(n13659), .X(n13657) );
  nand_x1_sg U42181 ( .A(n13662), .B(n13663), .X(n13661) );
  nand_x1_sg U42182 ( .A(n13666), .B(n13667), .X(n13665) );
  nand_x1_sg U42183 ( .A(n13670), .B(n13671), .X(n13669) );
  nand_x1_sg U42184 ( .A(n13674), .B(n13675), .X(n13673) );
  nand_x1_sg U42185 ( .A(n13678), .B(n13679), .X(n13677) );
  nand_x1_sg U42186 ( .A(n13682), .B(n13683), .X(n13681) );
  nand_x1_sg U42187 ( .A(n13686), .B(n13687), .X(n13685) );
  nand_x1_sg U42188 ( .A(n13690), .B(n13691), .X(n13689) );
  nand_x1_sg U42189 ( .A(n13694), .B(n13695), .X(n13693) );
  nand_x1_sg U42190 ( .A(n13704), .B(n13705), .X(n13703) );
  nand_x1_sg U42191 ( .A(n13708), .B(n13709), .X(n13707) );
  nand_x1_sg U42192 ( .A(n41523), .B(n13712), .X(n13711) );
  nand_x1_sg U42193 ( .A(n13715), .B(n13716), .X(n13714) );
  nand_x1_sg U42194 ( .A(n41522), .B(n13719), .X(n13718) );
  nand_x1_sg U42195 ( .A(n13722), .B(n13723), .X(n13721) );
  nand_x1_sg U42196 ( .A(n13726), .B(n13727), .X(n13725) );
  nand_x1_sg U42197 ( .A(n13730), .B(n13731), .X(n13729) );
  nand_x1_sg U42198 ( .A(n13734), .B(n13735), .X(n13733) );
  nand_x1_sg U42199 ( .A(n13738), .B(n13739), .X(n13737) );
  nand_x1_sg U42200 ( .A(n13742), .B(n13743), .X(n13741) );
  nand_x1_sg U42201 ( .A(n13746), .B(n13747), .X(n13745) );
  nand_x1_sg U42202 ( .A(n13750), .B(n13751), .X(n13749) );
  nand_x1_sg U42203 ( .A(n13754), .B(n13755), .X(n13753) );
  nand_x1_sg U42204 ( .A(n13758), .B(n13759), .X(n13757) );
  nand_x1_sg U42205 ( .A(n13762), .B(n13763), .X(n13761) );
  nand_x1_sg U42206 ( .A(n13766), .B(n13767), .X(n13765) );
  nand_x1_sg U42207 ( .A(n41521), .B(n13770), .X(n13769) );
  nand_x1_sg U42208 ( .A(n41520), .B(n13773), .X(n13772) );
  nand_x1_sg U42209 ( .A(n13776), .B(n13777), .X(n13775) );
  nand_x1_sg U42210 ( .A(n13785), .B(n13617), .X(n13784) );
  nand_x1_sg U42211 ( .A(n13823), .B(n13622), .X(n13822) );
  nand_x1_sg U42212 ( .A(n13854), .B(n13626), .X(n13853) );
  nand_x1_sg U42213 ( .A(n13885), .B(n13630), .X(n13884) );
  nand_x1_sg U42214 ( .A(n13916), .B(n13634), .X(n13915) );
  nand_x1_sg U42215 ( .A(n13947), .B(n13638), .X(n13946) );
  nand_x1_sg U42216 ( .A(n13978), .B(n13642), .X(n13977) );
  nand_x1_sg U42217 ( .A(n14009), .B(n13646), .X(n14008) );
  nand_x1_sg U42218 ( .A(n14040), .B(n13650), .X(n14039) );
  nand_x1_sg U42219 ( .A(n14071), .B(n13654), .X(n14070) );
  nand_x1_sg U42220 ( .A(n14102), .B(n13658), .X(n14101) );
  nand_x1_sg U42221 ( .A(n14133), .B(n13662), .X(n14132) );
  nand_x1_sg U42222 ( .A(n14164), .B(n13666), .X(n14163) );
  nand_x1_sg U42223 ( .A(n14195), .B(n13670), .X(n14194) );
  nand_x1_sg U42224 ( .A(n14226), .B(n13674), .X(n14225) );
  nand_x1_sg U42225 ( .A(n14257), .B(n13678), .X(n14256) );
  nand_x1_sg U42226 ( .A(n14288), .B(n13682), .X(n14287) );
  nand_x1_sg U42227 ( .A(n14319), .B(n13686), .X(n14318) );
  nand_x1_sg U42228 ( .A(n14350), .B(n13690), .X(n14349) );
  nand_x1_sg U42229 ( .A(n14381), .B(n13694), .X(n14380) );
  nand_x1_sg U42230 ( .A(n14413), .B(n13704), .X(n14412) );
  nand_x1_sg U42231 ( .A(n14444), .B(n13708), .X(n14443) );
  nand_x1_sg U42232 ( .A(n14475), .B(n41523), .X(n14474) );
  nand_x1_sg U42233 ( .A(n14508), .B(n13715), .X(n14507) );
  nand_x1_sg U42234 ( .A(n14539), .B(n41522), .X(n14538) );
  nand_x1_sg U42235 ( .A(n14570), .B(n13722), .X(n14569) );
  nand_x1_sg U42236 ( .A(n14601), .B(n13726), .X(n14600) );
  nand_x1_sg U42237 ( .A(n14632), .B(n13730), .X(n14631) );
  nand_x1_sg U42238 ( .A(n14663), .B(n13734), .X(n14662) );
  nand_x1_sg U42239 ( .A(n14694), .B(n13738), .X(n14693) );
  nand_x1_sg U42240 ( .A(n14725), .B(n13742), .X(n14724) );
  nand_x1_sg U42241 ( .A(n14756), .B(n13746), .X(n14755) );
  nand_x1_sg U42242 ( .A(n14787), .B(n13750), .X(n14786) );
  nand_x1_sg U42243 ( .A(n14818), .B(n13754), .X(n14817) );
  nand_x1_sg U42244 ( .A(n14849), .B(n13758), .X(n14848) );
  nand_x1_sg U42245 ( .A(n14880), .B(n13762), .X(n14879) );
  nand_x1_sg U42246 ( .A(n14911), .B(n13766), .X(n14910) );
  nand_x1_sg U42247 ( .A(n14942), .B(n41521), .X(n14941) );
  nand_x1_sg U42248 ( .A(n14973), .B(n41520), .X(n14972) );
  nand_x1_sg U42249 ( .A(n15004), .B(n13776), .X(n15003) );
  nand_x2_sg U42250 ( .A(n15058), .B(n15059), .X(n15057) );
  nand_x1_sg U42251 ( .A(n42404), .B(n15063), .X(n15062) );
  nand_x1_sg U42252 ( .A(n15080), .B(n15081), .X(n15079) );
  nand_x1_sg U42253 ( .A(n15082), .B(n15083), .X(n15081) );
  nand_x1_sg U42254 ( .A(n15074), .B(n15075), .X(n15070) );
  nand_x1_sg U42255 ( .A(n15077), .B(n15078), .X(n15076) );
  nand_x1_sg U42256 ( .A(n15156), .B(n15157), .X(n15155) );
  nand_x2_sg U42257 ( .A(n15159), .B(n15160), .X(n15158) );
  nand_x1_sg U42258 ( .A(n15163), .B(n15164), .X(n15162) );
  nand_x1_sg U42259 ( .A(n42390), .B(n15166), .X(n15165) );
  nand_x2_sg U42260 ( .A(n15194), .B(n15195), .X(n15193) );
  nand_x1_sg U42261 ( .A(n42397), .B(n15199), .X(n15198) );
  nand_x1_sg U42262 ( .A(n15210), .B(n15211), .X(n15206) );
  nand_x1_sg U42263 ( .A(n15213), .B(n15214), .X(n15212) );
  nand_x1_sg U42264 ( .A(n20910), .B(n20911), .X(n20909) );
  nand_x1_sg U42265 ( .A(n20917), .B(n20918), .X(n20910) );
  nand_x1_sg U42266 ( .A(n33718), .B(n35448), .X(n12778) );
  nand_x1_sg U42267 ( .A(n33717), .B(n35438), .X(n12826) );
  nand_x1_sg U42268 ( .A(n33798), .B(n35425), .X(n12908) );
  nand_x1_sg U42269 ( .A(n30013), .B(n35420), .X(n12956) );
  nand_x1_sg U42270 ( .A(n33735), .B(n13261), .X(n13260) );
  nand_x1_sg U42271 ( .A(n30994), .B(n13267), .X(n13266) );
  nand_x1_sg U42272 ( .A(n30001), .B(n13285), .X(n13284) );
  nand_x1_sg U42273 ( .A(n33636), .B(n13329), .X(n13328) );
  nand_x1_sg U42274 ( .A(n35621), .B(n13355), .X(n13354) );
  nand_x1_sg U42275 ( .A(n33742), .B(n13430), .X(n13429) );
  nand_x1_sg U42276 ( .A(n33743), .B(n13442), .X(n13441) );
  nand_x1_sg U42277 ( .A(n33742), .B(n13478), .X(n13477) );
  nand_x1_sg U42278 ( .A(n29997), .B(n13555), .X(n13554) );
  nand_x1_sg U42279 ( .A(n33721), .B(n13601), .X(n13600) );
  nand_x1_sg U42280 ( .A(n33737), .B(n13661), .X(n13660) );
  nand_x1_sg U42281 ( .A(n33738), .B(n13669), .X(n13668) );
  nand_x1_sg U42282 ( .A(n30993), .B(n13693), .X(n13692) );
  nand_x1_sg U42283 ( .A(n33726), .B(n13745), .X(n13744) );
  nand_x1_sg U42284 ( .A(n33726), .B(n13775), .X(n13774) );
  nand_x1_sg U42285 ( .A(n33633), .B(n14132), .X(n14131) );
  nand_x1_sg U42286 ( .A(n33632), .B(n14194), .X(n14193) );
  nand_x1_sg U42287 ( .A(n31001), .B(n14380), .X(n14379) );
  inv_x1_sg U42288 ( .A(n15069), .X(n42403) );
  inv_x1_sg U42289 ( .A(n11852), .X(n41647) );
  inv_x1_sg U42290 ( .A(n11830), .X(n41515) );
  inv_x1_sg U42291 ( .A(n11828), .X(n41514) );
  inv_x1_sg U42292 ( .A(n11824), .X(n41512) );
  nand_x1_sg U42293 ( .A(n30996), .B(n13753), .X(n13752) );
  nand_x1_sg U42294 ( .A(n30997), .B(n13567), .X(n13566) );
  inv_x1_sg U42295 ( .A(n13073), .X(n35601) );
  inv_x1_sg U42296 ( .A(n13037), .X(n35602) );
  inv_x1_sg U42297 ( .A(n13099), .X(n35603) );
  inv_x1_sg U42298 ( .A(n13001), .X(n35604) );
  nand_x1_sg U42299 ( .A(n29993), .B(n13335), .X(n13334) );
  nand_x1_sg U42300 ( .A(n33797), .B(n35427), .X(n12920) );
  nand_x1_sg U42301 ( .A(n35622), .B(n35441), .X(n12790) );
  inv_x1_sg U42302 ( .A(n35600), .X(n35606) );
  nand_x4_sg U42303 ( .A(n15035), .B(n19580), .X(n11535) );
  inv_x1_sg U42304 ( .A(n13085), .X(n35607) );
  inv_x1_sg U42305 ( .A(n13079), .X(n35608) );
  inv_x1_sg U42306 ( .A(n13067), .X(n35609) );
  inv_x1_sg U42307 ( .A(n13061), .X(n35610) );
  inv_x1_sg U42308 ( .A(n13049), .X(n35611) );
  inv_x1_sg U42309 ( .A(n13025), .X(n35612) );
  inv_x1_sg U42310 ( .A(n12989), .X(n35613) );
  inv_x1_sg U42311 ( .A(n12977), .X(n35614) );
  nand_x4_sg U42312 ( .A(n11688), .B(n11635), .X(n11667) );
  inv_x1_sg U42313 ( .A(n33631), .X(n41321) );
  nand_x1_sg U42314 ( .A(n32884), .B(n29667), .X(n28318) );
  nand_x1_sg U42315 ( .A(n15161), .B(n35273), .X(n15089) );
  inv_x1_sg U42316 ( .A(n11826), .X(n41513) );
  inv_x1_sg U42317 ( .A(n13055), .X(n35615) );
  inv_x1_sg U42318 ( .A(n13043), .X(n35616) );
  inv_x1_sg U42319 ( .A(n13031), .X(n35617) );
  inv_x1_sg U42320 ( .A(n13019), .X(n35618) );
  inv_x1_sg U42321 ( .A(n13007), .X(n35619) );
  nand_x1_sg U42322 ( .A(n15343), .B(n35273), .X(n15095) );
  nand_x1_sg U42323 ( .A(n34420), .B(n13700), .X(n35635) );
  nand_x1_sg U42324 ( .A(n30292), .B(n13856), .X(n13855) );
  nand_x1_sg U42325 ( .A(n34219), .B(n13825), .X(n13824) );
  nand_x1_sg U42326 ( .A(n34222), .B(n13788), .X(n13786) );
  nand_x1_sg U42327 ( .A(n15348), .B(n35273), .X(n15093) );
  inv_x1_sg U42328 ( .A(n13299), .X(n41708) );
  inv_x1_sg U42329 ( .A(n13306), .X(n41710) );
  inv_x1_sg U42330 ( .A(n13346), .X(n41723) );
  inv_x1_sg U42331 ( .A(n13350), .X(n41724) );
  inv_x1_sg U42332 ( .A(n15296), .X(n42369) );
  inv_x1_sg U42333 ( .A(n15311), .X(n42386) );
  nand_x1_sg U42334 ( .A(n21342), .B(n35484), .X(n21341) );
  nand_x1_sg U42335 ( .A(n20946), .B(n20938), .X(n20945) );
  inv_x1_sg U42336 ( .A(n21186), .X(n42546) );
  inv_x1_sg U42337 ( .A(n21686), .X(n42545) );
  nand_x1_sg U42338 ( .A(n20898), .B(n20899), .X(\shifter_0/n10240 ) );
  nand_x1_sg U42339 ( .A(n19595), .B(n19596), .X(\shifter_0/n10885 ) );
  inv_x1_sg U42340 ( .A(n21565), .X(n42534) );
  inv_x1_sg U42341 ( .A(n21378), .X(n42535) );
  nand_x1_sg U42342 ( .A(n19592), .B(n19593), .X(\shifter_0/n10886 ) );
  nand_x1_sg U42343 ( .A(n31019), .B(n32929), .X(n13367) );
  nand_x1_sg U42344 ( .A(n13118), .B(n13119), .X(\shifter_0/n7185 ) );
  nand_x1_sg U42345 ( .A(n13129), .B(n13130), .X(\shifter_0/n7177 ) );
  nand_x1_sg U42346 ( .A(n13206), .B(n13207), .X(\shifter_0/n7125 ) );
  nand_x1_sg U42347 ( .A(n13211), .B(n13212), .X(\shifter_0/n7121 ) );
  inv_x1_sg U42348 ( .A(n14442), .X(n41606) );
  inv_x1_sg U42349 ( .A(n14537), .X(n41609) );
  inv_x1_sg U42350 ( .A(n14630), .X(n41612) );
  inv_x1_sg U42351 ( .A(n12710), .X(n41563) );
  inv_x1_sg U42352 ( .A(n12724), .X(n41561) );
  inv_x1_sg U42353 ( .A(n12736), .X(n41559) );
  inv_x1_sg U42354 ( .A(n12748), .X(n41557) );
  inv_x1_sg U42355 ( .A(n12760), .X(n41555) );
  inv_x1_sg U42356 ( .A(n12772), .X(n41553) );
  inv_x1_sg U42357 ( .A(n12784), .X(n41551) );
  inv_x1_sg U42358 ( .A(n12796), .X(n41549) );
  inv_x1_sg U42359 ( .A(n12802), .X(n41548) );
  inv_x1_sg U42360 ( .A(n12808), .X(n41547) );
  inv_x1_sg U42361 ( .A(n12814), .X(n41546) );
  inv_x1_sg U42362 ( .A(n12820), .X(n41545) );
  inv_x1_sg U42363 ( .A(n12826), .X(n41544) );
  inv_x1_sg U42364 ( .A(n13360), .X(n41524) );
  inv_x1_sg U42365 ( .A(n13375), .X(n41526) );
  inv_x1_sg U42366 ( .A(n13387), .X(n41528) );
  inv_x1_sg U42367 ( .A(n13399), .X(n41530) );
  inv_x1_sg U42368 ( .A(n13411), .X(n41532) );
  inv_x1_sg U42369 ( .A(n13423), .X(n41534) );
  inv_x1_sg U42370 ( .A(n13435), .X(n41536) );
  inv_x1_sg U42371 ( .A(n13447), .X(n41538) );
  inv_x1_sg U42372 ( .A(n13453), .X(n41539) );
  inv_x1_sg U42373 ( .A(n13459), .X(n41540) );
  inv_x1_sg U42374 ( .A(n13465), .X(n41541) );
  inv_x1_sg U42375 ( .A(n13471), .X(n41542) );
  inv_x1_sg U42376 ( .A(n13477), .X(n41543) );
  inv_x1_sg U42377 ( .A(n12841), .X(n41665) );
  inv_x1_sg U42378 ( .A(n12854), .X(n41667) );
  inv_x1_sg U42379 ( .A(n12866), .X(n41669) );
  inv_x1_sg U42380 ( .A(n12878), .X(n41671) );
  inv_x1_sg U42381 ( .A(n12890), .X(n41673) );
  inv_x1_sg U42382 ( .A(n12902), .X(n41675) );
  inv_x1_sg U42383 ( .A(n12914), .X(n41677) );
  inv_x1_sg U42384 ( .A(n12926), .X(n41679) );
  inv_x1_sg U42385 ( .A(n12932), .X(n41680) );
  inv_x1_sg U42386 ( .A(n12938), .X(n41681) );
  inv_x1_sg U42387 ( .A(n12944), .X(n41682) );
  inv_x1_sg U42388 ( .A(n12950), .X(n41683) );
  inv_x1_sg U42389 ( .A(n12956), .X(n41684) );
  inv_x1_sg U42390 ( .A(n12718), .X(n41562) );
  inv_x1_sg U42391 ( .A(n12730), .X(n41560) );
  inv_x1_sg U42392 ( .A(n12742), .X(n41558) );
  inv_x1_sg U42393 ( .A(n12754), .X(n41556) );
  inv_x1_sg U42394 ( .A(n12766), .X(n41554) );
  inv_x1_sg U42395 ( .A(n12778), .X(n41552) );
  inv_x1_sg U42396 ( .A(n12790), .X(n41550) );
  inv_x1_sg U42397 ( .A(n13369), .X(n41525) );
  inv_x1_sg U42398 ( .A(n13381), .X(n41527) );
  inv_x1_sg U42399 ( .A(n13393), .X(n41529) );
  inv_x1_sg U42400 ( .A(n13405), .X(n41531) );
  inv_x1_sg U42401 ( .A(n13417), .X(n41533) );
  inv_x1_sg U42402 ( .A(n13429), .X(n41535) );
  inv_x1_sg U42403 ( .A(n13441), .X(n41537) );
  inv_x1_sg U42404 ( .A(n12848), .X(n41666) );
  inv_x1_sg U42405 ( .A(n12860), .X(n41668) );
  inv_x1_sg U42406 ( .A(n12872), .X(n41670) );
  inv_x1_sg U42407 ( .A(n12884), .X(n41672) );
  inv_x1_sg U42408 ( .A(n12896), .X(n41674) );
  inv_x1_sg U42409 ( .A(n12908), .X(n41676) );
  inv_x1_sg U42410 ( .A(n12920), .X(n41678) );
  inv_x1_sg U42411 ( .A(n14410), .X(n41605) );
  inv_x1_sg U42412 ( .A(n14506), .X(n41608) );
  inv_x1_sg U42413 ( .A(n14599), .X(n41611) );
  inv_x1_sg U42414 ( .A(n14692), .X(n41614) );
  inv_x1_sg U42415 ( .A(n14754), .X(n41616) );
  inv_x1_sg U42416 ( .A(n14816), .X(n41618) );
  inv_x1_sg U42417 ( .A(n14878), .X(n41620) );
  inv_x1_sg U42418 ( .A(n14940), .X(n41622) );
  inv_x1_sg U42419 ( .A(n15002), .X(n41624) );
  inv_x1_sg U42420 ( .A(n13489), .X(n41685) );
  inv_x1_sg U42421 ( .A(n13502), .X(n41687) );
  inv_x1_sg U42422 ( .A(n13513), .X(n41689) );
  inv_x1_sg U42423 ( .A(n13524), .X(n41691) );
  inv_x1_sg U42424 ( .A(n13536), .X(n41693) );
  inv_x1_sg U42425 ( .A(n13548), .X(n41695) );
  inv_x1_sg U42426 ( .A(n13560), .X(n41697) );
  inv_x1_sg U42427 ( .A(n13572), .X(n41699) );
  inv_x1_sg U42428 ( .A(n13578), .X(n41700) );
  inv_x1_sg U42429 ( .A(n13584), .X(n41701) );
  inv_x1_sg U42430 ( .A(n13590), .X(n41702) );
  inv_x1_sg U42431 ( .A(n13595), .X(n41703) );
  inv_x1_sg U42432 ( .A(n13600), .X(n41704) );
  inv_x1_sg U42433 ( .A(n13496), .X(n41686) );
  inv_x1_sg U42434 ( .A(n13507), .X(n41688) );
  inv_x1_sg U42435 ( .A(n13518), .X(n41690) );
  inv_x1_sg U42436 ( .A(n13530), .X(n41692) );
  inv_x1_sg U42437 ( .A(n13542), .X(n41694) );
  inv_x1_sg U42438 ( .A(n13554), .X(n41696) );
  inv_x1_sg U42439 ( .A(n13566), .X(n41698) );
  inv_x1_sg U42440 ( .A(n13782), .X(n41417) );
  inv_x1_sg U42441 ( .A(n13852), .X(n41409) );
  inv_x1_sg U42442 ( .A(n13914), .X(n41401) );
  inv_x1_sg U42443 ( .A(n13976), .X(n41393) );
  inv_x1_sg U42444 ( .A(n14038), .X(n41385) );
  inv_x1_sg U42445 ( .A(n14100), .X(n41377) );
  inv_x1_sg U42446 ( .A(n14162), .X(n41369) );
  inv_x1_sg U42447 ( .A(n14224), .X(n41361) );
  inv_x1_sg U42448 ( .A(n14255), .X(n41357) );
  inv_x1_sg U42449 ( .A(n14286), .X(n41353) );
  inv_x1_sg U42450 ( .A(n14317), .X(n41349) );
  inv_x1_sg U42451 ( .A(n14348), .X(n41345) );
  inv_x1_sg U42452 ( .A(n14379), .X(n41341) );
  inv_x1_sg U42453 ( .A(n14473), .X(n41607) );
  inv_x1_sg U42454 ( .A(n14568), .X(n41610) );
  inv_x1_sg U42455 ( .A(n14661), .X(n41613) );
  inv_x1_sg U42456 ( .A(n14723), .X(n41615) );
  inv_x1_sg U42457 ( .A(n14785), .X(n41617) );
  inv_x1_sg U42458 ( .A(n14847), .X(n41619) );
  inv_x1_sg U42459 ( .A(n14909), .X(n41621) );
  inv_x1_sg U42460 ( .A(n14971), .X(n41623) );
  inv_x1_sg U42461 ( .A(n13821), .X(n41413) );
  inv_x1_sg U42462 ( .A(n13883), .X(n41405) );
  inv_x1_sg U42463 ( .A(n13945), .X(n41397) );
  inv_x1_sg U42464 ( .A(n14007), .X(n41389) );
  inv_x1_sg U42465 ( .A(n14069), .X(n41381) );
  inv_x1_sg U42466 ( .A(n14131), .X(n41373) );
  inv_x1_sg U42467 ( .A(n14193), .X(n41365) );
  nand_x1_sg U42468 ( .A(n21337), .B(n21338), .X(\shifter_0/n10234 ) );
  nand_x1_sg U42469 ( .A(n20941), .B(n20942), .X(\shifter_0/n10237 ) );
  nand_x1_sg U42470 ( .A(n21324), .B(n21325), .X(\shifter_0/n10235 ) );
  nand_x1_sg U42471 ( .A(n21327), .B(n21328), .X(n21324) );
  nand_x1_sg U42472 ( .A(n20949), .B(n20950), .X(\shifter_0/n10236 ) );
  nand_x1_sg U42473 ( .A(n20906), .B(n20951), .X(n20950) );
  nand_x1_sg U42474 ( .A(n20952), .B(n20953), .X(n20951) );
  inv_x1_sg U42475 ( .A(n15307), .X(n42380) );
  inv_x1_sg U42476 ( .A(n15292), .X(n42385) );
  inv_x1_sg U42477 ( .A(n20930), .X(n42538) );
  nand_x1_sg U42478 ( .A(n21562), .B(n21563), .X(n21561) );
  nand_x1_sg U42479 ( .A(n21564), .B(n42534), .X(n21563) );
  nand_x1_sg U42480 ( .A(n21375), .B(n21376), .X(n21374) );
  nand_x1_sg U42481 ( .A(n21377), .B(n42535), .X(n21376) );
  nand_x1_sg U42482 ( .A(n21343), .B(n21344), .X(n21342) );
  nand_x1_sg U42483 ( .A(n20947), .B(n20948), .X(n20946) );
  nand_x1_sg U42484 ( .A(n35484), .B(n21350), .X(n21349) );
  nand_x1_sg U42485 ( .A(n26197), .B(n26205), .X(n26204) );
  nand_x1_sg U42486 ( .A(n13515), .B(n13308), .X(n13514) );
  nand_x1_sg U42487 ( .A(n13504), .B(n13301), .X(n13503) );
  nand_x1_sg U42488 ( .A(n13592), .B(n13348), .X(n13591) );
  nand_x1_sg U42489 ( .A(n13597), .B(n13352), .X(n13596) );
  inv_x1_sg U42490 ( .A(n15168), .X(n42390) );
  nand_x1_sg U42491 ( .A(n12449), .B(n12450), .X(\shifter_0/n7665 ) );
  nand_x1_sg U42492 ( .A(n12511), .B(n12512), .X(\shifter_0/n7605 ) );
  nand_x1_sg U42493 ( .A(n12516), .B(n12517), .X(\shifter_0/n7601 ) );
  nand_x1_sg U42494 ( .A(n13115), .B(n13116), .X(\shifter_0/n7186 ) );
  nand_x1_sg U42495 ( .A(n13126), .B(n13127), .X(\shifter_0/n7178 ) );
  nand_x1_sg U42496 ( .A(n13203), .B(n13204), .X(\shifter_0/n7126 ) );
  nand_x1_sg U42497 ( .A(n13208), .B(n13209), .X(\shifter_0/n7122 ) );
  nand_x1_sg U42498 ( .A(n12969), .B(n12970), .X(\shifter_0/n7274 ) );
  nand_x1_sg U42499 ( .A(n12978), .B(n12979), .X(\shifter_0/n7270 ) );
  nand_x1_sg U42500 ( .A(n12984), .B(n12985), .X(\shifter_0/n7266 ) );
  nand_x1_sg U42501 ( .A(n12990), .B(n12991), .X(\shifter_0/n7262 ) );
  nand_x1_sg U42502 ( .A(n12996), .B(n12997), .X(\shifter_0/n7258 ) );
  nand_x1_sg U42503 ( .A(n13002), .B(n13003), .X(\shifter_0/n7254 ) );
  nand_x1_sg U42504 ( .A(n13008), .B(n13009), .X(\shifter_0/n7250 ) );
  nand_x1_sg U42505 ( .A(n13014), .B(n13015), .X(\shifter_0/n7246 ) );
  nand_x1_sg U42506 ( .A(n13020), .B(n13021), .X(\shifter_0/n7242 ) );
  nand_x1_sg U42507 ( .A(n13026), .B(n13027), .X(\shifter_0/n7238 ) );
  nand_x1_sg U42508 ( .A(n13032), .B(n13033), .X(\shifter_0/n7234 ) );
  nand_x1_sg U42509 ( .A(n13038), .B(n13039), .X(\shifter_0/n7230 ) );
  nand_x1_sg U42510 ( .A(n13044), .B(n13045), .X(\shifter_0/n7226 ) );
  nand_x1_sg U42511 ( .A(n13050), .B(n13051), .X(\shifter_0/n7222 ) );
  nand_x1_sg U42512 ( .A(n13056), .B(n13057), .X(\shifter_0/n7218 ) );
  nand_x1_sg U42513 ( .A(n13062), .B(n13063), .X(\shifter_0/n7214 ) );
  nand_x1_sg U42514 ( .A(n13068), .B(n13069), .X(\shifter_0/n7210 ) );
  nand_x1_sg U42515 ( .A(n13074), .B(n13075), .X(\shifter_0/n7206 ) );
  nand_x1_sg U42516 ( .A(n13080), .B(n13081), .X(\shifter_0/n7202 ) );
  nand_x1_sg U42517 ( .A(n13086), .B(n13087), .X(\shifter_0/n7198 ) );
  nand_x1_sg U42518 ( .A(n13100), .B(n13101), .X(\shifter_0/n7194 ) );
  nand_x1_sg U42519 ( .A(n13109), .B(n13110), .X(\shifter_0/n7190 ) );
  nand_x1_sg U42520 ( .A(n13120), .B(n13121), .X(\shifter_0/n7182 ) );
  nand_x1_sg U42521 ( .A(n13131), .B(n13132), .X(\shifter_0/n7174 ) );
  nand_x1_sg U42522 ( .A(n13137), .B(n13138), .X(\shifter_0/n7170 ) );
  nand_x1_sg U42523 ( .A(n13143), .B(n13144), .X(\shifter_0/n7166 ) );
  nand_x1_sg U42524 ( .A(n13149), .B(n13150), .X(\shifter_0/n7162 ) );
  nand_x1_sg U42525 ( .A(n13155), .B(n13156), .X(\shifter_0/n7158 ) );
  nand_x1_sg U42526 ( .A(n13161), .B(n13162), .X(\shifter_0/n7154 ) );
  nand_x1_sg U42527 ( .A(n13167), .B(n13168), .X(\shifter_0/n7150 ) );
  nand_x1_sg U42528 ( .A(n13173), .B(n13174), .X(\shifter_0/n7146 ) );
  nand_x1_sg U42529 ( .A(n13179), .B(n13180), .X(\shifter_0/n7142 ) );
  nand_x1_sg U42530 ( .A(n13185), .B(n13186), .X(\shifter_0/n7138 ) );
  nand_x1_sg U42531 ( .A(n13191), .B(n13192), .X(\shifter_0/n7134 ) );
  nand_x1_sg U42532 ( .A(n13197), .B(n13198), .X(\shifter_0/n7130 ) );
  nand_x1_sg U42533 ( .A(n13213), .B(n13214), .X(\shifter_0/n7118 ) );
  nand_x1_sg U42534 ( .A(n34219), .B(n13887), .X(n13886) );
  nand_x1_sg U42535 ( .A(n30292), .B(n13918), .X(n13917) );
  nand_x1_sg U42536 ( .A(n31405), .B(n13949), .X(n13948) );
  inv_x1_sg U42537 ( .A(n13614), .X(n41416) );
  inv_x1_sg U42538 ( .A(n13624), .X(n41408) );
  inv_x1_sg U42539 ( .A(n13632), .X(n41400) );
  inv_x1_sg U42540 ( .A(n13640), .X(n41392) );
  inv_x1_sg U42541 ( .A(n13648), .X(n41384) );
  inv_x1_sg U42542 ( .A(n13656), .X(n41376) );
  inv_x1_sg U42543 ( .A(n13664), .X(n41368) );
  inv_x1_sg U42544 ( .A(n13672), .X(n41360) );
  inv_x1_sg U42545 ( .A(n13676), .X(n41356) );
  inv_x1_sg U42546 ( .A(n13680), .X(n41352) );
  inv_x1_sg U42547 ( .A(n13684), .X(n41348) );
  inv_x1_sg U42548 ( .A(n13688), .X(n41344) );
  inv_x1_sg U42549 ( .A(n13692), .X(n41340) );
  inv_x1_sg U42550 ( .A(n11799), .X(n41500) );
  inv_x1_sg U42551 ( .A(n11847), .X(n41645) );
  inv_x1_sg U42552 ( .A(n13620), .X(n41412) );
  inv_x1_sg U42553 ( .A(n13628), .X(n41404) );
  inv_x1_sg U42554 ( .A(n13636), .X(n41396) );
  inv_x1_sg U42555 ( .A(n13644), .X(n41388) );
  inv_x1_sg U42556 ( .A(n13652), .X(n41380) );
  inv_x1_sg U42557 ( .A(n13660), .X(n41372) );
  inv_x1_sg U42558 ( .A(n13668), .X(n41364) );
  inv_x1_sg U42559 ( .A(n13701), .X(n41625) );
  inv_x1_sg U42560 ( .A(n13710), .X(n41627) );
  inv_x1_sg U42561 ( .A(n13717), .X(n41629) );
  inv_x1_sg U42562 ( .A(n13724), .X(n41631) );
  inv_x1_sg U42563 ( .A(n13732), .X(n41633) );
  inv_x1_sg U42564 ( .A(n13740), .X(n41635) );
  inv_x1_sg U42565 ( .A(n13748), .X(n41637) );
  inv_x1_sg U42566 ( .A(n13756), .X(n41639) );
  inv_x1_sg U42567 ( .A(n13760), .X(n41640) );
  inv_x1_sg U42568 ( .A(n13764), .X(n41641) );
  inv_x1_sg U42569 ( .A(n13768), .X(n41642) );
  inv_x1_sg U42570 ( .A(n13771), .X(n41643) );
  inv_x1_sg U42571 ( .A(n13774), .X(n41644) );
  inv_x1_sg U42572 ( .A(n13706), .X(n41626) );
  inv_x1_sg U42573 ( .A(n13713), .X(n41628) );
  inv_x1_sg U42574 ( .A(n13720), .X(n41630) );
  inv_x1_sg U42575 ( .A(n13728), .X(n41632) );
  inv_x1_sg U42576 ( .A(n13736), .X(n41634) );
  inv_x1_sg U42577 ( .A(n13744), .X(n41636) );
  inv_x1_sg U42578 ( .A(n13752), .X(n41638) );
  inv_x1_sg U42579 ( .A(n13292), .X(n41706) );
  inv_x1_sg U42580 ( .A(n13313), .X(n41712) );
  inv_x1_sg U42581 ( .A(n13319), .X(n41714) );
  inv_x1_sg U42582 ( .A(n13325), .X(n41716) );
  inv_x1_sg U42583 ( .A(n13331), .X(n41718) );
  inv_x1_sg U42584 ( .A(n13337), .X(n41720) );
  inv_x1_sg U42585 ( .A(n13340), .X(n41721) );
  inv_x1_sg U42586 ( .A(n13343), .X(n41722) );
  inv_x1_sg U42587 ( .A(n13354), .X(n41725) );
  inv_x1_sg U42588 ( .A(n13296), .X(n41707) );
  inv_x1_sg U42589 ( .A(n13303), .X(n41709) );
  inv_x1_sg U42590 ( .A(n13310), .X(n41711) );
  inv_x1_sg U42591 ( .A(n13316), .X(n41713) );
  inv_x1_sg U42592 ( .A(n13322), .X(n41715) );
  inv_x1_sg U42593 ( .A(n13328), .X(n41717) );
  inv_x1_sg U42594 ( .A(n13334), .X(n41719) );
  inv_x1_sg U42595 ( .A(n11804), .X(n41502) );
  inv_x1_sg U42596 ( .A(n11808), .X(n41504) );
  inv_x1_sg U42597 ( .A(n11812), .X(n41506) );
  inv_x1_sg U42598 ( .A(n11816), .X(n41508) );
  inv_x1_sg U42599 ( .A(n11820), .X(n41510) );
  inv_x1_sg U42600 ( .A(n11832), .X(n41516) );
  inv_x1_sg U42601 ( .A(n11834), .X(n41517) );
  inv_x1_sg U42602 ( .A(n11836), .X(n41518) );
  inv_x1_sg U42603 ( .A(n11838), .X(n41519) );
  inv_x1_sg U42604 ( .A(n13226), .X(n41415) );
  inv_x1_sg U42605 ( .A(n13233), .X(n41407) );
  inv_x1_sg U42606 ( .A(n13239), .X(n41399) );
  inv_x1_sg U42607 ( .A(n13245), .X(n41391) );
  inv_x1_sg U42608 ( .A(n13251), .X(n41383) );
  inv_x1_sg U42609 ( .A(n13257), .X(n41375) );
  inv_x1_sg U42610 ( .A(n13263), .X(n41367) );
  inv_x1_sg U42611 ( .A(n13269), .X(n41359) );
  inv_x1_sg U42612 ( .A(n13272), .X(n41355) );
  inv_x1_sg U42613 ( .A(n13275), .X(n41351) );
  inv_x1_sg U42614 ( .A(n13278), .X(n41347) );
  inv_x1_sg U42615 ( .A(n13281), .X(n41343) );
  inv_x1_sg U42616 ( .A(n13284), .X(n41339) );
  inv_x1_sg U42617 ( .A(n11856), .X(n41649) );
  inv_x1_sg U42618 ( .A(n11860), .X(n41651) );
  inv_x1_sg U42619 ( .A(n11864), .X(n41653) );
  inv_x1_sg U42620 ( .A(n11868), .X(n41655) );
  inv_x1_sg U42621 ( .A(n11872), .X(n41657) );
  inv_x1_sg U42622 ( .A(n11876), .X(n41659) );
  inv_x1_sg U42623 ( .A(n11878), .X(n41660) );
  inv_x1_sg U42624 ( .A(n11880), .X(n41661) );
  inv_x1_sg U42625 ( .A(n11882), .X(n41662) );
  inv_x1_sg U42626 ( .A(n11884), .X(n41663) );
  inv_x1_sg U42627 ( .A(n11886), .X(n41664) );
  inv_x1_sg U42628 ( .A(n11802), .X(n41501) );
  inv_x1_sg U42629 ( .A(n11806), .X(n41503) );
  inv_x1_sg U42630 ( .A(n11810), .X(n41505) );
  inv_x1_sg U42631 ( .A(n11814), .X(n41507) );
  inv_x1_sg U42632 ( .A(n11818), .X(n41509) );
  inv_x1_sg U42633 ( .A(n11822), .X(n41511) );
  inv_x1_sg U42634 ( .A(n13230), .X(n41411) );
  inv_x1_sg U42635 ( .A(n13236), .X(n41403) );
  inv_x1_sg U42636 ( .A(n13242), .X(n41395) );
  inv_x1_sg U42637 ( .A(n13248), .X(n41387) );
  inv_x1_sg U42638 ( .A(n13254), .X(n41379) );
  inv_x1_sg U42639 ( .A(n13260), .X(n41371) );
  inv_x1_sg U42640 ( .A(n13266), .X(n41363) );
  inv_x1_sg U42641 ( .A(n11850), .X(n41646) );
  inv_x1_sg U42642 ( .A(n11854), .X(n41648) );
  inv_x1_sg U42643 ( .A(n11858), .X(n41650) );
  inv_x1_sg U42644 ( .A(n11862), .X(n41652) );
  inv_x1_sg U42645 ( .A(n11866), .X(n41654) );
  inv_x1_sg U42646 ( .A(n11870), .X(n41656) );
  inv_x1_sg U42647 ( .A(n11874), .X(n41658) );
  nand_x1_sg U42648 ( .A(n21954), .B(n21953), .X(\shifter_0/n10127 ) );
  nand_x1_sg U42649 ( .A(n21956), .B(n21955), .X(\shifter_0/n10126 ) );
  nand_x1_sg U42650 ( .A(n21958), .B(n21957), .X(\shifter_0/n10125 ) );
  nand_x1_sg U42651 ( .A(n18892), .B(n18891), .X(\shifter_0/n9935 ) );
  nand_x1_sg U42652 ( .A(n18894), .B(n18893), .X(\shifter_0/n9934 ) );
  nand_x1_sg U42653 ( .A(n18896), .B(n18895), .X(\shifter_0/n9933 ) );
  nand_x1_sg U42654 ( .A(n18956), .B(n18955), .X(\shifter_0/n9903 ) );
  nand_x1_sg U42655 ( .A(n18958), .B(n18957), .X(\shifter_0/n9902 ) );
  nand_x1_sg U42656 ( .A(n18960), .B(n18959), .X(\shifter_0/n9901 ) );
  nand_x1_sg U42657 ( .A(n19212), .B(n19211), .X(\shifter_0/n9775 ) );
  nand_x1_sg U42658 ( .A(n19214), .B(n19213), .X(\shifter_0/n9774 ) );
  nand_x1_sg U42659 ( .A(n19216), .B(n19215), .X(\shifter_0/n9773 ) );
  nand_x1_sg U42660 ( .A(n19486), .B(n19485), .X(\shifter_0/n9638 ) );
  nand_x1_sg U42661 ( .A(n19488), .B(n19487), .X(\shifter_0/n9637 ) );
  nand_x1_sg U42662 ( .A(n19490), .B(n19489), .X(\shifter_0/n9636 ) );
  nand_x1_sg U42663 ( .A(n21762), .B(n21761), .X(\shifter_0/n10223 ) );
  nand_x1_sg U42664 ( .A(n21764), .B(n21763), .X(\shifter_0/n10222 ) );
  nand_x1_sg U42665 ( .A(n21766), .B(n21765), .X(\shifter_0/n10221 ) );
  nand_x1_sg U42666 ( .A(n21850), .B(n21849), .X(\shifter_0/n10179 ) );
  nand_x1_sg U42667 ( .A(n21852), .B(n21851), .X(\shifter_0/n10178 ) );
  nand_x1_sg U42668 ( .A(n21854), .B(n21853), .X(\shifter_0/n10177 ) );
  nand_x1_sg U42669 ( .A(n18762), .B(n18761), .X(\shifter_0/n9999 ) );
  nand_x1_sg U42670 ( .A(n18766), .B(n18765), .X(\shifter_0/n9998 ) );
  nand_x1_sg U42671 ( .A(n18768), .B(n18767), .X(\shifter_0/n9997 ) );
  nand_x1_sg U42672 ( .A(n19340), .B(n19339), .X(\shifter_0/n9711 ) );
  nand_x1_sg U42673 ( .A(n19342), .B(n19341), .X(\shifter_0/n9710 ) );
  nand_x1_sg U42674 ( .A(n19344), .B(n19343), .X(\shifter_0/n9709 ) );
  nand_x1_sg U42675 ( .A(n21768), .B(n21767), .X(\shifter_0/n10220 ) );
  nand_x1_sg U42676 ( .A(n21770), .B(n21769), .X(\shifter_0/n10219 ) );
  nand_x1_sg U42677 ( .A(n21772), .B(n21771), .X(\shifter_0/n10218 ) );
  nand_x1_sg U42678 ( .A(n21774), .B(n21773), .X(\shifter_0/n10217 ) );
  nand_x1_sg U42679 ( .A(n21776), .B(n21775), .X(\shifter_0/n10216 ) );
  nand_x1_sg U42680 ( .A(n21778), .B(n21777), .X(\shifter_0/n10215 ) );
  nand_x1_sg U42681 ( .A(n21780), .B(n21779), .X(\shifter_0/n10214 ) );
  nand_x1_sg U42682 ( .A(n21782), .B(n21781), .X(\shifter_0/n10213 ) );
  nand_x1_sg U42683 ( .A(n21784), .B(n21783), .X(\shifter_0/n10212 ) );
  nand_x1_sg U42684 ( .A(n21786), .B(n21785), .X(\shifter_0/n10211 ) );
  nand_x1_sg U42685 ( .A(n21788), .B(n21787), .X(\shifter_0/n10210 ) );
  nand_x1_sg U42686 ( .A(n21790), .B(n21789), .X(\shifter_0/n10209 ) );
  nand_x1_sg U42687 ( .A(n21792), .B(n21791), .X(\shifter_0/n10208 ) );
  nand_x1_sg U42688 ( .A(n21794), .B(n21793), .X(\shifter_0/n10207 ) );
  nand_x1_sg U42689 ( .A(n21796), .B(n21795), .X(\shifter_0/n10206 ) );
  nand_x1_sg U42690 ( .A(n21798), .B(n21797), .X(\shifter_0/n10205 ) );
  nand_x1_sg U42691 ( .A(n21800), .B(n21799), .X(\shifter_0/n10204 ) );
  nand_x1_sg U42692 ( .A(n21802), .B(n21801), .X(\shifter_0/n10203 ) );
  nand_x1_sg U42693 ( .A(n21804), .B(n21803), .X(\shifter_0/n10202 ) );
  nand_x1_sg U42694 ( .A(n21806), .B(n21805), .X(\shifter_0/n10201 ) );
  nand_x1_sg U42695 ( .A(n21808), .B(n21807), .X(\shifter_0/n10200 ) );
  nand_x1_sg U42696 ( .A(n21810), .B(n21809), .X(\shifter_0/n10199 ) );
  nand_x1_sg U42697 ( .A(n21812), .B(n21811), .X(\shifter_0/n10198 ) );
  nand_x1_sg U42698 ( .A(n21814), .B(n21813), .X(\shifter_0/n10197 ) );
  nand_x1_sg U42699 ( .A(n21816), .B(n21815), .X(\shifter_0/n10196 ) );
  nand_x1_sg U42700 ( .A(n21818), .B(n21817), .X(\shifter_0/n10195 ) );
  nand_x1_sg U42701 ( .A(n21820), .B(n21819), .X(\shifter_0/n10194 ) );
  nand_x1_sg U42702 ( .A(n21822), .B(n21821), .X(\shifter_0/n10193 ) );
  nand_x1_sg U42703 ( .A(n21824), .B(n21823), .X(\shifter_0/n10192 ) );
  nand_x1_sg U42704 ( .A(n21856), .B(n21855), .X(\shifter_0/n10176 ) );
  nand_x1_sg U42705 ( .A(n21858), .B(n21857), .X(\shifter_0/n10175 ) );
  nand_x1_sg U42706 ( .A(n21860), .B(n21859), .X(\shifter_0/n10174 ) );
  nand_x1_sg U42707 ( .A(n21862), .B(n21861), .X(\shifter_0/n10173 ) );
  nand_x1_sg U42708 ( .A(n21864), .B(n21863), .X(\shifter_0/n10172 ) );
  nand_x1_sg U42709 ( .A(n21866), .B(n21865), .X(\shifter_0/n10171 ) );
  nand_x1_sg U42710 ( .A(n21868), .B(n21867), .X(\shifter_0/n10170 ) );
  nand_x1_sg U42711 ( .A(n21870), .B(n21869), .X(\shifter_0/n10169 ) );
  nand_x1_sg U42712 ( .A(n21872), .B(n21871), .X(\shifter_0/n10168 ) );
  nand_x1_sg U42713 ( .A(n21874), .B(n21873), .X(\shifter_0/n10167 ) );
  nand_x1_sg U42714 ( .A(n21876), .B(n21875), .X(\shifter_0/n10166 ) );
  nand_x1_sg U42715 ( .A(n21878), .B(n21877), .X(\shifter_0/n10165 ) );
  nand_x1_sg U42716 ( .A(n21880), .B(n21879), .X(\shifter_0/n10164 ) );
  nand_x1_sg U42717 ( .A(n21882), .B(n21881), .X(\shifter_0/n10163 ) );
  nand_x1_sg U42718 ( .A(n21884), .B(n21883), .X(\shifter_0/n10162 ) );
  nand_x1_sg U42719 ( .A(n21886), .B(n21885), .X(\shifter_0/n10161 ) );
  nand_x1_sg U42720 ( .A(n21888), .B(n21887), .X(\shifter_0/n10160 ) );
  nand_x1_sg U42721 ( .A(n21930), .B(n21929), .X(\shifter_0/n10139 ) );
  nand_x1_sg U42722 ( .A(n21932), .B(n21931), .X(\shifter_0/n10138 ) );
  nand_x1_sg U42723 ( .A(n21934), .B(n21933), .X(\shifter_0/n10137 ) );
  nand_x1_sg U42724 ( .A(n21936), .B(n21935), .X(\shifter_0/n10136 ) );
  nand_x1_sg U42725 ( .A(n21938), .B(n21937), .X(\shifter_0/n10135 ) );
  nand_x1_sg U42726 ( .A(n21940), .B(n21939), .X(\shifter_0/n10134 ) );
  nand_x1_sg U42727 ( .A(n21942), .B(n21941), .X(\shifter_0/n10133 ) );
  nand_x1_sg U42728 ( .A(n21944), .B(n21943), .X(\shifter_0/n10132 ) );
  nand_x1_sg U42729 ( .A(n21946), .B(n21945), .X(\shifter_0/n10131 ) );
  nand_x1_sg U42730 ( .A(n21948), .B(n21947), .X(\shifter_0/n10130 ) );
  nand_x1_sg U42731 ( .A(n21950), .B(n21949), .X(\shifter_0/n10129 ) );
  nand_x1_sg U42732 ( .A(n21952), .B(n21951), .X(\shifter_0/n10128 ) );
  nand_x1_sg U42733 ( .A(n22018), .B(n22017), .X(\shifter_0/n10095 ) );
  nand_x1_sg U42734 ( .A(n22020), .B(n22019), .X(\shifter_0/n10094 ) );
  nand_x1_sg U42735 ( .A(n22022), .B(n22021), .X(\shifter_0/n10093 ) );
  nand_x1_sg U42736 ( .A(n22024), .B(n22023), .X(\shifter_0/n10092 ) );
  nand_x1_sg U42737 ( .A(n22026), .B(n22025), .X(\shifter_0/n10091 ) );
  nand_x1_sg U42738 ( .A(n22028), .B(n22027), .X(\shifter_0/n10090 ) );
  nand_x1_sg U42739 ( .A(n22030), .B(n22029), .X(\shifter_0/n10089 ) );
  nand_x1_sg U42740 ( .A(n22032), .B(n22031), .X(\shifter_0/n10088 ) );
  nand_x1_sg U42741 ( .A(n22034), .B(n22033), .X(\shifter_0/n10087 ) );
  nand_x1_sg U42742 ( .A(n22036), .B(n22035), .X(\shifter_0/n10086 ) );
  nand_x1_sg U42743 ( .A(n22038), .B(n22037), .X(\shifter_0/n10085 ) );
  nand_x1_sg U42744 ( .A(n22040), .B(n22039), .X(\shifter_0/n10084 ) );
  nand_x1_sg U42745 ( .A(n22042), .B(n22041), .X(\shifter_0/n10083 ) );
  nand_x1_sg U42746 ( .A(n22044), .B(n22043), .X(\shifter_0/n10082 ) );
  nand_x1_sg U42747 ( .A(n22046), .B(n22045), .X(\shifter_0/n10081 ) );
  nand_x1_sg U42748 ( .A(n22048), .B(n22047), .X(\shifter_0/n10080 ) );
  nand_x1_sg U42749 ( .A(n22090), .B(n22089), .X(\shifter_0/n10059 ) );
  nand_x1_sg U42750 ( .A(n22092), .B(n22091), .X(\shifter_0/n10058 ) );
  nand_x1_sg U42751 ( .A(n22094), .B(n22093), .X(\shifter_0/n10057 ) );
  nand_x1_sg U42752 ( .A(n22096), .B(n22095), .X(\shifter_0/n10056 ) );
  nand_x1_sg U42753 ( .A(n22098), .B(n22097), .X(\shifter_0/n10055 ) );
  nand_x1_sg U42754 ( .A(n22100), .B(n22099), .X(\shifter_0/n10054 ) );
  nand_x1_sg U42755 ( .A(n22102), .B(n22101), .X(\shifter_0/n10053 ) );
  nand_x1_sg U42756 ( .A(n22104), .B(n22103), .X(\shifter_0/n10052 ) );
  nand_x1_sg U42757 ( .A(n22106), .B(n22105), .X(\shifter_0/n10051 ) );
  nand_x1_sg U42758 ( .A(n22108), .B(n22107), .X(\shifter_0/n10050 ) );
  nand_x1_sg U42759 ( .A(n22110), .B(n22109), .X(\shifter_0/n10049 ) );
  nand_x1_sg U42760 ( .A(n22112), .B(n22111), .X(\shifter_0/n10048 ) );
  nand_x1_sg U42761 ( .A(n22114), .B(n22113), .X(\shifter_0/n10047 ) );
  nand_x1_sg U42762 ( .A(n22116), .B(n22115), .X(\shifter_0/n10046 ) );
  nand_x1_sg U42763 ( .A(n22118), .B(n22117), .X(\shifter_0/n10045 ) );
  nand_x1_sg U42764 ( .A(n22120), .B(n22119), .X(\shifter_0/n10044 ) );
  nand_x1_sg U42765 ( .A(n22122), .B(n22121), .X(\shifter_0/n10043 ) );
  nand_x1_sg U42766 ( .A(n22124), .B(n22123), .X(\shifter_0/n10042 ) );
  nand_x1_sg U42767 ( .A(n22126), .B(n22125), .X(\shifter_0/n10041 ) );
  nand_x1_sg U42768 ( .A(n22128), .B(n22127), .X(\shifter_0/n10040 ) );
  nand_x1_sg U42769 ( .A(n22130), .B(n22129), .X(\shifter_0/n10039 ) );
  nand_x1_sg U42770 ( .A(n22132), .B(n22131), .X(\shifter_0/n10038 ) );
  nand_x1_sg U42771 ( .A(n22134), .B(n22133), .X(\shifter_0/n10037 ) );
  nand_x1_sg U42772 ( .A(n22136), .B(n22135), .X(\shifter_0/n10036 ) );
  nand_x1_sg U42773 ( .A(n22138), .B(n22137), .X(\shifter_0/n10035 ) );
  nand_x1_sg U42774 ( .A(n22140), .B(n22139), .X(\shifter_0/n10034 ) );
  nand_x1_sg U42775 ( .A(n22142), .B(n22141), .X(\shifter_0/n10033 ) );
  nand_x1_sg U42776 ( .A(n22144), .B(n22143), .X(\shifter_0/n10032 ) );
  nand_x1_sg U42777 ( .A(n22146), .B(n22145), .X(\shifter_0/n10031 ) );
  nand_x1_sg U42778 ( .A(n22148), .B(n22147), .X(\shifter_0/n10030 ) );
  nand_x1_sg U42779 ( .A(n22150), .B(n22149), .X(\shifter_0/n10029 ) );
  nand_x1_sg U42780 ( .A(n22152), .B(n22151), .X(\shifter_0/n10028 ) );
  nand_x1_sg U42781 ( .A(n22154), .B(n22153), .X(\shifter_0/n10027 ) );
  nand_x1_sg U42782 ( .A(n22156), .B(n22155), .X(\shifter_0/n10026 ) );
  nand_x1_sg U42783 ( .A(n22158), .B(n22157), .X(\shifter_0/n10025 ) );
  nand_x1_sg U42784 ( .A(n22160), .B(n22159), .X(\shifter_0/n10024 ) );
  nand_x1_sg U42785 ( .A(n22162), .B(n22161), .X(\shifter_0/n10023 ) );
  nand_x1_sg U42786 ( .A(n22164), .B(n22163), .X(\shifter_0/n10022 ) );
  nand_x1_sg U42787 ( .A(n22166), .B(n22165), .X(\shifter_0/n10021 ) );
  nand_x1_sg U42788 ( .A(n22168), .B(n22167), .X(\shifter_0/n10020 ) );
  nand_x1_sg U42789 ( .A(n22170), .B(n22169), .X(\shifter_0/n10019 ) );
  nand_x1_sg U42790 ( .A(n22172), .B(n22171), .X(\shifter_0/n10018 ) );
  nand_x1_sg U42791 ( .A(n22174), .B(n22173), .X(\shifter_0/n10017 ) );
  nand_x1_sg U42792 ( .A(n22176), .B(n22175), .X(\shifter_0/n10016 ) );
  nand_x1_sg U42793 ( .A(n22178), .B(n22177), .X(\shifter_0/n10015 ) );
  nand_x1_sg U42794 ( .A(n22180), .B(n22179), .X(\shifter_0/n10014 ) );
  nand_x1_sg U42795 ( .A(n22182), .B(n22181), .X(\shifter_0/n10013 ) );
  nand_x1_sg U42796 ( .A(n22184), .B(n22183), .X(\shifter_0/n10012 ) );
  nand_x1_sg U42797 ( .A(n22186), .B(n22185), .X(\shifter_0/n10011 ) );
  nand_x1_sg U42798 ( .A(n22188), .B(n22187), .X(\shifter_0/n10010 ) );
  nand_x1_sg U42799 ( .A(n22190), .B(n22189), .X(\shifter_0/n10009 ) );
  nand_x1_sg U42800 ( .A(n22192), .B(n22191), .X(\shifter_0/n10008 ) );
  nand_x1_sg U42801 ( .A(n22194), .B(n22193), .X(\shifter_0/n10007 ) );
  nand_x1_sg U42802 ( .A(n22196), .B(n22195), .X(\shifter_0/n10006 ) );
  nand_x1_sg U42803 ( .A(n22198), .B(n22197), .X(\shifter_0/n10005 ) );
  nand_x1_sg U42804 ( .A(n22200), .B(n22199), .X(\shifter_0/n10004 ) );
  nand_x1_sg U42805 ( .A(n22202), .B(n22201), .X(\shifter_0/n10003 ) );
  nand_x1_sg U42806 ( .A(n22204), .B(n22203), .X(\shifter_0/n10002 ) );
  nand_x1_sg U42807 ( .A(n22206), .B(n22205), .X(\shifter_0/n10001 ) );
  nand_x1_sg U42808 ( .A(n22208), .B(n22207), .X(\shifter_0/n10000 ) );
  nand_x1_sg U42809 ( .A(n18770), .B(n18769), .X(\shifter_0/n9996 ) );
  nand_x1_sg U42810 ( .A(n18772), .B(n18771), .X(\shifter_0/n9995 ) );
  nand_x1_sg U42811 ( .A(n18774), .B(n18773), .X(\shifter_0/n9994 ) );
  nand_x1_sg U42812 ( .A(n18776), .B(n18775), .X(\shifter_0/n9993 ) );
  nand_x1_sg U42813 ( .A(n18778), .B(n18777), .X(\shifter_0/n9992 ) );
  nand_x1_sg U42814 ( .A(n18780), .B(n18779), .X(\shifter_0/n9991 ) );
  nand_x1_sg U42815 ( .A(n18782), .B(n18781), .X(\shifter_0/n9990 ) );
  nand_x1_sg U42816 ( .A(n18784), .B(n18783), .X(\shifter_0/n9989 ) );
  nand_x1_sg U42817 ( .A(n18786), .B(n18785), .X(\shifter_0/n9988 ) );
  nand_x1_sg U42818 ( .A(n18788), .B(n18787), .X(\shifter_0/n9987 ) );
  nand_x1_sg U42819 ( .A(n18790), .B(n18789), .X(\shifter_0/n9986 ) );
  nand_x1_sg U42820 ( .A(n18792), .B(n18791), .X(\shifter_0/n9985 ) );
  nand_x1_sg U42821 ( .A(n18794), .B(n18793), .X(\shifter_0/n9984 ) );
  nand_x1_sg U42822 ( .A(n18796), .B(n18795), .X(\shifter_0/n9983 ) );
  nand_x1_sg U42823 ( .A(n18798), .B(n18797), .X(\shifter_0/n9982 ) );
  nand_x1_sg U42824 ( .A(n18800), .B(n18799), .X(\shifter_0/n9981 ) );
  nand_x1_sg U42825 ( .A(n18802), .B(n18801), .X(\shifter_0/n9980 ) );
  nand_x1_sg U42826 ( .A(n18844), .B(n18843), .X(\shifter_0/n9959 ) );
  nand_x1_sg U42827 ( .A(n18846), .B(n18845), .X(\shifter_0/n9958 ) );
  nand_x1_sg U42828 ( .A(n18848), .B(n18847), .X(\shifter_0/n9957 ) );
  nand_x1_sg U42829 ( .A(n18850), .B(n18849), .X(\shifter_0/n9956 ) );
  nand_x1_sg U42830 ( .A(n18852), .B(n18851), .X(\shifter_0/n9955 ) );
  nand_x1_sg U42831 ( .A(n18854), .B(n18853), .X(\shifter_0/n9954 ) );
  nand_x1_sg U42832 ( .A(n18856), .B(n18855), .X(\shifter_0/n9953 ) );
  nand_x1_sg U42833 ( .A(n18858), .B(n18857), .X(\shifter_0/n9952 ) );
  nand_x1_sg U42834 ( .A(n18860), .B(n18859), .X(\shifter_0/n9951 ) );
  nand_x1_sg U42835 ( .A(n18862), .B(n18861), .X(\shifter_0/n9950 ) );
  nand_x1_sg U42836 ( .A(n18864), .B(n18863), .X(\shifter_0/n9949 ) );
  nand_x1_sg U42837 ( .A(n18866), .B(n18865), .X(\shifter_0/n9948 ) );
  nand_x1_sg U42838 ( .A(n18868), .B(n18867), .X(\shifter_0/n9947 ) );
  nand_x1_sg U42839 ( .A(n18870), .B(n18869), .X(\shifter_0/n9946 ) );
  nand_x1_sg U42840 ( .A(n18872), .B(n18871), .X(\shifter_0/n9945 ) );
  nand_x1_sg U42841 ( .A(n18874), .B(n18873), .X(\shifter_0/n9944 ) );
  nand_x1_sg U42842 ( .A(n18876), .B(n18875), .X(\shifter_0/n9943 ) );
  nand_x1_sg U42843 ( .A(n18878), .B(n18877), .X(\shifter_0/n9942 ) );
  nand_x1_sg U42844 ( .A(n18880), .B(n18879), .X(\shifter_0/n9941 ) );
  nand_x1_sg U42845 ( .A(n18882), .B(n18881), .X(\shifter_0/n9940 ) );
  nand_x1_sg U42846 ( .A(n18884), .B(n18883), .X(\shifter_0/n9939 ) );
  nand_x1_sg U42847 ( .A(n18886), .B(n18885), .X(\shifter_0/n9938 ) );
  nand_x1_sg U42848 ( .A(n18888), .B(n18887), .X(\shifter_0/n9937 ) );
  nand_x1_sg U42849 ( .A(n18890), .B(n18889), .X(\shifter_0/n9936 ) );
  nand_x1_sg U42850 ( .A(n18950), .B(n18949), .X(\shifter_0/n9906 ) );
  nand_x1_sg U42851 ( .A(n18952), .B(n18951), .X(\shifter_0/n9905 ) );
  nand_x1_sg U42852 ( .A(n18954), .B(n18953), .X(\shifter_0/n9904 ) );
  nand_x1_sg U42853 ( .A(n19044), .B(n19043), .X(\shifter_0/n9859 ) );
  nand_x1_sg U42854 ( .A(n19046), .B(n19045), .X(\shifter_0/n9858 ) );
  nand_x1_sg U42855 ( .A(n19048), .B(n19047), .X(\shifter_0/n9857 ) );
  nand_x1_sg U42856 ( .A(n19050), .B(n19049), .X(\shifter_0/n9856 ) );
  nand_x1_sg U42857 ( .A(n19052), .B(n19051), .X(\shifter_0/n9855 ) );
  nand_x1_sg U42858 ( .A(n19054), .B(n19053), .X(\shifter_0/n9854 ) );
  nand_x1_sg U42859 ( .A(n19056), .B(n19055), .X(\shifter_0/n9853 ) );
  nand_x1_sg U42860 ( .A(n19058), .B(n19057), .X(\shifter_0/n9852 ) );
  nand_x1_sg U42861 ( .A(n19060), .B(n19059), .X(\shifter_0/n9851 ) );
  nand_x1_sg U42862 ( .A(n19062), .B(n19061), .X(\shifter_0/n9850 ) );
  nand_x1_sg U42863 ( .A(n19064), .B(n19063), .X(\shifter_0/n9849 ) );
  nand_x1_sg U42864 ( .A(n19066), .B(n19065), .X(\shifter_0/n9848 ) );
  nand_x1_sg U42865 ( .A(n19068), .B(n19067), .X(\shifter_0/n9847 ) );
  nand_x1_sg U42866 ( .A(n19070), .B(n19069), .X(\shifter_0/n9846 ) );
  nand_x1_sg U42867 ( .A(n19072), .B(n19071), .X(\shifter_0/n9845 ) );
  nand_x1_sg U42868 ( .A(n19074), .B(n19073), .X(\shifter_0/n9844 ) );
  nand_x1_sg U42869 ( .A(n19076), .B(n19075), .X(\shifter_0/n9843 ) );
  nand_x1_sg U42870 ( .A(n19078), .B(n19077), .X(\shifter_0/n9842 ) );
  nand_x1_sg U42871 ( .A(n19080), .B(n19079), .X(\shifter_0/n9841 ) );
  nand_x1_sg U42872 ( .A(n19082), .B(n19081), .X(\shifter_0/n9840 ) );
  nand_x1_sg U42873 ( .A(n19124), .B(n19123), .X(\shifter_0/n9819 ) );
  nand_x1_sg U42874 ( .A(n19126), .B(n19125), .X(\shifter_0/n9818 ) );
  nand_x1_sg U42875 ( .A(n19128), .B(n19127), .X(\shifter_0/n9817 ) );
  nand_x1_sg U42876 ( .A(n19130), .B(n19129), .X(\shifter_0/n9816 ) );
  nand_x1_sg U42877 ( .A(n19132), .B(n19131), .X(\shifter_0/n9815 ) );
  nand_x1_sg U42878 ( .A(n19134), .B(n19133), .X(\shifter_0/n9814 ) );
  nand_x1_sg U42879 ( .A(n19136), .B(n19135), .X(\shifter_0/n9813 ) );
  nand_x1_sg U42880 ( .A(n19138), .B(n19137), .X(\shifter_0/n9812 ) );
  nand_x1_sg U42881 ( .A(n19140), .B(n19139), .X(\shifter_0/n9811 ) );
  nand_x1_sg U42882 ( .A(n19142), .B(n19141), .X(\shifter_0/n9810 ) );
  nand_x1_sg U42883 ( .A(n19144), .B(n19143), .X(\shifter_0/n9809 ) );
  nand_x1_sg U42884 ( .A(n19146), .B(n19145), .X(\shifter_0/n9808 ) );
  nand_x1_sg U42885 ( .A(n19148), .B(n19147), .X(\shifter_0/n9807 ) );
  nand_x1_sg U42886 ( .A(n19150), .B(n19149), .X(\shifter_0/n9806 ) );
  nand_x1_sg U42887 ( .A(n19152), .B(n19151), .X(\shifter_0/n9805 ) );
  nand_x1_sg U42888 ( .A(n19154), .B(n19153), .X(\shifter_0/n9804 ) );
  nand_x1_sg U42889 ( .A(n19156), .B(n19155), .X(\shifter_0/n9803 ) );
  nand_x1_sg U42890 ( .A(n19158), .B(n19157), .X(\shifter_0/n9802 ) );
  nand_x1_sg U42891 ( .A(n19160), .B(n19159), .X(\shifter_0/n9801 ) );
  nand_x1_sg U42892 ( .A(n19162), .B(n19161), .X(\shifter_0/n9800 ) );
  nand_x1_sg U42893 ( .A(n19204), .B(n19203), .X(\shifter_0/n9779 ) );
  nand_x1_sg U42894 ( .A(n19206), .B(n19205), .X(\shifter_0/n9778 ) );
  nand_x1_sg U42895 ( .A(n19208), .B(n19207), .X(\shifter_0/n9777 ) );
  nand_x1_sg U42896 ( .A(n19210), .B(n19209), .X(\shifter_0/n9776 ) );
  nand_x1_sg U42897 ( .A(n19276), .B(n19275), .X(\shifter_0/n9743 ) );
  nand_x1_sg U42898 ( .A(n19278), .B(n19277), .X(\shifter_0/n9742 ) );
  nand_x1_sg U42899 ( .A(n19280), .B(n19279), .X(\shifter_0/n9741 ) );
  nand_x1_sg U42900 ( .A(n19282), .B(n19281), .X(\shifter_0/n9740 ) );
  nand_x1_sg U42901 ( .A(n19284), .B(n19283), .X(\shifter_0/n9739 ) );
  nand_x1_sg U42902 ( .A(n19286), .B(n19285), .X(\shifter_0/n9738 ) );
  nand_x1_sg U42903 ( .A(n19288), .B(n19287), .X(\shifter_0/n9737 ) );
  nand_x1_sg U42904 ( .A(n19290), .B(n19289), .X(\shifter_0/n9736 ) );
  nand_x1_sg U42905 ( .A(n19292), .B(n19291), .X(\shifter_0/n9735 ) );
  nand_x1_sg U42906 ( .A(n19294), .B(n19293), .X(\shifter_0/n9734 ) );
  nand_x1_sg U42907 ( .A(n19296), .B(n19295), .X(\shifter_0/n9733 ) );
  nand_x1_sg U42908 ( .A(n19298), .B(n19297), .X(\shifter_0/n9732 ) );
  nand_x1_sg U42909 ( .A(n19300), .B(n19299), .X(\shifter_0/n9731 ) );
  nand_x1_sg U42910 ( .A(n19302), .B(n19301), .X(\shifter_0/n9730 ) );
  nand_x1_sg U42911 ( .A(n19304), .B(n19303), .X(\shifter_0/n9729 ) );
  nand_x1_sg U42912 ( .A(n19306), .B(n19305), .X(\shifter_0/n9728 ) );
  nand_x1_sg U42913 ( .A(n19308), .B(n19307), .X(\shifter_0/n9727 ) );
  nand_x1_sg U42914 ( .A(n19310), .B(n19309), .X(\shifter_0/n9726 ) );
  nand_x1_sg U42915 ( .A(n19312), .B(n19311), .X(\shifter_0/n9725 ) );
  nand_x1_sg U42916 ( .A(n19314), .B(n19313), .X(\shifter_0/n9724 ) );
  nand_x1_sg U42917 ( .A(n19316), .B(n19315), .X(\shifter_0/n9723 ) );
  nand_x1_sg U42918 ( .A(n19318), .B(n19317), .X(\shifter_0/n9722 ) );
  nand_x1_sg U42919 ( .A(n19320), .B(n19319), .X(\shifter_0/n9721 ) );
  nand_x1_sg U42920 ( .A(n19322), .B(n19321), .X(\shifter_0/n9720 ) );
  nand_x1_sg U42921 ( .A(n19324), .B(n19323), .X(\shifter_0/n9719 ) );
  nand_x1_sg U42922 ( .A(n19326), .B(n19325), .X(\shifter_0/n9718 ) );
  nand_x1_sg U42923 ( .A(n19328), .B(n19327), .X(\shifter_0/n9717 ) );
  nand_x1_sg U42924 ( .A(n19330), .B(n19329), .X(\shifter_0/n9716 ) );
  nand_x1_sg U42925 ( .A(n19332), .B(n19331), .X(\shifter_0/n9715 ) );
  nand_x1_sg U42926 ( .A(n19334), .B(n19333), .X(\shifter_0/n9714 ) );
  nand_x1_sg U42927 ( .A(n19336), .B(n19335), .X(\shifter_0/n9713 ) );
  nand_x1_sg U42928 ( .A(n19338), .B(n19337), .X(\shifter_0/n9712 ) );
  nand_x1_sg U42929 ( .A(n19346), .B(n19345), .X(\shifter_0/n9708 ) );
  nand_x1_sg U42930 ( .A(n19348), .B(n19347), .X(\shifter_0/n9707 ) );
  nand_x1_sg U42931 ( .A(n19350), .B(n19349), .X(\shifter_0/n9706 ) );
  nand_x1_sg U42932 ( .A(n19352), .B(n19351), .X(\shifter_0/n9705 ) );
  nand_x1_sg U42933 ( .A(n19354), .B(n19353), .X(\shifter_0/n9704 ) );
  nand_x1_sg U42934 ( .A(n19356), .B(n19355), .X(\shifter_0/n9703 ) );
  nand_x1_sg U42935 ( .A(n19358), .B(n19357), .X(\shifter_0/n9702 ) );
  nand_x1_sg U42936 ( .A(n19360), .B(n19359), .X(\shifter_0/n9701 ) );
  nand_x1_sg U42937 ( .A(n19362), .B(n19361), .X(\shifter_0/n9700 ) );
  nand_x1_sg U42938 ( .A(n19404), .B(n19403), .X(\shifter_0/n9679 ) );
  nand_x1_sg U42939 ( .A(n19406), .B(n19405), .X(\shifter_0/n9678 ) );
  nand_x1_sg U42940 ( .A(n19408), .B(n19407), .X(\shifter_0/n9677 ) );
  nand_x1_sg U42941 ( .A(n19410), .B(n19409), .X(\shifter_0/n9676 ) );
  nand_x1_sg U42942 ( .A(n19412), .B(n19411), .X(\shifter_0/n9675 ) );
  nand_x1_sg U42943 ( .A(n19414), .B(n19413), .X(\shifter_0/n9674 ) );
  nand_x1_sg U42944 ( .A(n19416), .B(n19415), .X(\shifter_0/n9673 ) );
  nand_x1_sg U42945 ( .A(n19418), .B(n19417), .X(\shifter_0/n9672 ) );
  nand_x1_sg U42946 ( .A(n19420), .B(n19419), .X(\shifter_0/n9671 ) );
  nand_x1_sg U42947 ( .A(n19422), .B(n19421), .X(\shifter_0/n9670 ) );
  nand_x1_sg U42948 ( .A(n19424), .B(n19423), .X(\shifter_0/n9669 ) );
  nand_x1_sg U42949 ( .A(n19426), .B(n19425), .X(\shifter_0/n9668 ) );
  nand_x1_sg U42950 ( .A(n19428), .B(n19427), .X(\shifter_0/n9667 ) );
  nand_x1_sg U42951 ( .A(n19430), .B(n19429), .X(\shifter_0/n9666 ) );
  nand_x1_sg U42952 ( .A(n19432), .B(n19431), .X(\shifter_0/n9665 ) );
  nand_x1_sg U42953 ( .A(n19434), .B(n19433), .X(\shifter_0/n9664 ) );
  nand_x1_sg U42954 ( .A(n19436), .B(n19435), .X(\shifter_0/n9663 ) );
  nand_x1_sg U42955 ( .A(n19438), .B(n19437), .X(\shifter_0/n9662 ) );
  nand_x1_sg U42956 ( .A(n19440), .B(n19439), .X(\shifter_0/n9661 ) );
  nand_x1_sg U42957 ( .A(n19442), .B(n19441), .X(\shifter_0/n9660 ) );
  nand_x1_sg U42958 ( .A(n19484), .B(n19483), .X(\shifter_0/n9639 ) );
  nand_x1_sg U42959 ( .A(n21746), .B(n21745), .X(\shifter_0/n10231 ) );
  nand_x1_sg U42960 ( .A(n21748), .B(n21747), .X(\shifter_0/n10230 ) );
  nand_x1_sg U42961 ( .A(n21750), .B(n21749), .X(\shifter_0/n10229 ) );
  nand_x1_sg U42962 ( .A(n21752), .B(n21751), .X(\shifter_0/n10228 ) );
  nand_x1_sg U42963 ( .A(n21754), .B(n21753), .X(\shifter_0/n10227 ) );
  nand_x1_sg U42964 ( .A(n21756), .B(n21755), .X(\shifter_0/n10226 ) );
  nand_x1_sg U42965 ( .A(n21758), .B(n21757), .X(\shifter_0/n10225 ) );
  nand_x1_sg U42966 ( .A(n21760), .B(n21759), .X(\shifter_0/n10224 ) );
  nand_x1_sg U42967 ( .A(n21826), .B(n21825), .X(\shifter_0/n10191 ) );
  nand_x1_sg U42968 ( .A(n21828), .B(n21827), .X(\shifter_0/n10190 ) );
  nand_x1_sg U42969 ( .A(n21830), .B(n21829), .X(\shifter_0/n10189 ) );
  nand_x1_sg U42970 ( .A(n21832), .B(n21831), .X(\shifter_0/n10188 ) );
  nand_x1_sg U42971 ( .A(n21834), .B(n21833), .X(\shifter_0/n10187 ) );
  nand_x1_sg U42972 ( .A(n21836), .B(n21835), .X(\shifter_0/n10186 ) );
  nand_x1_sg U42973 ( .A(n21838), .B(n21837), .X(\shifter_0/n10185 ) );
  nand_x1_sg U42974 ( .A(n21840), .B(n21839), .X(\shifter_0/n10184 ) );
  nand_x1_sg U42975 ( .A(n21842), .B(n21841), .X(\shifter_0/n10183 ) );
  nand_x1_sg U42976 ( .A(n21844), .B(n21843), .X(\shifter_0/n10182 ) );
  nand_x1_sg U42977 ( .A(n21846), .B(n21845), .X(\shifter_0/n10181 ) );
  nand_x1_sg U42978 ( .A(n21848), .B(n21847), .X(\shifter_0/n10180 ) );
  nand_x1_sg U42979 ( .A(n21960), .B(n21959), .X(\shifter_0/n10124 ) );
  nand_x1_sg U42980 ( .A(n21962), .B(n21961), .X(\shifter_0/n10123 ) );
  nand_x1_sg U42981 ( .A(n21964), .B(n21963), .X(\shifter_0/n10122 ) );
  nand_x1_sg U42982 ( .A(n21966), .B(n21965), .X(\shifter_0/n10121 ) );
  nand_x1_sg U42983 ( .A(n21968), .B(n21967), .X(\shifter_0/n10120 ) );
  nand_x1_sg U42984 ( .A(n22010), .B(n22009), .X(\shifter_0/n10099 ) );
  nand_x1_sg U42985 ( .A(n22012), .B(n22011), .X(\shifter_0/n10098 ) );
  nand_x1_sg U42986 ( .A(n22014), .B(n22013), .X(\shifter_0/n10097 ) );
  nand_x1_sg U42987 ( .A(n22016), .B(n22015), .X(\shifter_0/n10096 ) );
  nand_x1_sg U42988 ( .A(n18898), .B(n18897), .X(\shifter_0/n9932 ) );
  nand_x1_sg U42989 ( .A(n18900), .B(n18899), .X(\shifter_0/n9931 ) );
  nand_x1_sg U42990 ( .A(n18902), .B(n18901), .X(\shifter_0/n9930 ) );
  nand_x1_sg U42991 ( .A(n18904), .B(n18903), .X(\shifter_0/n9929 ) );
  nand_x1_sg U42992 ( .A(n18906), .B(n18905), .X(\shifter_0/n9928 ) );
  nand_x1_sg U42993 ( .A(n18908), .B(n18907), .X(\shifter_0/n9927 ) );
  nand_x1_sg U42994 ( .A(n18910), .B(n18909), .X(\shifter_0/n9926 ) );
  nand_x1_sg U42995 ( .A(n18912), .B(n18911), .X(\shifter_0/n9925 ) );
  nand_x1_sg U42996 ( .A(n18914), .B(n18913), .X(\shifter_0/n9924 ) );
  nand_x1_sg U42997 ( .A(n18916), .B(n18915), .X(\shifter_0/n9923 ) );
  nand_x1_sg U42998 ( .A(n18918), .B(n18917), .X(\shifter_0/n9922 ) );
  nand_x1_sg U42999 ( .A(n18920), .B(n18919), .X(\shifter_0/n9921 ) );
  nand_x1_sg U43000 ( .A(n18922), .B(n18921), .X(\shifter_0/n9920 ) );
  nand_x1_sg U43001 ( .A(n18924), .B(n18923), .X(\shifter_0/n9919 ) );
  nand_x1_sg U43002 ( .A(n18926), .B(n18925), .X(\shifter_0/n9918 ) );
  nand_x1_sg U43003 ( .A(n18928), .B(n18927), .X(\shifter_0/n9917 ) );
  nand_x1_sg U43004 ( .A(n18930), .B(n18929), .X(\shifter_0/n9916 ) );
  nand_x1_sg U43005 ( .A(n18932), .B(n18931), .X(\shifter_0/n9915 ) );
  nand_x1_sg U43006 ( .A(n18934), .B(n18933), .X(\shifter_0/n9914 ) );
  nand_x1_sg U43007 ( .A(n18936), .B(n18935), .X(\shifter_0/n9913 ) );
  nand_x1_sg U43008 ( .A(n18938), .B(n18937), .X(\shifter_0/n9912 ) );
  nand_x1_sg U43009 ( .A(n18940), .B(n18939), .X(\shifter_0/n9911 ) );
  nand_x1_sg U43010 ( .A(n18942), .B(n18941), .X(\shifter_0/n9910 ) );
  nand_x1_sg U43011 ( .A(n18944), .B(n18943), .X(\shifter_0/n9909 ) );
  nand_x1_sg U43012 ( .A(n18946), .B(n18945), .X(\shifter_0/n9908 ) );
  nand_x1_sg U43013 ( .A(n18948), .B(n18947), .X(\shifter_0/n9907 ) );
  nand_x1_sg U43014 ( .A(n18962), .B(n18961), .X(\shifter_0/n9900 ) );
  nand_x1_sg U43015 ( .A(n18964), .B(n18963), .X(\shifter_0/n9899 ) );
  nand_x1_sg U43016 ( .A(n18966), .B(n18965), .X(\shifter_0/n9898 ) );
  nand_x1_sg U43017 ( .A(n18968), .B(n18967), .X(\shifter_0/n9897 ) );
  nand_x1_sg U43018 ( .A(n18970), .B(n18969), .X(\shifter_0/n9896 ) );
  nand_x1_sg U43019 ( .A(n18972), .B(n18971), .X(\shifter_0/n9895 ) );
  nand_x1_sg U43020 ( .A(n18974), .B(n18973), .X(\shifter_0/n9894 ) );
  nand_x1_sg U43021 ( .A(n18976), .B(n18975), .X(\shifter_0/n9893 ) );
  nand_x1_sg U43022 ( .A(n18978), .B(n18977), .X(\shifter_0/n9892 ) );
  nand_x1_sg U43023 ( .A(n18980), .B(n18979), .X(\shifter_0/n9891 ) );
  nand_x1_sg U43024 ( .A(n18982), .B(n18981), .X(\shifter_0/n9890 ) );
  nand_x1_sg U43025 ( .A(n18984), .B(n18983), .X(\shifter_0/n9889 ) );
  nand_x1_sg U43026 ( .A(n18986), .B(n18985), .X(\shifter_0/n9888 ) );
  nand_x1_sg U43027 ( .A(n18988), .B(n18987), .X(\shifter_0/n9887 ) );
  nand_x1_sg U43028 ( .A(n18990), .B(n18989), .X(\shifter_0/n9886 ) );
  nand_x1_sg U43029 ( .A(n18992), .B(n18991), .X(\shifter_0/n9885 ) );
  nand_x1_sg U43030 ( .A(n18994), .B(n18993), .X(\shifter_0/n9884 ) );
  nand_x1_sg U43031 ( .A(n18996), .B(n18995), .X(\shifter_0/n9883 ) );
  nand_x1_sg U43032 ( .A(n18998), .B(n18997), .X(\shifter_0/n9882 ) );
  nand_x1_sg U43033 ( .A(n19000), .B(n18999), .X(\shifter_0/n9881 ) );
  nand_x1_sg U43034 ( .A(n19002), .B(n19001), .X(\shifter_0/n9880 ) );
  nand_x1_sg U43035 ( .A(n19218), .B(n19217), .X(\shifter_0/n9772 ) );
  nand_x1_sg U43036 ( .A(n19220), .B(n19219), .X(\shifter_0/n9771 ) );
  nand_x1_sg U43037 ( .A(n19222), .B(n19221), .X(\shifter_0/n9770 ) );
  nand_x1_sg U43038 ( .A(n19224), .B(n19223), .X(\shifter_0/n9769 ) );
  nand_x1_sg U43039 ( .A(n19226), .B(n19225), .X(\shifter_0/n9768 ) );
  nand_x1_sg U43040 ( .A(n19228), .B(n19227), .X(\shifter_0/n9767 ) );
  nand_x1_sg U43041 ( .A(n19230), .B(n19229), .X(\shifter_0/n9766 ) );
  nand_x1_sg U43042 ( .A(n19232), .B(n19231), .X(\shifter_0/n9765 ) );
  nand_x1_sg U43043 ( .A(n19234), .B(n19233), .X(\shifter_0/n9764 ) );
  nand_x1_sg U43044 ( .A(n19236), .B(n19235), .X(\shifter_0/n9763 ) );
  nand_x1_sg U43045 ( .A(n19238), .B(n19237), .X(\shifter_0/n9762 ) );
  nand_x1_sg U43046 ( .A(n19240), .B(n19239), .X(\shifter_0/n9761 ) );
  nand_x1_sg U43047 ( .A(n19242), .B(n19241), .X(\shifter_0/n9760 ) );
  nand_x1_sg U43048 ( .A(n19244), .B(n19243), .X(\shifter_0/n9759 ) );
  nand_x1_sg U43049 ( .A(n19246), .B(n19245), .X(\shifter_0/n9758 ) );
  nand_x1_sg U43050 ( .A(n19248), .B(n19247), .X(\shifter_0/n9757 ) );
  nand_x1_sg U43051 ( .A(n19250), .B(n19249), .X(\shifter_0/n9756 ) );
  nand_x1_sg U43052 ( .A(n19252), .B(n19251), .X(\shifter_0/n9755 ) );
  nand_x1_sg U43053 ( .A(n19254), .B(n19253), .X(\shifter_0/n9754 ) );
  nand_x1_sg U43054 ( .A(n19256), .B(n19255), .X(\shifter_0/n9753 ) );
  nand_x1_sg U43055 ( .A(n19258), .B(n19257), .X(\shifter_0/n9752 ) );
  nand_x1_sg U43056 ( .A(n19260), .B(n19259), .X(\shifter_0/n9751 ) );
  nand_x1_sg U43057 ( .A(n19262), .B(n19261), .X(\shifter_0/n9750 ) );
  nand_x1_sg U43058 ( .A(n19264), .B(n19263), .X(\shifter_0/n9749 ) );
  nand_x1_sg U43059 ( .A(n19266), .B(n19265), .X(\shifter_0/n9748 ) );
  nand_x1_sg U43060 ( .A(n19268), .B(n19267), .X(\shifter_0/n9747 ) );
  nand_x1_sg U43061 ( .A(n19270), .B(n19269), .X(\shifter_0/n9746 ) );
  nand_x1_sg U43062 ( .A(n19272), .B(n19271), .X(\shifter_0/n9745 ) );
  nand_x1_sg U43063 ( .A(n19274), .B(n19273), .X(\shifter_0/n9744 ) );
  nand_x1_sg U43064 ( .A(n19492), .B(n19491), .X(\shifter_0/n9635 ) );
  nand_x1_sg U43065 ( .A(n19494), .B(n19493), .X(\shifter_0/n9634 ) );
  nand_x1_sg U43066 ( .A(n19496), .B(n19495), .X(\shifter_0/n9633 ) );
  nand_x1_sg U43067 ( .A(n19498), .B(n19497), .X(\shifter_0/n9632 ) );
  nand_x1_sg U43068 ( .A(n19500), .B(n19499), .X(\shifter_0/n9631 ) );
  nand_x1_sg U43069 ( .A(n19502), .B(n19501), .X(\shifter_0/n9630 ) );
  nand_x1_sg U43070 ( .A(n19504), .B(n19503), .X(\shifter_0/n9629 ) );
  nand_x1_sg U43071 ( .A(n19506), .B(n19505), .X(\shifter_0/n9628 ) );
  nand_x1_sg U43072 ( .A(n19508), .B(n19507), .X(\shifter_0/n9627 ) );
  nand_x1_sg U43073 ( .A(n19510), .B(n19509), .X(\shifter_0/n9626 ) );
  nand_x1_sg U43074 ( .A(n19512), .B(n19511), .X(\shifter_0/n9625 ) );
  nand_x1_sg U43075 ( .A(n19514), .B(n19513), .X(\shifter_0/n9624 ) );
  nand_x1_sg U43076 ( .A(n19516), .B(n19515), .X(\shifter_0/n9623 ) );
  nand_x1_sg U43077 ( .A(n19518), .B(n19517), .X(\shifter_0/n9622 ) );
  nand_x1_sg U43078 ( .A(n19520), .B(n19519), .X(\shifter_0/n9621 ) );
  nand_x1_sg U43079 ( .A(n19522), .B(n19521), .X(\shifter_0/n9620 ) );
  nand_x1_sg U43080 ( .A(n19564), .B(n19563), .X(\shifter_0/n9599 ) );
  nand_x1_sg U43081 ( .A(n19566), .B(n19565), .X(\shifter_0/n9598 ) );
  nand_x1_sg U43082 ( .A(n19568), .B(n19567), .X(\shifter_0/n9597 ) );
  nand_x1_sg U43083 ( .A(n19570), .B(n19569), .X(\shifter_0/n9596 ) );
  nand_x1_sg U43084 ( .A(n19572), .B(n19571), .X(\shifter_0/n9595 ) );
  nand_x1_sg U43085 ( .A(n19574), .B(n19573), .X(\shifter_0/n9594 ) );
  nand_x1_sg U43086 ( .A(n19576), .B(n19575), .X(\shifter_0/n9593 ) );
  nand_x1_sg U43087 ( .A(n19578), .B(n19577), .X(\shifter_0/n9592 ) );
  nand_x1_sg U43088 ( .A(n19532), .B(n19531), .X(\shifter_0/n9615 ) );
  nand_x1_sg U43089 ( .A(n19534), .B(n19533), .X(\shifter_0/n9614 ) );
  nand_x1_sg U43090 ( .A(n19536), .B(n19535), .X(\shifter_0/n9613 ) );
  nand_x1_sg U43091 ( .A(n22082), .B(n22081), .X(\shifter_0/n10063 ) );
  nand_x1_sg U43092 ( .A(n22084), .B(n22083), .X(\shifter_0/n10062 ) );
  nand_x1_sg U43093 ( .A(n22086), .B(n22085), .X(\shifter_0/n10061 ) );
  nand_x1_sg U43094 ( .A(n19020), .B(n19019), .X(\shifter_0/n9871 ) );
  nand_x1_sg U43095 ( .A(n19022), .B(n19021), .X(\shifter_0/n9870 ) );
  nand_x1_sg U43096 ( .A(n19024), .B(n19023), .X(\shifter_0/n9869 ) );
  nand_x1_sg U43097 ( .A(n19090), .B(n19089), .X(\shifter_0/n9836 ) );
  nand_x1_sg U43098 ( .A(n19092), .B(n19091), .X(\shifter_0/n9835 ) );
  nand_x1_sg U43099 ( .A(n19094), .B(n19093), .X(\shifter_0/n9834 ) );
  nand_x1_sg U43100 ( .A(n21890), .B(n21889), .X(\shifter_0/n10159 ) );
  nand_x1_sg U43101 ( .A(n21892), .B(n21891), .X(\shifter_0/n10158 ) );
  nand_x1_sg U43102 ( .A(n21894), .B(n21893), .X(\shifter_0/n10157 ) );
  nand_x1_sg U43103 ( .A(n21896), .B(n21895), .X(\shifter_0/n10156 ) );
  nand_x1_sg U43104 ( .A(n21898), .B(n21897), .X(\shifter_0/n10155 ) );
  nand_x1_sg U43105 ( .A(n21900), .B(n21899), .X(\shifter_0/n10154 ) );
  nand_x1_sg U43106 ( .A(n21902), .B(n21901), .X(\shifter_0/n10153 ) );
  nand_x1_sg U43107 ( .A(n21904), .B(n21903), .X(\shifter_0/n10152 ) );
  nand_x1_sg U43108 ( .A(n21906), .B(n21905), .X(\shifter_0/n10151 ) );
  nand_x1_sg U43109 ( .A(n21908), .B(n21907), .X(\shifter_0/n10150 ) );
  nand_x1_sg U43110 ( .A(n21910), .B(n21909), .X(\shifter_0/n10149 ) );
  nand_x1_sg U43111 ( .A(n21912), .B(n21911), .X(\shifter_0/n10148 ) );
  nand_x1_sg U43112 ( .A(n21914), .B(n21913), .X(\shifter_0/n10147 ) );
  nand_x1_sg U43113 ( .A(n21916), .B(n21915), .X(\shifter_0/n10146 ) );
  nand_x1_sg U43114 ( .A(n21918), .B(n21917), .X(\shifter_0/n10145 ) );
  nand_x1_sg U43115 ( .A(n21920), .B(n21919), .X(\shifter_0/n10144 ) );
  nand_x1_sg U43116 ( .A(n21922), .B(n21921), .X(\shifter_0/n10143 ) );
  nand_x1_sg U43117 ( .A(n21924), .B(n21923), .X(\shifter_0/n10142 ) );
  nand_x1_sg U43118 ( .A(n21926), .B(n21925), .X(\shifter_0/n10141 ) );
  nand_x1_sg U43119 ( .A(n21928), .B(n21927), .X(\shifter_0/n10140 ) );
  nand_x1_sg U43120 ( .A(n22050), .B(n22049), .X(\shifter_0/n10079 ) );
  nand_x1_sg U43121 ( .A(n22052), .B(n22051), .X(\shifter_0/n10078 ) );
  nand_x1_sg U43122 ( .A(n22054), .B(n22053), .X(\shifter_0/n10077 ) );
  nand_x1_sg U43123 ( .A(n22056), .B(n22055), .X(\shifter_0/n10076 ) );
  nand_x1_sg U43124 ( .A(n22058), .B(n22057), .X(\shifter_0/n10075 ) );
  nand_x1_sg U43125 ( .A(n22060), .B(n22059), .X(\shifter_0/n10074 ) );
  nand_x1_sg U43126 ( .A(n22062), .B(n22061), .X(\shifter_0/n10073 ) );
  nand_x1_sg U43127 ( .A(n22064), .B(n22063), .X(\shifter_0/n10072 ) );
  nand_x1_sg U43128 ( .A(n22066), .B(n22065), .X(\shifter_0/n10071 ) );
  nand_x1_sg U43129 ( .A(n22068), .B(n22067), .X(\shifter_0/n10070 ) );
  nand_x1_sg U43130 ( .A(n22070), .B(n22069), .X(\shifter_0/n10069 ) );
  nand_x1_sg U43131 ( .A(n22072), .B(n22071), .X(\shifter_0/n10068 ) );
  nand_x1_sg U43132 ( .A(n22074), .B(n22073), .X(\shifter_0/n10067 ) );
  nand_x1_sg U43133 ( .A(n22076), .B(n22075), .X(\shifter_0/n10066 ) );
  nand_x1_sg U43134 ( .A(n22078), .B(n22077), .X(\shifter_0/n10065 ) );
  nand_x1_sg U43135 ( .A(n22080), .B(n22079), .X(\shifter_0/n10064 ) );
  nand_x1_sg U43136 ( .A(n22088), .B(n22087), .X(\shifter_0/n10060 ) );
  nand_x1_sg U43137 ( .A(n18804), .B(n18803), .X(\shifter_0/n9979 ) );
  nand_x1_sg U43138 ( .A(n18806), .B(n18805), .X(\shifter_0/n9978 ) );
  nand_x1_sg U43139 ( .A(n18808), .B(n18807), .X(\shifter_0/n9977 ) );
  nand_x1_sg U43140 ( .A(n18810), .B(n18809), .X(\shifter_0/n9976 ) );
  nand_x1_sg U43141 ( .A(n18812), .B(n18811), .X(\shifter_0/n9975 ) );
  nand_x1_sg U43142 ( .A(n18814), .B(n18813), .X(\shifter_0/n9974 ) );
  nand_x1_sg U43143 ( .A(n18816), .B(n18815), .X(\shifter_0/n9973 ) );
  nand_x1_sg U43144 ( .A(n18818), .B(n18817), .X(\shifter_0/n9972 ) );
  nand_x1_sg U43145 ( .A(n18820), .B(n18819), .X(\shifter_0/n9971 ) );
  nand_x1_sg U43146 ( .A(n18822), .B(n18821), .X(\shifter_0/n9970 ) );
  nand_x1_sg U43147 ( .A(n18824), .B(n18823), .X(\shifter_0/n9969 ) );
  nand_x1_sg U43148 ( .A(n18826), .B(n18825), .X(\shifter_0/n9968 ) );
  nand_x1_sg U43149 ( .A(n18828), .B(n18827), .X(\shifter_0/n9967 ) );
  nand_x1_sg U43150 ( .A(n18830), .B(n18829), .X(\shifter_0/n9966 ) );
  nand_x1_sg U43151 ( .A(n18832), .B(n18831), .X(\shifter_0/n9965 ) );
  nand_x1_sg U43152 ( .A(n18834), .B(n18833), .X(\shifter_0/n9964 ) );
  nand_x1_sg U43153 ( .A(n18836), .B(n18835), .X(\shifter_0/n9963 ) );
  nand_x1_sg U43154 ( .A(n18838), .B(n18837), .X(\shifter_0/n9962 ) );
  nand_x1_sg U43155 ( .A(n18840), .B(n18839), .X(\shifter_0/n9961 ) );
  nand_x1_sg U43156 ( .A(n18842), .B(n18841), .X(\shifter_0/n9960 ) );
  nand_x1_sg U43157 ( .A(n19026), .B(n19025), .X(\shifter_0/n9868 ) );
  nand_x1_sg U43158 ( .A(n19028), .B(n19027), .X(\shifter_0/n9867 ) );
  nand_x1_sg U43159 ( .A(n19030), .B(n19029), .X(\shifter_0/n9866 ) );
  nand_x1_sg U43160 ( .A(n19032), .B(n19031), .X(\shifter_0/n9865 ) );
  nand_x1_sg U43161 ( .A(n19034), .B(n19033), .X(\shifter_0/n9864 ) );
  nand_x1_sg U43162 ( .A(n19036), .B(n19035), .X(\shifter_0/n9863 ) );
  nand_x1_sg U43163 ( .A(n19038), .B(n19037), .X(\shifter_0/n9862 ) );
  nand_x1_sg U43164 ( .A(n19040), .B(n19039), .X(\shifter_0/n9861 ) );
  nand_x1_sg U43165 ( .A(n19042), .B(n19041), .X(\shifter_0/n9860 ) );
  nand_x1_sg U43166 ( .A(n19096), .B(n19095), .X(\shifter_0/n9833 ) );
  nand_x1_sg U43167 ( .A(n19098), .B(n19097), .X(\shifter_0/n9832 ) );
  nand_x1_sg U43168 ( .A(n19100), .B(n19099), .X(\shifter_0/n9831 ) );
  nand_x1_sg U43169 ( .A(n19102), .B(n19101), .X(\shifter_0/n9830 ) );
  nand_x1_sg U43170 ( .A(n19104), .B(n19103), .X(\shifter_0/n9829 ) );
  nand_x1_sg U43171 ( .A(n19106), .B(n19105), .X(\shifter_0/n9828 ) );
  nand_x1_sg U43172 ( .A(n19108), .B(n19107), .X(\shifter_0/n9827 ) );
  nand_x1_sg U43173 ( .A(n19110), .B(n19109), .X(\shifter_0/n9826 ) );
  nand_x1_sg U43174 ( .A(n19112), .B(n19111), .X(\shifter_0/n9825 ) );
  nand_x1_sg U43175 ( .A(n19114), .B(n19113), .X(\shifter_0/n9824 ) );
  nand_x1_sg U43176 ( .A(n19116), .B(n19115), .X(\shifter_0/n9823 ) );
  nand_x1_sg U43177 ( .A(n19118), .B(n19117), .X(\shifter_0/n9822 ) );
  nand_x1_sg U43178 ( .A(n19120), .B(n19119), .X(\shifter_0/n9821 ) );
  nand_x1_sg U43179 ( .A(n19122), .B(n19121), .X(\shifter_0/n9820 ) );
  nand_x1_sg U43180 ( .A(n19164), .B(n19163), .X(\shifter_0/n9799 ) );
  nand_x1_sg U43181 ( .A(n19166), .B(n19165), .X(\shifter_0/n9798 ) );
  nand_x1_sg U43182 ( .A(n19168), .B(n19167), .X(\shifter_0/n9797 ) );
  nand_x1_sg U43183 ( .A(n19170), .B(n19169), .X(\shifter_0/n9796 ) );
  nand_x1_sg U43184 ( .A(n19172), .B(n19171), .X(\shifter_0/n9795 ) );
  nand_x1_sg U43185 ( .A(n19174), .B(n19173), .X(\shifter_0/n9794 ) );
  nand_x1_sg U43186 ( .A(n19176), .B(n19175), .X(\shifter_0/n9793 ) );
  nand_x1_sg U43187 ( .A(n19178), .B(n19177), .X(\shifter_0/n9792 ) );
  nand_x1_sg U43188 ( .A(n19180), .B(n19179), .X(\shifter_0/n9791 ) );
  nand_x1_sg U43189 ( .A(n19182), .B(n19181), .X(\shifter_0/n9790 ) );
  nand_x1_sg U43190 ( .A(n19184), .B(n19183), .X(\shifter_0/n9789 ) );
  nand_x1_sg U43191 ( .A(n19186), .B(n19185), .X(\shifter_0/n9788 ) );
  nand_x1_sg U43192 ( .A(n19188), .B(n19187), .X(\shifter_0/n9787 ) );
  nand_x1_sg U43193 ( .A(n19190), .B(n19189), .X(\shifter_0/n9786 ) );
  nand_x1_sg U43194 ( .A(n19192), .B(n19191), .X(\shifter_0/n9785 ) );
  nand_x1_sg U43195 ( .A(n19194), .B(n19193), .X(\shifter_0/n9784 ) );
  nand_x1_sg U43196 ( .A(n19196), .B(n19195), .X(\shifter_0/n9783 ) );
  nand_x1_sg U43197 ( .A(n19198), .B(n19197), .X(\shifter_0/n9782 ) );
  nand_x1_sg U43198 ( .A(n19200), .B(n19199), .X(\shifter_0/n9781 ) );
  nand_x1_sg U43199 ( .A(n19202), .B(n19201), .X(\shifter_0/n9780 ) );
  nand_x1_sg U43200 ( .A(n19364), .B(n19363), .X(\shifter_0/n9699 ) );
  nand_x1_sg U43201 ( .A(n19366), .B(n19365), .X(\shifter_0/n9698 ) );
  nand_x1_sg U43202 ( .A(n19368), .B(n19367), .X(\shifter_0/n9697 ) );
  nand_x1_sg U43203 ( .A(n19370), .B(n19369), .X(\shifter_0/n9696 ) );
  nand_x1_sg U43204 ( .A(n19372), .B(n19371), .X(\shifter_0/n9695 ) );
  nand_x1_sg U43205 ( .A(n19374), .B(n19373), .X(\shifter_0/n9694 ) );
  nand_x1_sg U43206 ( .A(n19376), .B(n19375), .X(\shifter_0/n9693 ) );
  nand_x1_sg U43207 ( .A(n19378), .B(n19377), .X(\shifter_0/n9692 ) );
  nand_x1_sg U43208 ( .A(n19380), .B(n19379), .X(\shifter_0/n9691 ) );
  nand_x1_sg U43209 ( .A(n19382), .B(n19381), .X(\shifter_0/n9690 ) );
  nand_x1_sg U43210 ( .A(n19384), .B(n19383), .X(\shifter_0/n9689 ) );
  nand_x1_sg U43211 ( .A(n19386), .B(n19385), .X(\shifter_0/n9688 ) );
  nand_x1_sg U43212 ( .A(n19388), .B(n19387), .X(\shifter_0/n9687 ) );
  nand_x1_sg U43213 ( .A(n19390), .B(n19389), .X(\shifter_0/n9686 ) );
  nand_x1_sg U43214 ( .A(n19392), .B(n19391), .X(\shifter_0/n9685 ) );
  nand_x1_sg U43215 ( .A(n19394), .B(n19393), .X(\shifter_0/n9684 ) );
  nand_x1_sg U43216 ( .A(n19396), .B(n19395), .X(\shifter_0/n9683 ) );
  nand_x1_sg U43217 ( .A(n19398), .B(n19397), .X(\shifter_0/n9682 ) );
  nand_x1_sg U43218 ( .A(n19400), .B(n19399), .X(\shifter_0/n9681 ) );
  nand_x1_sg U43219 ( .A(n19402), .B(n19401), .X(\shifter_0/n9680 ) );
  nand_x1_sg U43220 ( .A(n19444), .B(n19443), .X(\shifter_0/n9659 ) );
  nand_x1_sg U43221 ( .A(n19446), .B(n19445), .X(\shifter_0/n9658 ) );
  nand_x1_sg U43222 ( .A(n19448), .B(n19447), .X(\shifter_0/n9657 ) );
  nand_x1_sg U43223 ( .A(n19450), .B(n19449), .X(\shifter_0/n9656 ) );
  nand_x1_sg U43224 ( .A(n19452), .B(n19451), .X(\shifter_0/n9655 ) );
  nand_x1_sg U43225 ( .A(n19454), .B(n19453), .X(\shifter_0/n9654 ) );
  nand_x1_sg U43226 ( .A(n19456), .B(n19455), .X(\shifter_0/n9653 ) );
  nand_x1_sg U43227 ( .A(n19458), .B(n19457), .X(\shifter_0/n9652 ) );
  nand_x1_sg U43228 ( .A(n19460), .B(n19459), .X(\shifter_0/n9651 ) );
  nand_x1_sg U43229 ( .A(n19462), .B(n19461), .X(\shifter_0/n9650 ) );
  nand_x1_sg U43230 ( .A(n19464), .B(n19463), .X(\shifter_0/n9649 ) );
  nand_x1_sg U43231 ( .A(n19466), .B(n19465), .X(\shifter_0/n9648 ) );
  nand_x1_sg U43232 ( .A(n19468), .B(n19467), .X(\shifter_0/n9647 ) );
  nand_x1_sg U43233 ( .A(n19470), .B(n19469), .X(\shifter_0/n9646 ) );
  nand_x1_sg U43234 ( .A(n19472), .B(n19471), .X(\shifter_0/n9645 ) );
  nand_x1_sg U43235 ( .A(n19474), .B(n19473), .X(\shifter_0/n9644 ) );
  nand_x1_sg U43236 ( .A(n19476), .B(n19475), .X(\shifter_0/n9643 ) );
  nand_x1_sg U43237 ( .A(n19478), .B(n19477), .X(\shifter_0/n9642 ) );
  nand_x1_sg U43238 ( .A(n19480), .B(n19479), .X(\shifter_0/n9641 ) );
  nand_x1_sg U43239 ( .A(n19482), .B(n19481), .X(\shifter_0/n9640 ) );
  nand_x1_sg U43240 ( .A(n19526), .B(n19525), .X(\shifter_0/n9618 ) );
  nand_x1_sg U43241 ( .A(n19528), .B(n19527), .X(\shifter_0/n9617 ) );
  nand_x1_sg U43242 ( .A(n19530), .B(n19529), .X(\shifter_0/n9616 ) );
  nand_x1_sg U43243 ( .A(n21970), .B(n21969), .X(\shifter_0/n10119 ) );
  nand_x1_sg U43244 ( .A(n21972), .B(n21971), .X(\shifter_0/n10118 ) );
  nand_x1_sg U43245 ( .A(n21974), .B(n21973), .X(\shifter_0/n10117 ) );
  nand_x1_sg U43246 ( .A(n21976), .B(n21975), .X(\shifter_0/n10116 ) );
  nand_x1_sg U43247 ( .A(n21978), .B(n21977), .X(\shifter_0/n10115 ) );
  nand_x1_sg U43248 ( .A(n21980), .B(n21979), .X(\shifter_0/n10114 ) );
  nand_x1_sg U43249 ( .A(n21982), .B(n21981), .X(\shifter_0/n10113 ) );
  nand_x1_sg U43250 ( .A(n21984), .B(n21983), .X(\shifter_0/n10112 ) );
  nand_x1_sg U43251 ( .A(n21986), .B(n21985), .X(\shifter_0/n10111 ) );
  nand_x1_sg U43252 ( .A(n21988), .B(n21987), .X(\shifter_0/n10110 ) );
  nand_x1_sg U43253 ( .A(n21990), .B(n21989), .X(\shifter_0/n10109 ) );
  nand_x1_sg U43254 ( .A(n21992), .B(n21991), .X(\shifter_0/n10108 ) );
  nand_x1_sg U43255 ( .A(n21994), .B(n21993), .X(\shifter_0/n10107 ) );
  nand_x1_sg U43256 ( .A(n21996), .B(n21995), .X(\shifter_0/n10106 ) );
  nand_x1_sg U43257 ( .A(n21998), .B(n21997), .X(\shifter_0/n10105 ) );
  nand_x1_sg U43258 ( .A(n22000), .B(n21999), .X(\shifter_0/n10104 ) );
  nand_x1_sg U43259 ( .A(n22002), .B(n22001), .X(\shifter_0/n10103 ) );
  nand_x1_sg U43260 ( .A(n22004), .B(n22003), .X(\shifter_0/n10102 ) );
  nand_x1_sg U43261 ( .A(n22006), .B(n22005), .X(\shifter_0/n10101 ) );
  nand_x1_sg U43262 ( .A(n22008), .B(n22007), .X(\shifter_0/n10100 ) );
  nand_x1_sg U43263 ( .A(n19004), .B(n19003), .X(\shifter_0/n9879 ) );
  nand_x1_sg U43264 ( .A(n19006), .B(n19005), .X(\shifter_0/n9878 ) );
  nand_x1_sg U43265 ( .A(n19008), .B(n19007), .X(\shifter_0/n9877 ) );
  nand_x1_sg U43266 ( .A(n19010), .B(n19009), .X(\shifter_0/n9876 ) );
  nand_x1_sg U43267 ( .A(n19012), .B(n19011), .X(\shifter_0/n9875 ) );
  nand_x1_sg U43268 ( .A(n19014), .B(n19013), .X(\shifter_0/n9874 ) );
  nand_x1_sg U43269 ( .A(n19016), .B(n19015), .X(\shifter_0/n9873 ) );
  nand_x1_sg U43270 ( .A(n19018), .B(n19017), .X(\shifter_0/n9872 ) );
  nand_x1_sg U43271 ( .A(n19084), .B(n19083), .X(\shifter_0/n9839 ) );
  nand_x1_sg U43272 ( .A(n19086), .B(n19085), .X(\shifter_0/n9838 ) );
  nand_x1_sg U43273 ( .A(n19088), .B(n19087), .X(\shifter_0/n9837 ) );
  nand_x1_sg U43274 ( .A(n19524), .B(n19523), .X(\shifter_0/n9619 ) );
  nand_x1_sg U43275 ( .A(n19538), .B(n19537), .X(\shifter_0/n9612 ) );
  nand_x1_sg U43276 ( .A(n19540), .B(n19539), .X(\shifter_0/n9611 ) );
  nand_x1_sg U43277 ( .A(n19542), .B(n19541), .X(\shifter_0/n9610 ) );
  nand_x1_sg U43278 ( .A(n19544), .B(n19543), .X(\shifter_0/n9609 ) );
  nand_x1_sg U43279 ( .A(n19546), .B(n19545), .X(\shifter_0/n9608 ) );
  nand_x1_sg U43280 ( .A(n19548), .B(n19547), .X(\shifter_0/n9607 ) );
  nand_x1_sg U43281 ( .A(n19550), .B(n19549), .X(\shifter_0/n9606 ) );
  nand_x1_sg U43282 ( .A(n19552), .B(n19551), .X(\shifter_0/n9605 ) );
  nand_x1_sg U43283 ( .A(n19554), .B(n19553), .X(\shifter_0/n9604 ) );
  nand_x1_sg U43284 ( .A(n19556), .B(n19555), .X(\shifter_0/n9603 ) );
  nand_x1_sg U43285 ( .A(n19558), .B(n19557), .X(\shifter_0/n9602 ) );
  nand_x1_sg U43286 ( .A(n19560), .B(n19559), .X(\shifter_0/n9601 ) );
  nand_x1_sg U43287 ( .A(n19562), .B(n19561), .X(\shifter_0/n9600 ) );
  nand_x1_sg U43288 ( .A(n21345), .B(n21346), .X(\shifter_0/n10233 ) );
  nand_x1_sg U43289 ( .A(n21368), .B(n21369), .X(\shifter_0/n10232 ) );
  nand_x1_sg U43290 ( .A(n21372), .B(n21373), .X(n21371) );
  nand_x1_sg U43291 ( .A(n20902), .B(n20903), .X(\shifter_0/n10239 ) );
  nand_x1_sg U43292 ( .A(n20933), .B(n20934), .X(\shifter_0/n10238 ) );
  nand_x1_sg U43293 ( .A(n29076), .B(n29077), .X(\filter_0/n8517 ) );
  nand_x1_sg U43294 ( .A(n29078), .B(n29079), .X(\filter_0/n8516 ) );
  nand_x1_sg U43295 ( .A(n29080), .B(n29081), .X(\filter_0/n8515 ) );
  nand_x1_sg U43296 ( .A(n29082), .B(n29083), .X(\filter_0/n8514 ) );
  nand_x1_sg U43297 ( .A(n29084), .B(n29085), .X(\filter_0/n8513 ) );
  nand_x1_sg U43298 ( .A(n29086), .B(n29087), .X(\filter_0/n8512 ) );
  nand_x1_sg U43299 ( .A(n29088), .B(n29089), .X(\filter_0/n8511 ) );
  nand_x1_sg U43300 ( .A(n29090), .B(n29091), .X(\filter_0/n8510 ) );
  nand_x1_sg U43301 ( .A(n29092), .B(n29093), .X(\filter_0/n8509 ) );
  nand_x1_sg U43302 ( .A(n29094), .B(n29095), .X(\filter_0/n8508 ) );
  nand_x1_sg U43303 ( .A(n29096), .B(n29097), .X(\filter_0/n8507 ) );
  nand_x1_sg U43304 ( .A(n29098), .B(n29099), .X(\filter_0/n8506 ) );
  nand_x1_sg U43305 ( .A(n29100), .B(n29101), .X(\filter_0/n8505 ) );
  nand_x1_sg U43306 ( .A(n29102), .B(n29103), .X(\filter_0/n8504 ) );
  nand_x1_sg U43307 ( .A(n29289), .B(n29290), .X(\filter_0/n8417 ) );
  nand_x1_sg U43308 ( .A(n29291), .B(n29292), .X(\filter_0/n8416 ) );
  nand_x1_sg U43309 ( .A(n29293), .B(n29294), .X(\filter_0/n8415 ) );
  nand_x1_sg U43310 ( .A(n29295), .B(n29296), .X(\filter_0/n8414 ) );
  nand_x1_sg U43311 ( .A(n29297), .B(n29298), .X(\filter_0/n8413 ) );
  nand_x1_sg U43312 ( .A(n29299), .B(n29300), .X(\filter_0/n8412 ) );
  nand_x1_sg U43313 ( .A(n29301), .B(n29302), .X(\filter_0/n8411 ) );
  nand_x1_sg U43314 ( .A(n29303), .B(n29304), .X(\filter_0/n8410 ) );
  nand_x1_sg U43315 ( .A(n29305), .B(n29306), .X(\filter_0/n8409 ) );
  nand_x1_sg U43316 ( .A(n29307), .B(n29308), .X(\filter_0/n8408 ) );
  nand_x1_sg U43317 ( .A(n29309), .B(n29310), .X(\filter_0/n8407 ) );
  nand_x1_sg U43318 ( .A(n29311), .B(n29312), .X(\filter_0/n8406 ) );
  nand_x1_sg U43319 ( .A(n29313), .B(n29314), .X(\filter_0/n8405 ) );
  nand_x1_sg U43320 ( .A(n29315), .B(n29316), .X(\filter_0/n8404 ) );
  nand_x1_sg U43321 ( .A(n29072), .B(n29073), .X(\filter_0/n8519 ) );
  nand_x1_sg U43322 ( .A(n29985), .B(\filter_0/n8235 ), .X(n29073) );
  nand_x1_sg U43323 ( .A(n29074), .B(n29075), .X(\filter_0/n8518 ) );
  nand_x1_sg U43324 ( .A(n33466), .B(\filter_0/n8234 ), .X(n29075) );
  nand_x1_sg U43325 ( .A(n29285), .B(n29286), .X(\filter_0/n8419 ) );
  nand_x1_sg U43326 ( .A(n33405), .B(\filter_0/n8015 ), .X(n29286) );
  nand_x1_sg U43327 ( .A(n29287), .B(n29288), .X(\filter_0/n8418 ) );
  nand_x1_sg U43328 ( .A(n33406), .B(\filter_0/n8014 ), .X(n29288) );
  nand_x1_sg U43329 ( .A(n29033), .B(n29034), .X(\filter_0/n8537 ) );
  nand_x1_sg U43330 ( .A(n29035), .B(n29036), .X(\filter_0/n8536 ) );
  nand_x1_sg U43331 ( .A(n29037), .B(n29038), .X(\filter_0/n8535 ) );
  nand_x1_sg U43332 ( .A(n29039), .B(n29040), .X(\filter_0/n8534 ) );
  nand_x1_sg U43333 ( .A(n29041), .B(n29042), .X(\filter_0/n8533 ) );
  nand_x1_sg U43334 ( .A(n29043), .B(n29044), .X(\filter_0/n8532 ) );
  nand_x1_sg U43335 ( .A(n29045), .B(n29046), .X(\filter_0/n8531 ) );
  nand_x1_sg U43336 ( .A(n29047), .B(n29048), .X(\filter_0/n8530 ) );
  nand_x1_sg U43337 ( .A(n29049), .B(n29050), .X(\filter_0/n8529 ) );
  nand_x1_sg U43338 ( .A(n29051), .B(n29052), .X(\filter_0/n8528 ) );
  nand_x1_sg U43339 ( .A(n29053), .B(n29054), .X(\filter_0/n8527 ) );
  nand_x1_sg U43340 ( .A(n29055), .B(n29056), .X(\filter_0/n8526 ) );
  nand_x1_sg U43341 ( .A(n29057), .B(n29058), .X(\filter_0/n8525 ) );
  nand_x1_sg U43342 ( .A(n29059), .B(n29060), .X(\filter_0/n8524 ) );
  nand_x1_sg U43343 ( .A(n28990), .B(n28991), .X(\filter_0/n8557 ) );
  nand_x1_sg U43344 ( .A(n28992), .B(n28993), .X(\filter_0/n8556 ) );
  nand_x1_sg U43345 ( .A(n28994), .B(n28995), .X(\filter_0/n8555 ) );
  nand_x1_sg U43346 ( .A(n28996), .B(n28997), .X(\filter_0/n8554 ) );
  nand_x1_sg U43347 ( .A(n28998), .B(n28999), .X(\filter_0/n8553 ) );
  nand_x1_sg U43348 ( .A(n29000), .B(n29001), .X(\filter_0/n8552 ) );
  nand_x1_sg U43349 ( .A(n29002), .B(n29003), .X(\filter_0/n8551 ) );
  nand_x1_sg U43350 ( .A(n29004), .B(n29005), .X(\filter_0/n8550 ) );
  nand_x1_sg U43351 ( .A(n29006), .B(n29007), .X(\filter_0/n8549 ) );
  nand_x1_sg U43352 ( .A(n29008), .B(n29009), .X(\filter_0/n8548 ) );
  nand_x1_sg U43353 ( .A(n29010), .B(n29011), .X(\filter_0/n8547 ) );
  nand_x1_sg U43354 ( .A(n29012), .B(n29013), .X(\filter_0/n8546 ) );
  nand_x1_sg U43355 ( .A(n29014), .B(n29015), .X(\filter_0/n8545 ) );
  nand_x1_sg U43356 ( .A(n29016), .B(n29017), .X(\filter_0/n8544 ) );
  nand_x1_sg U43357 ( .A(n29205), .B(n29206), .X(\filter_0/n8457 ) );
  nand_x1_sg U43358 ( .A(n29207), .B(n29208), .X(\filter_0/n8456 ) );
  nand_x1_sg U43359 ( .A(n29209), .B(n29210), .X(\filter_0/n8455 ) );
  nand_x1_sg U43360 ( .A(n29211), .B(n29212), .X(\filter_0/n8454 ) );
  nand_x1_sg U43361 ( .A(n29213), .B(n29214), .X(\filter_0/n8453 ) );
  nand_x1_sg U43362 ( .A(n29215), .B(n29216), .X(\filter_0/n8452 ) );
  nand_x1_sg U43363 ( .A(n29217), .B(n29218), .X(\filter_0/n8451 ) );
  nand_x1_sg U43364 ( .A(n29219), .B(n29220), .X(\filter_0/n8450 ) );
  nand_x1_sg U43365 ( .A(n29221), .B(n29222), .X(\filter_0/n8449 ) );
  nand_x1_sg U43366 ( .A(n29223), .B(n29224), .X(\filter_0/n8448 ) );
  nand_x1_sg U43367 ( .A(n29225), .B(n29226), .X(\filter_0/n8447 ) );
  nand_x1_sg U43368 ( .A(n29227), .B(n29228), .X(\filter_0/n8446 ) );
  nand_x1_sg U43369 ( .A(n29229), .B(n29230), .X(\filter_0/n8445 ) );
  nand_x1_sg U43370 ( .A(n29231), .B(n29232), .X(\filter_0/n8444 ) );
  nand_x1_sg U43371 ( .A(n29163), .B(n29164), .X(\filter_0/n8477 ) );
  nand_x1_sg U43372 ( .A(n29165), .B(n29166), .X(\filter_0/n8476 ) );
  nand_x1_sg U43373 ( .A(n29167), .B(n29168), .X(\filter_0/n8475 ) );
  nand_x1_sg U43374 ( .A(n29169), .B(n29170), .X(\filter_0/n8474 ) );
  nand_x1_sg U43375 ( .A(n29171), .B(n29172), .X(\filter_0/n8473 ) );
  nand_x1_sg U43376 ( .A(n29173), .B(n29174), .X(\filter_0/n8472 ) );
  nand_x1_sg U43377 ( .A(n29175), .B(n29176), .X(\filter_0/n8471 ) );
  nand_x1_sg U43378 ( .A(n29177), .B(n29178), .X(\filter_0/n8470 ) );
  nand_x1_sg U43379 ( .A(n29179), .B(n29180), .X(\filter_0/n8469 ) );
  nand_x1_sg U43380 ( .A(n29181), .B(n29182), .X(\filter_0/n8468 ) );
  nand_x1_sg U43381 ( .A(n29183), .B(n29184), .X(\filter_0/n8467 ) );
  nand_x1_sg U43382 ( .A(n29185), .B(n29186), .X(\filter_0/n8466 ) );
  nand_x1_sg U43383 ( .A(n29187), .B(n29188), .X(\filter_0/n8465 ) );
  nand_x1_sg U43384 ( .A(n29189), .B(n29190), .X(\filter_0/n8464 ) );
  nand_x1_sg U43385 ( .A(n29332), .B(n29333), .X(\filter_0/n8397 ) );
  nand_x1_sg U43386 ( .A(n29334), .B(n29335), .X(\filter_0/n8396 ) );
  nand_x1_sg U43387 ( .A(n29336), .B(n29337), .X(\filter_0/n8395 ) );
  nand_x1_sg U43388 ( .A(n29338), .B(n29339), .X(\filter_0/n8394 ) );
  nand_x1_sg U43389 ( .A(n29340), .B(n29341), .X(\filter_0/n8393 ) );
  nand_x1_sg U43390 ( .A(n29342), .B(n29343), .X(\filter_0/n8392 ) );
  nand_x1_sg U43391 ( .A(n29344), .B(n29345), .X(\filter_0/n8391 ) );
  nand_x1_sg U43392 ( .A(n29346), .B(n29347), .X(\filter_0/n8390 ) );
  nand_x1_sg U43393 ( .A(n29348), .B(n29349), .X(\filter_0/n8389 ) );
  nand_x1_sg U43394 ( .A(n29350), .B(n29351), .X(\filter_0/n8388 ) );
  nand_x1_sg U43395 ( .A(n29352), .B(n29353), .X(\filter_0/n8387 ) );
  nand_x1_sg U43396 ( .A(n29354), .B(n29355), .X(\filter_0/n8386 ) );
  nand_x1_sg U43397 ( .A(n29356), .B(n29357), .X(\filter_0/n8385 ) );
  nand_x1_sg U43398 ( .A(n29358), .B(n29359), .X(\filter_0/n8384 ) );
  nand_x1_sg U43399 ( .A(n29374), .B(n29375), .X(\filter_0/n8377 ) );
  nand_x1_sg U43400 ( .A(n29376), .B(n29377), .X(\filter_0/n8376 ) );
  nand_x1_sg U43401 ( .A(n29378), .B(n29379), .X(\filter_0/n8375 ) );
  nand_x1_sg U43402 ( .A(n29380), .B(n29381), .X(\filter_0/n8374 ) );
  nand_x1_sg U43403 ( .A(n29382), .B(n29383), .X(\filter_0/n8373 ) );
  nand_x1_sg U43404 ( .A(n29384), .B(n29385), .X(\filter_0/n8372 ) );
  nand_x1_sg U43405 ( .A(n29386), .B(n29387), .X(\filter_0/n8371 ) );
  nand_x1_sg U43406 ( .A(n29388), .B(n29389), .X(\filter_0/n8370 ) );
  nand_x1_sg U43407 ( .A(n29390), .B(n29391), .X(\filter_0/n8369 ) );
  nand_x1_sg U43408 ( .A(n29392), .B(n29393), .X(\filter_0/n8368 ) );
  nand_x1_sg U43409 ( .A(n29394), .B(n29395), .X(\filter_0/n8367 ) );
  nand_x1_sg U43410 ( .A(n29396), .B(n29397), .X(\filter_0/n8366 ) );
  nand_x1_sg U43411 ( .A(n29398), .B(n29399), .X(\filter_0/n8365 ) );
  nand_x1_sg U43412 ( .A(n29400), .B(n29401), .X(\filter_0/n8364 ) );
  nand_x1_sg U43413 ( .A(n29062), .B(n29063), .X(\filter_0/n8523 ) );
  nand_x1_sg U43414 ( .A(n33467), .B(\filter_0/n8239 ), .X(n29063) );
  nand_x1_sg U43415 ( .A(n29066), .B(n29067), .X(\filter_0/n8522 ) );
  nand_x1_sg U43416 ( .A(n33468), .B(\filter_0/n8238 ), .X(n29067) );
  nand_x1_sg U43417 ( .A(n29068), .B(n29069), .X(\filter_0/n8521 ) );
  nand_x1_sg U43418 ( .A(n33467), .B(\filter_0/n8237 ), .X(n29069) );
  nand_x1_sg U43419 ( .A(n29070), .B(n29071), .X(\filter_0/n8520 ) );
  nand_x1_sg U43420 ( .A(n29985), .B(\filter_0/n8236 ), .X(n29071) );
  nand_x1_sg U43421 ( .A(n29275), .B(n29276), .X(\filter_0/n8423 ) );
  nand_x1_sg U43422 ( .A(n33408), .B(\filter_0/n8019 ), .X(n29276) );
  nand_x1_sg U43423 ( .A(n29279), .B(n29280), .X(\filter_0/n8422 ) );
  nand_x1_sg U43424 ( .A(n33406), .B(\filter_0/n8018 ), .X(n29280) );
  nand_x1_sg U43425 ( .A(n29281), .B(n29282), .X(\filter_0/n8421 ) );
  nand_x1_sg U43426 ( .A(n29961), .B(\filter_0/n8017 ), .X(n29282) );
  nand_x1_sg U43427 ( .A(n29283), .B(n29284), .X(\filter_0/n8420 ) );
  nand_x1_sg U43428 ( .A(n33408), .B(\filter_0/n8016 ), .X(n29284) );
  nand_x1_sg U43429 ( .A(n29255), .B(n29256), .X(\filter_0/n8433 ) );
  nand_x1_sg U43430 ( .A(n29267), .B(n29268), .X(\filter_0/n8427 ) );
  nand_x1_sg U43431 ( .A(n29251), .B(n29252), .X(\filter_0/n8435 ) );
  nand_x1_sg U43432 ( .A(n29263), .B(n29264), .X(\filter_0/n8429 ) );
  nand_x1_sg U43433 ( .A(n29247), .B(n29248), .X(\filter_0/n8437 ) );
  nand_x1_sg U43434 ( .A(n29259), .B(n29260), .X(\filter_0/n8431 ) );
  nand_x1_sg U43435 ( .A(n29271), .B(n29272), .X(\filter_0/n8425 ) );
  nand_x1_sg U43436 ( .A(n29467), .B(n29468), .X(\filter_0/n8333 ) );
  nand_x1_sg U43437 ( .A(n29479), .B(n29480), .X(\filter_0/n8327 ) );
  nand_x1_sg U43438 ( .A(n29463), .B(n29464), .X(\filter_0/n8335 ) );
  nand_x1_sg U43439 ( .A(n29475), .B(n29476), .X(\filter_0/n8329 ) );
  nand_x1_sg U43440 ( .A(n29459), .B(n29460), .X(\filter_0/n8337 ) );
  nand_x1_sg U43441 ( .A(n29471), .B(n29472), .X(\filter_0/n8331 ) );
  nand_x1_sg U43442 ( .A(n29483), .B(n29484), .X(\filter_0/n8325 ) );
  nand_x1_sg U43443 ( .A(n29029), .B(n29030), .X(\filter_0/n8539 ) );
  nand_x1_sg U43444 ( .A(n29925), .B(\filter_0/n8215 ), .X(n29030) );
  nand_x1_sg U43445 ( .A(n29031), .B(n29032), .X(\filter_0/n8538 ) );
  nand_x1_sg U43446 ( .A(n33316), .B(\filter_0/n8214 ), .X(n29032) );
  nand_x1_sg U43447 ( .A(n29201), .B(n29202), .X(\filter_0/n8459 ) );
  nand_x1_sg U43448 ( .A(n33435), .B(\filter_0/n8135 ), .X(n29202) );
  nand_x1_sg U43449 ( .A(n29203), .B(n29204), .X(\filter_0/n8458 ) );
  nand_x1_sg U43450 ( .A(n33437), .B(\filter_0/n8134 ), .X(n29204) );
  nand_x1_sg U43451 ( .A(n29328), .B(n29329), .X(\filter_0/n8399 ) );
  nand_x1_sg U43452 ( .A(n29923), .B(\filter_0/n8075 ), .X(n29329) );
  nand_x1_sg U43453 ( .A(n29330), .B(n29331), .X(\filter_0/n8398 ) );
  nand_x1_sg U43454 ( .A(n29923), .B(\filter_0/n8074 ), .X(n29331) );
  nand_x1_sg U43455 ( .A(n28986), .B(n28987), .X(\filter_0/n8559 ) );
  nand_x1_sg U43456 ( .A(n33306), .B(\filter_0/n8195 ), .X(n28987) );
  nand_x1_sg U43457 ( .A(n28988), .B(n28989), .X(\filter_0/n8558 ) );
  nand_x1_sg U43458 ( .A(n29921), .B(\filter_0/n8194 ), .X(n28989) );
  nand_x1_sg U43459 ( .A(n29159), .B(n29160), .X(\filter_0/n8479 ) );
  nand_x1_sg U43460 ( .A(n29983), .B(\filter_0/n8115 ), .X(n29160) );
  nand_x1_sg U43461 ( .A(n29161), .B(n29162), .X(\filter_0/n8478 ) );
  nand_x1_sg U43462 ( .A(n33462), .B(\filter_0/n8114 ), .X(n29162) );
  nand_x1_sg U43463 ( .A(n29370), .B(n29371), .X(\filter_0/n8379 ) );
  nand_x1_sg U43464 ( .A(n29975), .B(\filter_0/n8055 ), .X(n29371) );
  nand_x1_sg U43465 ( .A(n29372), .B(n29373), .X(\filter_0/n8378 ) );
  nand_x1_sg U43466 ( .A(n33442), .B(\filter_0/n8054 ), .X(n29373) );
  nand_x1_sg U43467 ( .A(n29249), .B(n29250), .X(\filter_0/n8436 ) );
  nand_x1_sg U43468 ( .A(n29261), .B(n29262), .X(\filter_0/n8430 ) );
  nand_x1_sg U43469 ( .A(n29273), .B(n29274), .X(\filter_0/n8424 ) );
  nand_x1_sg U43470 ( .A(n29257), .B(n29258), .X(\filter_0/n8432 ) );
  nand_x1_sg U43471 ( .A(n29269), .B(n29270), .X(\filter_0/n8426 ) );
  nand_x1_sg U43472 ( .A(n29253), .B(n29254), .X(\filter_0/n8434 ) );
  nand_x1_sg U43473 ( .A(n29265), .B(n29266), .X(\filter_0/n8428 ) );
  nand_x1_sg U43474 ( .A(n29243), .B(n29244), .X(\filter_0/n8439 ) );
  nand_x1_sg U43475 ( .A(n29957), .B(\filter_0/n8155 ), .X(n29244) );
  nand_x1_sg U43476 ( .A(n29019), .B(n29020), .X(\filter_0/n8543 ) );
  nand_x1_sg U43477 ( .A(n33315), .B(\filter_0/n8219 ), .X(n29020) );
  nand_x1_sg U43478 ( .A(n29023), .B(n29024), .X(\filter_0/n8542 ) );
  nand_x1_sg U43479 ( .A(n33318), .B(\filter_0/n8218 ), .X(n29024) );
  nand_x1_sg U43480 ( .A(n29025), .B(n29026), .X(\filter_0/n8541 ) );
  nand_x1_sg U43481 ( .A(n33315), .B(\filter_0/n8217 ), .X(n29026) );
  nand_x1_sg U43482 ( .A(n29027), .B(n29028), .X(\filter_0/n8540 ) );
  nand_x1_sg U43483 ( .A(n29925), .B(\filter_0/n8216 ), .X(n29028) );
  nand_x1_sg U43484 ( .A(n29191), .B(n29192), .X(\filter_0/n8463 ) );
  nand_x1_sg U43485 ( .A(n33436), .B(\filter_0/n8139 ), .X(n29192) );
  nand_x1_sg U43486 ( .A(n29195), .B(n29196), .X(\filter_0/n8462 ) );
  nand_x1_sg U43487 ( .A(n33437), .B(\filter_0/n8138 ), .X(n29196) );
  nand_x1_sg U43488 ( .A(n29197), .B(n29198), .X(\filter_0/n8461 ) );
  nand_x1_sg U43489 ( .A(n33436), .B(\filter_0/n8137 ), .X(n29198) );
  nand_x1_sg U43490 ( .A(n29199), .B(n29200), .X(\filter_0/n8460 ) );
  nand_x1_sg U43491 ( .A(n29973), .B(\filter_0/n8136 ), .X(n29200) );
  nand_x1_sg U43492 ( .A(n29318), .B(n29319), .X(\filter_0/n8403 ) );
  nand_x1_sg U43493 ( .A(n33313), .B(\filter_0/n8079 ), .X(n29319) );
  nand_x1_sg U43494 ( .A(n29322), .B(n29323), .X(\filter_0/n8402 ) );
  nand_x1_sg U43495 ( .A(n33310), .B(\filter_0/n8078 ), .X(n29323) );
  nand_x1_sg U43496 ( .A(n29324), .B(n29325), .X(\filter_0/n8401 ) );
  nand_x1_sg U43497 ( .A(n33311), .B(\filter_0/n8077 ), .X(n29325) );
  nand_x1_sg U43498 ( .A(n29326), .B(n29327), .X(\filter_0/n8400 ) );
  nand_x1_sg U43499 ( .A(n33311), .B(\filter_0/n8076 ), .X(n29327) );
  nand_x1_sg U43500 ( .A(n29461), .B(n29462), .X(\filter_0/n8336 ) );
  nand_x1_sg U43501 ( .A(n29465), .B(n29466), .X(\filter_0/n8334 ) );
  nand_x1_sg U43502 ( .A(n29469), .B(n29470), .X(\filter_0/n8332 ) );
  nand_x1_sg U43503 ( .A(n29473), .B(n29474), .X(\filter_0/n8330 ) );
  nand_x1_sg U43504 ( .A(n29477), .B(n29478), .X(\filter_0/n8328 ) );
  nand_x1_sg U43505 ( .A(n29481), .B(n29482), .X(\filter_0/n8326 ) );
  nand_x1_sg U43506 ( .A(n29485), .B(n29486), .X(\filter_0/n8324 ) );
  nand_x1_sg U43507 ( .A(n28976), .B(n28977), .X(\filter_0/n8563 ) );
  nand_x1_sg U43508 ( .A(n33306), .B(\filter_0/n8199 ), .X(n28977) );
  nand_x1_sg U43509 ( .A(n28980), .B(n28981), .X(\filter_0/n8562 ) );
  nand_x1_sg U43510 ( .A(n33305), .B(\filter_0/n8198 ), .X(n28981) );
  nand_x1_sg U43511 ( .A(n28982), .B(n28983), .X(\filter_0/n8561 ) );
  nand_x1_sg U43512 ( .A(n29921), .B(\filter_0/n8197 ), .X(n28983) );
  nand_x1_sg U43513 ( .A(n28984), .B(n28985), .X(\filter_0/n8560 ) );
  nand_x1_sg U43514 ( .A(n33307), .B(\filter_0/n8196 ), .X(n28985) );
  nand_x1_sg U43515 ( .A(n29149), .B(n29150), .X(\filter_0/n8483 ) );
  nand_x1_sg U43516 ( .A(n33463), .B(\filter_0/n8119 ), .X(n29150) );
  nand_x1_sg U43517 ( .A(n29153), .B(n29154), .X(\filter_0/n8482 ) );
  nand_x1_sg U43518 ( .A(n33460), .B(\filter_0/n8118 ), .X(n29154) );
  nand_x1_sg U43519 ( .A(n29155), .B(n29156), .X(\filter_0/n8481 ) );
  nand_x1_sg U43520 ( .A(n29983), .B(\filter_0/n8117 ), .X(n29156) );
  nand_x1_sg U43521 ( .A(n29157), .B(n29158), .X(\filter_0/n8480 ) );
  nand_x1_sg U43522 ( .A(n33461), .B(\filter_0/n8116 ), .X(n29158) );
  nand_x1_sg U43523 ( .A(n29360), .B(n29361), .X(\filter_0/n8383 ) );
  nand_x1_sg U43524 ( .A(n29975), .B(\filter_0/n8059 ), .X(n29361) );
  nand_x1_sg U43525 ( .A(n29364), .B(n29365), .X(\filter_0/n8382 ) );
  nand_x1_sg U43526 ( .A(n33442), .B(\filter_0/n8058 ), .X(n29365) );
  nand_x1_sg U43527 ( .A(n29366), .B(n29367), .X(\filter_0/n8381 ) );
  nand_x1_sg U43528 ( .A(n29975), .B(\filter_0/n8057 ), .X(n29367) );
  nand_x1_sg U43529 ( .A(n29368), .B(n29369), .X(\filter_0/n8380 ) );
  nand_x1_sg U43530 ( .A(n33442), .B(\filter_0/n8056 ), .X(n29369) );
  nand_x1_sg U43531 ( .A(n29455), .B(n29456), .X(\filter_0/n8339 ) );
  nand_x1_sg U43532 ( .A(n29959), .B(\filter_0/n7995 ), .X(n29456) );
  nand_x1_sg U43533 ( .A(n29504), .B(n29505), .X(\filter_0/n8317 ) );
  nand_x1_sg U43534 ( .A(n29508), .B(n29509), .X(\filter_0/n8315 ) );
  nand_x1_sg U43535 ( .A(n29512), .B(n29513), .X(\filter_0/n8313 ) );
  nand_x1_sg U43536 ( .A(n29516), .B(n29517), .X(\filter_0/n8311 ) );
  nand_x1_sg U43537 ( .A(n29520), .B(n29521), .X(\filter_0/n8309 ) );
  nand_x1_sg U43538 ( .A(n29524), .B(n29525), .X(\filter_0/n8307 ) );
  nand_x1_sg U43539 ( .A(n29528), .B(n29529), .X(\filter_0/n8305 ) );
  nand_x1_sg U43540 ( .A(n29548), .B(n29549), .X(\filter_0/n8297 ) );
  nand_x1_sg U43541 ( .A(n29552), .B(n29553), .X(\filter_0/n8295 ) );
  nand_x1_sg U43542 ( .A(n29556), .B(n29557), .X(\filter_0/n8293 ) );
  nand_x1_sg U43543 ( .A(n29560), .B(n29561), .X(\filter_0/n8291 ) );
  nand_x1_sg U43544 ( .A(n29564), .B(n29565), .X(\filter_0/n8289 ) );
  nand_x1_sg U43545 ( .A(n29568), .B(n29569), .X(\filter_0/n8287 ) );
  nand_x1_sg U43546 ( .A(n29572), .B(n29573), .X(\filter_0/n8285 ) );
  nand_x1_sg U43547 ( .A(n29233), .B(n29234), .X(\filter_0/n8443 ) );
  nand_x1_sg U43548 ( .A(n29957), .B(\filter_0/n8159 ), .X(n29234) );
  nand_x1_sg U43549 ( .A(n29239), .B(n29240), .X(\filter_0/n8441 ) );
  nand_x1_sg U43550 ( .A(n33398), .B(\filter_0/n8157 ), .X(n29240) );
  nand_x1_sg U43551 ( .A(n29451), .B(n29452), .X(\filter_0/n8341 ) );
  nand_x1_sg U43552 ( .A(n33400), .B(\filter_0/n7997 ), .X(n29452) );
  nand_x1_sg U43553 ( .A(n29245), .B(n29246), .X(\filter_0/n8438 ) );
  nand_x1_sg U43554 ( .A(n33395), .B(\filter_0/n8154 ), .X(n29246) );
  nand_x1_sg U43555 ( .A(n29445), .B(n29446), .X(\filter_0/n8343 ) );
  nand_x1_sg U43556 ( .A(n33400), .B(\filter_0/n7999 ), .X(n29446) );
  nand_x1_sg U43557 ( .A(n29550), .B(n29551), .X(\filter_0/n8296 ) );
  nand_x1_sg U43558 ( .A(n29554), .B(n29555), .X(\filter_0/n8294 ) );
  nand_x1_sg U43559 ( .A(n29558), .B(n29559), .X(\filter_0/n8292 ) );
  nand_x1_sg U43560 ( .A(n29562), .B(n29563), .X(\filter_0/n8290 ) );
  nand_x1_sg U43561 ( .A(n29566), .B(n29567), .X(\filter_0/n8288 ) );
  nand_x1_sg U43562 ( .A(n29570), .B(n29571), .X(\filter_0/n8286 ) );
  nand_x1_sg U43563 ( .A(n29574), .B(n29575), .X(\filter_0/n8284 ) );
  nand_x1_sg U43564 ( .A(n29457), .B(n29458), .X(\filter_0/n8338 ) );
  nand_x1_sg U43565 ( .A(n29959), .B(\filter_0/n7994 ), .X(n29458) );
  nand_x1_sg U43566 ( .A(n29506), .B(n29507), .X(\filter_0/n8316 ) );
  nand_x1_sg U43567 ( .A(n29510), .B(n29511), .X(\filter_0/n8314 ) );
  nand_x1_sg U43568 ( .A(n29514), .B(n29515), .X(\filter_0/n8312 ) );
  nand_x1_sg U43569 ( .A(n29518), .B(n29519), .X(\filter_0/n8310 ) );
  nand_x1_sg U43570 ( .A(n29522), .B(n29523), .X(\filter_0/n8308 ) );
  nand_x1_sg U43571 ( .A(n29526), .B(n29527), .X(\filter_0/n8306 ) );
  nand_x1_sg U43572 ( .A(n29530), .B(n29531), .X(\filter_0/n8304 ) );
  nand_x1_sg U43573 ( .A(n29237), .B(n29238), .X(\filter_0/n8442 ) );
  nand_x1_sg U43574 ( .A(n29957), .B(\filter_0/n8158 ), .X(n29238) );
  nand_x1_sg U43575 ( .A(n29241), .B(n29242), .X(\filter_0/n8440 ) );
  nand_x1_sg U43576 ( .A(n33397), .B(\filter_0/n8156 ), .X(n29242) );
  nand_x1_sg U43577 ( .A(n29500), .B(n29501), .X(\filter_0/n8319 ) );
  nand_x1_sg U43578 ( .A(n29919), .B(\filter_0/n7975 ), .X(n29501) );
  nand_x1_sg U43579 ( .A(n29544), .B(n29545), .X(\filter_0/n8299 ) );
  nand_x1_sg U43580 ( .A(n29917), .B(\filter_0/n7955 ), .X(n29545) );
  nand_x1_sg U43581 ( .A(n29449), .B(n29450), .X(\filter_0/n8342 ) );
  nand_x1_sg U43582 ( .A(n33403), .B(\filter_0/n7998 ), .X(n29450) );
  nand_x1_sg U43583 ( .A(n29453), .B(n29454), .X(\filter_0/n8340 ) );
  nand_x1_sg U43584 ( .A(n33403), .B(\filter_0/n7996 ), .X(n29454) );
  nand_x1_sg U43585 ( .A(n29496), .B(n29497), .X(\filter_0/n8321 ) );
  nand_x1_sg U43586 ( .A(n33300), .B(\filter_0/n7977 ), .X(n29497) );
  nand_x1_sg U43587 ( .A(n29540), .B(n29541), .X(\filter_0/n8301 ) );
  nand_x1_sg U43588 ( .A(n33295), .B(\filter_0/n7957 ), .X(n29541) );
  nand_x1_sg U43589 ( .A(n29490), .B(n29491), .X(\filter_0/n8323 ) );
  nand_x1_sg U43590 ( .A(n33301), .B(\filter_0/n7979 ), .X(n29491) );
  nand_x1_sg U43591 ( .A(n29534), .B(n29535), .X(\filter_0/n8303 ) );
  nand_x1_sg U43592 ( .A(n33297), .B(\filter_0/n7959 ), .X(n29535) );
  nand_x1_sg U43593 ( .A(n29546), .B(n29547), .X(\filter_0/n8298 ) );
  nand_x1_sg U43594 ( .A(n33298), .B(\filter_0/n7954 ), .X(n29547) );
  nand_x1_sg U43595 ( .A(n29502), .B(n29503), .X(\filter_0/n8318 ) );
  nand_x1_sg U43596 ( .A(n33303), .B(\filter_0/n7974 ), .X(n29503) );
  nand_x1_sg U43597 ( .A(n19603), .B(n19604), .X(\shifter_0/n10883 ) );
  nand_x1_sg U43598 ( .A(n29494), .B(n29495), .X(\filter_0/n8322 ) );
  nand_x1_sg U43599 ( .A(n33301), .B(\filter_0/n7978 ), .X(n29495) );
  nand_x1_sg U43600 ( .A(n29538), .B(n29539), .X(\filter_0/n8302 ) );
  nand_x1_sg U43601 ( .A(n33298), .B(\filter_0/n7958 ), .X(n29539) );
  nand_x1_sg U43602 ( .A(n29498), .B(n29499), .X(\filter_0/n8320 ) );
  nand_x1_sg U43603 ( .A(n29919), .B(\filter_0/n7976 ), .X(n29499) );
  nand_x1_sg U43604 ( .A(n29542), .B(n29543), .X(\filter_0/n8300 ) );
  nand_x1_sg U43605 ( .A(n33296), .B(\filter_0/n7956 ), .X(n29543) );
  nand_x1_sg U43606 ( .A(n26036), .B(n26037), .X(n4074) );
  nand_x1_sg U43607 ( .A(n26040), .B(n26041), .X(n4072) );
  nand_x1_sg U43608 ( .A(n26042), .B(n26043), .X(n4071) );
  nand_x1_sg U43609 ( .A(n26046), .B(n26047), .X(n4069) );
  nand_x1_sg U43610 ( .A(n26048), .B(n26049), .X(n4068) );
  nand_x1_sg U43611 ( .A(n26052), .B(n26053), .X(n4066) );
  nand_x1_sg U43612 ( .A(n26054), .B(n26055), .X(n4065) );
  nand_x1_sg U43613 ( .A(n26058), .B(n26059), .X(n4063) );
  nand_x1_sg U43614 ( .A(n26060), .B(n26061), .X(n4062) );
  nand_x1_sg U43615 ( .A(n26064), .B(n26065), .X(n4060) );
  nand_x1_sg U43616 ( .A(n26130), .B(n26131), .X(n4027) );
  nand_x1_sg U43617 ( .A(n26132), .B(n26133), .X(n4026) );
  nand_x1_sg U43618 ( .A(n26136), .B(n26137), .X(n4024) );
  nand_x1_sg U43619 ( .A(n26138), .B(n26139), .X(n4023) );
  nand_x1_sg U43620 ( .A(n26142), .B(n26143), .X(n4021) );
  nand_x1_sg U43621 ( .A(n26144), .B(n26145), .X(n4020) );
  nand_x1_sg U43622 ( .A(n26148), .B(n26149), .X(n4018) );
  nand_x1_sg U43623 ( .A(n26150), .B(n26151), .X(n4017) );
  nand_x1_sg U43624 ( .A(n25428), .B(n25429), .X(n4378) );
  nand_x1_sg U43625 ( .A(n25430), .B(n25431), .X(n4377) );
  nand_x1_sg U43626 ( .A(n25434), .B(n25435), .X(n4375) );
  nand_x1_sg U43627 ( .A(n25436), .B(n25437), .X(n4374) );
  nand_x1_sg U43628 ( .A(n25482), .B(n25483), .X(n4351) );
  nand_x1_sg U43629 ( .A(n25484), .B(n25485), .X(n4350) );
  nand_x1_sg U43630 ( .A(n25488), .B(n25489), .X(n4348) );
  nand_x1_sg U43631 ( .A(n25560), .B(n25561), .X(n4312) );
  nand_x1_sg U43632 ( .A(n25562), .B(n25563), .X(n4311) );
  nand_x1_sg U43633 ( .A(n25566), .B(n25567), .X(n4309) );
  nand_x1_sg U43634 ( .A(n25568), .B(n25569), .X(n4308) );
  nand_x1_sg U43635 ( .A(n25572), .B(n25573), .X(n4306) );
  nand_x1_sg U43636 ( .A(n25574), .B(n25575), .X(n4305) );
  nand_x1_sg U43637 ( .A(n25578), .B(n25579), .X(n4303) );
  nand_x1_sg U43638 ( .A(n25580), .B(n25581), .X(n4302) );
  nand_x1_sg U43639 ( .A(n25584), .B(n25585), .X(n4300) );
  nand_x1_sg U43640 ( .A(n25586), .B(n25587), .X(n4299) );
  nand_x1_sg U43641 ( .A(n25590), .B(n25591), .X(n4297) );
  nand_x1_sg U43642 ( .A(n25592), .B(n25593), .X(n4296) );
  nand_x1_sg U43643 ( .A(n25596), .B(n25597), .X(n4294) );
  nand_x1_sg U43644 ( .A(n25598), .B(n25599), .X(n4293) );
  nand_x1_sg U43645 ( .A(n25722), .B(n25723), .X(n4231) );
  nand_x1_sg U43646 ( .A(n25724), .B(n25725), .X(n4230) );
  nand_x1_sg U43647 ( .A(n25728), .B(n25729), .X(n4228) );
  nand_x1_sg U43648 ( .A(n25730), .B(n25731), .X(n4227) );
  nand_x1_sg U43649 ( .A(n25734), .B(n25735), .X(n4225) );
  nand_x1_sg U43650 ( .A(n25736), .B(n25737), .X(n4224) );
  nand_x1_sg U43651 ( .A(n25740), .B(n25741), .X(n4222) );
  nand_x1_sg U43652 ( .A(n25742), .B(n25743), .X(n4221) );
  nand_x1_sg U43653 ( .A(n25002), .B(n25003), .X(n4591) );
  nand_x1_sg U43654 ( .A(n25004), .B(n25005), .X(n4590) );
  nand_x1_sg U43655 ( .A(n25008), .B(n25009), .X(n4588) );
  nand_x1_sg U43656 ( .A(n25010), .B(n25011), .X(n4587) );
  nand_x1_sg U43657 ( .A(n25014), .B(n25015), .X(n4585) );
  nand_x1_sg U43658 ( .A(n25016), .B(n25017), .X(n4584) );
  nand_x1_sg U43659 ( .A(n25020), .B(n25021), .X(n4582) );
  nand_x1_sg U43660 ( .A(n25022), .B(n25023), .X(n4581) );
  nand_x1_sg U43661 ( .A(n25026), .B(n25027), .X(n4579) );
  nand_x1_sg U43662 ( .A(n25028), .B(n25029), .X(n4578) );
  nand_x1_sg U43663 ( .A(n25032), .B(n25033), .X(n4576) );
  nand_x1_sg U43664 ( .A(n25034), .B(n25035), .X(n4575) );
  nand_x1_sg U43665 ( .A(n25038), .B(n25039), .X(n4573) );
  nand_x1_sg U43666 ( .A(n25040), .B(n25041), .X(n4572) );
  nand_x1_sg U43667 ( .A(n25106), .B(n25107), .X(n4539) );
  nand_x1_sg U43668 ( .A(n25110), .B(n25111), .X(n4537) );
  nand_x1_sg U43669 ( .A(n25112), .B(n25113), .X(n4536) );
  nand_x1_sg U43670 ( .A(n25116), .B(n25117), .X(n4534) );
  nand_x1_sg U43671 ( .A(n25118), .B(n25119), .X(n4533) );
  nand_x1_sg U43672 ( .A(n25122), .B(n25123), .X(n4531) );
  nand_x1_sg U43673 ( .A(n25164), .B(n25165), .X(n4510) );
  nand_x1_sg U43674 ( .A(n25166), .B(n25167), .X(n4509) );
  nand_x1_sg U43675 ( .A(n24852), .B(n24853), .X(n4666) );
  nand_x1_sg U43676 ( .A(n24854), .B(n24855), .X(n4665) );
  nand_x1_sg U43677 ( .A(n24858), .B(n24859), .X(n4663) );
  nand_x1_sg U43678 ( .A(n24860), .B(n24861), .X(n4662) );
  nand_x1_sg U43679 ( .A(n24864), .B(n24865), .X(n4660) );
  nand_x1_sg U43680 ( .A(n24866), .B(n24867), .X(n4659) );
  nand_x1_sg U43681 ( .A(n24870), .B(n24871), .X(n4657) );
  nand_x1_sg U43682 ( .A(n24872), .B(n24873), .X(n4656) );
  nand_x1_sg U43683 ( .A(n24876), .B(n24877), .X(n4654) );
  nand_x1_sg U43684 ( .A(n24878), .B(n24879), .X(n4653) );
  nand_x1_sg U43685 ( .A(n24882), .B(n24883), .X(n4651) );
  nand_x1_sg U43686 ( .A(n24884), .B(n24885), .X(n4650) );
  nand_x1_sg U43687 ( .A(n24294), .B(n24295), .X(n4945) );
  nand_x1_sg U43688 ( .A(n24296), .B(n24297), .X(n4944) );
  nand_x1_sg U43689 ( .A(n24300), .B(n24301), .X(n4942) );
  nand_x1_sg U43690 ( .A(n24302), .B(n24303), .X(n4941) );
  nand_x1_sg U43691 ( .A(n24306), .B(n24307), .X(n4939) );
  nand_x1_sg U43692 ( .A(n24308), .B(n24309), .X(n4938) );
  nand_x1_sg U43693 ( .A(n24312), .B(n24313), .X(n4936) );
  nand_x1_sg U43694 ( .A(n24314), .B(n24315), .X(n4935) );
  nand_x1_sg U43695 ( .A(n24318), .B(n24319), .X(n4933) );
  nand_x1_sg U43696 ( .A(n24320), .B(n24321), .X(n4932) );
  nand_x1_sg U43697 ( .A(n24324), .B(n24325), .X(n4930) );
  nand_x1_sg U43698 ( .A(n24326), .B(n24327), .X(n4929) );
  nand_x1_sg U43699 ( .A(n24330), .B(n24331), .X(n4927) );
  nand_x1_sg U43700 ( .A(n24402), .B(n24403), .X(n4891) );
  nand_x1_sg U43701 ( .A(n24404), .B(n24405), .X(n4890) );
  nand_x1_sg U43702 ( .A(n24408), .B(n24409), .X(n4888) );
  nand_x1_sg U43703 ( .A(n24410), .B(n24411), .X(n4887) );
  nand_x1_sg U43704 ( .A(n24452), .B(n24453), .X(n4866) );
  nand_x1_sg U43705 ( .A(n24456), .B(n24457), .X(n4864) );
  nand_x1_sg U43706 ( .A(n24458), .B(n24459), .X(n4863) );
  nand_x1_sg U43707 ( .A(n24462), .B(n24463), .X(n4861) );
  nand_x1_sg U43708 ( .A(n24464), .B(n24465), .X(n4860) );
  nand_x1_sg U43709 ( .A(n24534), .B(n24535), .X(n4825) );
  nand_x1_sg U43710 ( .A(n24536), .B(n24537), .X(n4824) );
  nand_x1_sg U43711 ( .A(n24540), .B(n24541), .X(n4822) );
  nand_x1_sg U43712 ( .A(n24542), .B(n24543), .X(n4821) );
  nand_x1_sg U43713 ( .A(n24546), .B(n24547), .X(n4819) );
  nand_x1_sg U43714 ( .A(n24548), .B(n24549), .X(n4818) );
  nand_x1_sg U43715 ( .A(n24552), .B(n24553), .X(n4816) );
  nand_x1_sg U43716 ( .A(n24554), .B(n24555), .X(n4815) );
  nand_x1_sg U43717 ( .A(n24558), .B(n24559), .X(n4813) );
  nand_x1_sg U43718 ( .A(n24560), .B(n24561), .X(n4812) );
  nand_x1_sg U43719 ( .A(n23826), .B(n23827), .X(n5179) );
  nand_x1_sg U43720 ( .A(n23828), .B(n23829), .X(n5178) );
  nand_x1_sg U43721 ( .A(n23832), .B(n23833), .X(n5176) );
  nand_x1_sg U43722 ( .A(n23834), .B(n23835), .X(n5175) );
  nand_x1_sg U43723 ( .A(n23838), .B(n23839), .X(n5173) );
  nand_x1_sg U43724 ( .A(n23840), .B(n23841), .X(n5172) );
  nand_x1_sg U43725 ( .A(n23844), .B(n23845), .X(n5170) );
  nand_x1_sg U43726 ( .A(n23846), .B(n23847), .X(n5169) );
  nand_x1_sg U43727 ( .A(n23850), .B(n23851), .X(n5167) );
  nand_x1_sg U43728 ( .A(n23852), .B(n23853), .X(n5166) );
  nand_x1_sg U43729 ( .A(n23976), .B(n23977), .X(n5104) );
  nand_x1_sg U43730 ( .A(n23978), .B(n23979), .X(n5103) );
  nand_x1_sg U43731 ( .A(n23982), .B(n23983), .X(n5101) );
  nand_x1_sg U43732 ( .A(n23984), .B(n23985), .X(n5100) );
  nand_x1_sg U43733 ( .A(n23988), .B(n23989), .X(n5098) );
  nand_x1_sg U43734 ( .A(n23990), .B(n23991), .X(n5097) );
  nand_x1_sg U43735 ( .A(n23994), .B(n23995), .X(n5095) );
  nand_x1_sg U43736 ( .A(n23996), .B(n23997), .X(n5094) );
  nand_x1_sg U43737 ( .A(n24000), .B(n24001), .X(n5092) );
  nand_x1_sg U43738 ( .A(n24002), .B(n24003), .X(n5091) );
  nand_x1_sg U43739 ( .A(n24006), .B(n24007), .X(n5089) );
  nand_x1_sg U43740 ( .A(n24008), .B(n24009), .X(n5088) );
  nand_x1_sg U43741 ( .A(n24012), .B(n24013), .X(n5086) );
  nand_x1_sg U43742 ( .A(n24014), .B(n24015), .X(n5085) );
  nand_x1_sg U43743 ( .A(n23726), .B(n23727), .X(n5229) );
  nand_x1_sg U43744 ( .A(n23730), .B(n23731), .X(n5227) );
  nand_x1_sg U43745 ( .A(n23732), .B(n23733), .X(n5226) );
  nand_x1_sg U43746 ( .A(n23736), .B(n23737), .X(n5224) );
  nand_x1_sg U43747 ( .A(n23738), .B(n23739), .X(n5223) );
  nand_x1_sg U43748 ( .A(n23742), .B(n23743), .X(n5221) );
  nand_x1_sg U43749 ( .A(n23744), .B(n23745), .X(n5220) );
  nand_x1_sg U43750 ( .A(n23748), .B(n23749), .X(n5218) );
  nand_x1_sg U43751 ( .A(n23750), .B(n23751), .X(n5217) );
  nand_x1_sg U43752 ( .A(n23754), .B(n23755), .X(n5215) );
  nand_x1_sg U43753 ( .A(n23756), .B(n23757), .X(n5214) );
  nand_x1_sg U43754 ( .A(n23760), .B(n23761), .X(n5212) );
  nand_x1_sg U43755 ( .A(n26038), .B(n26039), .X(n4073) );
  nand_x1_sg U43756 ( .A(n26044), .B(n26045), .X(n4070) );
  nand_x1_sg U43757 ( .A(n26050), .B(n26051), .X(n4067) );
  nand_x1_sg U43758 ( .A(n26056), .B(n26057), .X(n4064) );
  nand_x1_sg U43759 ( .A(n26062), .B(n26063), .X(n4061) );
  nand_x1_sg U43760 ( .A(n26134), .B(n26135), .X(n4025) );
  nand_x1_sg U43761 ( .A(n26140), .B(n26141), .X(n4022) );
  nand_x1_sg U43762 ( .A(n26146), .B(n26147), .X(n4019) );
  nand_x1_sg U43763 ( .A(n26152), .B(n26153), .X(n4016) );
  nand_x1_sg U43764 ( .A(n25426), .B(n25427), .X(n4379) );
  nand_x1_sg U43765 ( .A(n25432), .B(n25433), .X(n4376) );
  nand_x1_sg U43766 ( .A(n25438), .B(n25439), .X(n4373) );
  nand_x1_sg U43767 ( .A(n25480), .B(n25481), .X(n4352) );
  nand_x1_sg U43768 ( .A(n25486), .B(n25487), .X(n4349) );
  nand_x1_sg U43769 ( .A(n25564), .B(n25565), .X(n4310) );
  nand_x1_sg U43770 ( .A(n25570), .B(n25571), .X(n4307) );
  nand_x1_sg U43771 ( .A(n25576), .B(n25577), .X(n4304) );
  nand_x1_sg U43772 ( .A(n25582), .B(n25583), .X(n4301) );
  nand_x1_sg U43773 ( .A(n25588), .B(n25589), .X(n4298) );
  nand_x1_sg U43774 ( .A(n25594), .B(n25595), .X(n4295) );
  nand_x1_sg U43775 ( .A(n25720), .B(n25721), .X(n4232) );
  nand_x1_sg U43776 ( .A(n25726), .B(n25727), .X(n4229) );
  nand_x1_sg U43777 ( .A(n25732), .B(n25733), .X(n4226) );
  nand_x1_sg U43778 ( .A(n25738), .B(n25739), .X(n4223) );
  nand_x1_sg U43779 ( .A(n25744), .B(n25745), .X(n4220) );
  nand_x1_sg U43780 ( .A(n25000), .B(n25001), .X(n4592) );
  nand_x1_sg U43781 ( .A(n25006), .B(n25007), .X(n4589) );
  nand_x1_sg U43782 ( .A(n25012), .B(n25013), .X(n4586) );
  nand_x1_sg U43783 ( .A(n25018), .B(n25019), .X(n4583) );
  nand_x1_sg U43784 ( .A(n25024), .B(n25025), .X(n4580) );
  nand_x1_sg U43785 ( .A(n25030), .B(n25031), .X(n4577) );
  nand_x1_sg U43786 ( .A(n25036), .B(n25037), .X(n4574) );
  nand_x1_sg U43787 ( .A(n25108), .B(n25109), .X(n4538) );
  nand_x1_sg U43788 ( .A(n25114), .B(n25115), .X(n4535) );
  nand_x1_sg U43789 ( .A(n25120), .B(n25121), .X(n4532) );
  nand_x1_sg U43790 ( .A(n25168), .B(n25169), .X(n4508) );
  nand_x1_sg U43791 ( .A(n24850), .B(n24851), .X(n4667) );
  nand_x1_sg U43792 ( .A(n24856), .B(n24857), .X(n4664) );
  nand_x1_sg U43793 ( .A(n24862), .B(n24863), .X(n4661) );
  nand_x1_sg U43794 ( .A(n24868), .B(n24869), .X(n4658) );
  nand_x1_sg U43795 ( .A(n24874), .B(n24875), .X(n4655) );
  nand_x1_sg U43796 ( .A(n24880), .B(n24881), .X(n4652) );
  nand_x1_sg U43797 ( .A(n24886), .B(n24887), .X(n4649) );
  nand_x1_sg U43798 ( .A(n24292), .B(n24293), .X(n4946) );
  nand_x1_sg U43799 ( .A(n24298), .B(n24299), .X(n4943) );
  nand_x1_sg U43800 ( .A(n24304), .B(n24305), .X(n4940) );
  nand_x1_sg U43801 ( .A(n24310), .B(n24311), .X(n4937) );
  nand_x1_sg U43802 ( .A(n24316), .B(n24317), .X(n4934) );
  nand_x1_sg U43803 ( .A(n24322), .B(n24323), .X(n4931) );
  nand_x1_sg U43804 ( .A(n24328), .B(n24329), .X(n4928) );
  nand_x1_sg U43805 ( .A(n24406), .B(n24407), .X(n4889) );
  nand_x1_sg U43806 ( .A(n24454), .B(n24455), .X(n4865) );
  nand_x1_sg U43807 ( .A(n24460), .B(n24461), .X(n4862) );
  nand_x1_sg U43808 ( .A(n24532), .B(n24533), .X(n4826) );
  nand_x1_sg U43809 ( .A(n24538), .B(n24539), .X(n4823) );
  nand_x1_sg U43810 ( .A(n24544), .B(n24545), .X(n4820) );
  nand_x1_sg U43811 ( .A(n24550), .B(n24551), .X(n4817) );
  nand_x1_sg U43812 ( .A(n24556), .B(n24557), .X(n4814) );
  nand_x1_sg U43813 ( .A(n23830), .B(n23831), .X(n5177) );
  nand_x1_sg U43814 ( .A(n23836), .B(n23837), .X(n5174) );
  nand_x1_sg U43815 ( .A(n23842), .B(n23843), .X(n5171) );
  nand_x1_sg U43816 ( .A(n23848), .B(n23849), .X(n5168) );
  nand_x1_sg U43817 ( .A(n23854), .B(n23855), .X(n5165) );
  nand_x1_sg U43818 ( .A(n23980), .B(n23981), .X(n5102) );
  nand_x1_sg U43819 ( .A(n23986), .B(n23987), .X(n5099) );
  nand_x1_sg U43820 ( .A(n23992), .B(n23993), .X(n5096) );
  nand_x1_sg U43821 ( .A(n23998), .B(n23999), .X(n5093) );
  nand_x1_sg U43822 ( .A(n24004), .B(n24005), .X(n5090) );
  nand_x1_sg U43823 ( .A(n24010), .B(n24011), .X(n5087) );
  nand_x1_sg U43824 ( .A(n23728), .B(n23729), .X(n5228) );
  nand_x1_sg U43825 ( .A(n23734), .B(n23735), .X(n5225) );
  nand_x1_sg U43826 ( .A(n23740), .B(n23741), .X(n5222) );
  nand_x1_sg U43827 ( .A(n23746), .B(n23747), .X(n5219) );
  nand_x1_sg U43828 ( .A(n23752), .B(n23753), .X(n5216) );
  nand_x1_sg U43829 ( .A(n23758), .B(n23759), .X(n5213) );
  inv_x1_sg U43830 ( .A(n15345), .X(n42388) );
  nand_x1_sg U43831 ( .A(n26004), .B(n26005), .X(n4090) );
  nand_x1_sg U43832 ( .A(n26006), .B(n26007), .X(n4089) );
  nand_x1_sg U43833 ( .A(n26010), .B(n26011), .X(n4087) );
  nand_x1_sg U43834 ( .A(n26012), .B(n26013), .X(n4086) );
  nand_x1_sg U43835 ( .A(n26016), .B(n26017), .X(n4084) );
  nand_x1_sg U43836 ( .A(n26018), .B(n26019), .X(n4083) );
  nand_x1_sg U43837 ( .A(n26022), .B(n26023), .X(n4081) );
  nand_x1_sg U43838 ( .A(n26024), .B(n26025), .X(n4080) );
  nand_x1_sg U43839 ( .A(n26028), .B(n26029), .X(n4078) );
  nand_x1_sg U43840 ( .A(n26030), .B(n26031), .X(n4077) );
  nand_x1_sg U43841 ( .A(n26034), .B(n26035), .X(n4075) );
  nand_x1_sg U43842 ( .A(n26154), .B(n26155), .X(n4015) );
  nand_x1_sg U43843 ( .A(n26156), .B(n26157), .X(n4014) );
  nand_x1_sg U43844 ( .A(n26160), .B(n26161), .X(n4012) );
  nand_x1_sg U43845 ( .A(n26162), .B(n26163), .X(n4011) );
  nand_x1_sg U43846 ( .A(n26166), .B(n26167), .X(n4009) );
  nand_x1_sg U43847 ( .A(n26168), .B(n26169), .X(n4008) );
  nand_x1_sg U43848 ( .A(n26172), .B(n26173), .X(n4006) );
  nand_x1_sg U43849 ( .A(n26174), .B(n26175), .X(n4005) );
  nand_x1_sg U43850 ( .A(n26178), .B(n26179), .X(n4003) );
  nand_x1_sg U43851 ( .A(n26180), .B(n26181), .X(n4002) );
  nand_x1_sg U43852 ( .A(n26184), .B(n26185), .X(n4000) );
  nand_x1_sg U43853 ( .A(n26186), .B(n26187), .X(n3999) );
  nand_x1_sg U43854 ( .A(n26190), .B(n26191), .X(n3997) );
  nand_x1_sg U43855 ( .A(n26192), .B(n26193), .X(n3996) );
  nand_x1_sg U43856 ( .A(n25440), .B(n25441), .X(n4372) );
  nand_x1_sg U43857 ( .A(n25442), .B(n25443), .X(n4371) );
  nand_x1_sg U43858 ( .A(n25446), .B(n25447), .X(n4369) );
  nand_x1_sg U43859 ( .A(n25448), .B(n25449), .X(n4368) );
  nand_x1_sg U43860 ( .A(n25452), .B(n25453), .X(n4366) );
  nand_x1_sg U43861 ( .A(n25454), .B(n25455), .X(n4365) );
  nand_x1_sg U43862 ( .A(n25458), .B(n25459), .X(n4363) );
  nand_x1_sg U43863 ( .A(n25460), .B(n25461), .X(n4362) );
  nand_x1_sg U43864 ( .A(n25464), .B(n25465), .X(n4360) );
  nand_x1_sg U43865 ( .A(n25466), .B(n25467), .X(n4359) );
  nand_x1_sg U43866 ( .A(n25470), .B(n25471), .X(n4357) );
  nand_x1_sg U43867 ( .A(n25472), .B(n25473), .X(n4356) );
  nand_x1_sg U43868 ( .A(n25476), .B(n25477), .X(n4354) );
  nand_x1_sg U43869 ( .A(n25478), .B(n25479), .X(n4353) );
  nand_x1_sg U43870 ( .A(n25554), .B(n25555), .X(n4315) );
  nand_x1_sg U43871 ( .A(n25556), .B(n25557), .X(n4314) );
  nand_x1_sg U43872 ( .A(n25602), .B(n25603), .X(n4291) );
  nand_x1_sg U43873 ( .A(n25604), .B(n25605), .X(n4290) );
  nand_x1_sg U43874 ( .A(n25608), .B(n25609), .X(n4288) );
  nand_x1_sg U43875 ( .A(n25610), .B(n25611), .X(n4287) );
  nand_x1_sg U43876 ( .A(n25614), .B(n25615), .X(n4285) );
  nand_x1_sg U43877 ( .A(n25616), .B(n25617), .X(n4284) );
  nand_x1_sg U43878 ( .A(n25682), .B(n25683), .X(n4251) );
  nand_x1_sg U43879 ( .A(n25686), .B(n25687), .X(n4249) );
  nand_x1_sg U43880 ( .A(n25688), .B(n25689), .X(n4248) );
  nand_x1_sg U43881 ( .A(n25692), .B(n25693), .X(n4246) );
  nand_x1_sg U43882 ( .A(n25694), .B(n25695), .X(n4245) );
  nand_x1_sg U43883 ( .A(n25698), .B(n25699), .X(n4243) );
  nand_x1_sg U43884 ( .A(n25700), .B(n25701), .X(n4242) );
  nand_x1_sg U43885 ( .A(n25704), .B(n25705), .X(n4240) );
  nand_x1_sg U43886 ( .A(n25706), .B(n25707), .X(n4239) );
  nand_x1_sg U43887 ( .A(n25710), .B(n25711), .X(n4237) );
  nand_x1_sg U43888 ( .A(n25712), .B(n25713), .X(n4236) );
  nand_x1_sg U43889 ( .A(n25716), .B(n25717), .X(n4234) );
  nand_x1_sg U43890 ( .A(n25718), .B(n25719), .X(n4233) );
  nand_x1_sg U43891 ( .A(n25124), .B(n25125), .X(n4530) );
  nand_x1_sg U43892 ( .A(n25128), .B(n25129), .X(n4528) );
  nand_x1_sg U43893 ( .A(n25130), .B(n25131), .X(n4527) );
  nand_x1_sg U43894 ( .A(n25134), .B(n25135), .X(n4525) );
  nand_x1_sg U43895 ( .A(n25136), .B(n25137), .X(n4524) );
  nand_x1_sg U43896 ( .A(n25140), .B(n25141), .X(n4522) );
  nand_x1_sg U43897 ( .A(n25142), .B(n25143), .X(n4521) );
  nand_x1_sg U43898 ( .A(n25146), .B(n25147), .X(n4519) );
  nand_x1_sg U43899 ( .A(n25148), .B(n25149), .X(n4518) );
  nand_x1_sg U43900 ( .A(n25152), .B(n25153), .X(n4516) );
  nand_x1_sg U43901 ( .A(n25154), .B(n25155), .X(n4515) );
  nand_x1_sg U43902 ( .A(n25158), .B(n25159), .X(n4513) );
  nand_x1_sg U43903 ( .A(n25160), .B(n25161), .X(n4512) );
  nand_x1_sg U43904 ( .A(n24888), .B(n24889), .X(n4648) );
  nand_x1_sg U43905 ( .A(n24890), .B(n24891), .X(n4647) );
  nand_x1_sg U43906 ( .A(n24894), .B(n24895), .X(n4645) );
  nand_x1_sg U43907 ( .A(n24896), .B(n24897), .X(n4644) );
  nand_x1_sg U43908 ( .A(n24900), .B(n24901), .X(n4642) );
  nand_x1_sg U43909 ( .A(n24902), .B(n24903), .X(n4641) );
  nand_x1_sg U43910 ( .A(n24906), .B(n24907), .X(n4639) );
  nand_x1_sg U43911 ( .A(n24908), .B(n24909), .X(n4638) );
  nand_x1_sg U43912 ( .A(n24912), .B(n24913), .X(n4636) );
  nand_x1_sg U43913 ( .A(n24978), .B(n24979), .X(n4603) );
  nand_x1_sg U43914 ( .A(n24980), .B(n24981), .X(n4602) );
  nand_x1_sg U43915 ( .A(n24984), .B(n24985), .X(n4600) );
  nand_x1_sg U43916 ( .A(n24986), .B(n24987), .X(n4599) );
  nand_x1_sg U43917 ( .A(n24990), .B(n24991), .X(n4597) );
  nand_x1_sg U43918 ( .A(n24992), .B(n24993), .X(n4596) );
  nand_x1_sg U43919 ( .A(n24996), .B(n24997), .X(n4594) );
  nand_x1_sg U43920 ( .A(n24998), .B(n24999), .X(n4593) );
  nand_x1_sg U43921 ( .A(n24276), .B(n24277), .X(n4954) );
  nand_x1_sg U43922 ( .A(n24278), .B(n24279), .X(n4953) );
  nand_x1_sg U43923 ( .A(n24282), .B(n24283), .X(n4951) );
  nand_x1_sg U43924 ( .A(n24284), .B(n24285), .X(n4950) );
  nand_x1_sg U43925 ( .A(n24288), .B(n24289), .X(n4948) );
  nand_x1_sg U43926 ( .A(n24290), .B(n24291), .X(n4947) );
  nand_x1_sg U43927 ( .A(n24332), .B(n24333), .X(n4926) );
  nand_x1_sg U43928 ( .A(n24336), .B(n24337), .X(n4924) );
  nand_x1_sg U43929 ( .A(n24414), .B(n24415), .X(n4885) );
  nand_x1_sg U43930 ( .A(n24416), .B(n24417), .X(n4884) );
  nand_x1_sg U43931 ( .A(n24420), .B(n24421), .X(n4882) );
  nand_x1_sg U43932 ( .A(n24422), .B(n24423), .X(n4881) );
  nand_x1_sg U43933 ( .A(n24426), .B(n24427), .X(n4879) );
  nand_x1_sg U43934 ( .A(n24428), .B(n24429), .X(n4878) );
  nand_x1_sg U43935 ( .A(n24432), .B(n24433), .X(n4876) );
  nand_x1_sg U43936 ( .A(n24434), .B(n24435), .X(n4875) );
  nand_x1_sg U43937 ( .A(n24438), .B(n24439), .X(n4873) );
  nand_x1_sg U43938 ( .A(n24440), .B(n24441), .X(n4872) );
  nand_x1_sg U43939 ( .A(n24444), .B(n24445), .X(n4870) );
  nand_x1_sg U43940 ( .A(n24446), .B(n24447), .X(n4869) );
  nand_x1_sg U43941 ( .A(n24450), .B(n24451), .X(n4867) );
  nand_x1_sg U43942 ( .A(n24530), .B(n24531), .X(n4827) );
  nand_x1_sg U43943 ( .A(n24564), .B(n24565), .X(n4810) );
  nand_x1_sg U43944 ( .A(n24566), .B(n24567), .X(n4809) );
  nand_x1_sg U43945 ( .A(n24570), .B(n24571), .X(n4807) );
  nand_x1_sg U43946 ( .A(n24572), .B(n24573), .X(n4806) );
  nand_x1_sg U43947 ( .A(n24576), .B(n24577), .X(n4804) );
  nand_x1_sg U43948 ( .A(n24578), .B(n24579), .X(n4803) );
  nand_x1_sg U43949 ( .A(n24582), .B(n24583), .X(n4801) );
  nand_x1_sg U43950 ( .A(n24584), .B(n24585), .X(n4800) );
  nand_x1_sg U43951 ( .A(n24588), .B(n24589), .X(n4798) );
  nand_x1_sg U43952 ( .A(n24590), .B(n24591), .X(n4797) );
  nand_x1_sg U43953 ( .A(n23856), .B(n23857), .X(n5164) );
  nand_x1_sg U43954 ( .A(n23858), .B(n23859), .X(n5163) );
  nand_x1_sg U43955 ( .A(n23862), .B(n23863), .X(n5161) );
  nand_x1_sg U43956 ( .A(n23864), .B(n23865), .X(n5160) );
  nand_x1_sg U43957 ( .A(n23868), .B(n23869), .X(n5158) );
  nand_x1_sg U43958 ( .A(n23870), .B(n23871), .X(n5157) );
  nand_x1_sg U43959 ( .A(n23874), .B(n23875), .X(n5155) );
  nand_x1_sg U43960 ( .A(n23876), .B(n23877), .X(n5154) );
  nand_x1_sg U43961 ( .A(n23880), .B(n23881), .X(n5152) );
  nand_x1_sg U43962 ( .A(n23882), .B(n23883), .X(n5151) );
  nand_x1_sg U43963 ( .A(n23886), .B(n23887), .X(n5149) );
  nand_x1_sg U43964 ( .A(n23888), .B(n23889), .X(n5148) );
  nand_x1_sg U43965 ( .A(n23954), .B(n23955), .X(n5115) );
  nand_x1_sg U43966 ( .A(n23958), .B(n23959), .X(n5113) );
  nand_x1_sg U43967 ( .A(n23960), .B(n23961), .X(n5112) );
  nand_x1_sg U43968 ( .A(n23964), .B(n23965), .X(n5110) );
  nand_x1_sg U43969 ( .A(n23966), .B(n23967), .X(n5109) );
  nand_x1_sg U43970 ( .A(n23970), .B(n23971), .X(n5107) );
  nand_x1_sg U43971 ( .A(n23972), .B(n23973), .X(n5106) );
  nand_x1_sg U43972 ( .A(n23700), .B(n23701), .X(n5242) );
  nand_x1_sg U43973 ( .A(n23702), .B(n23703), .X(n5241) );
  nand_x1_sg U43974 ( .A(n23706), .B(n23707), .X(n5239) );
  nand_x1_sg U43975 ( .A(n23708), .B(n23709), .X(n5238) );
  nand_x1_sg U43976 ( .A(n23712), .B(n23713), .X(n5236) );
  nand_x1_sg U43977 ( .A(n23714), .B(n23715), .X(n5235) );
  nand_x1_sg U43978 ( .A(n23718), .B(n23719), .X(n5233) );
  nand_x1_sg U43979 ( .A(n23720), .B(n23721), .X(n5232) );
  nand_x1_sg U43980 ( .A(n23724), .B(n23725), .X(n5230) );
  nand_x1_sg U43981 ( .A(n26002), .B(n26003), .X(n4091) );
  nand_x1_sg U43982 ( .A(n26008), .B(n26009), .X(n4088) );
  nand_x1_sg U43983 ( .A(n26014), .B(n26015), .X(n4085) );
  nand_x1_sg U43984 ( .A(n26020), .B(n26021), .X(n4082) );
  nand_x1_sg U43985 ( .A(n26026), .B(n26027), .X(n4079) );
  nand_x1_sg U43986 ( .A(n26032), .B(n26033), .X(n4076) );
  nand_x1_sg U43987 ( .A(n26158), .B(n26159), .X(n4013) );
  nand_x1_sg U43988 ( .A(n26164), .B(n26165), .X(n4010) );
  nand_x1_sg U43989 ( .A(n26170), .B(n26171), .X(n4007) );
  nand_x1_sg U43990 ( .A(n26176), .B(n26177), .X(n4004) );
  nand_x1_sg U43991 ( .A(n26182), .B(n26183), .X(n4001) );
  nand_x1_sg U43992 ( .A(n26188), .B(n26189), .X(n3998) );
  nand_x1_sg U43993 ( .A(n25444), .B(n25445), .X(n4370) );
  nand_x1_sg U43994 ( .A(n25450), .B(n25451), .X(n4367) );
  nand_x1_sg U43995 ( .A(n25456), .B(n25457), .X(n4364) );
  nand_x1_sg U43996 ( .A(n25462), .B(n25463), .X(n4361) );
  nand_x1_sg U43997 ( .A(n25468), .B(n25469), .X(n4358) );
  nand_x1_sg U43998 ( .A(n25474), .B(n25475), .X(n4355) );
  nand_x1_sg U43999 ( .A(n25558), .B(n25559), .X(n4313) );
  nand_x1_sg U44000 ( .A(n25600), .B(n25601), .X(n4292) );
  nand_x1_sg U44001 ( .A(n25606), .B(n25607), .X(n4289) );
  nand_x1_sg U44002 ( .A(n25612), .B(n25613), .X(n4286) );
  nand_x1_sg U44003 ( .A(n25684), .B(n25685), .X(n4250) );
  nand_x1_sg U44004 ( .A(n25690), .B(n25691), .X(n4247) );
  nand_x1_sg U44005 ( .A(n25696), .B(n25697), .X(n4244) );
  nand_x1_sg U44006 ( .A(n25702), .B(n25703), .X(n4241) );
  nand_x1_sg U44007 ( .A(n25708), .B(n25709), .X(n4238) );
  nand_x1_sg U44008 ( .A(n25714), .B(n25715), .X(n4235) );
  nand_x1_sg U44009 ( .A(n25126), .B(n25127), .X(n4529) );
  nand_x1_sg U44010 ( .A(n25132), .B(n25133), .X(n4526) );
  nand_x1_sg U44011 ( .A(n25138), .B(n25139), .X(n4523) );
  nand_x1_sg U44012 ( .A(n25144), .B(n25145), .X(n4520) );
  nand_x1_sg U44013 ( .A(n25150), .B(n25151), .X(n4517) );
  nand_x1_sg U44014 ( .A(n25156), .B(n25157), .X(n4514) );
  nand_x1_sg U44015 ( .A(n25162), .B(n25163), .X(n4511) );
  nand_x1_sg U44016 ( .A(n24892), .B(n24893), .X(n4646) );
  nand_x1_sg U44017 ( .A(n24898), .B(n24899), .X(n4643) );
  nand_x1_sg U44018 ( .A(n24904), .B(n24905), .X(n4640) );
  nand_x1_sg U44019 ( .A(n24910), .B(n24911), .X(n4637) );
  nand_x1_sg U44020 ( .A(n24982), .B(n24983), .X(n4601) );
  nand_x1_sg U44021 ( .A(n24988), .B(n24989), .X(n4598) );
  nand_x1_sg U44022 ( .A(n24994), .B(n24995), .X(n4595) );
  nand_x1_sg U44023 ( .A(n24274), .B(n24275), .X(n4955) );
  nand_x1_sg U44024 ( .A(n24280), .B(n24281), .X(n4952) );
  nand_x1_sg U44025 ( .A(n24286), .B(n24287), .X(n4949) );
  nand_x1_sg U44026 ( .A(n24334), .B(n24335), .X(n4925) );
  nand_x1_sg U44027 ( .A(n24412), .B(n24413), .X(n4886) );
  nand_x1_sg U44028 ( .A(n24418), .B(n24419), .X(n4883) );
  nand_x1_sg U44029 ( .A(n24424), .B(n24425), .X(n4880) );
  nand_x1_sg U44030 ( .A(n24430), .B(n24431), .X(n4877) );
  nand_x1_sg U44031 ( .A(n24436), .B(n24437), .X(n4874) );
  nand_x1_sg U44032 ( .A(n24442), .B(n24443), .X(n4871) );
  nand_x1_sg U44033 ( .A(n24448), .B(n24449), .X(n4868) );
  nand_x1_sg U44034 ( .A(n24562), .B(n24563), .X(n4811) );
  nand_x1_sg U44035 ( .A(n24568), .B(n24569), .X(n4808) );
  nand_x1_sg U44036 ( .A(n24574), .B(n24575), .X(n4805) );
  nand_x1_sg U44037 ( .A(n24580), .B(n24581), .X(n4802) );
  nand_x1_sg U44038 ( .A(n24586), .B(n24587), .X(n4799) );
  nand_x1_sg U44039 ( .A(n24592), .B(n24593), .X(n4796) );
  nand_x1_sg U44040 ( .A(n23860), .B(n23861), .X(n5162) );
  nand_x1_sg U44041 ( .A(n23866), .B(n23867), .X(n5159) );
  nand_x1_sg U44042 ( .A(n23872), .B(n23873), .X(n5156) );
  nand_x1_sg U44043 ( .A(n23878), .B(n23879), .X(n5153) );
  nand_x1_sg U44044 ( .A(n23884), .B(n23885), .X(n5150) );
  nand_x1_sg U44045 ( .A(n23956), .B(n23957), .X(n5114) );
  nand_x1_sg U44046 ( .A(n23962), .B(n23963), .X(n5111) );
  nand_x1_sg U44047 ( .A(n23968), .B(n23969), .X(n5108) );
  nand_x1_sg U44048 ( .A(n23974), .B(n23975), .X(n5105) );
  nand_x1_sg U44049 ( .A(n24016), .B(n24017), .X(n5084) );
  nand_x1_sg U44050 ( .A(n23698), .B(n23699), .X(n5243) );
  nand_x1_sg U44051 ( .A(n23704), .B(n23705), .X(n5240) );
  nand_x1_sg U44052 ( .A(n23710), .B(n23711), .X(n5237) );
  nand_x1_sg U44053 ( .A(n23716), .B(n23717), .X(n5234) );
  nand_x1_sg U44054 ( .A(n23722), .B(n23723), .X(n5231) );
  nand_x1_sg U44055 ( .A(n25796), .B(n25797), .X(n4194) );
  nand_x1_sg U44056 ( .A(n25800), .B(n25801), .X(n4192) );
  nand_x1_sg U44057 ( .A(n25802), .B(n25803), .X(n4191) );
  nand_x1_sg U44058 ( .A(n25806), .B(n25807), .X(n4189) );
  nand_x1_sg U44059 ( .A(n25808), .B(n25809), .X(n4188) );
  nand_x1_sg U44060 ( .A(n25812), .B(n25813), .X(n4186) );
  nand_x1_sg U44061 ( .A(n25814), .B(n25815), .X(n4185) );
  nand_x1_sg U44062 ( .A(n25818), .B(n25819), .X(n4183) );
  nand_x1_sg U44063 ( .A(n25820), .B(n25821), .X(n4182) );
  nand_x1_sg U44064 ( .A(n25824), .B(n25825), .X(n4180) );
  nand_x1_sg U44065 ( .A(n25826), .B(n25827), .X(n4179) );
  nand_x1_sg U44066 ( .A(n25830), .B(n25831), .X(n4177) );
  nand_x1_sg U44067 ( .A(n25832), .B(n25833), .X(n4176) );
  nand_x1_sg U44068 ( .A(n25878), .B(n25879), .X(n4153) );
  nand_x1_sg U44069 ( .A(n25880), .B(n25881), .X(n4152) );
  nand_x1_sg U44070 ( .A(n25884), .B(n25885), .X(n4150) );
  nand_x1_sg U44071 ( .A(n25886), .B(n25887), .X(n4149) );
  nand_x1_sg U44072 ( .A(n25890), .B(n25891), .X(n4147) );
  nand_x1_sg U44073 ( .A(n25892), .B(n25893), .X(n4146) );
  nand_x1_sg U44074 ( .A(n25896), .B(n25897), .X(n4144) );
  nand_x1_sg U44075 ( .A(n25898), .B(n25899), .X(n4143) );
  nand_x1_sg U44076 ( .A(n25902), .B(n25903), .X(n4141) );
  nand_x1_sg U44077 ( .A(n25904), .B(n25905), .X(n4140) );
  nand_x1_sg U44078 ( .A(n25908), .B(n25909), .X(n4138) );
  nand_x1_sg U44079 ( .A(n25910), .B(n25911), .X(n4137) );
  nand_x1_sg U44080 ( .A(n25914), .B(n25915), .X(n4135) );
  nand_x1_sg U44081 ( .A(n25956), .B(n25957), .X(n4114) );
  nand_x1_sg U44082 ( .A(n25958), .B(n25959), .X(n4113) );
  nand_x1_sg U44083 ( .A(n25962), .B(n25963), .X(n4111) );
  nand_x1_sg U44084 ( .A(n25964), .B(n25965), .X(n4110) );
  nand_x1_sg U44085 ( .A(n25968), .B(n25969), .X(n4108) );
  nand_x1_sg U44086 ( .A(n25970), .B(n25971), .X(n4107) );
  nand_x1_sg U44087 ( .A(n25974), .B(n25975), .X(n4105) );
  nand_x1_sg U44088 ( .A(n25976), .B(n25977), .X(n4104) );
  nand_x1_sg U44089 ( .A(n25980), .B(n25981), .X(n4102) );
  nand_x1_sg U44090 ( .A(n25982), .B(n25983), .X(n4101) );
  nand_x1_sg U44091 ( .A(n25986), .B(n25987), .X(n4099) );
  nand_x1_sg U44092 ( .A(n25988), .B(n25989), .X(n4098) );
  nand_x1_sg U44093 ( .A(n25992), .B(n25993), .X(n4096) );
  nand_x1_sg U44094 ( .A(n25994), .B(n25995), .X(n4095) );
  nand_x1_sg U44095 ( .A(n26066), .B(n26067), .X(n4059) );
  nand_x1_sg U44096 ( .A(n26070), .B(n26071), .X(n4057) );
  nand_x1_sg U44097 ( .A(n26072), .B(n26073), .X(n4056) );
  nand_x1_sg U44098 ( .A(n26118), .B(n26119), .X(n4033) );
  nand_x1_sg U44099 ( .A(n26120), .B(n26121), .X(n4032) );
  nand_x1_sg U44100 ( .A(n26124), .B(n26125), .X(n4030) );
  nand_x1_sg U44101 ( .A(n26126), .B(n26127), .X(n4029) );
  nand_x1_sg U44102 ( .A(n25398), .B(n25399), .X(n4393) );
  nand_x1_sg U44103 ( .A(n25400), .B(n25401), .X(n4392) );
  nand_x1_sg U44104 ( .A(n25404), .B(n25405), .X(n4390) );
  nand_x1_sg U44105 ( .A(n25406), .B(n25407), .X(n4389) );
  nand_x1_sg U44106 ( .A(n25410), .B(n25411), .X(n4387) );
  nand_x1_sg U44107 ( .A(n25412), .B(n25413), .X(n4386) );
  nand_x1_sg U44108 ( .A(n25416), .B(n25417), .X(n4384) );
  nand_x1_sg U44109 ( .A(n25418), .B(n25419), .X(n4383) );
  nand_x1_sg U44110 ( .A(n25422), .B(n25423), .X(n4381) );
  nand_x1_sg U44111 ( .A(n25424), .B(n25425), .X(n4380) );
  nand_x1_sg U44112 ( .A(n25490), .B(n25491), .X(n4347) );
  nand_x1_sg U44113 ( .A(n25494), .B(n25495), .X(n4345) );
  nand_x1_sg U44114 ( .A(n25496), .B(n25497), .X(n4344) );
  nand_x1_sg U44115 ( .A(n25500), .B(n25501), .X(n4342) );
  nand_x1_sg U44116 ( .A(n25502), .B(n25503), .X(n4341) );
  nand_x1_sg U44117 ( .A(n25506), .B(n25507), .X(n4339) );
  nand_x1_sg U44118 ( .A(n25508), .B(n25509), .X(n4338) );
  nand_x1_sg U44119 ( .A(n25512), .B(n25513), .X(n4336) );
  nand_x1_sg U44120 ( .A(n25514), .B(n25515), .X(n4335) );
  nand_x1_sg U44121 ( .A(n25518), .B(n25519), .X(n4333) );
  nand_x1_sg U44122 ( .A(n25640), .B(n25641), .X(n4272) );
  nand_x1_sg U44123 ( .A(n25644), .B(n25645), .X(n4270) );
  nand_x1_sg U44124 ( .A(n25646), .B(n25647), .X(n4269) );
  nand_x1_sg U44125 ( .A(n25650), .B(n25651), .X(n4267) );
  nand_x1_sg U44126 ( .A(n25652), .B(n25653), .X(n4266) );
  nand_x1_sg U44127 ( .A(n25656), .B(n25657), .X(n4264) );
  nand_x1_sg U44128 ( .A(n25658), .B(n25659), .X(n4263) );
  nand_x1_sg U44129 ( .A(n25662), .B(n25663), .X(n4261) );
  nand_x1_sg U44130 ( .A(n25664), .B(n25665), .X(n4260) );
  nand_x1_sg U44131 ( .A(n25668), .B(n25669), .X(n4258) );
  nand_x1_sg U44132 ( .A(n25670), .B(n25671), .X(n4257) );
  nand_x1_sg U44133 ( .A(n25674), .B(n25675), .X(n4255) );
  nand_x1_sg U44134 ( .A(n25676), .B(n25677), .X(n4254) );
  nand_x1_sg U44135 ( .A(n25746), .B(n25747), .X(n4219) );
  nand_x1_sg U44136 ( .A(n25748), .B(n25749), .X(n4218) );
  nand_x1_sg U44137 ( .A(n25752), .B(n25753), .X(n4216) );
  nand_x1_sg U44138 ( .A(n25754), .B(n25755), .X(n4215) );
  nand_x1_sg U44139 ( .A(n25086), .B(n25087), .X(n4549) );
  nand_x1_sg U44140 ( .A(n25088), .B(n25089), .X(n4548) );
  nand_x1_sg U44141 ( .A(n25092), .B(n25093), .X(n4546) );
  nand_x1_sg U44142 ( .A(n25094), .B(n25095), .X(n4545) );
  nand_x1_sg U44143 ( .A(n25098), .B(n25099), .X(n4543) );
  nand_x1_sg U44144 ( .A(n25100), .B(n25101), .X(n4542) );
  nand_x1_sg U44145 ( .A(n25104), .B(n25105), .X(n4540) );
  nand_x1_sg U44146 ( .A(n25170), .B(n25171), .X(n4507) );
  nand_x1_sg U44147 ( .A(n25172), .B(n25173), .X(n4506) );
  nand_x1_sg U44148 ( .A(n25176), .B(n25177), .X(n4504) );
  nand_x1_sg U44149 ( .A(n25178), .B(n25179), .X(n4503) );
  nand_x1_sg U44150 ( .A(n25182), .B(n25183), .X(n4501) );
  nand_x1_sg U44151 ( .A(n25184), .B(n25185), .X(n4500) );
  nand_x1_sg U44152 ( .A(n25188), .B(n25189), .X(n4498) );
  nand_x1_sg U44153 ( .A(n25190), .B(n25191), .X(n4497) );
  nand_x1_sg U44154 ( .A(n25194), .B(n25195), .X(n4495) );
  nand_x1_sg U44155 ( .A(n25196), .B(n25197), .X(n4494) );
  nand_x1_sg U44156 ( .A(n25200), .B(n25201), .X(n4492) );
  nand_x1_sg U44157 ( .A(n25202), .B(n25203), .X(n4491) );
  nand_x1_sg U44158 ( .A(n25244), .B(n25245), .X(n4470) );
  nand_x1_sg U44159 ( .A(n25248), .B(n25249), .X(n4468) );
  nand_x1_sg U44160 ( .A(n25250), .B(n25251), .X(n4467) );
  nand_x1_sg U44161 ( .A(n25254), .B(n25255), .X(n4465) );
  nand_x1_sg U44162 ( .A(n25256), .B(n25257), .X(n4464) );
  nand_x1_sg U44163 ( .A(n25260), .B(n25261), .X(n4462) );
  nand_x1_sg U44164 ( .A(n25262), .B(n25263), .X(n4461) );
  nand_x1_sg U44165 ( .A(n25266), .B(n25267), .X(n4459) );
  nand_x1_sg U44166 ( .A(n25268), .B(n25269), .X(n4458) );
  nand_x1_sg U44167 ( .A(n25272), .B(n25273), .X(n4456) );
  nand_x1_sg U44168 ( .A(n25274), .B(n25275), .X(n4455) );
  nand_x1_sg U44169 ( .A(n25278), .B(n25279), .X(n4453) );
  nand_x1_sg U44170 ( .A(n25280), .B(n25281), .X(n4452) );
  nand_x1_sg U44171 ( .A(n25326), .B(n25327), .X(n4429) );
  nand_x1_sg U44172 ( .A(n25328), .B(n25329), .X(n4428) );
  nand_x1_sg U44173 ( .A(n25332), .B(n25333), .X(n4426) );
  nand_x1_sg U44174 ( .A(n25334), .B(n25335), .X(n4425) );
  nand_x1_sg U44175 ( .A(n25338), .B(n25339), .X(n4423) );
  nand_x1_sg U44176 ( .A(n25340), .B(n25341), .X(n4422) );
  nand_x1_sg U44177 ( .A(n25344), .B(n25345), .X(n4420) );
  nand_x1_sg U44178 ( .A(n25346), .B(n25347), .X(n4419) );
  nand_x1_sg U44179 ( .A(n25350), .B(n25351), .X(n4417) );
  nand_x1_sg U44180 ( .A(n25352), .B(n25353), .X(n4416) );
  nand_x1_sg U44181 ( .A(n25356), .B(n25357), .X(n4414) );
  nand_x1_sg U44182 ( .A(n24602), .B(n24603), .X(n4791) );
  nand_x1_sg U44183 ( .A(n24606), .B(n24607), .X(n4789) );
  nand_x1_sg U44184 ( .A(n24608), .B(n24609), .X(n4788) );
  nand_x1_sg U44185 ( .A(n24612), .B(n24613), .X(n4786) );
  nand_x1_sg U44186 ( .A(n24614), .B(n24615), .X(n4785) );
  nand_x1_sg U44187 ( .A(n24618), .B(n24619), .X(n4783) );
  nand_x1_sg U44188 ( .A(n24620), .B(n24621), .X(n4782) );
  nand_x1_sg U44189 ( .A(n24624), .B(n24625), .X(n4780) );
  nand_x1_sg U44190 ( .A(n24626), .B(n24627), .X(n4779) );
  nand_x1_sg U44191 ( .A(n24630), .B(n24631), .X(n4777) );
  nand_x1_sg U44192 ( .A(n24632), .B(n24633), .X(n4776) );
  nand_x1_sg U44193 ( .A(n24636), .B(n24637), .X(n4774) );
  nand_x1_sg U44194 ( .A(n24638), .B(n24639), .X(n4773) );
  nand_x1_sg U44195 ( .A(n24642), .B(n24643), .X(n4771) );
  nand_x1_sg U44196 ( .A(n24644), .B(n24645), .X(n4770) );
  nand_x1_sg U44197 ( .A(n24690), .B(n24691), .X(n4747) );
  nand_x1_sg U44198 ( .A(n24692), .B(n24693), .X(n4746) );
  nand_x1_sg U44199 ( .A(n24696), .B(n24697), .X(n4744) );
  nand_x1_sg U44200 ( .A(n24698), .B(n24699), .X(n4743) );
  nand_x1_sg U44201 ( .A(n24702), .B(n24703), .X(n4741) );
  nand_x1_sg U44202 ( .A(n24704), .B(n24705), .X(n4740) );
  nand_x1_sg U44203 ( .A(n24708), .B(n24709), .X(n4738) );
  nand_x1_sg U44204 ( .A(n24710), .B(n24711), .X(n4737) );
  nand_x1_sg U44205 ( .A(n24714), .B(n24715), .X(n4735) );
  nand_x1_sg U44206 ( .A(n24716), .B(n24717), .X(n4734) );
  nand_x1_sg U44207 ( .A(n24720), .B(n24721), .X(n4732) );
  nand_x1_sg U44208 ( .A(n24722), .B(n24723), .X(n4731) );
  nand_x1_sg U44209 ( .A(n24726), .B(n24727), .X(n4729) );
  nand_x1_sg U44210 ( .A(n24768), .B(n24769), .X(n4708) );
  nand_x1_sg U44211 ( .A(n24770), .B(n24771), .X(n4707) );
  nand_x1_sg U44212 ( .A(n24774), .B(n24775), .X(n4705) );
  nand_x1_sg U44213 ( .A(n24776), .B(n24777), .X(n4704) );
  nand_x1_sg U44214 ( .A(n24780), .B(n24781), .X(n4702) );
  nand_x1_sg U44215 ( .A(n24782), .B(n24783), .X(n4701) );
  nand_x1_sg U44216 ( .A(n24786), .B(n24787), .X(n4699) );
  nand_x1_sg U44217 ( .A(n24788), .B(n24789), .X(n4698) );
  nand_x1_sg U44218 ( .A(n24792), .B(n24793), .X(n4696) );
  nand_x1_sg U44219 ( .A(n24794), .B(n24795), .X(n4695) );
  nand_x1_sg U44220 ( .A(n24798), .B(n24799), .X(n4693) );
  nand_x1_sg U44221 ( .A(n24800), .B(n24801), .X(n4692) );
  nand_x1_sg U44222 ( .A(n24804), .B(n24805), .X(n4690) );
  nand_x1_sg U44223 ( .A(n24806), .B(n24807), .X(n4689) );
  nand_x1_sg U44224 ( .A(n24848), .B(n24849), .X(n4668) );
  nand_x1_sg U44225 ( .A(n24930), .B(n24931), .X(n4627) );
  nand_x1_sg U44226 ( .A(n24932), .B(n24933), .X(n4626) );
  nand_x1_sg U44227 ( .A(n24936), .B(n24937), .X(n4624) );
  nand_x1_sg U44228 ( .A(n24938), .B(n24939), .X(n4623) );
  nand_x1_sg U44229 ( .A(n24942), .B(n24943), .X(n4621) );
  nand_x1_sg U44230 ( .A(n24944), .B(n24945), .X(n4620) );
  nand_x1_sg U44231 ( .A(n24948), .B(n24949), .X(n4618) );
  nand_x1_sg U44232 ( .A(n24950), .B(n24951), .X(n4617) );
  nand_x1_sg U44233 ( .A(n24954), .B(n24955), .X(n4615) );
  nand_x1_sg U44234 ( .A(n24956), .B(n24957), .X(n4614) );
  nand_x1_sg U44235 ( .A(n24204), .B(n24205), .X(n4990) );
  nand_x1_sg U44236 ( .A(n24206), .B(n24207), .X(n4989) );
  nand_x1_sg U44237 ( .A(n24210), .B(n24211), .X(n4987) );
  nand_x1_sg U44238 ( .A(n24212), .B(n24213), .X(n4986) );
  nand_x1_sg U44239 ( .A(n24216), .B(n24217), .X(n4984) );
  nand_x1_sg U44240 ( .A(n24218), .B(n24219), .X(n4983) );
  nand_x1_sg U44241 ( .A(n24222), .B(n24223), .X(n4981) );
  nand_x1_sg U44242 ( .A(n24224), .B(n24225), .X(n4980) );
  nand_x1_sg U44243 ( .A(n24228), .B(n24229), .X(n4978) );
  nand_x1_sg U44244 ( .A(n24230), .B(n24231), .X(n4977) );
  nand_x1_sg U44245 ( .A(n24234), .B(n24235), .X(n4975) );
  nand_x1_sg U44246 ( .A(n24236), .B(n24237), .X(n4974) );
  nand_x1_sg U44247 ( .A(n24240), .B(n24241), .X(n4972) );
  nand_x1_sg U44248 ( .A(n24242), .B(n24243), .X(n4971) );
  nand_x1_sg U44249 ( .A(n24246), .B(n24247), .X(n4969) );
  nand_x1_sg U44250 ( .A(n24248), .B(n24249), .X(n4968) );
  nand_x1_sg U44251 ( .A(n24372), .B(n24373), .X(n4906) );
  nand_x1_sg U44252 ( .A(n24374), .B(n24375), .X(n4905) );
  nand_x1_sg U44253 ( .A(n24378), .B(n24379), .X(n4903) );
  nand_x1_sg U44254 ( .A(n24380), .B(n24381), .X(n4902) );
  nand_x1_sg U44255 ( .A(n24384), .B(n24385), .X(n4900) );
  nand_x1_sg U44256 ( .A(n24386), .B(n24387), .X(n4899) );
  nand_x1_sg U44257 ( .A(n24390), .B(n24391), .X(n4897) );
  nand_x1_sg U44258 ( .A(n24392), .B(n24393), .X(n4896) );
  nand_x1_sg U44259 ( .A(n24396), .B(n24397), .X(n4894) );
  nand_x1_sg U44260 ( .A(n24398), .B(n24399), .X(n4893) );
  nand_x1_sg U44261 ( .A(n24468), .B(n24469), .X(n4858) );
  nand_x1_sg U44262 ( .A(n24470), .B(n24471), .X(n4857) );
  nand_x1_sg U44263 ( .A(n24474), .B(n24475), .X(n4855) );
  nand_x1_sg U44264 ( .A(n24476), .B(n24477), .X(n4854) );
  nand_x1_sg U44265 ( .A(n24480), .B(n24481), .X(n4852) );
  nand_x1_sg U44266 ( .A(n24482), .B(n24483), .X(n4851) );
  nand_x1_sg U44267 ( .A(n24486), .B(n24487), .X(n4849) );
  nand_x1_sg U44268 ( .A(n24488), .B(n24489), .X(n4848) );
  nand_x1_sg U44269 ( .A(n23808), .B(n23809), .X(n5188) );
  nand_x1_sg U44270 ( .A(n23810), .B(n23811), .X(n5187) );
  nand_x1_sg U44271 ( .A(n23814), .B(n23815), .X(n5185) );
  nand_x1_sg U44272 ( .A(n23816), .B(n23817), .X(n5184) );
  nand_x1_sg U44273 ( .A(n23820), .B(n23821), .X(n5182) );
  nand_x1_sg U44274 ( .A(n23822), .B(n23823), .X(n5181) );
  nand_x1_sg U44275 ( .A(n23898), .B(n23899), .X(n5143) );
  nand_x1_sg U44276 ( .A(n23900), .B(n23901), .X(n5142) );
  nand_x1_sg U44277 ( .A(n23904), .B(n23905), .X(n5140) );
  nand_x1_sg U44278 ( .A(n23906), .B(n23907), .X(n5139) );
  nand_x1_sg U44279 ( .A(n23910), .B(n23911), .X(n5137) );
  nand_x1_sg U44280 ( .A(n23912), .B(n23913), .X(n5136) );
  nand_x1_sg U44281 ( .A(n23916), .B(n23917), .X(n5134) );
  nand_x1_sg U44282 ( .A(n23918), .B(n23919), .X(n5133) );
  nand_x1_sg U44283 ( .A(n23922), .B(n23923), .X(n5131) );
  nand_x1_sg U44284 ( .A(n23924), .B(n23925), .X(n5130) );
  nand_x1_sg U44285 ( .A(n23928), .B(n23929), .X(n5128) );
  nand_x1_sg U44286 ( .A(n23930), .B(n23931), .X(n5127) );
  nand_x1_sg U44287 ( .A(n23934), .B(n23935), .X(n5125) );
  nand_x1_sg U44288 ( .A(n24056), .B(n24057), .X(n5064) );
  nand_x1_sg U44289 ( .A(n24060), .B(n24061), .X(n5062) );
  nand_x1_sg U44290 ( .A(n24062), .B(n24063), .X(n5061) );
  nand_x1_sg U44291 ( .A(n24066), .B(n24067), .X(n5059) );
  nand_x1_sg U44292 ( .A(n24068), .B(n24069), .X(n5058) );
  nand_x1_sg U44293 ( .A(n24072), .B(n24073), .X(n5056) );
  nand_x1_sg U44294 ( .A(n24074), .B(n24075), .X(n5055) );
  nand_x1_sg U44295 ( .A(n24078), .B(n24079), .X(n5053) );
  nand_x1_sg U44296 ( .A(n24080), .B(n24081), .X(n5052) );
  nand_x1_sg U44297 ( .A(n24084), .B(n24085), .X(n5050) );
  nand_x1_sg U44298 ( .A(n24086), .B(n24087), .X(n5049) );
  nand_x1_sg U44299 ( .A(n24090), .B(n24091), .X(n5047) );
  nand_x1_sg U44300 ( .A(n24092), .B(n24093), .X(n5046) );
  nand_x1_sg U44301 ( .A(n24138), .B(n24139), .X(n5023) );
  nand_x1_sg U44302 ( .A(n24140), .B(n24141), .X(n5022) );
  nand_x1_sg U44303 ( .A(n24144), .B(n24145), .X(n5020) );
  nand_x1_sg U44304 ( .A(n24146), .B(n24147), .X(n5019) );
  nand_x1_sg U44305 ( .A(n24150), .B(n24151), .X(n5017) );
  nand_x1_sg U44306 ( .A(n24152), .B(n24153), .X(n5016) );
  nand_x1_sg U44307 ( .A(n24156), .B(n24157), .X(n5014) );
  nand_x1_sg U44308 ( .A(n24158), .B(n24159), .X(n5013) );
  nand_x1_sg U44309 ( .A(n24162), .B(n24163), .X(n5011) );
  nand_x1_sg U44310 ( .A(n23633), .B(n23634), .X(n5275) );
  nand_x1_sg U44311 ( .A(n23636), .B(n23637), .X(n5274) );
  nand_x1_sg U44312 ( .A(n23640), .B(n23641), .X(n5272) );
  nand_x1_sg U44313 ( .A(n23642), .B(n23643), .X(n5271) );
  nand_x1_sg U44314 ( .A(n23646), .B(n23647), .X(n5269) );
  nand_x1_sg U44315 ( .A(n23648), .B(n23649), .X(n5268) );
  nand_x1_sg U44316 ( .A(n23652), .B(n23653), .X(n5266) );
  nand_x1_sg U44317 ( .A(n23654), .B(n23655), .X(n5265) );
  nand_x1_sg U44318 ( .A(n23658), .B(n23659), .X(n5263) );
  nand_x1_sg U44319 ( .A(n23660), .B(n23661), .X(n5262) );
  nand_x1_sg U44320 ( .A(n23664), .B(n23665), .X(n5260) );
  nand_x1_sg U44321 ( .A(n23666), .B(n23667), .X(n5259) );
  nand_x1_sg U44322 ( .A(n23670), .B(n23671), .X(n5257) );
  nand_x1_sg U44323 ( .A(n23672), .B(n23673), .X(n5256) );
  nand_x1_sg U44324 ( .A(n23676), .B(n23677), .X(n5254) );
  nand_x1_sg U44325 ( .A(n23678), .B(n23679), .X(n5253) );
  nand_x1_sg U44326 ( .A(n23682), .B(n23683), .X(n5251) );
  nand_x1_sg U44327 ( .A(n23684), .B(n23685), .X(n5250) );
  nand_x1_sg U44328 ( .A(n23762), .B(n23763), .X(n5211) );
  nand_x1_sg U44329 ( .A(n25798), .B(n25799), .X(n4193) );
  nand_x1_sg U44330 ( .A(n25804), .B(n25805), .X(n4190) );
  nand_x1_sg U44331 ( .A(n25810), .B(n25811), .X(n4187) );
  nand_x1_sg U44332 ( .A(n25816), .B(n25817), .X(n4184) );
  nand_x1_sg U44333 ( .A(n25822), .B(n25823), .X(n4181) );
  nand_x1_sg U44334 ( .A(n25828), .B(n25829), .X(n4178) );
  nand_x1_sg U44335 ( .A(n25834), .B(n25835), .X(n4175) );
  nand_x1_sg U44336 ( .A(n25876), .B(n25877), .X(n4154) );
  nand_x1_sg U44337 ( .A(n25882), .B(n25883), .X(n4151) );
  nand_x1_sg U44338 ( .A(n25888), .B(n25889), .X(n4148) );
  nand_x1_sg U44339 ( .A(n25894), .B(n25895), .X(n4145) );
  nand_x1_sg U44340 ( .A(n25900), .B(n25901), .X(n4142) );
  nand_x1_sg U44341 ( .A(n25906), .B(n25907), .X(n4139) );
  nand_x1_sg U44342 ( .A(n25912), .B(n25913), .X(n4136) );
  nand_x1_sg U44343 ( .A(n25960), .B(n25961), .X(n4112) );
  nand_x1_sg U44344 ( .A(n25966), .B(n25967), .X(n4109) );
  nand_x1_sg U44345 ( .A(n25972), .B(n25973), .X(n4106) );
  nand_x1_sg U44346 ( .A(n25978), .B(n25979), .X(n4103) );
  nand_x1_sg U44347 ( .A(n25984), .B(n25985), .X(n4100) );
  nand_x1_sg U44348 ( .A(n25990), .B(n25991), .X(n4097) );
  nand_x1_sg U44349 ( .A(n26068), .B(n26069), .X(n4058) );
  nand_x1_sg U44350 ( .A(n26074), .B(n26075), .X(n4055) );
  nand_x1_sg U44351 ( .A(n26116), .B(n26117), .X(n4034) );
  nand_x1_sg U44352 ( .A(n26122), .B(n26123), .X(n4031) );
  nand_x1_sg U44353 ( .A(n26128), .B(n26129), .X(n4028) );
  nand_x1_sg U44354 ( .A(n25402), .B(n25403), .X(n4391) );
  nand_x1_sg U44355 ( .A(n25408), .B(n25409), .X(n4388) );
  nand_x1_sg U44356 ( .A(n25414), .B(n25415), .X(n4385) );
  nand_x1_sg U44357 ( .A(n25420), .B(n25421), .X(n4382) );
  nand_x1_sg U44358 ( .A(n25492), .B(n25493), .X(n4346) );
  nand_x1_sg U44359 ( .A(n25498), .B(n25499), .X(n4343) );
  nand_x1_sg U44360 ( .A(n25504), .B(n25505), .X(n4340) );
  nand_x1_sg U44361 ( .A(n25510), .B(n25511), .X(n4337) );
  nand_x1_sg U44362 ( .A(n25516), .B(n25517), .X(n4334) );
  nand_x1_sg U44363 ( .A(n25642), .B(n25643), .X(n4271) );
  nand_x1_sg U44364 ( .A(n25648), .B(n25649), .X(n4268) );
  nand_x1_sg U44365 ( .A(n25654), .B(n25655), .X(n4265) );
  nand_x1_sg U44366 ( .A(n25660), .B(n25661), .X(n4262) );
  nand_x1_sg U44367 ( .A(n25666), .B(n25667), .X(n4259) );
  nand_x1_sg U44368 ( .A(n25672), .B(n25673), .X(n4256) );
  nand_x1_sg U44369 ( .A(n25678), .B(n25679), .X(n4253) );
  nand_x1_sg U44370 ( .A(n25750), .B(n25751), .X(n4217) );
  nand_x1_sg U44371 ( .A(n25042), .B(n25043), .X(n4571) );
  nand_x1_sg U44372 ( .A(n25084), .B(n25085), .X(n4550) );
  nand_x1_sg U44373 ( .A(n25090), .B(n25091), .X(n4547) );
  nand_x1_sg U44374 ( .A(n25096), .B(n25097), .X(n4544) );
  nand_x1_sg U44375 ( .A(n25102), .B(n25103), .X(n4541) );
  nand_x1_sg U44376 ( .A(n25174), .B(n25175), .X(n4505) );
  nand_x1_sg U44377 ( .A(n25180), .B(n25181), .X(n4502) );
  nand_x1_sg U44378 ( .A(n25186), .B(n25187), .X(n4499) );
  nand_x1_sg U44379 ( .A(n25192), .B(n25193), .X(n4496) );
  nand_x1_sg U44380 ( .A(n25198), .B(n25199), .X(n4493) );
  nand_x1_sg U44381 ( .A(n25246), .B(n25247), .X(n4469) );
  nand_x1_sg U44382 ( .A(n25252), .B(n25253), .X(n4466) );
  nand_x1_sg U44383 ( .A(n25258), .B(n25259), .X(n4463) );
  nand_x1_sg U44384 ( .A(n25264), .B(n25265), .X(n4460) );
  nand_x1_sg U44385 ( .A(n25270), .B(n25271), .X(n4457) );
  nand_x1_sg U44386 ( .A(n25276), .B(n25277), .X(n4454) );
  nand_x1_sg U44387 ( .A(n25282), .B(n25283), .X(n4451) );
  nand_x1_sg U44388 ( .A(n25324), .B(n25325), .X(n4430) );
  nand_x1_sg U44389 ( .A(n25330), .B(n25331), .X(n4427) );
  nand_x1_sg U44390 ( .A(n25336), .B(n25337), .X(n4424) );
  nand_x1_sg U44391 ( .A(n25342), .B(n25343), .X(n4421) );
  nand_x1_sg U44392 ( .A(n25348), .B(n25349), .X(n4418) );
  nand_x1_sg U44393 ( .A(n25354), .B(n25355), .X(n4415) );
  nand_x1_sg U44394 ( .A(n24604), .B(n24605), .X(n4790) );
  nand_x1_sg U44395 ( .A(n24610), .B(n24611), .X(n4787) );
  nand_x1_sg U44396 ( .A(n24616), .B(n24617), .X(n4784) );
  nand_x1_sg U44397 ( .A(n24622), .B(n24623), .X(n4781) );
  nand_x1_sg U44398 ( .A(n24628), .B(n24629), .X(n4778) );
  nand_x1_sg U44399 ( .A(n24634), .B(n24635), .X(n4775) );
  nand_x1_sg U44400 ( .A(n24640), .B(n24641), .X(n4772) );
  nand_x1_sg U44401 ( .A(n24646), .B(n24647), .X(n4769) );
  nand_x1_sg U44402 ( .A(n24688), .B(n24689), .X(n4748) );
  nand_x1_sg U44403 ( .A(n24694), .B(n24695), .X(n4745) );
  nand_x1_sg U44404 ( .A(n24700), .B(n24701), .X(n4742) );
  nand_x1_sg U44405 ( .A(n24706), .B(n24707), .X(n4739) );
  nand_x1_sg U44406 ( .A(n24712), .B(n24713), .X(n4736) );
  nand_x1_sg U44407 ( .A(n24718), .B(n24719), .X(n4733) );
  nand_x1_sg U44408 ( .A(n24724), .B(n24725), .X(n4730) );
  nand_x1_sg U44409 ( .A(n24772), .B(n24773), .X(n4706) );
  nand_x1_sg U44410 ( .A(n24778), .B(n24779), .X(n4703) );
  nand_x1_sg U44411 ( .A(n24784), .B(n24785), .X(n4700) );
  nand_x1_sg U44412 ( .A(n24790), .B(n24791), .X(n4697) );
  nand_x1_sg U44413 ( .A(n24796), .B(n24797), .X(n4694) );
  nand_x1_sg U44414 ( .A(n24802), .B(n24803), .X(n4691) );
  nand_x1_sg U44415 ( .A(n24928), .B(n24929), .X(n4628) );
  nand_x1_sg U44416 ( .A(n24934), .B(n24935), .X(n4625) );
  nand_x1_sg U44417 ( .A(n24940), .B(n24941), .X(n4622) );
  nand_x1_sg U44418 ( .A(n24946), .B(n24947), .X(n4619) );
  nand_x1_sg U44419 ( .A(n24952), .B(n24953), .X(n4616) );
  nand_x1_sg U44420 ( .A(n24958), .B(n24959), .X(n4613) );
  nand_x1_sg U44421 ( .A(n24208), .B(n24209), .X(n4988) );
  nand_x1_sg U44422 ( .A(n24214), .B(n24215), .X(n4985) );
  nand_x1_sg U44423 ( .A(n24220), .B(n24221), .X(n4982) );
  nand_x1_sg U44424 ( .A(n24226), .B(n24227), .X(n4979) );
  nand_x1_sg U44425 ( .A(n24232), .B(n24233), .X(n4976) );
  nand_x1_sg U44426 ( .A(n24238), .B(n24239), .X(n4973) );
  nand_x1_sg U44427 ( .A(n24244), .B(n24245), .X(n4970) );
  nand_x1_sg U44428 ( .A(n24250), .B(n24251), .X(n4967) );
  nand_x1_sg U44429 ( .A(n24376), .B(n24377), .X(n4904) );
  nand_x1_sg U44430 ( .A(n24382), .B(n24383), .X(n4901) );
  nand_x1_sg U44431 ( .A(n24388), .B(n24389), .X(n4898) );
  nand_x1_sg U44432 ( .A(n24394), .B(n24395), .X(n4895) );
  nand_x1_sg U44433 ( .A(n24400), .B(n24401), .X(n4892) );
  nand_x1_sg U44434 ( .A(n24466), .B(n24467), .X(n4859) );
  nand_x1_sg U44435 ( .A(n24472), .B(n24473), .X(n4856) );
  nand_x1_sg U44436 ( .A(n24478), .B(n24479), .X(n4853) );
  nand_x1_sg U44437 ( .A(n24484), .B(n24485), .X(n4850) );
  nand_x1_sg U44438 ( .A(n24490), .B(n24491), .X(n4847) );
  nand_x1_sg U44439 ( .A(n23806), .B(n23807), .X(n5189) );
  nand_x1_sg U44440 ( .A(n23812), .B(n23813), .X(n5186) );
  nand_x1_sg U44441 ( .A(n23818), .B(n23819), .X(n5183) );
  nand_x1_sg U44442 ( .A(n23824), .B(n23825), .X(n5180) );
  nand_x1_sg U44443 ( .A(n23896), .B(n23897), .X(n5144) );
  nand_x1_sg U44444 ( .A(n23902), .B(n23903), .X(n5141) );
  nand_x1_sg U44445 ( .A(n23908), .B(n23909), .X(n5138) );
  nand_x1_sg U44446 ( .A(n23914), .B(n23915), .X(n5135) );
  nand_x1_sg U44447 ( .A(n23920), .B(n23921), .X(n5132) );
  nand_x1_sg U44448 ( .A(n23926), .B(n23927), .X(n5129) );
  nand_x1_sg U44449 ( .A(n23932), .B(n23933), .X(n5126) );
  nand_x1_sg U44450 ( .A(n24058), .B(n24059), .X(n5063) );
  nand_x1_sg U44451 ( .A(n24064), .B(n24065), .X(n5060) );
  nand_x1_sg U44452 ( .A(n24070), .B(n24071), .X(n5057) );
  nand_x1_sg U44453 ( .A(n24076), .B(n24077), .X(n5054) );
  nand_x1_sg U44454 ( .A(n24082), .B(n24083), .X(n5051) );
  nand_x1_sg U44455 ( .A(n24088), .B(n24089), .X(n5048) );
  nand_x1_sg U44456 ( .A(n24094), .B(n24095), .X(n5045) );
  nand_x1_sg U44457 ( .A(n24136), .B(n24137), .X(n5024) );
  nand_x1_sg U44458 ( .A(n24142), .B(n24143), .X(n5021) );
  nand_x1_sg U44459 ( .A(n24148), .B(n24149), .X(n5018) );
  nand_x1_sg U44460 ( .A(n24154), .B(n24155), .X(n5015) );
  nand_x1_sg U44461 ( .A(n24160), .B(n24161), .X(n5012) );
  nand_x1_sg U44462 ( .A(n23638), .B(n23639), .X(n5273) );
  nand_x1_sg U44463 ( .A(n23644), .B(n23645), .X(n5270) );
  nand_x1_sg U44464 ( .A(n23650), .B(n23651), .X(n5267) );
  nand_x1_sg U44465 ( .A(n23656), .B(n23657), .X(n5264) );
  nand_x1_sg U44466 ( .A(n23662), .B(n23663), .X(n5261) );
  nand_x1_sg U44467 ( .A(n23668), .B(n23669), .X(n5258) );
  nand_x1_sg U44468 ( .A(n23674), .B(n23675), .X(n5255) );
  nand_x1_sg U44469 ( .A(n23680), .B(n23681), .X(n5252) );
  nand_x1_sg U44470 ( .A(n23764), .B(n23765), .X(n5210) );
  inv_x1_sg U44471 ( .A(n15329), .X(n42370) );
  nand_x1_sg U44472 ( .A(n29635), .B(n29636), .X(\filter_0/n8257 ) );
  nand_x1_sg U44473 ( .A(n29637), .B(n29638), .X(\filter_0/n8256 ) );
  nand_x1_sg U44474 ( .A(n29639), .B(n29640), .X(\filter_0/n8255 ) );
  nand_x1_sg U44475 ( .A(n29641), .B(n29642), .X(\filter_0/n8254 ) );
  nand_x1_sg U44476 ( .A(n29643), .B(n29644), .X(\filter_0/n8253 ) );
  nand_x1_sg U44477 ( .A(n29645), .B(n29646), .X(\filter_0/n8252 ) );
  nand_x1_sg U44478 ( .A(n29647), .B(n29648), .X(\filter_0/n8251 ) );
  nand_x1_sg U44479 ( .A(n29649), .B(n29650), .X(\filter_0/n8250 ) );
  nand_x1_sg U44480 ( .A(n29651), .B(n29652), .X(\filter_0/n8249 ) );
  nand_x1_sg U44481 ( .A(n29653), .B(n29654), .X(\filter_0/n8248 ) );
  nand_x1_sg U44482 ( .A(n29655), .B(n29656), .X(\filter_0/n8247 ) );
  nand_x1_sg U44483 ( .A(n29657), .B(n29658), .X(\filter_0/n8246 ) );
  nand_x1_sg U44484 ( .A(n29659), .B(n29660), .X(\filter_0/n8245 ) );
  nand_x1_sg U44485 ( .A(n29661), .B(n29662), .X(\filter_0/n8244 ) );
  nand_x1_sg U44486 ( .A(n29119), .B(n29120), .X(\filter_0/n8497 ) );
  nand_x1_sg U44487 ( .A(n29121), .B(n29122), .X(\filter_0/n8496 ) );
  nand_x1_sg U44488 ( .A(n29123), .B(n29124), .X(\filter_0/n8495 ) );
  nand_x1_sg U44489 ( .A(n29125), .B(n29126), .X(\filter_0/n8494 ) );
  nand_x1_sg U44490 ( .A(n29127), .B(n29128), .X(\filter_0/n8493 ) );
  nand_x1_sg U44491 ( .A(n29129), .B(n29130), .X(\filter_0/n8492 ) );
  nand_x1_sg U44492 ( .A(n29131), .B(n29132), .X(\filter_0/n8491 ) );
  nand_x1_sg U44493 ( .A(n29133), .B(n29134), .X(\filter_0/n8490 ) );
  nand_x1_sg U44494 ( .A(n29135), .B(n29136), .X(\filter_0/n8489 ) );
  nand_x1_sg U44495 ( .A(n29137), .B(n29138), .X(\filter_0/n8488 ) );
  nand_x1_sg U44496 ( .A(n29139), .B(n29140), .X(\filter_0/n8487 ) );
  nand_x1_sg U44497 ( .A(n29141), .B(n29142), .X(\filter_0/n8486 ) );
  nand_x1_sg U44498 ( .A(n29143), .B(n29144), .X(\filter_0/n8485 ) );
  nand_x1_sg U44499 ( .A(n29145), .B(n29146), .X(\filter_0/n8484 ) );
  nand_x1_sg U44500 ( .A(n28936), .B(n28937), .X(\filter_0/n8581 ) );
  nand_x1_sg U44501 ( .A(n28938), .B(n28939), .X(\filter_0/n8580 ) );
  nand_x1_sg U44502 ( .A(n28940), .B(n28941), .X(\filter_0/n8579 ) );
  nand_x1_sg U44503 ( .A(n28942), .B(n28943), .X(\filter_0/n8578 ) );
  nand_x1_sg U44504 ( .A(n28944), .B(n28945), .X(\filter_0/n8577 ) );
  nand_x1_sg U44505 ( .A(n28946), .B(n28947), .X(\filter_0/n8576 ) );
  nand_x1_sg U44506 ( .A(n28948), .B(n28949), .X(\filter_0/n8575 ) );
  nand_x1_sg U44507 ( .A(n28950), .B(n28951), .X(\filter_0/n8574 ) );
  nand_x1_sg U44508 ( .A(n28952), .B(n28953), .X(\filter_0/n8573 ) );
  nand_x1_sg U44509 ( .A(n28954), .B(n28955), .X(\filter_0/n8572 ) );
  nand_x1_sg U44510 ( .A(n28956), .B(n28957), .X(\filter_0/n8571 ) );
  nand_x1_sg U44511 ( .A(n28958), .B(n28959), .X(\filter_0/n8570 ) );
  nand_x1_sg U44512 ( .A(n28960), .B(n28961), .X(\filter_0/n8569 ) );
  nand_x1_sg U44513 ( .A(n28962), .B(n28963), .X(\filter_0/n8568 ) );
  nand_x1_sg U44514 ( .A(n28420), .B(n28421), .X(\filter_0/n8821 ) );
  nand_x1_sg U44515 ( .A(n28422), .B(n28423), .X(\filter_0/n8820 ) );
  nand_x1_sg U44516 ( .A(n28424), .B(n28425), .X(\filter_0/n8819 ) );
  nand_x1_sg U44517 ( .A(n28426), .B(n28427), .X(\filter_0/n8818 ) );
  nand_x1_sg U44518 ( .A(n28428), .B(n28429), .X(\filter_0/n8817 ) );
  nand_x1_sg U44519 ( .A(n28430), .B(n28431), .X(\filter_0/n8816 ) );
  nand_x1_sg U44520 ( .A(n28432), .B(n28433), .X(\filter_0/n8815 ) );
  nand_x1_sg U44521 ( .A(n28434), .B(n28435), .X(\filter_0/n8814 ) );
  nand_x1_sg U44522 ( .A(n28436), .B(n28437), .X(\filter_0/n8813 ) );
  nand_x1_sg U44523 ( .A(n28438), .B(n28439), .X(\filter_0/n8812 ) );
  nand_x1_sg U44524 ( .A(n28440), .B(n28441), .X(\filter_0/n8811 ) );
  nand_x1_sg U44525 ( .A(n28442), .B(n28443), .X(\filter_0/n8810 ) );
  nand_x1_sg U44526 ( .A(n28444), .B(n28445), .X(\filter_0/n8809 ) );
  nand_x1_sg U44527 ( .A(n28446), .B(n28447), .X(\filter_0/n8808 ) );
  nand_x1_sg U44528 ( .A(n25874), .B(n25875), .X(n4155) );
  nand_x1_sg U44529 ( .A(n25916), .B(n25917), .X(n4134) );
  nand_x1_sg U44530 ( .A(n25918), .B(n25919), .X(n4133) );
  nand_x1_sg U44531 ( .A(n25920), .B(n25921), .X(n4132) );
  nand_x1_sg U44532 ( .A(n25922), .B(n25923), .X(n4131) );
  nand_x1_sg U44533 ( .A(n25924), .B(n25925), .X(n4130) );
  nand_x1_sg U44534 ( .A(n25926), .B(n25927), .X(n4129) );
  nand_x1_sg U44535 ( .A(n25928), .B(n25929), .X(n4128) );
  nand_x1_sg U44536 ( .A(n25930), .B(n25931), .X(n4127) );
  nand_x1_sg U44537 ( .A(n25932), .B(n25933), .X(n4126) );
  nand_x1_sg U44538 ( .A(n25934), .B(n25935), .X(n4125) );
  nand_x1_sg U44539 ( .A(n25936), .B(n25937), .X(n4124) );
  nand_x1_sg U44540 ( .A(n25938), .B(n25939), .X(n4123) );
  nand_x1_sg U44541 ( .A(n25940), .B(n25941), .X(n4122) );
  nand_x1_sg U44542 ( .A(n25942), .B(n25943), .X(n4121) );
  nand_x1_sg U44543 ( .A(n25944), .B(n25945), .X(n4120) );
  nand_x1_sg U44544 ( .A(n25946), .B(n25947), .X(n4119) );
  nand_x1_sg U44545 ( .A(n25948), .B(n25949), .X(n4118) );
  nand_x1_sg U44546 ( .A(n25950), .B(n25951), .X(n4117) );
  nand_x1_sg U44547 ( .A(n25952), .B(n25953), .X(n4116) );
  nand_x1_sg U44548 ( .A(n25954), .B(n25955), .X(n4115) );
  nand_x1_sg U44549 ( .A(n25996), .B(n25997), .X(n4094) );
  nand_x1_sg U44550 ( .A(n25998), .B(n25999), .X(n4093) );
  nand_x1_sg U44551 ( .A(n26000), .B(n26001), .X(n4092) );
  nand_x1_sg U44552 ( .A(n25618), .B(n25619), .X(n4283) );
  nand_x1_sg U44553 ( .A(n25620), .B(n25621), .X(n4282) );
  nand_x1_sg U44554 ( .A(n25622), .B(n25623), .X(n4281) );
  nand_x1_sg U44555 ( .A(n25624), .B(n25625), .X(n4280) );
  nand_x1_sg U44556 ( .A(n25626), .B(n25627), .X(n4279) );
  nand_x1_sg U44557 ( .A(n25628), .B(n25629), .X(n4278) );
  nand_x1_sg U44558 ( .A(n25630), .B(n25631), .X(n4277) );
  nand_x1_sg U44559 ( .A(n25632), .B(n25633), .X(n4276) );
  nand_x1_sg U44560 ( .A(n25634), .B(n25635), .X(n4275) );
  nand_x1_sg U44561 ( .A(n25636), .B(n25637), .X(n4274) );
  nand_x1_sg U44562 ( .A(n25638), .B(n25639), .X(n4273) );
  nand_x1_sg U44563 ( .A(n25680), .B(n25681), .X(n4252) );
  nand_x1_sg U44564 ( .A(n25044), .B(n25045), .X(n4570) );
  nand_x1_sg U44565 ( .A(n25046), .B(n25047), .X(n4569) );
  nand_x1_sg U44566 ( .A(n25048), .B(n25049), .X(n4568) );
  nand_x1_sg U44567 ( .A(n25050), .B(n25051), .X(n4567) );
  nand_x1_sg U44568 ( .A(n25052), .B(n25053), .X(n4566) );
  nand_x1_sg U44569 ( .A(n25054), .B(n25055), .X(n4565) );
  nand_x1_sg U44570 ( .A(n25056), .B(n25057), .X(n4564) );
  nand_x1_sg U44571 ( .A(n25058), .B(n25059), .X(n4563) );
  nand_x1_sg U44572 ( .A(n25060), .B(n25061), .X(n4562) );
  nand_x1_sg U44573 ( .A(n25062), .B(n25063), .X(n4561) );
  nand_x1_sg U44574 ( .A(n25064), .B(n25065), .X(n4560) );
  nand_x1_sg U44575 ( .A(n25066), .B(n25067), .X(n4559) );
  nand_x1_sg U44576 ( .A(n25068), .B(n25069), .X(n4558) );
  nand_x1_sg U44577 ( .A(n25070), .B(n25071), .X(n4557) );
  nand_x1_sg U44578 ( .A(n25072), .B(n25073), .X(n4556) );
  nand_x1_sg U44579 ( .A(n25074), .B(n25075), .X(n4555) );
  nand_x1_sg U44580 ( .A(n25076), .B(n25077), .X(n4554) );
  nand_x1_sg U44581 ( .A(n25078), .B(n25079), .X(n4553) );
  nand_x1_sg U44582 ( .A(n25080), .B(n25081), .X(n4552) );
  nand_x1_sg U44583 ( .A(n25082), .B(n25083), .X(n4551) );
  nand_x1_sg U44584 ( .A(n25298), .B(n25299), .X(n4443) );
  nand_x1_sg U44585 ( .A(n25300), .B(n25301), .X(n4442) );
  nand_x1_sg U44586 ( .A(n25302), .B(n25303), .X(n4441) );
  nand_x1_sg U44587 ( .A(n25304), .B(n25305), .X(n4440) );
  nand_x1_sg U44588 ( .A(n25306), .B(n25307), .X(n4439) );
  nand_x1_sg U44589 ( .A(n25308), .B(n25309), .X(n4438) );
  nand_x1_sg U44590 ( .A(n25310), .B(n25311), .X(n4437) );
  nand_x1_sg U44591 ( .A(n25312), .B(n25313), .X(n4436) );
  nand_x1_sg U44592 ( .A(n25314), .B(n25315), .X(n4435) );
  nand_x1_sg U44593 ( .A(n25316), .B(n25317), .X(n4434) );
  nand_x1_sg U44594 ( .A(n25318), .B(n25319), .X(n4433) );
  nand_x1_sg U44595 ( .A(n25320), .B(n25321), .X(n4432) );
  nand_x1_sg U44596 ( .A(n25322), .B(n25323), .X(n4431) );
  nand_x1_sg U44597 ( .A(n25358), .B(n25359), .X(n4413) );
  nand_x1_sg U44598 ( .A(n25360), .B(n25361), .X(n4412) );
  nand_x1_sg U44599 ( .A(n25362), .B(n25363), .X(n4411) );
  nand_x1_sg U44600 ( .A(n25364), .B(n25365), .X(n4410) );
  nand_x1_sg U44601 ( .A(n25366), .B(n25367), .X(n4409) );
  nand_x1_sg U44602 ( .A(n25368), .B(n25369), .X(n4408) );
  nand_x1_sg U44603 ( .A(n25370), .B(n25371), .X(n4407) );
  nand_x1_sg U44604 ( .A(n25372), .B(n25373), .X(n4406) );
  nand_x1_sg U44605 ( .A(n25374), .B(n25375), .X(n4405) );
  nand_x1_sg U44606 ( .A(n25376), .B(n25377), .X(n4404) );
  nand_x1_sg U44607 ( .A(n25378), .B(n25379), .X(n4403) );
  nand_x1_sg U44608 ( .A(n25380), .B(n25381), .X(n4402) );
  nand_x1_sg U44609 ( .A(n25382), .B(n25383), .X(n4401) );
  nand_x1_sg U44610 ( .A(n25384), .B(n25385), .X(n4400) );
  nand_x1_sg U44611 ( .A(n25386), .B(n25387), .X(n4399) );
  nand_x1_sg U44612 ( .A(n25388), .B(n25389), .X(n4398) );
  nand_x1_sg U44613 ( .A(n25390), .B(n25391), .X(n4397) );
  nand_x1_sg U44614 ( .A(n25392), .B(n25393), .X(n4396) );
  nand_x1_sg U44615 ( .A(n25394), .B(n25395), .X(n4395) );
  nand_x1_sg U44616 ( .A(n25396), .B(n25397), .X(n4394) );
  nand_x1_sg U44617 ( .A(n24728), .B(n24729), .X(n4728) );
  nand_x1_sg U44618 ( .A(n24730), .B(n24731), .X(n4727) );
  nand_x1_sg U44619 ( .A(n24732), .B(n24733), .X(n4726) );
  nand_x1_sg U44620 ( .A(n24734), .B(n24735), .X(n4725) );
  nand_x1_sg U44621 ( .A(n24736), .B(n24737), .X(n4724) );
  nand_x1_sg U44622 ( .A(n24738), .B(n24739), .X(n4723) );
  nand_x1_sg U44623 ( .A(n24740), .B(n24741), .X(n4722) );
  nand_x1_sg U44624 ( .A(n24742), .B(n24743), .X(n4721) );
  nand_x1_sg U44625 ( .A(n24744), .B(n24745), .X(n4720) );
  nand_x1_sg U44626 ( .A(n24746), .B(n24747), .X(n4719) );
  nand_x1_sg U44627 ( .A(n24748), .B(n24749), .X(n4718) );
  nand_x1_sg U44628 ( .A(n24750), .B(n24751), .X(n4717) );
  nand_x1_sg U44629 ( .A(n24752), .B(n24753), .X(n4716) );
  nand_x1_sg U44630 ( .A(n24754), .B(n24755), .X(n4715) );
  nand_x1_sg U44631 ( .A(n24756), .B(n24757), .X(n4714) );
  nand_x1_sg U44632 ( .A(n24758), .B(n24759), .X(n4713) );
  nand_x1_sg U44633 ( .A(n24760), .B(n24761), .X(n4712) );
  nand_x1_sg U44634 ( .A(n24762), .B(n24763), .X(n4711) );
  nand_x1_sg U44635 ( .A(n24764), .B(n24765), .X(n4710) );
  nand_x1_sg U44636 ( .A(n24766), .B(n24767), .X(n4709) );
  nand_x1_sg U44637 ( .A(n24808), .B(n24809), .X(n4688) );
  nand_x1_sg U44638 ( .A(n24810), .B(n24811), .X(n4687) );
  nand_x1_sg U44639 ( .A(n24812), .B(n24813), .X(n4686) );
  nand_x1_sg U44640 ( .A(n24814), .B(n24815), .X(n4685) );
  nand_x1_sg U44641 ( .A(n24816), .B(n24817), .X(n4684) );
  nand_x1_sg U44642 ( .A(n24818), .B(n24819), .X(n4683) );
  nand_x1_sg U44643 ( .A(n24820), .B(n24821), .X(n4682) );
  nand_x1_sg U44644 ( .A(n24822), .B(n24823), .X(n4681) );
  nand_x1_sg U44645 ( .A(n24824), .B(n24825), .X(n4680) );
  nand_x1_sg U44646 ( .A(n24826), .B(n24827), .X(n4679) );
  nand_x1_sg U44647 ( .A(n24828), .B(n24829), .X(n4678) );
  nand_x1_sg U44648 ( .A(n24830), .B(n24831), .X(n4677) );
  nand_x1_sg U44649 ( .A(n24832), .B(n24833), .X(n4676) );
  nand_x1_sg U44650 ( .A(n24834), .B(n24835), .X(n4675) );
  nand_x1_sg U44651 ( .A(n24836), .B(n24837), .X(n4674) );
  nand_x1_sg U44652 ( .A(n24838), .B(n24839), .X(n4673) );
  nand_x1_sg U44653 ( .A(n24840), .B(n24841), .X(n4672) );
  nand_x1_sg U44654 ( .A(n24842), .B(n24843), .X(n4671) );
  nand_x1_sg U44655 ( .A(n24844), .B(n24845), .X(n4670) );
  nand_x1_sg U44656 ( .A(n24846), .B(n24847), .X(n4669) );
  nand_x1_sg U44657 ( .A(n24252), .B(n24253), .X(n4966) );
  nand_x1_sg U44658 ( .A(n24254), .B(n24255), .X(n4965) );
  nand_x1_sg U44659 ( .A(n24256), .B(n24257), .X(n4964) );
  nand_x1_sg U44660 ( .A(n24258), .B(n24259), .X(n4963) );
  nand_x1_sg U44661 ( .A(n24260), .B(n24261), .X(n4962) );
  nand_x1_sg U44662 ( .A(n24262), .B(n24263), .X(n4961) );
  nand_x1_sg U44663 ( .A(n24264), .B(n24265), .X(n4960) );
  nand_x1_sg U44664 ( .A(n24266), .B(n24267), .X(n4959) );
  nand_x1_sg U44665 ( .A(n24268), .B(n24269), .X(n4958) );
  nand_x1_sg U44666 ( .A(n24270), .B(n24271), .X(n4957) );
  nand_x1_sg U44667 ( .A(n24272), .B(n24273), .X(n4956) );
  nand_x1_sg U44668 ( .A(n24492), .B(n24493), .X(n4846) );
  nand_x1_sg U44669 ( .A(n24494), .B(n24495), .X(n4845) );
  nand_x1_sg U44670 ( .A(n24496), .B(n24497), .X(n4844) );
  nand_x1_sg U44671 ( .A(n24498), .B(n24499), .X(n4843) );
  nand_x1_sg U44672 ( .A(n24500), .B(n24501), .X(n4842) );
  nand_x1_sg U44673 ( .A(n24502), .B(n24503), .X(n4841) );
  nand_x1_sg U44674 ( .A(n24504), .B(n24505), .X(n4840) );
  nand_x1_sg U44675 ( .A(n24506), .B(n24507), .X(n4839) );
  nand_x1_sg U44676 ( .A(n24508), .B(n24509), .X(n4838) );
  nand_x1_sg U44677 ( .A(n24510), .B(n24511), .X(n4837) );
  nand_x1_sg U44678 ( .A(n24512), .B(n24513), .X(n4836) );
  nand_x1_sg U44679 ( .A(n24514), .B(n24515), .X(n4835) );
  nand_x1_sg U44680 ( .A(n24516), .B(n24517), .X(n4834) );
  nand_x1_sg U44681 ( .A(n24518), .B(n24519), .X(n4833) );
  nand_x1_sg U44682 ( .A(n24520), .B(n24521), .X(n4832) );
  nand_x1_sg U44683 ( .A(n24522), .B(n24523), .X(n4831) );
  nand_x1_sg U44684 ( .A(n24524), .B(n24525), .X(n4830) );
  nand_x1_sg U44685 ( .A(n24526), .B(n24527), .X(n4829) );
  nand_x1_sg U44686 ( .A(n24528), .B(n24529), .X(n4828) );
  nand_x1_sg U44687 ( .A(n23890), .B(n23891), .X(n5147) );
  nand_x1_sg U44688 ( .A(n23892), .B(n23893), .X(n5146) );
  nand_x1_sg U44689 ( .A(n23894), .B(n23895), .X(n5145) );
  nand_x1_sg U44690 ( .A(n23936), .B(n23937), .X(n5124) );
  nand_x1_sg U44691 ( .A(n23938), .B(n23939), .X(n5123) );
  nand_x1_sg U44692 ( .A(n23940), .B(n23941), .X(n5122) );
  nand_x1_sg U44693 ( .A(n23942), .B(n23943), .X(n5121) );
  nand_x1_sg U44694 ( .A(n23944), .B(n23945), .X(n5120) );
  nand_x1_sg U44695 ( .A(n23946), .B(n23947), .X(n5119) );
  nand_x1_sg U44696 ( .A(n23948), .B(n23949), .X(n5118) );
  nand_x1_sg U44697 ( .A(n23950), .B(n23951), .X(n5117) );
  nand_x1_sg U44698 ( .A(n23952), .B(n23953), .X(n5116) );
  nand_x1_sg U44699 ( .A(n24164), .B(n24165), .X(n5010) );
  nand_x1_sg U44700 ( .A(n24166), .B(n24167), .X(n5009) );
  nand_x1_sg U44701 ( .A(n24168), .B(n24169), .X(n5008) );
  nand_x1_sg U44702 ( .A(n24170), .B(n24171), .X(n5007) );
  nand_x1_sg U44703 ( .A(n24172), .B(n24173), .X(n5006) );
  nand_x1_sg U44704 ( .A(n24174), .B(n24175), .X(n5005) );
  nand_x1_sg U44705 ( .A(n24176), .B(n24177), .X(n5004) );
  nand_x1_sg U44706 ( .A(n24178), .B(n24179), .X(n5003) );
  nand_x1_sg U44707 ( .A(n24180), .B(n24181), .X(n5002) );
  nand_x1_sg U44708 ( .A(n24182), .B(n24183), .X(n5001) );
  nand_x1_sg U44709 ( .A(n24184), .B(n24185), .X(n5000) );
  nand_x1_sg U44710 ( .A(n24186), .B(n24187), .X(n4999) );
  nand_x1_sg U44711 ( .A(n24188), .B(n24189), .X(n4998) );
  nand_x1_sg U44712 ( .A(n24190), .B(n24191), .X(n4997) );
  nand_x1_sg U44713 ( .A(n24192), .B(n24193), .X(n4996) );
  nand_x1_sg U44714 ( .A(n24194), .B(n24195), .X(n4995) );
  nand_x1_sg U44715 ( .A(n24196), .B(n24197), .X(n4994) );
  nand_x1_sg U44716 ( .A(n24198), .B(n24199), .X(n4993) );
  nand_x1_sg U44717 ( .A(n24200), .B(n24201), .X(n4992) );
  nand_x1_sg U44718 ( .A(n24202), .B(n24203), .X(n4991) );
  nand_x1_sg U44719 ( .A(n23686), .B(n23687), .X(n5249) );
  nand_x1_sg U44720 ( .A(n23688), .B(n23689), .X(n5248) );
  nand_x1_sg U44721 ( .A(n23690), .B(n23691), .X(n5247) );
  nand_x1_sg U44722 ( .A(n23692), .B(n23693), .X(n5246) );
  nand_x1_sg U44723 ( .A(n23694), .B(n23695), .X(n5245) );
  nand_x1_sg U44724 ( .A(n23696), .B(n23697), .X(n5244) );
  inv_x1_sg U44725 ( .A(n15340), .X(n42382) );
  nand_x1_sg U44726 ( .A(n25836), .B(n25837), .X(n4174) );
  nand_x1_sg U44727 ( .A(n25838), .B(n25839), .X(n4173) );
  nand_x1_sg U44728 ( .A(n25840), .B(n25841), .X(n4172) );
  nand_x1_sg U44729 ( .A(n25842), .B(n25843), .X(n4171) );
  nand_x1_sg U44730 ( .A(n25844), .B(n25845), .X(n4170) );
  nand_x1_sg U44731 ( .A(n25846), .B(n25847), .X(n4169) );
  nand_x1_sg U44732 ( .A(n25848), .B(n25849), .X(n4168) );
  nand_x1_sg U44733 ( .A(n25850), .B(n25851), .X(n4167) );
  nand_x1_sg U44734 ( .A(n25852), .B(n25853), .X(n4166) );
  nand_x1_sg U44735 ( .A(n25854), .B(n25855), .X(n4165) );
  nand_x1_sg U44736 ( .A(n25856), .B(n25857), .X(n4164) );
  nand_x1_sg U44737 ( .A(n25858), .B(n25859), .X(n4163) );
  nand_x1_sg U44738 ( .A(n25860), .B(n25861), .X(n4162) );
  nand_x1_sg U44739 ( .A(n25862), .B(n25863), .X(n4161) );
  nand_x1_sg U44740 ( .A(n25864), .B(n25865), .X(n4160) );
  nand_x1_sg U44741 ( .A(n25866), .B(n25867), .X(n4159) );
  nand_x1_sg U44742 ( .A(n25868), .B(n25869), .X(n4158) );
  nand_x1_sg U44743 ( .A(n25870), .B(n25871), .X(n4157) );
  nand_x1_sg U44744 ( .A(n25872), .B(n25873), .X(n4156) );
  nand_x1_sg U44745 ( .A(n26076), .B(n26077), .X(n4054) );
  nand_x1_sg U44746 ( .A(n26078), .B(n26079), .X(n4053) );
  nand_x1_sg U44747 ( .A(n26080), .B(n26081), .X(n4052) );
  nand_x1_sg U44748 ( .A(n26082), .B(n26083), .X(n4051) );
  nand_x1_sg U44749 ( .A(n26084), .B(n26085), .X(n4050) );
  nand_x1_sg U44750 ( .A(n26086), .B(n26087), .X(n4049) );
  nand_x1_sg U44751 ( .A(n26088), .B(n26089), .X(n4048) );
  nand_x1_sg U44752 ( .A(n26090), .B(n26091), .X(n4047) );
  nand_x1_sg U44753 ( .A(n26092), .B(n26093), .X(n4046) );
  nand_x1_sg U44754 ( .A(n26094), .B(n26095), .X(n4045) );
  nand_x1_sg U44755 ( .A(n26096), .B(n26097), .X(n4044) );
  nand_x1_sg U44756 ( .A(n26098), .B(n26099), .X(n4043) );
  nand_x1_sg U44757 ( .A(n26100), .B(n26101), .X(n4042) );
  nand_x1_sg U44758 ( .A(n26102), .B(n26103), .X(n4041) );
  nand_x1_sg U44759 ( .A(n26104), .B(n26105), .X(n4040) );
  nand_x1_sg U44760 ( .A(n26106), .B(n26107), .X(n4039) );
  nand_x1_sg U44761 ( .A(n26108), .B(n26109), .X(n4038) );
  nand_x1_sg U44762 ( .A(n26110), .B(n26111), .X(n4037) );
  nand_x1_sg U44763 ( .A(n26112), .B(n26113), .X(n4036) );
  nand_x1_sg U44764 ( .A(n26114), .B(n26115), .X(n4035) );
  nand_x1_sg U44765 ( .A(n25520), .B(n25521), .X(n4332) );
  nand_x1_sg U44766 ( .A(n25522), .B(n25523), .X(n4331) );
  nand_x1_sg U44767 ( .A(n25524), .B(n25525), .X(n4330) );
  nand_x1_sg U44768 ( .A(n25526), .B(n25527), .X(n4329) );
  nand_x1_sg U44769 ( .A(n25528), .B(n25529), .X(n4328) );
  nand_x1_sg U44770 ( .A(n25530), .B(n25531), .X(n4327) );
  nand_x1_sg U44771 ( .A(n25532), .B(n25533), .X(n4326) );
  nand_x1_sg U44772 ( .A(n25534), .B(n25535), .X(n4325) );
  nand_x1_sg U44773 ( .A(n25536), .B(n25537), .X(n4324) );
  nand_x1_sg U44774 ( .A(n25538), .B(n25539), .X(n4323) );
  nand_x1_sg U44775 ( .A(n25540), .B(n25541), .X(n4322) );
  nand_x1_sg U44776 ( .A(n25542), .B(n25543), .X(n4321) );
  nand_x1_sg U44777 ( .A(n25544), .B(n25545), .X(n4320) );
  nand_x1_sg U44778 ( .A(n25546), .B(n25547), .X(n4319) );
  nand_x1_sg U44779 ( .A(n25548), .B(n25549), .X(n4318) );
  nand_x1_sg U44780 ( .A(n25550), .B(n25551), .X(n4317) );
  nand_x1_sg U44781 ( .A(n25552), .B(n25553), .X(n4316) );
  nand_x1_sg U44782 ( .A(n25756), .B(n25757), .X(n4214) );
  nand_x1_sg U44783 ( .A(n25758), .B(n25759), .X(n4213) );
  nand_x1_sg U44784 ( .A(n25760), .B(n25761), .X(n4212) );
  nand_x1_sg U44785 ( .A(n25762), .B(n25763), .X(n4211) );
  nand_x1_sg U44786 ( .A(n25764), .B(n25765), .X(n4210) );
  nand_x1_sg U44787 ( .A(n25766), .B(n25767), .X(n4209) );
  nand_x1_sg U44788 ( .A(n25768), .B(n25769), .X(n4208) );
  nand_x1_sg U44789 ( .A(n25770), .B(n25771), .X(n4207) );
  nand_x1_sg U44790 ( .A(n25772), .B(n25773), .X(n4206) );
  nand_x1_sg U44791 ( .A(n25774), .B(n25775), .X(n4205) );
  nand_x1_sg U44792 ( .A(n25776), .B(n25777), .X(n4204) );
  nand_x1_sg U44793 ( .A(n25778), .B(n25779), .X(n4203) );
  nand_x1_sg U44794 ( .A(n25780), .B(n25781), .X(n4202) );
  nand_x1_sg U44795 ( .A(n25782), .B(n25783), .X(n4201) );
  nand_x1_sg U44796 ( .A(n25784), .B(n25785), .X(n4200) );
  nand_x1_sg U44797 ( .A(n25786), .B(n25787), .X(n4199) );
  nand_x1_sg U44798 ( .A(n25788), .B(n25789), .X(n4198) );
  nand_x1_sg U44799 ( .A(n25790), .B(n25791), .X(n4197) );
  nand_x1_sg U44800 ( .A(n25792), .B(n25793), .X(n4196) );
  nand_x1_sg U44801 ( .A(n25794), .B(n25795), .X(n4195) );
  nand_x1_sg U44802 ( .A(n25204), .B(n25205), .X(n4490) );
  nand_x1_sg U44803 ( .A(n25206), .B(n25207), .X(n4489) );
  nand_x1_sg U44804 ( .A(n25208), .B(n25209), .X(n4488) );
  nand_x1_sg U44805 ( .A(n25210), .B(n25211), .X(n4487) );
  nand_x1_sg U44806 ( .A(n25212), .B(n25213), .X(n4486) );
  nand_x1_sg U44807 ( .A(n25214), .B(n25215), .X(n4485) );
  nand_x1_sg U44808 ( .A(n25216), .B(n25217), .X(n4484) );
  nand_x1_sg U44809 ( .A(n25218), .B(n25219), .X(n4483) );
  nand_x1_sg U44810 ( .A(n25220), .B(n25221), .X(n4482) );
  nand_x1_sg U44811 ( .A(n25222), .B(n25223), .X(n4481) );
  nand_x1_sg U44812 ( .A(n25224), .B(n25225), .X(n4480) );
  nand_x1_sg U44813 ( .A(n25226), .B(n25227), .X(n4479) );
  nand_x1_sg U44814 ( .A(n25228), .B(n25229), .X(n4478) );
  nand_x1_sg U44815 ( .A(n25230), .B(n25231), .X(n4477) );
  nand_x1_sg U44816 ( .A(n25232), .B(n25233), .X(n4476) );
  nand_x1_sg U44817 ( .A(n25234), .B(n25235), .X(n4475) );
  nand_x1_sg U44818 ( .A(n25236), .B(n25237), .X(n4474) );
  nand_x1_sg U44819 ( .A(n25238), .B(n25239), .X(n4473) );
  nand_x1_sg U44820 ( .A(n25240), .B(n25241), .X(n4472) );
  nand_x1_sg U44821 ( .A(n25242), .B(n25243), .X(n4471) );
  nand_x1_sg U44822 ( .A(n25284), .B(n25285), .X(n4450) );
  nand_x1_sg U44823 ( .A(n25286), .B(n25287), .X(n4449) );
  nand_x1_sg U44824 ( .A(n25288), .B(n25289), .X(n4448) );
  nand_x1_sg U44825 ( .A(n25290), .B(n25291), .X(n4447) );
  nand_x1_sg U44826 ( .A(n25292), .B(n25293), .X(n4446) );
  nand_x1_sg U44827 ( .A(n25294), .B(n25295), .X(n4445) );
  nand_x1_sg U44828 ( .A(n25296), .B(n25297), .X(n4444) );
  nand_x1_sg U44829 ( .A(n24648), .B(n24649), .X(n4768) );
  nand_x1_sg U44830 ( .A(n24650), .B(n24651), .X(n4767) );
  nand_x1_sg U44831 ( .A(n24652), .B(n24653), .X(n4766) );
  nand_x1_sg U44832 ( .A(n24654), .B(n24655), .X(n4765) );
  nand_x1_sg U44833 ( .A(n24656), .B(n24657), .X(n4764) );
  nand_x1_sg U44834 ( .A(n24658), .B(n24659), .X(n4763) );
  nand_x1_sg U44835 ( .A(n24660), .B(n24661), .X(n4762) );
  nand_x1_sg U44836 ( .A(n24662), .B(n24663), .X(n4761) );
  nand_x1_sg U44837 ( .A(n24664), .B(n24665), .X(n4760) );
  nand_x1_sg U44838 ( .A(n24666), .B(n24667), .X(n4759) );
  nand_x1_sg U44839 ( .A(n24668), .B(n24669), .X(n4758) );
  nand_x1_sg U44840 ( .A(n24670), .B(n24671), .X(n4757) );
  nand_x1_sg U44841 ( .A(n24672), .B(n24673), .X(n4756) );
  nand_x1_sg U44842 ( .A(n24674), .B(n24675), .X(n4755) );
  nand_x1_sg U44843 ( .A(n24676), .B(n24677), .X(n4754) );
  nand_x1_sg U44844 ( .A(n24678), .B(n24679), .X(n4753) );
  nand_x1_sg U44845 ( .A(n24680), .B(n24681), .X(n4752) );
  nand_x1_sg U44846 ( .A(n24682), .B(n24683), .X(n4751) );
  nand_x1_sg U44847 ( .A(n24684), .B(n24685), .X(n4750) );
  nand_x1_sg U44848 ( .A(n24686), .B(n24687), .X(n4749) );
  nand_x1_sg U44849 ( .A(n24914), .B(n24915), .X(n4635) );
  nand_x1_sg U44850 ( .A(n24916), .B(n24917), .X(n4634) );
  nand_x1_sg U44851 ( .A(n24918), .B(n24919), .X(n4633) );
  nand_x1_sg U44852 ( .A(n24920), .B(n24921), .X(n4632) );
  nand_x1_sg U44853 ( .A(n24922), .B(n24923), .X(n4631) );
  nand_x1_sg U44854 ( .A(n24924), .B(n24925), .X(n4630) );
  nand_x1_sg U44855 ( .A(n24926), .B(n24927), .X(n4629) );
  nand_x1_sg U44856 ( .A(n24960), .B(n24961), .X(n4612) );
  nand_x1_sg U44857 ( .A(n24962), .B(n24963), .X(n4611) );
  nand_x1_sg U44858 ( .A(n24964), .B(n24965), .X(n4610) );
  nand_x1_sg U44859 ( .A(n24966), .B(n24967), .X(n4609) );
  nand_x1_sg U44860 ( .A(n24968), .B(n24969), .X(n4608) );
  nand_x1_sg U44861 ( .A(n24970), .B(n24971), .X(n4607) );
  nand_x1_sg U44862 ( .A(n24972), .B(n24973), .X(n4606) );
  nand_x1_sg U44863 ( .A(n24974), .B(n24975), .X(n4605) );
  nand_x1_sg U44864 ( .A(n24976), .B(n24977), .X(n4604) );
  nand_x1_sg U44865 ( .A(n24338), .B(n24339), .X(n4923) );
  nand_x1_sg U44866 ( .A(n24340), .B(n24341), .X(n4922) );
  nand_x1_sg U44867 ( .A(n24342), .B(n24343), .X(n4921) );
  nand_x1_sg U44868 ( .A(n24344), .B(n24345), .X(n4920) );
  nand_x1_sg U44869 ( .A(n24346), .B(n24347), .X(n4919) );
  nand_x1_sg U44870 ( .A(n24348), .B(n24349), .X(n4918) );
  nand_x1_sg U44871 ( .A(n24350), .B(n24351), .X(n4917) );
  nand_x1_sg U44872 ( .A(n24352), .B(n24353), .X(n4916) );
  nand_x1_sg U44873 ( .A(n24354), .B(n24355), .X(n4915) );
  nand_x1_sg U44874 ( .A(n24356), .B(n24357), .X(n4914) );
  nand_x1_sg U44875 ( .A(n24358), .B(n24359), .X(n4913) );
  nand_x1_sg U44876 ( .A(n24360), .B(n24361), .X(n4912) );
  nand_x1_sg U44877 ( .A(n24362), .B(n24363), .X(n4911) );
  nand_x1_sg U44878 ( .A(n24364), .B(n24365), .X(n4910) );
  nand_x1_sg U44879 ( .A(n24366), .B(n24367), .X(n4909) );
  nand_x1_sg U44880 ( .A(n24368), .B(n24369), .X(n4908) );
  nand_x1_sg U44881 ( .A(n24370), .B(n24371), .X(n4907) );
  nand_x1_sg U44882 ( .A(n24594), .B(n24595), .X(n4795) );
  nand_x1_sg U44883 ( .A(n24596), .B(n24597), .X(n4794) );
  nand_x1_sg U44884 ( .A(n24598), .B(n24599), .X(n4793) );
  nand_x1_sg U44885 ( .A(n24600), .B(n24601), .X(n4792) );
  nand_x1_sg U44886 ( .A(n24018), .B(n24019), .X(n5083) );
  nand_x1_sg U44887 ( .A(n24020), .B(n24021), .X(n5082) );
  nand_x1_sg U44888 ( .A(n24022), .B(n24023), .X(n5081) );
  nand_x1_sg U44889 ( .A(n24024), .B(n24025), .X(n5080) );
  nand_x1_sg U44890 ( .A(n24026), .B(n24027), .X(n5079) );
  nand_x1_sg U44891 ( .A(n24028), .B(n24029), .X(n5078) );
  nand_x1_sg U44892 ( .A(n24030), .B(n24031), .X(n5077) );
  nand_x1_sg U44893 ( .A(n24032), .B(n24033), .X(n5076) );
  nand_x1_sg U44894 ( .A(n24034), .B(n24035), .X(n5075) );
  nand_x1_sg U44895 ( .A(n24036), .B(n24037), .X(n5074) );
  nand_x1_sg U44896 ( .A(n24038), .B(n24039), .X(n5073) );
  nand_x1_sg U44897 ( .A(n24040), .B(n24041), .X(n5072) );
  nand_x1_sg U44898 ( .A(n24042), .B(n24043), .X(n5071) );
  nand_x1_sg U44899 ( .A(n24044), .B(n24045), .X(n5070) );
  nand_x1_sg U44900 ( .A(n24046), .B(n24047), .X(n5069) );
  nand_x1_sg U44901 ( .A(n24048), .B(n24049), .X(n5068) );
  nand_x1_sg U44902 ( .A(n24050), .B(n24051), .X(n5067) );
  nand_x1_sg U44903 ( .A(n24052), .B(n24053), .X(n5066) );
  nand_x1_sg U44904 ( .A(n24054), .B(n24055), .X(n5065) );
  nand_x1_sg U44905 ( .A(n24096), .B(n24097), .X(n5044) );
  nand_x1_sg U44906 ( .A(n24098), .B(n24099), .X(n5043) );
  nand_x1_sg U44907 ( .A(n24100), .B(n24101), .X(n5042) );
  nand_x1_sg U44908 ( .A(n24102), .B(n24103), .X(n5041) );
  nand_x1_sg U44909 ( .A(n24104), .B(n24105), .X(n5040) );
  nand_x1_sg U44910 ( .A(n24106), .B(n24107), .X(n5039) );
  nand_x1_sg U44911 ( .A(n24108), .B(n24109), .X(n5038) );
  nand_x1_sg U44912 ( .A(n24110), .B(n24111), .X(n5037) );
  nand_x1_sg U44913 ( .A(n24112), .B(n24113), .X(n5036) );
  nand_x1_sg U44914 ( .A(n24114), .B(n24115), .X(n5035) );
  nand_x1_sg U44915 ( .A(n24116), .B(n24117), .X(n5034) );
  nand_x1_sg U44916 ( .A(n24118), .B(n24119), .X(n5033) );
  nand_x1_sg U44917 ( .A(n24120), .B(n24121), .X(n5032) );
  nand_x1_sg U44918 ( .A(n24122), .B(n24123), .X(n5031) );
  nand_x1_sg U44919 ( .A(n24124), .B(n24125), .X(n5030) );
  nand_x1_sg U44920 ( .A(n24126), .B(n24127), .X(n5029) );
  nand_x1_sg U44921 ( .A(n24128), .B(n24129), .X(n5028) );
  nand_x1_sg U44922 ( .A(n24130), .B(n24131), .X(n5027) );
  nand_x1_sg U44923 ( .A(n24132), .B(n24133), .X(n5026) );
  nand_x1_sg U44924 ( .A(n24134), .B(n24135), .X(n5025) );
  nand_x1_sg U44925 ( .A(n23766), .B(n23767), .X(n5209) );
  nand_x1_sg U44926 ( .A(n23768), .B(n23769), .X(n5208) );
  nand_x1_sg U44927 ( .A(n23770), .B(n23771), .X(n5207) );
  nand_x1_sg U44928 ( .A(n23772), .B(n23773), .X(n5206) );
  nand_x1_sg U44929 ( .A(n23774), .B(n23775), .X(n5205) );
  nand_x1_sg U44930 ( .A(n23776), .B(n23777), .X(n5204) );
  nand_x1_sg U44931 ( .A(n23778), .B(n23779), .X(n5203) );
  nand_x1_sg U44932 ( .A(n23780), .B(n23781), .X(n5202) );
  nand_x1_sg U44933 ( .A(n23782), .B(n23783), .X(n5201) );
  nand_x1_sg U44934 ( .A(n23784), .B(n23785), .X(n5200) );
  nand_x1_sg U44935 ( .A(n23786), .B(n23787), .X(n5199) );
  nand_x1_sg U44936 ( .A(n23788), .B(n23789), .X(n5198) );
  nand_x1_sg U44937 ( .A(n23790), .B(n23791), .X(n5197) );
  nand_x1_sg U44938 ( .A(n23792), .B(n23793), .X(n5196) );
  nand_x1_sg U44939 ( .A(n23794), .B(n23795), .X(n5195) );
  nand_x1_sg U44940 ( .A(n23796), .B(n23797), .X(n5194) );
  nand_x1_sg U44941 ( .A(n23798), .B(n23799), .X(n5193) );
  nand_x1_sg U44942 ( .A(n23800), .B(n23801), .X(n5192) );
  nand_x1_sg U44943 ( .A(n23802), .B(n23803), .X(n5191) );
  nand_x1_sg U44944 ( .A(n23804), .B(n23805), .X(n5190) );
  nand_x1_sg U44945 ( .A(n28377), .B(n28378), .X(\filter_0/n8841 ) );
  nand_x1_sg U44946 ( .A(n28379), .B(n28380), .X(\filter_0/n8840 ) );
  nand_x1_sg U44947 ( .A(n28381), .B(n28382), .X(\filter_0/n8839 ) );
  nand_x1_sg U44948 ( .A(n28383), .B(n28384), .X(\filter_0/n8838 ) );
  nand_x1_sg U44949 ( .A(n28385), .B(n28386), .X(\filter_0/n8837 ) );
  nand_x1_sg U44950 ( .A(n28387), .B(n28388), .X(\filter_0/n8836 ) );
  nand_x1_sg U44951 ( .A(n28389), .B(n28390), .X(\filter_0/n8835 ) );
  nand_x1_sg U44952 ( .A(n28391), .B(n28392), .X(\filter_0/n8834 ) );
  nand_x1_sg U44953 ( .A(n28393), .B(n28394), .X(\filter_0/n8833 ) );
  nand_x1_sg U44954 ( .A(n28395), .B(n28396), .X(\filter_0/n8832 ) );
  nand_x1_sg U44955 ( .A(n28397), .B(n28398), .X(\filter_0/n8831 ) );
  nand_x1_sg U44956 ( .A(n28399), .B(n28400), .X(\filter_0/n8830 ) );
  nand_x1_sg U44957 ( .A(n28401), .B(n28402), .X(\filter_0/n8829 ) );
  nand_x1_sg U44958 ( .A(n28403), .B(n28404), .X(\filter_0/n8828 ) );
  nand_x1_sg U44959 ( .A(n28590), .B(n28591), .X(\filter_0/n8741 ) );
  nand_x1_sg U44960 ( .A(n28592), .B(n28593), .X(\filter_0/n8740 ) );
  nand_x1_sg U44961 ( .A(n28594), .B(n28595), .X(\filter_0/n8739 ) );
  nand_x1_sg U44962 ( .A(n28596), .B(n28597), .X(\filter_0/n8738 ) );
  nand_x1_sg U44963 ( .A(n28598), .B(n28599), .X(\filter_0/n8737 ) );
  nand_x1_sg U44964 ( .A(n28600), .B(n28601), .X(\filter_0/n8736 ) );
  nand_x1_sg U44965 ( .A(n28602), .B(n28603), .X(\filter_0/n8735 ) );
  nand_x1_sg U44966 ( .A(n28604), .B(n28605), .X(\filter_0/n8734 ) );
  nand_x1_sg U44967 ( .A(n28606), .B(n28607), .X(\filter_0/n8733 ) );
  nand_x1_sg U44968 ( .A(n28608), .B(n28609), .X(\filter_0/n8732 ) );
  nand_x1_sg U44969 ( .A(n28610), .B(n28611), .X(\filter_0/n8731 ) );
  nand_x1_sg U44970 ( .A(n28612), .B(n28613), .X(\filter_0/n8730 ) );
  nand_x1_sg U44971 ( .A(n28614), .B(n28615), .X(\filter_0/n8729 ) );
  nand_x1_sg U44972 ( .A(n28616), .B(n28617), .X(\filter_0/n8728 ) );
  nand_x1_sg U44973 ( .A(n28760), .B(n28761), .X(\filter_0/n8661 ) );
  nand_x1_sg U44974 ( .A(n28762), .B(n28763), .X(\filter_0/n8660 ) );
  nand_x1_sg U44975 ( .A(n28764), .B(n28765), .X(\filter_0/n8659 ) );
  nand_x1_sg U44976 ( .A(n28766), .B(n28767), .X(\filter_0/n8658 ) );
  nand_x1_sg U44977 ( .A(n28768), .B(n28769), .X(\filter_0/n8657 ) );
  nand_x1_sg U44978 ( .A(n28770), .B(n28771), .X(\filter_0/n8656 ) );
  nand_x1_sg U44979 ( .A(n28772), .B(n28773), .X(\filter_0/n8655 ) );
  nand_x1_sg U44980 ( .A(n28774), .B(n28775), .X(\filter_0/n8654 ) );
  nand_x1_sg U44981 ( .A(n28776), .B(n28777), .X(\filter_0/n8653 ) );
  nand_x1_sg U44982 ( .A(n28778), .B(n28779), .X(\filter_0/n8652 ) );
  nand_x1_sg U44983 ( .A(n28780), .B(n28781), .X(\filter_0/n8651 ) );
  nand_x1_sg U44984 ( .A(n28782), .B(n28783), .X(\filter_0/n8650 ) );
  nand_x1_sg U44985 ( .A(n28784), .B(n28785), .X(\filter_0/n8649 ) );
  nand_x1_sg U44986 ( .A(n28786), .B(n28787), .X(\filter_0/n8648 ) );
  nand_x1_sg U44987 ( .A(n29631), .B(n29632), .X(\filter_0/n8259 ) );
  nand_x1_sg U44988 ( .A(n33390), .B(\filter_0/n8175 ), .X(n29632) );
  nand_x1_sg U44989 ( .A(n29633), .B(n29634), .X(\filter_0/n8258 ) );
  nand_x1_sg U44990 ( .A(n33391), .B(\filter_0/n8174 ), .X(n29634) );
  nand_x1_sg U44991 ( .A(n29115), .B(n29116), .X(\filter_0/n8499 ) );
  nand_x1_sg U44992 ( .A(n33456), .B(\filter_0/n8095 ), .X(n29116) );
  nand_x1_sg U44993 ( .A(n29117), .B(n29118), .X(\filter_0/n8498 ) );
  nand_x1_sg U44994 ( .A(n33456), .B(\filter_0/n8094 ), .X(n29118) );
  nand_x1_sg U44995 ( .A(n28932), .B(n28933), .X(\filter_0/n8583 ) );
  nand_x1_sg U44996 ( .A(n33450), .B(\filter_0/n7846 ), .X(n28933) );
  nand_x1_sg U44997 ( .A(n28934), .B(n28935), .X(\filter_0/n8582 ) );
  nand_x1_sg U44998 ( .A(n29979), .B(\filter_0/n7845 ), .X(n28935) );
  nand_x1_sg U44999 ( .A(n28416), .B(n28417), .X(\filter_0/n8823 ) );
  nand_x1_sg U45000 ( .A(n33387), .B(\filter_0/n7766 ), .X(n28417) );
  nand_x1_sg U45001 ( .A(n28418), .B(n28419), .X(\filter_0/n8822 ) );
  nand_x1_sg U45002 ( .A(n29953), .B(\filter_0/n7765 ), .X(n28419) );
  inv_x1_sg U45003 ( .A(n15325), .X(n42387) );
  nand_x1_sg U45004 ( .A(n28373), .B(n28374), .X(\filter_0/n8843 ) );
  nand_x1_sg U45005 ( .A(n33448), .B(\filter_0/n7906 ), .X(n28374) );
  nand_x1_sg U45006 ( .A(n28375), .B(n28376), .X(\filter_0/n8842 ) );
  nand_x1_sg U45007 ( .A(n29977), .B(\filter_0/n7905 ), .X(n28376) );
  nand_x1_sg U45008 ( .A(n28586), .B(n28587), .X(\filter_0/n8743 ) );
  nand_x1_sg U45009 ( .A(n33380), .B(\filter_0/n7686 ), .X(n28587) );
  nand_x1_sg U45010 ( .A(n28588), .B(n28589), .X(\filter_0/n8742 ) );
  nand_x1_sg U45011 ( .A(n33381), .B(\filter_0/n7685 ), .X(n28589) );
  nand_x1_sg U45012 ( .A(n28756), .B(n28757), .X(\filter_0/n8663 ) );
  nand_x1_sg U45013 ( .A(n33377), .B(\filter_0/n7666 ), .X(n28757) );
  nand_x1_sg U45014 ( .A(n28758), .B(n28759), .X(\filter_0/n8662 ) );
  nand_x1_sg U45015 ( .A(n33378), .B(\filter_0/n7665 ), .X(n28759) );
  nand_x1_sg U45016 ( .A(n28334), .B(n28335), .X(\filter_0/n8861 ) );
  nand_x1_sg U45017 ( .A(n28336), .B(n28337), .X(\filter_0/n8860 ) );
  nand_x1_sg U45018 ( .A(n28338), .B(n28339), .X(\filter_0/n8859 ) );
  nand_x1_sg U45019 ( .A(n28340), .B(n28341), .X(\filter_0/n8858 ) );
  nand_x1_sg U45020 ( .A(n28342), .B(n28343), .X(\filter_0/n8857 ) );
  nand_x1_sg U45021 ( .A(n28344), .B(n28345), .X(\filter_0/n8856 ) );
  nand_x1_sg U45022 ( .A(n28346), .B(n28347), .X(\filter_0/n8855 ) );
  nand_x1_sg U45023 ( .A(n28348), .B(n28349), .X(\filter_0/n8854 ) );
  nand_x1_sg U45024 ( .A(n28350), .B(n28351), .X(\filter_0/n8853 ) );
  nand_x1_sg U45025 ( .A(n28352), .B(n28353), .X(\filter_0/n8852 ) );
  nand_x1_sg U45026 ( .A(n28354), .B(n28355), .X(\filter_0/n8851 ) );
  nand_x1_sg U45027 ( .A(n28356), .B(n28357), .X(\filter_0/n8850 ) );
  nand_x1_sg U45028 ( .A(n28358), .B(n28359), .X(\filter_0/n8849 ) );
  nand_x1_sg U45029 ( .A(n28360), .B(n28361), .X(\filter_0/n8848 ) );
  nand_x1_sg U45030 ( .A(n28290), .B(n28291), .X(\filter_0/n8881 ) );
  nand_x1_sg U45031 ( .A(n28292), .B(n28293), .X(\filter_0/n8880 ) );
  nand_x1_sg U45032 ( .A(n28294), .B(n28295), .X(\filter_0/n8879 ) );
  nand_x1_sg U45033 ( .A(n28296), .B(n28297), .X(\filter_0/n8878 ) );
  nand_x1_sg U45034 ( .A(n28298), .B(n28299), .X(\filter_0/n8877 ) );
  nand_x1_sg U45035 ( .A(n28300), .B(n28301), .X(\filter_0/n8876 ) );
  nand_x1_sg U45036 ( .A(n28302), .B(n28303), .X(\filter_0/n8875 ) );
  nand_x1_sg U45037 ( .A(n28304), .B(n28305), .X(\filter_0/n8874 ) );
  nand_x1_sg U45038 ( .A(n28306), .B(n28307), .X(\filter_0/n8873 ) );
  nand_x1_sg U45039 ( .A(n28308), .B(n28309), .X(\filter_0/n8872 ) );
  nand_x1_sg U45040 ( .A(n28310), .B(n28311), .X(\filter_0/n8871 ) );
  nand_x1_sg U45041 ( .A(n28312), .B(n28313), .X(\filter_0/n8870 ) );
  nand_x1_sg U45042 ( .A(n28314), .B(n28315), .X(\filter_0/n8869 ) );
  nand_x1_sg U45043 ( .A(n28316), .B(n28317), .X(\filter_0/n8868 ) );
  nand_x1_sg U45044 ( .A(n28506), .B(n28507), .X(\filter_0/n8781 ) );
  nand_x1_sg U45045 ( .A(n28508), .B(n28509), .X(\filter_0/n8780 ) );
  nand_x1_sg U45046 ( .A(n28510), .B(n28511), .X(\filter_0/n8779 ) );
  nand_x1_sg U45047 ( .A(n28512), .B(n28513), .X(\filter_0/n8778 ) );
  nand_x1_sg U45048 ( .A(n28514), .B(n28515), .X(\filter_0/n8777 ) );
  nand_x1_sg U45049 ( .A(n28516), .B(n28517), .X(\filter_0/n8776 ) );
  nand_x1_sg U45050 ( .A(n28518), .B(n28519), .X(\filter_0/n8775 ) );
  nand_x1_sg U45051 ( .A(n28520), .B(n28521), .X(\filter_0/n8774 ) );
  nand_x1_sg U45052 ( .A(n28522), .B(n28523), .X(\filter_0/n8773 ) );
  nand_x1_sg U45053 ( .A(n28524), .B(n28525), .X(\filter_0/n8772 ) );
  nand_x1_sg U45054 ( .A(n28526), .B(n28527), .X(\filter_0/n8771 ) );
  nand_x1_sg U45055 ( .A(n28528), .B(n28529), .X(\filter_0/n8770 ) );
  nand_x1_sg U45056 ( .A(n28530), .B(n28531), .X(\filter_0/n8769 ) );
  nand_x1_sg U45057 ( .A(n28532), .B(n28533), .X(\filter_0/n8768 ) );
  nand_x1_sg U45058 ( .A(n28464), .B(n28465), .X(\filter_0/n8801 ) );
  nand_x1_sg U45059 ( .A(n28466), .B(n28467), .X(\filter_0/n8800 ) );
  nand_x1_sg U45060 ( .A(n28468), .B(n28469), .X(\filter_0/n8799 ) );
  nand_x1_sg U45061 ( .A(n28470), .B(n28471), .X(\filter_0/n8798 ) );
  nand_x1_sg U45062 ( .A(n28472), .B(n28473), .X(\filter_0/n8797 ) );
  nand_x1_sg U45063 ( .A(n28474), .B(n28475), .X(\filter_0/n8796 ) );
  nand_x1_sg U45064 ( .A(n28476), .B(n28477), .X(\filter_0/n8795 ) );
  nand_x1_sg U45065 ( .A(n28478), .B(n28479), .X(\filter_0/n8794 ) );
  nand_x1_sg U45066 ( .A(n28480), .B(n28481), .X(\filter_0/n8793 ) );
  nand_x1_sg U45067 ( .A(n28482), .B(n28483), .X(\filter_0/n8792 ) );
  nand_x1_sg U45068 ( .A(n28484), .B(n28485), .X(\filter_0/n8791 ) );
  nand_x1_sg U45069 ( .A(n28486), .B(n28487), .X(\filter_0/n8790 ) );
  nand_x1_sg U45070 ( .A(n28488), .B(n28489), .X(\filter_0/n8789 ) );
  nand_x1_sg U45071 ( .A(n28490), .B(n28491), .X(\filter_0/n8788 ) );
  nand_x1_sg U45072 ( .A(n28633), .B(n28634), .X(\filter_0/n8721 ) );
  nand_x1_sg U45073 ( .A(n28635), .B(n28636), .X(\filter_0/n8720 ) );
  nand_x1_sg U45074 ( .A(n28637), .B(n28638), .X(\filter_0/n8719 ) );
  nand_x1_sg U45075 ( .A(n28639), .B(n28640), .X(\filter_0/n8718 ) );
  nand_x1_sg U45076 ( .A(n28641), .B(n28642), .X(\filter_0/n8717 ) );
  nand_x1_sg U45077 ( .A(n28643), .B(n28644), .X(\filter_0/n8716 ) );
  nand_x1_sg U45078 ( .A(n28645), .B(n28646), .X(\filter_0/n8715 ) );
  nand_x1_sg U45079 ( .A(n28647), .B(n28648), .X(\filter_0/n8714 ) );
  nand_x1_sg U45080 ( .A(n28649), .B(n28650), .X(\filter_0/n8713 ) );
  nand_x1_sg U45081 ( .A(n28651), .B(n28652), .X(\filter_0/n8712 ) );
  nand_x1_sg U45082 ( .A(n28653), .B(n28654), .X(\filter_0/n8711 ) );
  nand_x1_sg U45083 ( .A(n28655), .B(n28656), .X(\filter_0/n8710 ) );
  nand_x1_sg U45084 ( .A(n28657), .B(n28658), .X(\filter_0/n8709 ) );
  nand_x1_sg U45085 ( .A(n28659), .B(n28660), .X(\filter_0/n8708 ) );
  nand_x1_sg U45086 ( .A(n28675), .B(n28676), .X(\filter_0/n8701 ) );
  nand_x1_sg U45087 ( .A(n28677), .B(n28678), .X(\filter_0/n8700 ) );
  nand_x1_sg U45088 ( .A(n28679), .B(n28680), .X(\filter_0/n8699 ) );
  nand_x1_sg U45089 ( .A(n28681), .B(n28682), .X(\filter_0/n8698 ) );
  nand_x1_sg U45090 ( .A(n28683), .B(n28684), .X(\filter_0/n8697 ) );
  nand_x1_sg U45091 ( .A(n28685), .B(n28686), .X(\filter_0/n8696 ) );
  nand_x1_sg U45092 ( .A(n28687), .B(n28688), .X(\filter_0/n8695 ) );
  nand_x1_sg U45093 ( .A(n28689), .B(n28690), .X(\filter_0/n8694 ) );
  nand_x1_sg U45094 ( .A(n28691), .B(n28692), .X(\filter_0/n8693 ) );
  nand_x1_sg U45095 ( .A(n28693), .B(n28694), .X(\filter_0/n8692 ) );
  nand_x1_sg U45096 ( .A(n28695), .B(n28696), .X(\filter_0/n8691 ) );
  nand_x1_sg U45097 ( .A(n28697), .B(n28698), .X(\filter_0/n8690 ) );
  nand_x1_sg U45098 ( .A(n28699), .B(n28700), .X(\filter_0/n8689 ) );
  nand_x1_sg U45099 ( .A(n28701), .B(n28702), .X(\filter_0/n8688 ) );
  nand_x1_sg U45100 ( .A(n28805), .B(n28806), .X(\filter_0/n8641 ) );
  nand_x1_sg U45101 ( .A(n28807), .B(n28808), .X(\filter_0/n8640 ) );
  nand_x1_sg U45102 ( .A(n28809), .B(n28810), .X(\filter_0/n8639 ) );
  nand_x1_sg U45103 ( .A(n28811), .B(n28812), .X(\filter_0/n8638 ) );
  nand_x1_sg U45104 ( .A(n28813), .B(n28814), .X(\filter_0/n8637 ) );
  nand_x1_sg U45105 ( .A(n28815), .B(n28816), .X(\filter_0/n8636 ) );
  nand_x1_sg U45106 ( .A(n28817), .B(n28818), .X(\filter_0/n8635 ) );
  nand_x1_sg U45107 ( .A(n28819), .B(n28820), .X(\filter_0/n8634 ) );
  nand_x1_sg U45108 ( .A(n28821), .B(n28822), .X(\filter_0/n8633 ) );
  nand_x1_sg U45109 ( .A(n28823), .B(n28824), .X(\filter_0/n8632 ) );
  nand_x1_sg U45110 ( .A(n28825), .B(n28826), .X(\filter_0/n8631 ) );
  nand_x1_sg U45111 ( .A(n28827), .B(n28828), .X(\filter_0/n8630 ) );
  nand_x1_sg U45112 ( .A(n28829), .B(n28830), .X(\filter_0/n8629 ) );
  nand_x1_sg U45113 ( .A(n28831), .B(n28832), .X(\filter_0/n8628 ) );
  nand_x1_sg U45114 ( .A(n28849), .B(n28850), .X(\filter_0/n8621 ) );
  nand_x1_sg U45115 ( .A(n28851), .B(n28852), .X(\filter_0/n8620 ) );
  nand_x1_sg U45116 ( .A(n28853), .B(n28854), .X(\filter_0/n8619 ) );
  nand_x1_sg U45117 ( .A(n28855), .B(n28856), .X(\filter_0/n8618 ) );
  nand_x1_sg U45118 ( .A(n28857), .B(n28858), .X(\filter_0/n8617 ) );
  nand_x1_sg U45119 ( .A(n28859), .B(n28860), .X(\filter_0/n8616 ) );
  nand_x1_sg U45120 ( .A(n28861), .B(n28862), .X(\filter_0/n8615 ) );
  nand_x1_sg U45121 ( .A(n28863), .B(n28864), .X(\filter_0/n8614 ) );
  nand_x1_sg U45122 ( .A(n28865), .B(n28866), .X(\filter_0/n8613 ) );
  nand_x1_sg U45123 ( .A(n28867), .B(n28868), .X(\filter_0/n8612 ) );
  nand_x1_sg U45124 ( .A(n28869), .B(n28870), .X(\filter_0/n8611 ) );
  nand_x1_sg U45125 ( .A(n28871), .B(n28872), .X(\filter_0/n8610 ) );
  nand_x1_sg U45126 ( .A(n28873), .B(n28874), .X(\filter_0/n8609 ) );
  nand_x1_sg U45127 ( .A(n28875), .B(n28876), .X(\filter_0/n8608 ) );
  nand_x1_sg U45128 ( .A(n29621), .B(n29622), .X(\filter_0/n8263 ) );
  nand_x1_sg U45129 ( .A(n29955), .B(\filter_0/n8179 ), .X(n29622) );
  nand_x1_sg U45130 ( .A(n29625), .B(n29626), .X(\filter_0/n8262 ) );
  nand_x1_sg U45131 ( .A(n33393), .B(\filter_0/n8178 ), .X(n29626) );
  nand_x1_sg U45132 ( .A(n29627), .B(n29628), .X(\filter_0/n8261 ) );
  nand_x1_sg U45133 ( .A(n33390), .B(\filter_0/n8177 ), .X(n29628) );
  nand_x1_sg U45134 ( .A(n29629), .B(n29630), .X(\filter_0/n8260 ) );
  nand_x1_sg U45135 ( .A(n33393), .B(\filter_0/n8176 ), .X(n29630) );
  nand_x1_sg U45136 ( .A(n29105), .B(n29106), .X(\filter_0/n8503 ) );
  nand_x1_sg U45137 ( .A(n33458), .B(\filter_0/n8099 ), .X(n29106) );
  nand_x1_sg U45138 ( .A(n29109), .B(n29110), .X(\filter_0/n8502 ) );
  nand_x1_sg U45139 ( .A(n29981), .B(\filter_0/n8098 ), .X(n29110) );
  nand_x1_sg U45140 ( .A(n29111), .B(n29112), .X(\filter_0/n8501 ) );
  nand_x1_sg U45141 ( .A(n33455), .B(\filter_0/n8097 ), .X(n29112) );
  nand_x1_sg U45142 ( .A(n29113), .B(n29114), .X(\filter_0/n8500 ) );
  nand_x1_sg U45143 ( .A(n33457), .B(\filter_0/n8096 ), .X(n29114) );
  nand_x1_sg U45144 ( .A(n28922), .B(n28923), .X(\filter_0/n8587 ) );
  nand_x1_sg U45145 ( .A(n33452), .B(\filter_0/n7850 ), .X(n28923) );
  nand_x1_sg U45146 ( .A(n28926), .B(n28927), .X(\filter_0/n8586 ) );
  nand_x1_sg U45147 ( .A(n33450), .B(\filter_0/n7849 ), .X(n28927) );
  nand_x1_sg U45148 ( .A(n28928), .B(n28929), .X(\filter_0/n8585 ) );
  nand_x1_sg U45149 ( .A(n33451), .B(\filter_0/n7848 ), .X(n28929) );
  nand_x1_sg U45150 ( .A(n28930), .B(n28931), .X(\filter_0/n8584 ) );
  nand_x1_sg U45151 ( .A(n33452), .B(\filter_0/n7847 ), .X(n28931) );
  nand_x1_sg U45152 ( .A(n28406), .B(n28407), .X(\filter_0/n8827 ) );
  nand_x1_sg U45153 ( .A(n33387), .B(\filter_0/n7770 ), .X(n28407) );
  nand_x1_sg U45154 ( .A(n28410), .B(n28411), .X(\filter_0/n8826 ) );
  nand_x1_sg U45155 ( .A(n33385), .B(\filter_0/n7769 ), .X(n28411) );
  nand_x1_sg U45156 ( .A(n28412), .B(n28413), .X(\filter_0/n8825 ) );
  nand_x1_sg U45157 ( .A(n33386), .B(\filter_0/n7768 ), .X(n28413) );
  nand_x1_sg U45158 ( .A(n28414), .B(n28415), .X(\filter_0/n8824 ) );
  nand_x1_sg U45159 ( .A(n33387), .B(\filter_0/n7767 ), .X(n28415) );
  nand_x1_sg U45160 ( .A(n29424), .B(n29425), .X(\filter_0/n8353 ) );
  nand_x1_sg U45161 ( .A(n29436), .B(n29437), .X(\filter_0/n8347 ) );
  nand_x1_sg U45162 ( .A(n29600), .B(n29601), .X(\filter_0/n8273 ) );
  nand_x1_sg U45163 ( .A(n29612), .B(n29613), .X(\filter_0/n8267 ) );
  nand_x1_sg U45164 ( .A(n28725), .B(n28726), .X(\filter_0/n8677 ) );
  nand_x1_sg U45165 ( .A(n28737), .B(n28738), .X(\filter_0/n8671 ) );
  nand_x1_sg U45166 ( .A(n28901), .B(n28902), .X(\filter_0/n8597 ) );
  nand_x1_sg U45167 ( .A(n28913), .B(n28914), .X(\filter_0/n8591 ) );
  nand_x1_sg U45168 ( .A(n29420), .B(n29421), .X(\filter_0/n8355 ) );
  nand_x1_sg U45169 ( .A(n29432), .B(n29433), .X(\filter_0/n8349 ) );
  nand_x1_sg U45170 ( .A(n29596), .B(n29597), .X(\filter_0/n8275 ) );
  nand_x1_sg U45171 ( .A(n29608), .B(n29609), .X(\filter_0/n8269 ) );
  nand_x1_sg U45172 ( .A(n28721), .B(n28722), .X(\filter_0/n8679 ) );
  nand_x1_sg U45173 ( .A(n28733), .B(n28734), .X(\filter_0/n8673 ) );
  nand_x1_sg U45174 ( .A(n28897), .B(n28898), .X(\filter_0/n8599 ) );
  nand_x1_sg U45175 ( .A(n28909), .B(n28910), .X(\filter_0/n8593 ) );
  nand_x1_sg U45176 ( .A(n29416), .B(n29417), .X(\filter_0/n8357 ) );
  nand_x1_sg U45177 ( .A(n29428), .B(n29429), .X(\filter_0/n8351 ) );
  nand_x1_sg U45178 ( .A(n29440), .B(n29441), .X(\filter_0/n8345 ) );
  nand_x1_sg U45179 ( .A(n29592), .B(n29593), .X(\filter_0/n8277 ) );
  nand_x1_sg U45180 ( .A(n29604), .B(n29605), .X(\filter_0/n8271 ) );
  nand_x1_sg U45181 ( .A(n29616), .B(n29617), .X(\filter_0/n8265 ) );
  nand_x1_sg U45182 ( .A(n28717), .B(n28718), .X(\filter_0/n8681 ) );
  nand_x1_sg U45183 ( .A(n28729), .B(n28730), .X(\filter_0/n8675 ) );
  nand_x1_sg U45184 ( .A(n28741), .B(n28742), .X(\filter_0/n8669 ) );
  nand_x1_sg U45185 ( .A(n28893), .B(n28894), .X(\filter_0/n8601 ) );
  nand_x1_sg U45186 ( .A(n28905), .B(n28906), .X(\filter_0/n8595 ) );
  nand_x1_sg U45187 ( .A(n28917), .B(n28918), .X(\filter_0/n8589 ) );
  nand_x1_sg U45188 ( .A(n28363), .B(n28364), .X(\filter_0/n8847 ) );
  nand_x1_sg U45189 ( .A(n29977), .B(\filter_0/n7910 ), .X(n28364) );
  nand_x1_sg U45190 ( .A(n28367), .B(n28368), .X(\filter_0/n8846 ) );
  nand_x1_sg U45191 ( .A(n33447), .B(\filter_0/n7909 ), .X(n28368) );
  nand_x1_sg U45192 ( .A(n28369), .B(n28370), .X(\filter_0/n8845 ) );
  nand_x1_sg U45193 ( .A(n33446), .B(\filter_0/n7908 ), .X(n28370) );
  nand_x1_sg U45194 ( .A(n28371), .B(n28372), .X(\filter_0/n8844 ) );
  nand_x1_sg U45195 ( .A(n33445), .B(\filter_0/n7907 ), .X(n28372) );
  nand_x1_sg U45196 ( .A(n28576), .B(n28577), .X(\filter_0/n8747 ) );
  nand_x1_sg U45197 ( .A(n33382), .B(\filter_0/n7690 ), .X(n28577) );
  nand_x1_sg U45198 ( .A(n28580), .B(n28581), .X(\filter_0/n8746 ) );
  nand_x1_sg U45199 ( .A(n29951), .B(\filter_0/n7689 ), .X(n28581) );
  nand_x1_sg U45200 ( .A(n28582), .B(n28583), .X(\filter_0/n8745 ) );
  nand_x1_sg U45201 ( .A(n33380), .B(\filter_0/n7688 ), .X(n28583) );
  nand_x1_sg U45202 ( .A(n28584), .B(n28585), .X(\filter_0/n8744 ) );
  nand_x1_sg U45203 ( .A(n33380), .B(\filter_0/n7687 ), .X(n28585) );
  nand_x1_sg U45204 ( .A(n28746), .B(n28747), .X(\filter_0/n8667 ) );
  nand_x1_sg U45205 ( .A(n33378), .B(\filter_0/n7670 ), .X(n28747) );
  nand_x1_sg U45206 ( .A(n28750), .B(n28751), .X(\filter_0/n8666 ) );
  nand_x1_sg U45207 ( .A(n29949), .B(\filter_0/n7669 ), .X(n28751) );
  nand_x1_sg U45208 ( .A(n28752), .B(n28753), .X(\filter_0/n8665 ) );
  nand_x1_sg U45209 ( .A(n29949), .B(\filter_0/n7668 ), .X(n28753) );
  nand_x1_sg U45210 ( .A(n28754), .B(n28755), .X(\filter_0/n8664 ) );
  nand_x1_sg U45211 ( .A(n33376), .B(\filter_0/n7667 ), .X(n28755) );
  nand_x1_sg U45212 ( .A(n28330), .B(n28331), .X(\filter_0/n8863 ) );
  nand_x1_sg U45213 ( .A(n29945), .B(\filter_0/n7886 ), .X(n28331) );
  nand_x1_sg U45214 ( .A(n28332), .B(n28333), .X(\filter_0/n8862 ) );
  nand_x1_sg U45215 ( .A(n33367), .B(\filter_0/n7885 ), .X(n28333) );
  nand_x1_sg U45216 ( .A(n28286), .B(n28287), .X(\filter_0/n8883 ) );
  nand_x1_sg U45217 ( .A(n33351), .B(\filter_0/n7866 ), .X(n28287) );
  nand_x1_sg U45218 ( .A(n28288), .B(n28289), .X(\filter_0/n8882 ) );
  nand_x1_sg U45219 ( .A(n33350), .B(\filter_0/n7865 ), .X(n28289) );
  nand_x1_sg U45220 ( .A(n28502), .B(n28503), .X(\filter_0/n8783 ) );
  nand_x1_sg U45221 ( .A(n33470), .B(\filter_0/n7806 ), .X(n28503) );
  nand_x1_sg U45222 ( .A(n28504), .B(n28505), .X(\filter_0/n8782 ) );
  nand_x1_sg U45223 ( .A(n29987), .B(\filter_0/n7805 ), .X(n28505) );
  nand_x1_sg U45224 ( .A(n28460), .B(n28461), .X(\filter_0/n8803 ) );
  nand_x1_sg U45225 ( .A(n33348), .B(\filter_0/n7786 ), .X(n28461) );
  nand_x1_sg U45226 ( .A(n28462), .B(n28463), .X(\filter_0/n8802 ) );
  nand_x1_sg U45227 ( .A(n29937), .B(\filter_0/n7785 ), .X(n28463) );
  nand_x1_sg U45228 ( .A(n28629), .B(n28630), .X(\filter_0/n8723 ) );
  nand_x1_sg U45229 ( .A(n33362), .B(\filter_0/n7746 ), .X(n28630) );
  nand_x1_sg U45230 ( .A(n28631), .B(n28632), .X(\filter_0/n8722 ) );
  nand_x1_sg U45231 ( .A(n33362), .B(\filter_0/n7745 ), .X(n28632) );
  nand_x1_sg U45232 ( .A(n28671), .B(n28672), .X(\filter_0/n8703 ) );
  nand_x1_sg U45233 ( .A(n33340), .B(\filter_0/n7726 ), .X(n28672) );
  nand_x1_sg U45234 ( .A(n28673), .B(n28674), .X(\filter_0/n8702 ) );
  nand_x1_sg U45235 ( .A(n33341), .B(\filter_0/n7725 ), .X(n28674) );
  nand_x1_sg U45236 ( .A(n28801), .B(n28802), .X(\filter_0/n8643 ) );
  nand_x1_sg U45237 ( .A(n33357), .B(\filter_0/n7646 ), .X(n28802) );
  nand_x1_sg U45238 ( .A(n28803), .B(n28804), .X(\filter_0/n8642 ) );
  nand_x1_sg U45239 ( .A(n33355), .B(\filter_0/n7645 ), .X(n28804) );
  nand_x1_sg U45240 ( .A(n28845), .B(n28846), .X(\filter_0/n8623 ) );
  nand_x1_sg U45241 ( .A(n33337), .B(\filter_0/n7626 ), .X(n28846) );
  nand_x1_sg U45242 ( .A(n28847), .B(n28848), .X(\filter_0/n8622 ) );
  nand_x1_sg U45243 ( .A(n33336), .B(\filter_0/n7625 ), .X(n28848) );
  nand_x1_sg U45244 ( .A(n28556), .B(n28557), .X(\filter_0/n8757 ) );
  nand_x1_sg U45245 ( .A(n28568), .B(n28569), .X(\filter_0/n8751 ) );
  nand_x1_sg U45246 ( .A(n28552), .B(n28553), .X(\filter_0/n8759 ) );
  nand_x1_sg U45247 ( .A(n28564), .B(n28565), .X(\filter_0/n8753 ) );
  nand_x1_sg U45248 ( .A(n28548), .B(n28549), .X(\filter_0/n8761 ) );
  nand_x1_sg U45249 ( .A(n28560), .B(n28561), .X(\filter_0/n8755 ) );
  nand_x1_sg U45250 ( .A(n28572), .B(n28573), .X(\filter_0/n8749 ) );
  nand_x1_sg U45251 ( .A(n29418), .B(n29419), .X(\filter_0/n8356 ) );
  nand_x1_sg U45252 ( .A(n29430), .B(n29431), .X(\filter_0/n8350 ) );
  nand_x1_sg U45253 ( .A(n29442), .B(n29443), .X(\filter_0/n8344 ) );
  nand_x1_sg U45254 ( .A(n29594), .B(n29595), .X(\filter_0/n8276 ) );
  nand_x1_sg U45255 ( .A(n29606), .B(n29607), .X(\filter_0/n8270 ) );
  nand_x1_sg U45256 ( .A(n29618), .B(n29619), .X(\filter_0/n8264 ) );
  nand_x1_sg U45257 ( .A(n28719), .B(n28720), .X(\filter_0/n8680 ) );
  nand_x1_sg U45258 ( .A(n28731), .B(n28732), .X(\filter_0/n8674 ) );
  nand_x1_sg U45259 ( .A(n28743), .B(n28744), .X(\filter_0/n8668 ) );
  nand_x1_sg U45260 ( .A(n28895), .B(n28896), .X(\filter_0/n8600 ) );
  nand_x1_sg U45261 ( .A(n28907), .B(n28908), .X(\filter_0/n8594 ) );
  nand_x1_sg U45262 ( .A(n28919), .B(n28920), .X(\filter_0/n8588 ) );
  nand_x1_sg U45263 ( .A(n29426), .B(n29427), .X(\filter_0/n8352 ) );
  nand_x1_sg U45264 ( .A(n29438), .B(n29439), .X(\filter_0/n8346 ) );
  nand_x1_sg U45265 ( .A(n29602), .B(n29603), .X(\filter_0/n8272 ) );
  nand_x1_sg U45266 ( .A(n29614), .B(n29615), .X(\filter_0/n8266 ) );
  nand_x1_sg U45267 ( .A(n28727), .B(n28728), .X(\filter_0/n8676 ) );
  nand_x1_sg U45268 ( .A(n28739), .B(n28740), .X(\filter_0/n8670 ) );
  nand_x1_sg U45269 ( .A(n28903), .B(n28904), .X(\filter_0/n8596 ) );
  nand_x1_sg U45270 ( .A(n28915), .B(n28916), .X(\filter_0/n8590 ) );
  nand_x1_sg U45271 ( .A(n29422), .B(n29423), .X(\filter_0/n8354 ) );
  nand_x1_sg U45272 ( .A(n29434), .B(n29435), .X(\filter_0/n8348 ) );
  nand_x1_sg U45273 ( .A(n29598), .B(n29599), .X(\filter_0/n8274 ) );
  nand_x1_sg U45274 ( .A(n29610), .B(n29611), .X(\filter_0/n8268 ) );
  nand_x1_sg U45275 ( .A(n28723), .B(n28724), .X(\filter_0/n8678 ) );
  nand_x1_sg U45276 ( .A(n28735), .B(n28736), .X(\filter_0/n8672 ) );
  nand_x1_sg U45277 ( .A(n28899), .B(n28900), .X(\filter_0/n8598 ) );
  nand_x1_sg U45278 ( .A(n28911), .B(n28912), .X(\filter_0/n8592 ) );
  nand_x1_sg U45279 ( .A(n29412), .B(n29413), .X(\filter_0/n8359 ) );
  nand_x1_sg U45280 ( .A(n33332), .B(\filter_0/n8035 ), .X(n29413) );
  nand_x1_sg U45281 ( .A(n29588), .B(n29589), .X(\filter_0/n8279 ) );
  nand_x1_sg U45282 ( .A(n33325), .B(\filter_0/n7935 ), .X(n29589) );
  nand_x1_sg U45283 ( .A(n28713), .B(n28714), .X(\filter_0/n8683 ) );
  nand_x1_sg U45284 ( .A(n29947), .B(\filter_0/n7706 ), .X(n28714) );
  nand_x1_sg U45285 ( .A(n28889), .B(n28890), .X(\filter_0/n8603 ) );
  nand_x1_sg U45286 ( .A(n33322), .B(\filter_0/n7606 ), .X(n28890) );
  nand_x1_sg U45287 ( .A(n28320), .B(n28321), .X(\filter_0/n8867 ) );
  nand_x1_sg U45288 ( .A(n33368), .B(\filter_0/n7890 ), .X(n28321) );
  nand_x1_sg U45289 ( .A(n28324), .B(n28325), .X(\filter_0/n8866 ) );
  nand_x1_sg U45290 ( .A(n29945), .B(\filter_0/n7889 ), .X(n28325) );
  nand_x1_sg U45291 ( .A(n28326), .B(n28327), .X(\filter_0/n8865 ) );
  nand_x1_sg U45292 ( .A(n33365), .B(\filter_0/n7888 ), .X(n28327) );
  nand_x1_sg U45293 ( .A(n28328), .B(n28329), .X(\filter_0/n8864 ) );
  nand_x1_sg U45294 ( .A(n33368), .B(\filter_0/n7887 ), .X(n28329) );
  nand_x1_sg U45295 ( .A(n28276), .B(n28277), .X(\filter_0/n8887 ) );
  nand_x1_sg U45296 ( .A(n29939), .B(\filter_0/n7870 ), .X(n28277) );
  nand_x1_sg U45297 ( .A(n28280), .B(n28281), .X(\filter_0/n8886 ) );
  nand_x1_sg U45298 ( .A(n29939), .B(\filter_0/n7869 ), .X(n28281) );
  nand_x1_sg U45299 ( .A(n28282), .B(n28283), .X(\filter_0/n8885 ) );
  nand_x1_sg U45300 ( .A(n33350), .B(\filter_0/n7868 ), .X(n28283) );
  nand_x1_sg U45301 ( .A(n28284), .B(n28285), .X(\filter_0/n8884 ) );
  nand_x1_sg U45302 ( .A(n33352), .B(\filter_0/n7867 ), .X(n28285) );
  nand_x1_sg U45303 ( .A(n28492), .B(n28493), .X(\filter_0/n8787 ) );
  nand_x1_sg U45304 ( .A(n33472), .B(\filter_0/n7810 ), .X(n28493) );
  nand_x1_sg U45305 ( .A(n28496), .B(n28497), .X(\filter_0/n8786 ) );
  nand_x1_sg U45306 ( .A(n33473), .B(\filter_0/n7809 ), .X(n28497) );
  nand_x1_sg U45307 ( .A(n28498), .B(n28499), .X(\filter_0/n8785 ) );
  nand_x1_sg U45308 ( .A(n33471), .B(\filter_0/n7808 ), .X(n28499) );
  nand_x1_sg U45309 ( .A(n28500), .B(n28501), .X(\filter_0/n8784 ) );
  nand_x1_sg U45310 ( .A(n29987), .B(\filter_0/n7807 ), .X(n28501) );
  nand_x1_sg U45311 ( .A(n28450), .B(n28451), .X(\filter_0/n8807 ) );
  nand_x1_sg U45312 ( .A(n33346), .B(\filter_0/n7790 ), .X(n28451) );
  nand_x1_sg U45313 ( .A(n28454), .B(n28455), .X(\filter_0/n8806 ) );
  nand_x1_sg U45314 ( .A(n33348), .B(\filter_0/n7789 ), .X(n28455) );
  nand_x1_sg U45315 ( .A(n28456), .B(n28457), .X(\filter_0/n8805 ) );
  nand_x1_sg U45316 ( .A(n33346), .B(\filter_0/n7788 ), .X(n28457) );
  nand_x1_sg U45317 ( .A(n28458), .B(n28459), .X(\filter_0/n8804 ) );
  nand_x1_sg U45318 ( .A(n33347), .B(\filter_0/n7787 ), .X(n28459) );
  nand_x1_sg U45319 ( .A(n28619), .B(n28620), .X(\filter_0/n8727 ) );
  nand_x1_sg U45320 ( .A(n29943), .B(\filter_0/n7750 ), .X(n28620) );
  nand_x1_sg U45321 ( .A(n28623), .B(n28624), .X(\filter_0/n8726 ) );
  nand_x1_sg U45322 ( .A(n33361), .B(\filter_0/n7749 ), .X(n28624) );
  nand_x1_sg U45323 ( .A(n28625), .B(n28626), .X(\filter_0/n8725 ) );
  nand_x1_sg U45324 ( .A(n33361), .B(\filter_0/n7748 ), .X(n28626) );
  nand_x1_sg U45325 ( .A(n28627), .B(n28628), .X(\filter_0/n8724 ) );
  nand_x1_sg U45326 ( .A(n29943), .B(\filter_0/n7747 ), .X(n28628) );
  nand_x1_sg U45327 ( .A(n28661), .B(n28662), .X(\filter_0/n8707 ) );
  nand_x1_sg U45328 ( .A(n33343), .B(\filter_0/n7730 ), .X(n28662) );
  nand_x1_sg U45329 ( .A(n28665), .B(n28666), .X(\filter_0/n8706 ) );
  nand_x1_sg U45330 ( .A(n33341), .B(\filter_0/n7729 ), .X(n28666) );
  nand_x1_sg U45331 ( .A(n28667), .B(n28668), .X(\filter_0/n8705 ) );
  nand_x1_sg U45332 ( .A(n33342), .B(\filter_0/n7728 ), .X(n28668) );
  nand_x1_sg U45333 ( .A(n28669), .B(n28670), .X(\filter_0/n8704 ) );
  nand_x1_sg U45334 ( .A(n29935), .B(\filter_0/n7727 ), .X(n28670) );
  nand_x1_sg U45335 ( .A(n28791), .B(n28792), .X(\filter_0/n8647 ) );
  nand_x1_sg U45336 ( .A(n29941), .B(\filter_0/n7650 ), .X(n28792) );
  nand_x1_sg U45337 ( .A(n28795), .B(n28796), .X(\filter_0/n8646 ) );
  nand_x1_sg U45338 ( .A(n33358), .B(\filter_0/n7649 ), .X(n28796) );
  nand_x1_sg U45339 ( .A(n28797), .B(n28798), .X(\filter_0/n8645 ) );
  nand_x1_sg U45340 ( .A(n33356), .B(\filter_0/n7648 ), .X(n28798) );
  nand_x1_sg U45341 ( .A(n28799), .B(n28800), .X(\filter_0/n8644 ) );
  nand_x1_sg U45342 ( .A(n33357), .B(\filter_0/n7647 ), .X(n28800) );
  nand_x1_sg U45343 ( .A(n28835), .B(n28836), .X(\filter_0/n8627 ) );
  nand_x1_sg U45344 ( .A(n33338), .B(\filter_0/n7630 ), .X(n28836) );
  nand_x1_sg U45345 ( .A(n28839), .B(n28840), .X(\filter_0/n8626 ) );
  nand_x1_sg U45346 ( .A(n29933), .B(\filter_0/n7629 ), .X(n28840) );
  nand_x1_sg U45347 ( .A(n28841), .B(n28842), .X(\filter_0/n8625 ) );
  nand_x1_sg U45348 ( .A(n33336), .B(\filter_0/n7628 ), .X(n28842) );
  nand_x1_sg U45349 ( .A(n28843), .B(n28844), .X(\filter_0/n8624 ) );
  nand_x1_sg U45350 ( .A(n29933), .B(\filter_0/n7627 ), .X(n28844) );
  nand_x1_sg U45351 ( .A(n28550), .B(n28551), .X(\filter_0/n8760 ) );
  nand_x1_sg U45352 ( .A(n28562), .B(n28563), .X(\filter_0/n8754 ) );
  nand_x1_sg U45353 ( .A(n28574), .B(n28575), .X(\filter_0/n8748 ) );
  nand_x1_sg U45354 ( .A(n28558), .B(n28559), .X(\filter_0/n8756 ) );
  nand_x1_sg U45355 ( .A(n28570), .B(n28571), .X(\filter_0/n8750 ) );
  nand_x1_sg U45356 ( .A(n28554), .B(n28555), .X(\filter_0/n8758 ) );
  nand_x1_sg U45357 ( .A(n28566), .B(n28567), .X(\filter_0/n8752 ) );
  nand_x1_sg U45358 ( .A(n29402), .B(n29403), .X(\filter_0/n8363 ) );
  nand_x1_sg U45359 ( .A(n33330), .B(\filter_0/n8039 ), .X(n29403) );
  nand_x1_sg U45360 ( .A(n29408), .B(n29409), .X(\filter_0/n8361 ) );
  nand_x1_sg U45361 ( .A(n33330), .B(\filter_0/n8037 ), .X(n29409) );
  nand_x1_sg U45362 ( .A(n29578), .B(n29579), .X(\filter_0/n8283 ) );
  nand_x1_sg U45363 ( .A(n33326), .B(\filter_0/n7939 ), .X(n29579) );
  nand_x1_sg U45364 ( .A(n29584), .B(n29585), .X(\filter_0/n8281 ) );
  nand_x1_sg U45365 ( .A(n29929), .B(\filter_0/n7937 ), .X(n29585) );
  nand_x1_sg U45366 ( .A(n28703), .B(n28704), .X(\filter_0/n8687 ) );
  nand_x1_sg U45367 ( .A(n33372), .B(\filter_0/n7710 ), .X(n28704) );
  nand_x1_sg U45368 ( .A(n28709), .B(n28710), .X(\filter_0/n8685 ) );
  nand_x1_sg U45369 ( .A(n33371), .B(\filter_0/n7708 ), .X(n28710) );
  nand_x1_sg U45370 ( .A(n28879), .B(n28880), .X(\filter_0/n8607 ) );
  nand_x1_sg U45371 ( .A(n33323), .B(\filter_0/n7610 ), .X(n28880) );
  nand_x1_sg U45372 ( .A(n28885), .B(n28886), .X(\filter_0/n8605 ) );
  nand_x1_sg U45373 ( .A(n29927), .B(\filter_0/n7608 ), .X(n28886) );
  nand_x1_sg U45374 ( .A(n28544), .B(n28545), .X(\filter_0/n8763 ) );
  nand_x1_sg U45375 ( .A(n33431), .B(\filter_0/n7826 ), .X(n28545) );
  nand_x1_sg U45376 ( .A(n29414), .B(n29415), .X(\filter_0/n8358 ) );
  nand_x1_sg U45377 ( .A(n29931), .B(\filter_0/n8034 ), .X(n29415) );
  nand_x1_sg U45378 ( .A(n29590), .B(n29591), .X(\filter_0/n8278 ) );
  nand_x1_sg U45379 ( .A(n33328), .B(\filter_0/n7934 ), .X(n29591) );
  nand_x1_sg U45380 ( .A(n28715), .B(n28716), .X(\filter_0/n8682 ) );
  nand_x1_sg U45381 ( .A(n33370), .B(\filter_0/n7705 ), .X(n28716) );
  nand_x1_sg U45382 ( .A(n28891), .B(n28892), .X(\filter_0/n8602 ) );
  nand_x1_sg U45383 ( .A(n29927), .B(\filter_0/n7605 ), .X(n28892) );
  nand_x1_sg U45384 ( .A(n28534), .B(n28535), .X(\filter_0/n8767 ) );
  nand_x1_sg U45385 ( .A(n33430), .B(\filter_0/n7830 ), .X(n28535) );
  nand_x1_sg U45386 ( .A(n28540), .B(n28541), .X(\filter_0/n8765 ) );
  nand_x1_sg U45387 ( .A(n33430), .B(\filter_0/n7828 ), .X(n28541) );
  nand_x1_sg U45388 ( .A(n29406), .B(n29407), .X(\filter_0/n8362 ) );
  nand_x1_sg U45389 ( .A(n33333), .B(\filter_0/n8038 ), .X(n29407) );
  nand_x1_sg U45390 ( .A(n29582), .B(n29583), .X(\filter_0/n8282 ) );
  nand_x1_sg U45391 ( .A(n29929), .B(\filter_0/n7938 ), .X(n29583) );
  nand_x1_sg U45392 ( .A(n28707), .B(n28708), .X(\filter_0/n8686 ) );
  nand_x1_sg U45393 ( .A(n29947), .B(\filter_0/n7709 ), .X(n28708) );
  nand_x1_sg U45394 ( .A(n28883), .B(n28884), .X(\filter_0/n8606 ) );
  nand_x1_sg U45395 ( .A(n33321), .B(\filter_0/n7609 ), .X(n28884) );
  nand_x1_sg U45396 ( .A(n28546), .B(n28547), .X(\filter_0/n8762 ) );
  nand_x1_sg U45397 ( .A(n29971), .B(\filter_0/n7825 ), .X(n28547) );
  nand_x1_sg U45398 ( .A(n29410), .B(n29411), .X(\filter_0/n8360 ) );
  nand_x1_sg U45399 ( .A(n29931), .B(\filter_0/n8036 ), .X(n29411) );
  nand_x1_sg U45400 ( .A(n29586), .B(n29587), .X(\filter_0/n8280 ) );
  nand_x1_sg U45401 ( .A(n33328), .B(\filter_0/n7936 ), .X(n29587) );
  nand_x1_sg U45402 ( .A(n28711), .B(n28712), .X(\filter_0/n8684 ) );
  nand_x1_sg U45403 ( .A(n33372), .B(\filter_0/n7707 ), .X(n28712) );
  nand_x1_sg U45404 ( .A(n28887), .B(n28888), .X(\filter_0/n8604 ) );
  nand_x1_sg U45405 ( .A(n29927), .B(\filter_0/n7607 ), .X(n28888) );
  nand_x1_sg U45406 ( .A(n28538), .B(n28539), .X(\filter_0/n8766 ) );
  nand_x1_sg U45407 ( .A(n33431), .B(\filter_0/n7829 ), .X(n28539) );
  nand_x1_sg U45408 ( .A(n28542), .B(n28543), .X(\filter_0/n8764 ) );
  nand_x1_sg U45409 ( .A(n33432), .B(\filter_0/n7827 ), .X(n28543) );
  nand_x1_sg U45410 ( .A(n28145), .B(n28146), .X(\filter_0/n8918 ) );
  nand_x1_sg U45411 ( .A(n28140), .B(n28141), .X(\filter_0/n8919 ) );
  nand_x1_sg U45412 ( .A(n28135), .B(n28136), .X(\filter_0/n8920 ) );
  nand_x1_sg U45413 ( .A(n28130), .B(n28131), .X(\filter_0/n8921 ) );
  nand_x1_sg U45414 ( .A(n28125), .B(n28126), .X(\filter_0/n8922 ) );
  nand_x1_sg U45415 ( .A(n28120), .B(n28121), .X(\filter_0/n8923 ) );
  nand_x1_sg U45416 ( .A(n28115), .B(n28116), .X(\filter_0/n8924 ) );
  nand_x1_sg U45417 ( .A(n28110), .B(n28111), .X(\filter_0/n8925 ) );
  nand_x1_sg U45418 ( .A(n28105), .B(n28106), .X(\filter_0/n8926 ) );
  nand_x1_sg U45419 ( .A(n28100), .B(n28101), .X(\filter_0/n8927 ) );
  nand_x1_sg U45420 ( .A(n28095), .B(n28096), .X(\filter_0/n8928 ) );
  nand_x1_sg U45421 ( .A(n28090), .B(n28091), .X(\filter_0/n8929 ) );
  nand_x1_sg U45422 ( .A(n28085), .B(n28086), .X(\filter_0/n8930 ) );
  nand_x1_sg U45423 ( .A(n28080), .B(n28081), .X(\filter_0/n8931 ) );
  nand_x1_sg U45424 ( .A(n28075), .B(n28076), .X(\filter_0/n8932 ) );
  nand_x1_sg U45425 ( .A(n28070), .B(n28071), .X(\filter_0/n8933 ) );
  nand_x1_sg U45426 ( .A(n28065), .B(n28066), .X(\filter_0/n8934 ) );
  nand_x1_sg U45427 ( .A(n28060), .B(n28061), .X(\filter_0/n8935 ) );
  nand_x1_sg U45428 ( .A(n28055), .B(n28056), .X(\filter_0/n8936 ) );
  nand_x1_sg U45429 ( .A(n28050), .B(n28051), .X(\filter_0/n8937 ) );
  nand_x1_sg U45430 ( .A(n28045), .B(n28046), .X(\filter_0/n8938 ) );
  nand_x1_sg U45431 ( .A(n28030), .B(n28031), .X(\filter_0/n8941 ) );
  nand_x1_sg U45432 ( .A(n28025), .B(n28026), .X(\filter_0/n8942 ) );
  nand_x1_sg U45433 ( .A(n28020), .B(n28021), .X(\filter_0/n8943 ) );
  nand_x1_sg U45434 ( .A(n28015), .B(n28016), .X(\filter_0/n8944 ) );
  nand_x1_sg U45435 ( .A(n28010), .B(n28011), .X(\filter_0/n8945 ) );
  nand_x1_sg U45436 ( .A(n28005), .B(n28006), .X(\filter_0/n8946 ) );
  nand_x1_sg U45437 ( .A(n28000), .B(n28001), .X(\filter_0/n8947 ) );
  nand_x1_sg U45438 ( .A(n27995), .B(n27996), .X(\filter_0/n8948 ) );
  nand_x1_sg U45439 ( .A(n27990), .B(n27991), .X(\filter_0/n8949 ) );
  nand_x1_sg U45440 ( .A(n27985), .B(n27986), .X(\filter_0/n8950 ) );
  nand_x1_sg U45441 ( .A(n27980), .B(n27981), .X(\filter_0/n8951 ) );
  nand_x1_sg U45442 ( .A(n27975), .B(n27976), .X(\filter_0/n8952 ) );
  nand_x1_sg U45443 ( .A(n27970), .B(n27971), .X(\filter_0/n8953 ) );
  nand_x1_sg U45444 ( .A(n27965), .B(n27966), .X(\filter_0/n8954 ) );
  nand_x1_sg U45445 ( .A(n27960), .B(n27961), .X(\filter_0/n8955 ) );
  nand_x1_sg U45446 ( .A(n27955), .B(n27956), .X(\filter_0/n8956 ) );
  nand_x1_sg U45447 ( .A(n27950), .B(n27951), .X(\filter_0/n8957 ) );
  nand_x1_sg U45448 ( .A(n27945), .B(n27946), .X(\filter_0/n8958 ) );
  nand_x1_sg U45449 ( .A(n28250), .B(n28251), .X(\filter_0/n8897 ) );
  nand_x1_sg U45450 ( .A(n27893), .B(n27894), .X(\filter_0/n8981 ) );
  nand_x1_sg U45451 ( .A(n27887), .B(n27888), .X(\filter_0/n8984 ) );
  nand_x1_sg U45452 ( .A(n27881), .B(n27882), .X(\filter_0/n8987 ) );
  nand_x1_sg U45453 ( .A(n27875), .B(n27876), .X(\filter_0/n8990 ) );
  nand_x1_sg U45454 ( .A(n27869), .B(n27870), .X(\filter_0/n8993 ) );
  nand_x1_sg U45455 ( .A(n27863), .B(n27864), .X(\filter_0/n8996 ) );
  nand_x1_sg U45456 ( .A(n27857), .B(n27858), .X(\filter_0/n8999 ) );
  nand_x1_sg U45457 ( .A(n27851), .B(n27852), .X(\filter_0/n9002 ) );
  nand_x1_sg U45458 ( .A(n27809), .B(n27810), .X(\filter_0/n9023 ) );
  nand_x1_sg U45459 ( .A(n27803), .B(n27804), .X(\filter_0/n9026 ) );
  nand_x1_sg U45460 ( .A(n27797), .B(n27798), .X(\filter_0/n9029 ) );
  nand_x1_sg U45461 ( .A(n27791), .B(n27792), .X(\filter_0/n9032 ) );
  nand_x1_sg U45462 ( .A(n27785), .B(n27786), .X(\filter_0/n9035 ) );
  nand_x1_sg U45463 ( .A(n27779), .B(n27780), .X(\filter_0/n9038 ) );
  nand_x1_sg U45464 ( .A(n27773), .B(n27774), .X(\filter_0/n9041 ) );
  nand_x1_sg U45465 ( .A(n27731), .B(n27732), .X(\filter_0/n9062 ) );
  nand_x1_sg U45466 ( .A(n27725), .B(n27726), .X(\filter_0/n9065 ) );
  nand_x1_sg U45467 ( .A(n27719), .B(n27720), .X(\filter_0/n9068 ) );
  nand_x1_sg U45468 ( .A(n27713), .B(n27714), .X(\filter_0/n9071 ) );
  nand_x1_sg U45469 ( .A(n27707), .B(n27708), .X(\filter_0/n9074 ) );
  nand_x1_sg U45470 ( .A(n27701), .B(n27702), .X(\filter_0/n9077 ) );
  nand_x1_sg U45471 ( .A(n27695), .B(n27696), .X(\filter_0/n9080 ) );
  nand_x1_sg U45472 ( .A(n27689), .B(n27690), .X(\filter_0/n9083 ) );
  nand_x1_sg U45473 ( .A(n27683), .B(n27684), .X(\filter_0/n9086 ) );
  nand_x1_sg U45474 ( .A(n27677), .B(n27678), .X(\filter_0/n9089 ) );
  nand_x1_sg U45475 ( .A(n27671), .B(n27672), .X(\filter_0/n9092 ) );
  nand_x1_sg U45476 ( .A(n27665), .B(n27666), .X(\filter_0/n9095 ) );
  nand_x1_sg U45477 ( .A(n27659), .B(n27660), .X(\filter_0/n9098 ) );
  nand_x1_sg U45478 ( .A(n27653), .B(n27654), .X(\filter_0/n9101 ) );
  nand_x1_sg U45479 ( .A(n27647), .B(n27648), .X(\filter_0/n9104 ) );
  nand_x1_sg U45480 ( .A(n27641), .B(n27642), .X(\filter_0/n9107 ) );
  nand_x1_sg U45481 ( .A(n27635), .B(n27636), .X(\filter_0/n9110 ) );
  nand_x1_sg U45482 ( .A(n27629), .B(n27630), .X(\filter_0/n9113 ) );
  nand_x1_sg U45483 ( .A(n27623), .B(n27624), .X(\filter_0/n9116 ) );
  nand_x1_sg U45484 ( .A(n27617), .B(n27618), .X(\filter_0/n9119 ) );
  nand_x1_sg U45485 ( .A(n27611), .B(n27612), .X(\filter_0/n9122 ) );
  nand_x1_sg U45486 ( .A(n27593), .B(n27594), .X(\filter_0/n9131 ) );
  nand_x1_sg U45487 ( .A(n27587), .B(n27588), .X(\filter_0/n9134 ) );
  nand_x1_sg U45488 ( .A(n27581), .B(n27582), .X(\filter_0/n9137 ) );
  nand_x1_sg U45489 ( .A(n27575), .B(n27576), .X(\filter_0/n9140 ) );
  nand_x1_sg U45490 ( .A(n27569), .B(n27570), .X(\filter_0/n9143 ) );
  nand_x1_sg U45491 ( .A(n27563), .B(n27564), .X(\filter_0/n9146 ) );
  nand_x1_sg U45492 ( .A(n27527), .B(n27528), .X(\filter_0/n9164 ) );
  nand_x1_sg U45493 ( .A(n27521), .B(n27522), .X(\filter_0/n9167 ) );
  nand_x1_sg U45494 ( .A(n27515), .B(n27516), .X(\filter_0/n9170 ) );
  nand_x1_sg U45495 ( .A(n27509), .B(n27510), .X(\filter_0/n9173 ) );
  nand_x1_sg U45496 ( .A(n27503), .B(n27504), .X(\filter_0/n9176 ) );
  nand_x1_sg U45497 ( .A(n27497), .B(n27498), .X(\filter_0/n9179 ) );
  nand_x1_sg U45498 ( .A(n27491), .B(n27492), .X(\filter_0/n9182 ) );
  nand_x1_sg U45499 ( .A(n27485), .B(n27486), .X(\filter_0/n9185 ) );
  nand_x1_sg U45500 ( .A(n27479), .B(n27480), .X(\filter_0/n9188 ) );
  nand_x1_sg U45501 ( .A(n27473), .B(n27474), .X(\filter_0/n9191 ) );
  nand_x1_sg U45502 ( .A(n27467), .B(n27468), .X(\filter_0/n9194 ) );
  nand_x1_sg U45503 ( .A(n27461), .B(n27462), .X(\filter_0/n9197 ) );
  nand_x1_sg U45504 ( .A(n27431), .B(n27432), .X(\filter_0/n9212 ) );
  nand_x1_sg U45505 ( .A(n27425), .B(n27426), .X(\filter_0/n9215 ) );
  nand_x1_sg U45506 ( .A(n27419), .B(n27420), .X(\filter_0/n9218 ) );
  nand_x1_sg U45507 ( .A(n27413), .B(n27414), .X(\filter_0/n9221 ) );
  nand_x1_sg U45508 ( .A(n27407), .B(n27408), .X(\filter_0/n9224 ) );
  nand_x1_sg U45509 ( .A(n27365), .B(n27366), .X(\filter_0/n9245 ) );
  nand_x1_sg U45510 ( .A(n27359), .B(n27360), .X(\filter_0/n9248 ) );
  nand_x1_sg U45511 ( .A(n27353), .B(n27354), .X(\filter_0/n9251 ) );
  nand_x1_sg U45512 ( .A(n27347), .B(n27348), .X(\filter_0/n9254 ) );
  nand_x1_sg U45513 ( .A(n27329), .B(n27330), .X(\filter_0/n9263 ) );
  nand_x1_sg U45514 ( .A(n27323), .B(n27324), .X(\filter_0/n9266 ) );
  nand_x1_sg U45515 ( .A(n27317), .B(n27318), .X(\filter_0/n9269 ) );
  nand_x1_sg U45516 ( .A(n27311), .B(n27312), .X(\filter_0/n9272 ) );
  nand_x1_sg U45517 ( .A(n27305), .B(n27306), .X(\filter_0/n9275 ) );
  nand_x1_sg U45518 ( .A(n27299), .B(n27300), .X(\filter_0/n9278 ) );
  nand_x1_sg U45519 ( .A(n27293), .B(n27294), .X(\filter_0/n9281 ) );
  nand_x1_sg U45520 ( .A(n27287), .B(n27288), .X(\filter_0/n9284 ) );
  nand_x1_sg U45521 ( .A(n27281), .B(n27282), .X(\filter_0/n9287 ) );
  nand_x1_sg U45522 ( .A(n27275), .B(n27276), .X(\filter_0/n9290 ) );
  nand_x1_sg U45523 ( .A(n27269), .B(n27270), .X(\filter_0/n9293 ) );
  nand_x1_sg U45524 ( .A(n27263), .B(n27264), .X(\filter_0/n9296 ) );
  nand_x1_sg U45525 ( .A(n27257), .B(n27258), .X(\filter_0/n9299 ) );
  nand_x1_sg U45526 ( .A(n27251), .B(n27252), .X(\filter_0/n9302 ) );
  nand_x1_sg U45527 ( .A(n27245), .B(n27246), .X(\filter_0/n9305 ) );
  nand_x1_sg U45528 ( .A(n27215), .B(n27216), .X(\filter_0/n9320 ) );
  nand_x1_sg U45529 ( .A(n27209), .B(n27210), .X(\filter_0/n9323 ) );
  nand_x1_sg U45530 ( .A(n27203), .B(n27204), .X(\filter_0/n9326 ) );
  nand_x1_sg U45531 ( .A(n27197), .B(n27198), .X(\filter_0/n9329 ) );
  nand_x1_sg U45532 ( .A(n27191), .B(n27192), .X(\filter_0/n9332 ) );
  nand_x1_sg U45533 ( .A(n27185), .B(n27186), .X(\filter_0/n9335 ) );
  nand_x1_sg U45534 ( .A(n27161), .B(n27162), .X(\filter_0/n9347 ) );
  nand_x1_sg U45535 ( .A(n27155), .B(n27156), .X(\filter_0/n9350 ) );
  nand_x1_sg U45536 ( .A(n27149), .B(n27150), .X(\filter_0/n9353 ) );
  nand_x1_sg U45537 ( .A(n27143), .B(n27144), .X(\filter_0/n9356 ) );
  nand_x1_sg U45538 ( .A(n27137), .B(n27138), .X(\filter_0/n9359 ) );
  nand_x1_sg U45539 ( .A(n27131), .B(n27132), .X(\filter_0/n9362 ) );
  nand_x1_sg U45540 ( .A(n27125), .B(n27126), .X(\filter_0/n9365 ) );
  nand_x1_sg U45541 ( .A(n27119), .B(n27120), .X(\filter_0/n9368 ) );
  nand_x1_sg U45542 ( .A(n27113), .B(n27114), .X(\filter_0/n9371 ) );
  nand_x1_sg U45543 ( .A(n27107), .B(n27108), .X(\filter_0/n9374 ) );
  nand_x1_sg U45544 ( .A(n27101), .B(n27102), .X(\filter_0/n9377 ) );
  nand_x1_sg U45545 ( .A(n27095), .B(n27096), .X(\filter_0/n9380 ) );
  nand_x1_sg U45546 ( .A(n27089), .B(n27090), .X(\filter_0/n9383 ) );
  nand_x1_sg U45547 ( .A(n27083), .B(n27084), .X(\filter_0/n9386 ) );
  nand_x1_sg U45548 ( .A(n27077), .B(n27078), .X(\filter_0/n9389 ) );
  nand_x1_sg U45549 ( .A(n27071), .B(n27072), .X(\filter_0/n9392 ) );
  nand_x1_sg U45550 ( .A(n27053), .B(n27054), .X(\filter_0/n9401 ) );
  nand_x1_sg U45551 ( .A(n27047), .B(n27048), .X(\filter_0/n9404 ) );
  nand_x1_sg U45552 ( .A(n27041), .B(n27042), .X(\filter_0/n9407 ) );
  nand_x1_sg U45553 ( .A(n26999), .B(n27000), .X(\filter_0/n9428 ) );
  nand_x1_sg U45554 ( .A(n26993), .B(n26994), .X(\filter_0/n9431 ) );
  nand_x1_sg U45555 ( .A(n26987), .B(n26988), .X(\filter_0/n9434 ) );
  nand_x1_sg U45556 ( .A(n26981), .B(n26982), .X(\filter_0/n9437 ) );
  nand_x1_sg U45557 ( .A(n26975), .B(n26976), .X(\filter_0/n9440 ) );
  nand_x1_sg U45558 ( .A(n26969), .B(n26970), .X(\filter_0/n9443 ) );
  nand_x1_sg U45559 ( .A(n26939), .B(n26940), .X(\filter_0/n9458 ) );
  nand_x1_sg U45560 ( .A(n26933), .B(n26934), .X(\filter_0/n9461 ) );
  nand_x1_sg U45561 ( .A(n26927), .B(n26928), .X(\filter_0/n9464 ) );
  nand_x1_sg U45562 ( .A(n26921), .B(n26922), .X(\filter_0/n9467 ) );
  nand_x1_sg U45563 ( .A(n26915), .B(n26916), .X(\filter_0/n9470 ) );
  nand_x1_sg U45564 ( .A(n26909), .B(n26910), .X(\filter_0/n9473 ) );
  nand_x1_sg U45565 ( .A(n26903), .B(n26904), .X(\filter_0/n9476 ) );
  nand_x1_sg U45566 ( .A(n26897), .B(n26898), .X(\filter_0/n9479 ) );
  nand_x1_sg U45567 ( .A(n26891), .B(n26892), .X(\filter_0/n9482 ) );
  nand_x1_sg U45568 ( .A(n26885), .B(n26886), .X(\filter_0/n9485 ) );
  nand_x1_sg U45569 ( .A(n26879), .B(n26880), .X(\filter_0/n9488 ) );
  nand_x1_sg U45570 ( .A(n26837), .B(n26838), .X(\filter_0/n9509 ) );
  nand_x1_sg U45571 ( .A(n26831), .B(n26832), .X(\filter_0/n9512 ) );
  nand_x1_sg U45572 ( .A(n26825), .B(n26826), .X(\filter_0/n9515 ) );
  nand_x1_sg U45573 ( .A(n26819), .B(n26820), .X(\filter_0/n9518 ) );
  nand_x1_sg U45574 ( .A(n26813), .B(n26814), .X(\filter_0/n9521 ) );
  nand_x1_sg U45575 ( .A(n26807), .B(n26808), .X(\filter_0/n9524 ) );
  nand_x1_sg U45576 ( .A(n26795), .B(n26796), .X(\filter_0/n9530 ) );
  nand_x1_sg U45577 ( .A(n26789), .B(n26790), .X(\filter_0/n9533 ) );
  nand_x1_sg U45578 ( .A(n26783), .B(n26784), .X(\filter_0/n9536 ) );
  nand_x1_sg U45579 ( .A(n26777), .B(n26778), .X(\filter_0/n9539 ) );
  nand_x1_sg U45580 ( .A(n26771), .B(n26772), .X(\filter_0/n9542 ) );
  nand_x1_sg U45581 ( .A(n26765), .B(n26766), .X(\filter_0/n9545 ) );
  nand_x1_sg U45582 ( .A(n26759), .B(n26760), .X(\filter_0/n9548 ) );
  nand_x1_sg U45583 ( .A(n26753), .B(n26754), .X(\filter_0/n9551 ) );
  nand_x1_sg U45584 ( .A(n26747), .B(n26748), .X(\filter_0/n9554 ) );
  nand_x1_sg U45585 ( .A(n26741), .B(n26742), .X(\filter_0/n9557 ) );
  nand_x1_sg U45586 ( .A(n26735), .B(n26736), .X(\filter_0/n9560 ) );
  nand_x1_sg U45587 ( .A(n26729), .B(n26730), .X(\filter_0/n9563 ) );
  nand_x1_sg U45588 ( .A(n26723), .B(n26724), .X(\filter_0/n9566 ) );
  nand_x1_sg U45589 ( .A(n26717), .B(n26718), .X(\filter_0/n9569 ) );
  nand_x1_sg U45590 ( .A(n26711), .B(n26712), .X(\filter_0/n9572 ) );
  nand_x1_sg U45591 ( .A(n26705), .B(n26706), .X(\filter_0/n9575 ) );
  nand_x1_sg U45592 ( .A(n26699), .B(n26700), .X(\filter_0/n9578 ) );
  nand_x1_sg U45593 ( .A(n26693), .B(n26694), .X(\filter_0/n9581 ) );
  nand_x1_sg U45594 ( .A(n26687), .B(n26688), .X(\filter_0/n9584 ) );
  nand_x1_sg U45595 ( .A(n26681), .B(n26682), .X(\filter_0/n9587 ) );
  nand_x1_sg U45596 ( .A(n26675), .B(n26676), .X(\filter_0/n9590 ) );
  nand_x1_sg U45597 ( .A(n26633), .B(n26634), .X(\filter_0/n9611 ) );
  nand_x1_sg U45598 ( .A(n26627), .B(n26628), .X(\filter_0/n9614 ) );
  nand_x1_sg U45599 ( .A(n26621), .B(n26622), .X(\filter_0/n9617 ) );
  nand_x1_sg U45600 ( .A(n26615), .B(n26616), .X(\filter_0/n9620 ) );
  nand_x1_sg U45601 ( .A(n26609), .B(n26610), .X(\filter_0/n9623 ) );
  nand_x1_sg U45602 ( .A(n26603), .B(n26604), .X(\filter_0/n9626 ) );
  nand_x1_sg U45603 ( .A(n26597), .B(n26598), .X(\filter_0/n9629 ) );
  nand_x1_sg U45604 ( .A(n26591), .B(n26592), .X(\filter_0/n9632 ) );
  nand_x1_sg U45605 ( .A(n28245), .B(n28246), .X(\filter_0/n8898 ) );
  nand_x1_sg U45606 ( .A(n28240), .B(n28241), .X(\filter_0/n8899 ) );
  nand_x1_sg U45607 ( .A(n27897), .B(n27898), .X(\filter_0/n8979 ) );
  nand_x1_sg U45608 ( .A(n27895), .B(n27896), .X(\filter_0/n8980 ) );
  nand_x1_sg U45609 ( .A(n27891), .B(n27892), .X(\filter_0/n8982 ) );
  nand_x1_sg U45610 ( .A(n27889), .B(n27890), .X(\filter_0/n8983 ) );
  nand_x1_sg U45611 ( .A(n27885), .B(n27886), .X(\filter_0/n8985 ) );
  nand_x1_sg U45612 ( .A(n27883), .B(n27884), .X(\filter_0/n8986 ) );
  nand_x1_sg U45613 ( .A(n27879), .B(n27880), .X(\filter_0/n8988 ) );
  nand_x1_sg U45614 ( .A(n27877), .B(n27878), .X(\filter_0/n8989 ) );
  nand_x1_sg U45615 ( .A(n27873), .B(n27874), .X(\filter_0/n8991 ) );
  nand_x1_sg U45616 ( .A(n27871), .B(n27872), .X(\filter_0/n8992 ) );
  nand_x1_sg U45617 ( .A(n27867), .B(n27868), .X(\filter_0/n8994 ) );
  nand_x1_sg U45618 ( .A(n27865), .B(n27866), .X(\filter_0/n8995 ) );
  nand_x1_sg U45619 ( .A(n27861), .B(n27862), .X(\filter_0/n8997 ) );
  nand_x1_sg U45620 ( .A(n27859), .B(n27860), .X(\filter_0/n8998 ) );
  nand_x1_sg U45621 ( .A(n27855), .B(n27856), .X(\filter_0/n9000 ) );
  nand_x1_sg U45622 ( .A(n27853), .B(n27854), .X(\filter_0/n9001 ) );
  nand_x1_sg U45623 ( .A(n27849), .B(n27850), .X(\filter_0/n9003 ) );
  nand_x1_sg U45624 ( .A(n27847), .B(n27848), .X(\filter_0/n9004 ) );
  nand_x1_sg U45625 ( .A(n27807), .B(n27808), .X(\filter_0/n9024 ) );
  nand_x1_sg U45626 ( .A(n27805), .B(n27806), .X(\filter_0/n9025 ) );
  nand_x1_sg U45627 ( .A(n27801), .B(n27802), .X(\filter_0/n9027 ) );
  nand_x1_sg U45628 ( .A(n27799), .B(n27800), .X(\filter_0/n9028 ) );
  nand_x1_sg U45629 ( .A(n27795), .B(n27796), .X(\filter_0/n9030 ) );
  nand_x1_sg U45630 ( .A(n27793), .B(n27794), .X(\filter_0/n9031 ) );
  nand_x1_sg U45631 ( .A(n27789), .B(n27790), .X(\filter_0/n9033 ) );
  nand_x1_sg U45632 ( .A(n27787), .B(n27788), .X(\filter_0/n9034 ) );
  nand_x1_sg U45633 ( .A(n27783), .B(n27784), .X(\filter_0/n9036 ) );
  nand_x1_sg U45634 ( .A(n27781), .B(n27782), .X(\filter_0/n9037 ) );
  nand_x1_sg U45635 ( .A(n27777), .B(n27778), .X(\filter_0/n9039 ) );
  nand_x1_sg U45636 ( .A(n27775), .B(n27776), .X(\filter_0/n9040 ) );
  nand_x1_sg U45637 ( .A(n27733), .B(n27734), .X(\filter_0/n9061 ) );
  nand_x1_sg U45638 ( .A(n27729), .B(n27730), .X(\filter_0/n9063 ) );
  nand_x1_sg U45639 ( .A(n27727), .B(n27728), .X(\filter_0/n9064 ) );
  nand_x1_sg U45640 ( .A(n27723), .B(n27724), .X(\filter_0/n9066 ) );
  nand_x1_sg U45641 ( .A(n27717), .B(n27718), .X(\filter_0/n9069 ) );
  nand_x1_sg U45642 ( .A(n27715), .B(n27716), .X(\filter_0/n9070 ) );
  nand_x1_sg U45643 ( .A(n27711), .B(n27712), .X(\filter_0/n9072 ) );
  nand_x1_sg U45644 ( .A(n27709), .B(n27710), .X(\filter_0/n9073 ) );
  nand_x1_sg U45645 ( .A(n27705), .B(n27706), .X(\filter_0/n9075 ) );
  nand_x1_sg U45646 ( .A(n27703), .B(n27704), .X(\filter_0/n9076 ) );
  nand_x1_sg U45647 ( .A(n27699), .B(n27700), .X(\filter_0/n9078 ) );
  nand_x1_sg U45648 ( .A(n27697), .B(n27698), .X(\filter_0/n9079 ) );
  nand_x1_sg U45649 ( .A(n27693), .B(n27694), .X(\filter_0/n9081 ) );
  nand_x1_sg U45650 ( .A(n27691), .B(n27692), .X(\filter_0/n9082 ) );
  nand_x1_sg U45651 ( .A(n27687), .B(n27688), .X(\filter_0/n9084 ) );
  nand_x1_sg U45652 ( .A(n27685), .B(n27686), .X(\filter_0/n9085 ) );
  nand_x1_sg U45653 ( .A(n27681), .B(n27682), .X(\filter_0/n9087 ) );
  nand_x1_sg U45654 ( .A(n27679), .B(n27680), .X(\filter_0/n9088 ) );
  nand_x1_sg U45655 ( .A(n27675), .B(n27676), .X(\filter_0/n9090 ) );
  nand_x1_sg U45656 ( .A(n27673), .B(n27674), .X(\filter_0/n9091 ) );
  nand_x1_sg U45657 ( .A(n27669), .B(n27670), .X(\filter_0/n9093 ) );
  nand_x1_sg U45658 ( .A(n27667), .B(n27668), .X(\filter_0/n9094 ) );
  nand_x1_sg U45659 ( .A(n27663), .B(n27664), .X(\filter_0/n9096 ) );
  nand_x1_sg U45660 ( .A(n27661), .B(n27662), .X(\filter_0/n9097 ) );
  nand_x1_sg U45661 ( .A(n27657), .B(n27658), .X(\filter_0/n9099 ) );
  nand_x1_sg U45662 ( .A(n27655), .B(n27656), .X(\filter_0/n9100 ) );
  nand_x1_sg U45663 ( .A(n27651), .B(n27652), .X(\filter_0/n9102 ) );
  nand_x1_sg U45664 ( .A(n27649), .B(n27650), .X(\filter_0/n9103 ) );
  nand_x1_sg U45665 ( .A(n27645), .B(n27646), .X(\filter_0/n9105 ) );
  nand_x1_sg U45666 ( .A(n27643), .B(n27644), .X(\filter_0/n9106 ) );
  nand_x1_sg U45667 ( .A(n27639), .B(n27640), .X(\filter_0/n9108 ) );
  nand_x1_sg U45668 ( .A(n27637), .B(n27638), .X(\filter_0/n9109 ) );
  nand_x1_sg U45669 ( .A(n27633), .B(n27634), .X(\filter_0/n9111 ) );
  nand_x1_sg U45670 ( .A(n27631), .B(n27632), .X(\filter_0/n9112 ) );
  nand_x1_sg U45671 ( .A(n27627), .B(n27628), .X(\filter_0/n9114 ) );
  nand_x1_sg U45672 ( .A(n27625), .B(n27626), .X(\filter_0/n9115 ) );
  nand_x1_sg U45673 ( .A(n27621), .B(n27622), .X(\filter_0/n9117 ) );
  nand_x1_sg U45674 ( .A(n27619), .B(n27620), .X(\filter_0/n9118 ) );
  nand_x1_sg U45675 ( .A(n27615), .B(n27616), .X(\filter_0/n9120 ) );
  nand_x1_sg U45676 ( .A(n27613), .B(n27614), .X(\filter_0/n9121 ) );
  nand_x1_sg U45677 ( .A(n27609), .B(n27610), .X(\filter_0/n9123 ) );
  nand_x1_sg U45678 ( .A(n27595), .B(n27596), .X(\filter_0/n9130 ) );
  nand_x1_sg U45679 ( .A(n27591), .B(n27592), .X(\filter_0/n9132 ) );
  nand_x1_sg U45680 ( .A(n27589), .B(n27590), .X(\filter_0/n9133 ) );
  nand_x1_sg U45681 ( .A(n27585), .B(n27586), .X(\filter_0/n9135 ) );
  nand_x1_sg U45682 ( .A(n27583), .B(n27584), .X(\filter_0/n9136 ) );
  nand_x1_sg U45683 ( .A(n27579), .B(n27580), .X(\filter_0/n9138 ) );
  nand_x1_sg U45684 ( .A(n27577), .B(n27578), .X(\filter_0/n9139 ) );
  nand_x1_sg U45685 ( .A(n27573), .B(n27574), .X(\filter_0/n9141 ) );
  nand_x1_sg U45686 ( .A(n27571), .B(n27572), .X(\filter_0/n9142 ) );
  nand_x1_sg U45687 ( .A(n27567), .B(n27568), .X(\filter_0/n9144 ) );
  nand_x1_sg U45688 ( .A(n27565), .B(n27566), .X(\filter_0/n9145 ) );
  nand_x1_sg U45689 ( .A(n27561), .B(n27562), .X(\filter_0/n9147 ) );
  nand_x1_sg U45690 ( .A(n27559), .B(n27560), .X(\filter_0/n9148 ) );
  nand_x1_sg U45691 ( .A(n27531), .B(n27532), .X(\filter_0/n9162 ) );
  nand_x1_sg U45692 ( .A(n27529), .B(n27530), .X(\filter_0/n9163 ) );
  nand_x1_sg U45693 ( .A(n27525), .B(n27526), .X(\filter_0/n9165 ) );
  nand_x1_sg U45694 ( .A(n27523), .B(n27524), .X(\filter_0/n9166 ) );
  nand_x1_sg U45695 ( .A(n27519), .B(n27520), .X(\filter_0/n9168 ) );
  nand_x1_sg U45696 ( .A(n27517), .B(n27518), .X(\filter_0/n9169 ) );
  nand_x1_sg U45697 ( .A(n27513), .B(n27514), .X(\filter_0/n9171 ) );
  nand_x1_sg U45698 ( .A(n27511), .B(n27512), .X(\filter_0/n9172 ) );
  nand_x1_sg U45699 ( .A(n27507), .B(n27508), .X(\filter_0/n9174 ) );
  nand_x1_sg U45700 ( .A(n27505), .B(n27506), .X(\filter_0/n9175 ) );
  nand_x1_sg U45701 ( .A(n27501), .B(n27502), .X(\filter_0/n9177 ) );
  nand_x1_sg U45702 ( .A(n27499), .B(n27500), .X(\filter_0/n9178 ) );
  nand_x1_sg U45703 ( .A(n27495), .B(n27496), .X(\filter_0/n9180 ) );
  nand_x1_sg U45704 ( .A(n27493), .B(n27494), .X(\filter_0/n9181 ) );
  nand_x1_sg U45705 ( .A(n27489), .B(n27490), .X(\filter_0/n9183 ) );
  nand_x1_sg U45706 ( .A(n27487), .B(n27488), .X(\filter_0/n9184 ) );
  nand_x1_sg U45707 ( .A(n27483), .B(n27484), .X(\filter_0/n9186 ) );
  nand_x1_sg U45708 ( .A(n27481), .B(n27482), .X(\filter_0/n9187 ) );
  nand_x1_sg U45709 ( .A(n27477), .B(n27478), .X(\filter_0/n9189 ) );
  nand_x1_sg U45710 ( .A(n27475), .B(n27476), .X(\filter_0/n9190 ) );
  nand_x1_sg U45711 ( .A(n27471), .B(n27472), .X(\filter_0/n9192 ) );
  nand_x1_sg U45712 ( .A(n27469), .B(n27470), .X(\filter_0/n9193 ) );
  nand_x1_sg U45713 ( .A(n27465), .B(n27466), .X(\filter_0/n9195 ) );
  nand_x1_sg U45714 ( .A(n27463), .B(n27464), .X(\filter_0/n9196 ) );
  nand_x1_sg U45715 ( .A(n27459), .B(n27460), .X(\filter_0/n9198 ) );
  nand_x1_sg U45716 ( .A(n27457), .B(n27458), .X(\filter_0/n9199 ) );
  nand_x1_sg U45717 ( .A(n27429), .B(n27430), .X(\filter_0/n9213 ) );
  nand_x1_sg U45718 ( .A(n27427), .B(n27428), .X(\filter_0/n9214 ) );
  nand_x1_sg U45719 ( .A(n27423), .B(n27424), .X(\filter_0/n9216 ) );
  nand_x1_sg U45720 ( .A(n27421), .B(n27422), .X(\filter_0/n9217 ) );
  nand_x1_sg U45721 ( .A(n27417), .B(n27418), .X(\filter_0/n9219 ) );
  nand_x1_sg U45722 ( .A(n27415), .B(n27416), .X(\filter_0/n9220 ) );
  nand_x1_sg U45723 ( .A(n27411), .B(n27412), .X(\filter_0/n9222 ) );
  nand_x1_sg U45724 ( .A(n27409), .B(n27410), .X(\filter_0/n9223 ) );
  nand_x1_sg U45725 ( .A(n27367), .B(n27368), .X(\filter_0/n9244 ) );
  nand_x1_sg U45726 ( .A(n27363), .B(n27364), .X(\filter_0/n9246 ) );
  nand_x1_sg U45727 ( .A(n27361), .B(n27362), .X(\filter_0/n9247 ) );
  nand_x1_sg U45728 ( .A(n27357), .B(n27358), .X(\filter_0/n9249 ) );
  nand_x1_sg U45729 ( .A(n27355), .B(n27356), .X(\filter_0/n9250 ) );
  nand_x1_sg U45730 ( .A(n27351), .B(n27352), .X(\filter_0/n9252 ) );
  nand_x1_sg U45731 ( .A(n27349), .B(n27350), .X(\filter_0/n9253 ) );
  nand_x1_sg U45732 ( .A(n27345), .B(n27346), .X(\filter_0/n9255 ) );
  nand_x1_sg U45733 ( .A(n27327), .B(n27328), .X(\filter_0/n9264 ) );
  nand_x1_sg U45734 ( .A(n27325), .B(n27326), .X(\filter_0/n9265 ) );
  nand_x1_sg U45735 ( .A(n27321), .B(n27322), .X(\filter_0/n9267 ) );
  nand_x1_sg U45736 ( .A(n27319), .B(n27320), .X(\filter_0/n9268 ) );
  nand_x1_sg U45737 ( .A(n27315), .B(n27316), .X(\filter_0/n9270 ) );
  nand_x1_sg U45738 ( .A(n27313), .B(n27314), .X(\filter_0/n9271 ) );
  nand_x1_sg U45739 ( .A(n27309), .B(n27310), .X(\filter_0/n9273 ) );
  nand_x1_sg U45740 ( .A(n27307), .B(n27308), .X(\filter_0/n9274 ) );
  nand_x1_sg U45741 ( .A(n27303), .B(n27304), .X(\filter_0/n9276 ) );
  nand_x1_sg U45742 ( .A(n27301), .B(n27302), .X(\filter_0/n9277 ) );
  nand_x1_sg U45743 ( .A(n27297), .B(n27298), .X(\filter_0/n9279 ) );
  nand_x1_sg U45744 ( .A(n27295), .B(n27296), .X(\filter_0/n9280 ) );
  nand_x1_sg U45745 ( .A(n27291), .B(n27292), .X(\filter_0/n9282 ) );
  nand_x1_sg U45746 ( .A(n27289), .B(n27290), .X(\filter_0/n9283 ) );
  nand_x1_sg U45747 ( .A(n27285), .B(n27286), .X(\filter_0/n9285 ) );
  nand_x1_sg U45748 ( .A(n27283), .B(n27284), .X(\filter_0/n9286 ) );
  nand_x1_sg U45749 ( .A(n27279), .B(n27280), .X(\filter_0/n9288 ) );
  nand_x1_sg U45750 ( .A(n27277), .B(n27278), .X(\filter_0/n9289 ) );
  nand_x1_sg U45751 ( .A(n27273), .B(n27274), .X(\filter_0/n9291 ) );
  nand_x1_sg U45752 ( .A(n27271), .B(n27272), .X(\filter_0/n9292 ) );
  nand_x1_sg U45753 ( .A(n27267), .B(n27268), .X(\filter_0/n9294 ) );
  nand_x1_sg U45754 ( .A(n27265), .B(n27266), .X(\filter_0/n9295 ) );
  nand_x1_sg U45755 ( .A(n27261), .B(n27262), .X(\filter_0/n9297 ) );
  nand_x1_sg U45756 ( .A(n27259), .B(n27260), .X(\filter_0/n9298 ) );
  nand_x1_sg U45757 ( .A(n27255), .B(n27256), .X(\filter_0/n9300 ) );
  nand_x1_sg U45758 ( .A(n27253), .B(n27254), .X(\filter_0/n9301 ) );
  nand_x1_sg U45759 ( .A(n27249), .B(n27250), .X(\filter_0/n9303 ) );
  nand_x1_sg U45760 ( .A(n27247), .B(n27248), .X(\filter_0/n9304 ) );
  nand_x1_sg U45761 ( .A(n27243), .B(n27244), .X(\filter_0/n9306 ) );
  nand_x1_sg U45762 ( .A(n27217), .B(n27218), .X(\filter_0/n9319 ) );
  nand_x1_sg U45763 ( .A(n27213), .B(n27214), .X(\filter_0/n9321 ) );
  nand_x1_sg U45764 ( .A(n27211), .B(n27212), .X(\filter_0/n9322 ) );
  nand_x1_sg U45765 ( .A(n27207), .B(n27208), .X(\filter_0/n9324 ) );
  nand_x1_sg U45766 ( .A(n27205), .B(n27206), .X(\filter_0/n9325 ) );
  nand_x1_sg U45767 ( .A(n27201), .B(n27202), .X(\filter_0/n9327 ) );
  nand_x1_sg U45768 ( .A(n27199), .B(n27200), .X(\filter_0/n9328 ) );
  nand_x1_sg U45769 ( .A(n27195), .B(n27196), .X(\filter_0/n9330 ) );
  nand_x1_sg U45770 ( .A(n27193), .B(n27194), .X(\filter_0/n9331 ) );
  nand_x1_sg U45771 ( .A(n27189), .B(n27190), .X(\filter_0/n9333 ) );
  nand_x1_sg U45772 ( .A(n27187), .B(n27188), .X(\filter_0/n9334 ) );
  nand_x1_sg U45773 ( .A(n27183), .B(n27184), .X(\filter_0/n9336 ) );
  nand_x1_sg U45774 ( .A(n27181), .B(n27182), .X(\filter_0/n9337 ) );
  nand_x1_sg U45775 ( .A(n27165), .B(n27166), .X(\filter_0/n9345 ) );
  nand_x1_sg U45776 ( .A(n27163), .B(n27164), .X(\filter_0/n9346 ) );
  nand_x1_sg U45777 ( .A(n27159), .B(n27160), .X(\filter_0/n9348 ) );
  nand_x1_sg U45778 ( .A(n27157), .B(n27158), .X(\filter_0/n9349 ) );
  nand_x1_sg U45779 ( .A(n27153), .B(n27154), .X(\filter_0/n9351 ) );
  nand_x1_sg U45780 ( .A(n27151), .B(n27152), .X(\filter_0/n9352 ) );
  nand_x1_sg U45781 ( .A(n27147), .B(n27148), .X(\filter_0/n9354 ) );
  nand_x1_sg U45782 ( .A(n27145), .B(n27146), .X(\filter_0/n9355 ) );
  nand_x1_sg U45783 ( .A(n27141), .B(n27142), .X(\filter_0/n9357 ) );
  nand_x1_sg U45784 ( .A(n27139), .B(n27140), .X(\filter_0/n9358 ) );
  nand_x1_sg U45785 ( .A(n27135), .B(n27136), .X(\filter_0/n9360 ) );
  nand_x1_sg U45786 ( .A(n27133), .B(n27134), .X(\filter_0/n9361 ) );
  nand_x1_sg U45787 ( .A(n27129), .B(n27130), .X(\filter_0/n9363 ) );
  nand_x1_sg U45788 ( .A(n27127), .B(n27128), .X(\filter_0/n9364 ) );
  nand_x1_sg U45789 ( .A(n27123), .B(n27124), .X(\filter_0/n9366 ) );
  nand_x1_sg U45790 ( .A(n27121), .B(n27122), .X(\filter_0/n9367 ) );
  nand_x1_sg U45791 ( .A(n27117), .B(n27118), .X(\filter_0/n9369 ) );
  nand_x1_sg U45792 ( .A(n27115), .B(n27116), .X(\filter_0/n9370 ) );
  nand_x1_sg U45793 ( .A(n27111), .B(n27112), .X(\filter_0/n9372 ) );
  nand_x1_sg U45794 ( .A(n27109), .B(n27110), .X(\filter_0/n9373 ) );
  nand_x1_sg U45795 ( .A(n27105), .B(n27106), .X(\filter_0/n9375 ) );
  nand_x1_sg U45796 ( .A(n27103), .B(n27104), .X(\filter_0/n9376 ) );
  nand_x1_sg U45797 ( .A(n27099), .B(n27100), .X(\filter_0/n9378 ) );
  nand_x1_sg U45798 ( .A(n27097), .B(n27098), .X(\filter_0/n9379 ) );
  nand_x1_sg U45799 ( .A(n27093), .B(n27094), .X(\filter_0/n9381 ) );
  nand_x1_sg U45800 ( .A(n27091), .B(n27092), .X(\filter_0/n9382 ) );
  nand_x1_sg U45801 ( .A(n27087), .B(n27088), .X(\filter_0/n9384 ) );
  nand_x1_sg U45802 ( .A(n27085), .B(n27086), .X(\filter_0/n9385 ) );
  nand_x1_sg U45803 ( .A(n27081), .B(n27082), .X(\filter_0/n9387 ) );
  nand_x1_sg U45804 ( .A(n27079), .B(n27080), .X(\filter_0/n9388 ) );
  nand_x1_sg U45805 ( .A(n27075), .B(n27076), .X(\filter_0/n9390 ) );
  nand_x1_sg U45806 ( .A(n27073), .B(n27074), .X(\filter_0/n9391 ) );
  nand_x1_sg U45807 ( .A(n27069), .B(n27070), .X(\filter_0/n9393 ) );
  nand_x1_sg U45808 ( .A(n27067), .B(n27068), .X(\filter_0/n9394 ) );
  nand_x1_sg U45809 ( .A(n27051), .B(n27052), .X(\filter_0/n9402 ) );
  nand_x1_sg U45810 ( .A(n27049), .B(n27050), .X(\filter_0/n9403 ) );
  nand_x1_sg U45811 ( .A(n27045), .B(n27046), .X(\filter_0/n9405 ) );
  nand_x1_sg U45812 ( .A(n27043), .B(n27044), .X(\filter_0/n9406 ) );
  nand_x1_sg U45813 ( .A(n27001), .B(n27002), .X(\filter_0/n9427 ) );
  nand_x1_sg U45814 ( .A(n26997), .B(n26998), .X(\filter_0/n9429 ) );
  nand_x1_sg U45815 ( .A(n26995), .B(n26996), .X(\filter_0/n9430 ) );
  nand_x1_sg U45816 ( .A(n26991), .B(n26992), .X(\filter_0/n9432 ) );
  nand_x1_sg U45817 ( .A(n26989), .B(n26990), .X(\filter_0/n9433 ) );
  nand_x1_sg U45818 ( .A(n26985), .B(n26986), .X(\filter_0/n9435 ) );
  nand_x1_sg U45819 ( .A(n26983), .B(n26984), .X(\filter_0/n9436 ) );
  nand_x1_sg U45820 ( .A(n26979), .B(n26980), .X(\filter_0/n9438 ) );
  nand_x1_sg U45821 ( .A(n26977), .B(n26978), .X(\filter_0/n9439 ) );
  nand_x1_sg U45822 ( .A(n26973), .B(n26974), .X(\filter_0/n9441 ) );
  nand_x1_sg U45823 ( .A(n26971), .B(n26972), .X(\filter_0/n9442 ) );
  nand_x1_sg U45824 ( .A(n26967), .B(n26968), .X(\filter_0/n9444 ) );
  nand_x1_sg U45825 ( .A(n26937), .B(n26938), .X(\filter_0/n9459 ) );
  nand_x1_sg U45826 ( .A(n26935), .B(n26936), .X(\filter_0/n9460 ) );
  nand_x1_sg U45827 ( .A(n26931), .B(n26932), .X(\filter_0/n9462 ) );
  nand_x1_sg U45828 ( .A(n26929), .B(n26930), .X(\filter_0/n9463 ) );
  nand_x1_sg U45829 ( .A(n26925), .B(n26926), .X(\filter_0/n9465 ) );
  nand_x1_sg U45830 ( .A(n26923), .B(n26924), .X(\filter_0/n9466 ) );
  nand_x1_sg U45831 ( .A(n26919), .B(n26920), .X(\filter_0/n9468 ) );
  nand_x1_sg U45832 ( .A(n26917), .B(n26918), .X(\filter_0/n9469 ) );
  nand_x1_sg U45833 ( .A(n26913), .B(n26914), .X(\filter_0/n9471 ) );
  nand_x1_sg U45834 ( .A(n26911), .B(n26912), .X(\filter_0/n9472 ) );
  nand_x1_sg U45835 ( .A(n26907), .B(n26908), .X(\filter_0/n9474 ) );
  nand_x1_sg U45836 ( .A(n26905), .B(n26906), .X(\filter_0/n9475 ) );
  nand_x1_sg U45837 ( .A(n26901), .B(n26902), .X(\filter_0/n9477 ) );
  nand_x1_sg U45838 ( .A(n26899), .B(n26900), .X(\filter_0/n9478 ) );
  nand_x1_sg U45839 ( .A(n26895), .B(n26896), .X(\filter_0/n9480 ) );
  nand_x1_sg U45840 ( .A(n26893), .B(n26894), .X(\filter_0/n9481 ) );
  nand_x1_sg U45841 ( .A(n26889), .B(n26890), .X(\filter_0/n9483 ) );
  nand_x1_sg U45842 ( .A(n26887), .B(n26888), .X(\filter_0/n9484 ) );
  nand_x1_sg U45843 ( .A(n26883), .B(n26884), .X(\filter_0/n9486 ) );
  nand_x1_sg U45844 ( .A(n26881), .B(n26882), .X(\filter_0/n9487 ) );
  nand_x1_sg U45845 ( .A(n26877), .B(n26878), .X(\filter_0/n9489 ) );
  nand_x1_sg U45846 ( .A(n26839), .B(n26840), .X(\filter_0/n9508 ) );
  nand_x1_sg U45847 ( .A(n26835), .B(n26836), .X(\filter_0/n9510 ) );
  nand_x1_sg U45848 ( .A(n26833), .B(n26834), .X(\filter_0/n9511 ) );
  nand_x1_sg U45849 ( .A(n26829), .B(n26830), .X(\filter_0/n9513 ) );
  nand_x1_sg U45850 ( .A(n26827), .B(n26828), .X(\filter_0/n9514 ) );
  nand_x1_sg U45851 ( .A(n26823), .B(n26824), .X(\filter_0/n9516 ) );
  nand_x1_sg U45852 ( .A(n26821), .B(n26822), .X(\filter_0/n9517 ) );
  nand_x1_sg U45853 ( .A(n26817), .B(n26818), .X(\filter_0/n9519 ) );
  nand_x1_sg U45854 ( .A(n26815), .B(n26816), .X(\filter_0/n9520 ) );
  nand_x1_sg U45855 ( .A(n26811), .B(n26812), .X(\filter_0/n9522 ) );
  nand_x1_sg U45856 ( .A(n26809), .B(n26810), .X(\filter_0/n9523 ) );
  nand_x1_sg U45857 ( .A(n26805), .B(n26806), .X(\filter_0/n9525 ) );
  nand_x1_sg U45858 ( .A(n26803), .B(n26804), .X(\filter_0/n9526 ) );
  nand_x1_sg U45859 ( .A(n26799), .B(n26800), .X(\filter_0/n9528 ) );
  nand_x1_sg U45860 ( .A(n26797), .B(n26798), .X(\filter_0/n9529 ) );
  nand_x1_sg U45861 ( .A(n26793), .B(n26794), .X(\filter_0/n9531 ) );
  nand_x1_sg U45862 ( .A(n26791), .B(n26792), .X(\filter_0/n9532 ) );
  nand_x1_sg U45863 ( .A(n26787), .B(n26788), .X(\filter_0/n9534 ) );
  nand_x1_sg U45864 ( .A(n26785), .B(n26786), .X(\filter_0/n9535 ) );
  nand_x1_sg U45865 ( .A(n26781), .B(n26782), .X(\filter_0/n9537 ) );
  nand_x1_sg U45866 ( .A(n26779), .B(n26780), .X(\filter_0/n9538 ) );
  nand_x1_sg U45867 ( .A(n26775), .B(n26776), .X(\filter_0/n9540 ) );
  nand_x1_sg U45868 ( .A(n26773), .B(n26774), .X(\filter_0/n9541 ) );
  nand_x1_sg U45869 ( .A(n26769), .B(n26770), .X(\filter_0/n9543 ) );
  nand_x1_sg U45870 ( .A(n26767), .B(n26768), .X(\filter_0/n9544 ) );
  nand_x1_sg U45871 ( .A(n26763), .B(n26764), .X(\filter_0/n9546 ) );
  nand_x1_sg U45872 ( .A(n26761), .B(n26762), .X(\filter_0/n9547 ) );
  nand_x1_sg U45873 ( .A(n26757), .B(n26758), .X(\filter_0/n9549 ) );
  nand_x1_sg U45874 ( .A(n26755), .B(n26756), .X(\filter_0/n9550 ) );
  nand_x1_sg U45875 ( .A(n26751), .B(n26752), .X(\filter_0/n9552 ) );
  nand_x1_sg U45876 ( .A(n26749), .B(n26750), .X(\filter_0/n9553 ) );
  nand_x1_sg U45877 ( .A(n26745), .B(n26746), .X(\filter_0/n9555 ) );
  nand_x1_sg U45878 ( .A(n26743), .B(n26744), .X(\filter_0/n9556 ) );
  nand_x1_sg U45879 ( .A(n26739), .B(n26740), .X(\filter_0/n9558 ) );
  nand_x1_sg U45880 ( .A(n26737), .B(n26738), .X(\filter_0/n9559 ) );
  nand_x1_sg U45881 ( .A(n26733), .B(n26734), .X(\filter_0/n9561 ) );
  nand_x1_sg U45882 ( .A(n26731), .B(n26732), .X(\filter_0/n9562 ) );
  nand_x1_sg U45883 ( .A(n26727), .B(n26728), .X(\filter_0/n9564 ) );
  nand_x1_sg U45884 ( .A(n26725), .B(n26726), .X(\filter_0/n9565 ) );
  nand_x1_sg U45885 ( .A(n26721), .B(n26722), .X(\filter_0/n9567 ) );
  nand_x1_sg U45886 ( .A(n26719), .B(n26720), .X(\filter_0/n9568 ) );
  nand_x1_sg U45887 ( .A(n26715), .B(n26716), .X(\filter_0/n9570 ) );
  nand_x1_sg U45888 ( .A(n26713), .B(n26714), .X(\filter_0/n9571 ) );
  nand_x1_sg U45889 ( .A(n26709), .B(n26710), .X(\filter_0/n9573 ) );
  nand_x1_sg U45890 ( .A(n26707), .B(n26708), .X(\filter_0/n9574 ) );
  nand_x1_sg U45891 ( .A(n26703), .B(n26704), .X(\filter_0/n9576 ) );
  nand_x1_sg U45892 ( .A(n26701), .B(n26702), .X(\filter_0/n9577 ) );
  nand_x1_sg U45893 ( .A(n26697), .B(n26698), .X(\filter_0/n9579 ) );
  nand_x1_sg U45894 ( .A(n26695), .B(n26696), .X(\filter_0/n9580 ) );
  nand_x1_sg U45895 ( .A(n26691), .B(n26692), .X(\filter_0/n9582 ) );
  nand_x1_sg U45896 ( .A(n26689), .B(n26690), .X(\filter_0/n9583 ) );
  nand_x1_sg U45897 ( .A(n26685), .B(n26686), .X(\filter_0/n9585 ) );
  nand_x1_sg U45898 ( .A(n26683), .B(n26684), .X(\filter_0/n9586 ) );
  nand_x1_sg U45899 ( .A(n26679), .B(n26680), .X(\filter_0/n9588 ) );
  nand_x1_sg U45900 ( .A(n26677), .B(n26678), .X(\filter_0/n9589 ) );
  nand_x1_sg U45901 ( .A(n26635), .B(n26636), .X(\filter_0/n9610 ) );
  nand_x1_sg U45902 ( .A(n26631), .B(n26632), .X(\filter_0/n9612 ) );
  nand_x1_sg U45903 ( .A(n26629), .B(n26630), .X(\filter_0/n9613 ) );
  nand_x1_sg U45904 ( .A(n26625), .B(n26626), .X(\filter_0/n9615 ) );
  nand_x1_sg U45905 ( .A(n26623), .B(n26624), .X(\filter_0/n9616 ) );
  nand_x1_sg U45906 ( .A(n26619), .B(n26620), .X(\filter_0/n9618 ) );
  nand_x1_sg U45907 ( .A(n26617), .B(n26618), .X(\filter_0/n9619 ) );
  nand_x1_sg U45908 ( .A(n26613), .B(n26614), .X(\filter_0/n9621 ) );
  nand_x1_sg U45909 ( .A(n26611), .B(n26612), .X(\filter_0/n9622 ) );
  nand_x1_sg U45910 ( .A(n26607), .B(n26608), .X(\filter_0/n9624 ) );
  nand_x1_sg U45911 ( .A(n26605), .B(n26606), .X(\filter_0/n9625 ) );
  nand_x1_sg U45912 ( .A(n26601), .B(n26602), .X(\filter_0/n9627 ) );
  nand_x1_sg U45913 ( .A(n26599), .B(n26600), .X(\filter_0/n9628 ) );
  nand_x1_sg U45914 ( .A(n26595), .B(n26596), .X(\filter_0/n9630 ) );
  nand_x1_sg U45915 ( .A(n26593), .B(n26594), .X(\filter_0/n9631 ) );
  nand_x1_sg U45916 ( .A(n28235), .B(n28236), .X(\filter_0/n8900 ) );
  nand_x1_sg U45917 ( .A(n28230), .B(n28231), .X(\filter_0/n8901 ) );
  nand_x1_sg U45918 ( .A(n28225), .B(n28226), .X(\filter_0/n8902 ) );
  nand_x1_sg U45919 ( .A(n28220), .B(n28221), .X(\filter_0/n8903 ) );
  nand_x1_sg U45920 ( .A(n28215), .B(n28216), .X(\filter_0/n8904 ) );
  nand_x1_sg U45921 ( .A(n28210), .B(n28211), .X(\filter_0/n8905 ) );
  nand_x1_sg U45922 ( .A(n28205), .B(n28206), .X(\filter_0/n8906 ) );
  nand_x1_sg U45923 ( .A(n28200), .B(n28201), .X(\filter_0/n8907 ) );
  nand_x1_sg U45924 ( .A(n28195), .B(n28196), .X(\filter_0/n8908 ) );
  nand_x1_sg U45925 ( .A(n28190), .B(n28191), .X(\filter_0/n8909 ) );
  nand_x1_sg U45926 ( .A(n28185), .B(n28186), .X(\filter_0/n8910 ) );
  nand_x1_sg U45927 ( .A(n28180), .B(n28181), .X(\filter_0/n8911 ) );
  nand_x1_sg U45928 ( .A(n28175), .B(n28176), .X(\filter_0/n8912 ) );
  nand_x1_sg U45929 ( .A(n28170), .B(n28171), .X(\filter_0/n8913 ) );
  nand_x1_sg U45930 ( .A(n28165), .B(n28166), .X(\filter_0/n8914 ) );
  nand_x1_sg U45931 ( .A(n28160), .B(n28161), .X(\filter_0/n8915 ) );
  nand_x1_sg U45932 ( .A(n28155), .B(n28156), .X(\filter_0/n8916 ) );
  nand_x1_sg U45933 ( .A(n28150), .B(n28151), .X(\filter_0/n8917 ) );
  nand_x1_sg U45934 ( .A(n28040), .B(n28041), .X(\filter_0/n8939 ) );
  nand_x1_sg U45935 ( .A(n28035), .B(n28036), .X(\filter_0/n8940 ) );
  nand_x1_sg U45936 ( .A(n27940), .B(n27941), .X(\filter_0/n8959 ) );
  nand_x1_sg U45937 ( .A(n27935), .B(n27936), .X(\filter_0/n8960 ) );
  nand_x1_sg U45938 ( .A(n27929), .B(n27930), .X(\filter_0/n8963 ) );
  nand_x1_sg U45939 ( .A(n27923), .B(n27924), .X(\filter_0/n8966 ) );
  nand_x1_sg U45940 ( .A(n27917), .B(n27918), .X(\filter_0/n8969 ) );
  nand_x1_sg U45941 ( .A(n27911), .B(n27912), .X(\filter_0/n8972 ) );
  nand_x1_sg U45942 ( .A(n27905), .B(n27906), .X(\filter_0/n8975 ) );
  nand_x1_sg U45943 ( .A(n27899), .B(n27900), .X(\filter_0/n8978 ) );
  nand_x1_sg U45944 ( .A(n27845), .B(n27846), .X(\filter_0/n9005 ) );
  nand_x1_sg U45945 ( .A(n27839), .B(n27840), .X(\filter_0/n9008 ) );
  nand_x1_sg U45946 ( .A(n27833), .B(n27834), .X(\filter_0/n9011 ) );
  nand_x1_sg U45947 ( .A(n27827), .B(n27828), .X(\filter_0/n9014 ) );
  nand_x1_sg U45948 ( .A(n27821), .B(n27822), .X(\filter_0/n9017 ) );
  nand_x1_sg U45949 ( .A(n27815), .B(n27816), .X(\filter_0/n9020 ) );
  nand_x1_sg U45950 ( .A(n27767), .B(n27768), .X(\filter_0/n9044 ) );
  nand_x1_sg U45951 ( .A(n27761), .B(n27762), .X(\filter_0/n9047 ) );
  nand_x1_sg U45952 ( .A(n27755), .B(n27756), .X(\filter_0/n9050 ) );
  nand_x1_sg U45953 ( .A(n27749), .B(n27750), .X(\filter_0/n9053 ) );
  nand_x1_sg U45954 ( .A(n27743), .B(n27744), .X(\filter_0/n9056 ) );
  nand_x1_sg U45955 ( .A(n27737), .B(n27738), .X(\filter_0/n9059 ) );
  nand_x1_sg U45956 ( .A(n27605), .B(n27606), .X(\filter_0/n9125 ) );
  nand_x1_sg U45957 ( .A(n27599), .B(n27600), .X(\filter_0/n9128 ) );
  nand_x1_sg U45958 ( .A(n27557), .B(n27558), .X(\filter_0/n9149 ) );
  nand_x1_sg U45959 ( .A(n27551), .B(n27552), .X(\filter_0/n9152 ) );
  nand_x1_sg U45960 ( .A(n27545), .B(n27546), .X(\filter_0/n9155 ) );
  nand_x1_sg U45961 ( .A(n27539), .B(n27540), .X(\filter_0/n9158 ) );
  nand_x1_sg U45962 ( .A(n27533), .B(n27534), .X(\filter_0/n9161 ) );
  nand_x1_sg U45963 ( .A(n27455), .B(n27456), .X(\filter_0/n9200 ) );
  nand_x1_sg U45964 ( .A(n27449), .B(n27450), .X(\filter_0/n9203 ) );
  nand_x1_sg U45965 ( .A(n27443), .B(n27444), .X(\filter_0/n9206 ) );
  nand_x1_sg U45966 ( .A(n27437), .B(n27438), .X(\filter_0/n9209 ) );
  nand_x1_sg U45967 ( .A(n27401), .B(n27402), .X(\filter_0/n9227 ) );
  nand_x1_sg U45968 ( .A(n27395), .B(n27396), .X(\filter_0/n9230 ) );
  nand_x1_sg U45969 ( .A(n27389), .B(n27390), .X(\filter_0/n9233 ) );
  nand_x1_sg U45970 ( .A(n27383), .B(n27384), .X(\filter_0/n9236 ) );
  nand_x1_sg U45971 ( .A(n27377), .B(n27378), .X(\filter_0/n9239 ) );
  nand_x1_sg U45972 ( .A(n27371), .B(n27372), .X(\filter_0/n9242 ) );
  nand_x1_sg U45973 ( .A(n27341), .B(n27342), .X(\filter_0/n9257 ) );
  nand_x1_sg U45974 ( .A(n27335), .B(n27336), .X(\filter_0/n9260 ) );
  nand_x1_sg U45975 ( .A(n27239), .B(n27240), .X(\filter_0/n9308 ) );
  nand_x1_sg U45976 ( .A(n27233), .B(n27234), .X(\filter_0/n9311 ) );
  nand_x1_sg U45977 ( .A(n27227), .B(n27228), .X(\filter_0/n9314 ) );
  nand_x1_sg U45978 ( .A(n27221), .B(n27222), .X(\filter_0/n9317 ) );
  nand_x1_sg U45979 ( .A(n27179), .B(n27180), .X(\filter_0/n9338 ) );
  nand_x1_sg U45980 ( .A(n27173), .B(n27174), .X(\filter_0/n9341 ) );
  nand_x1_sg U45981 ( .A(n27167), .B(n27168), .X(\filter_0/n9344 ) );
  nand_x1_sg U45982 ( .A(n27065), .B(n27066), .X(\filter_0/n9395 ) );
  nand_x1_sg U45983 ( .A(n27059), .B(n27060), .X(\filter_0/n9398 ) );
  nand_x1_sg U45984 ( .A(n27035), .B(n27036), .X(\filter_0/n9410 ) );
  nand_x1_sg U45985 ( .A(n27029), .B(n27030), .X(\filter_0/n9413 ) );
  nand_x1_sg U45986 ( .A(n27023), .B(n27024), .X(\filter_0/n9416 ) );
  nand_x1_sg U45987 ( .A(n27017), .B(n27018), .X(\filter_0/n9419 ) );
  nand_x1_sg U45988 ( .A(n27011), .B(n27012), .X(\filter_0/n9422 ) );
  nand_x1_sg U45989 ( .A(n27005), .B(n27006), .X(\filter_0/n9425 ) );
  nand_x1_sg U45990 ( .A(n26963), .B(n26964), .X(\filter_0/n9446 ) );
  nand_x1_sg U45991 ( .A(n26957), .B(n26958), .X(\filter_0/n9449 ) );
  nand_x1_sg U45992 ( .A(n26951), .B(n26952), .X(\filter_0/n9452 ) );
  nand_x1_sg U45993 ( .A(n26945), .B(n26946), .X(\filter_0/n9455 ) );
  nand_x1_sg U45994 ( .A(n26873), .B(n26874), .X(\filter_0/n9491 ) );
  nand_x1_sg U45995 ( .A(n26867), .B(n26868), .X(\filter_0/n9494 ) );
  nand_x1_sg U45996 ( .A(n26861), .B(n26862), .X(\filter_0/n9497 ) );
  nand_x1_sg U45997 ( .A(n26855), .B(n26856), .X(\filter_0/n9500 ) );
  nand_x1_sg U45998 ( .A(n26849), .B(n26850), .X(\filter_0/n9503 ) );
  nand_x1_sg U45999 ( .A(n26843), .B(n26844), .X(\filter_0/n9506 ) );
  nand_x1_sg U46000 ( .A(n26801), .B(n26802), .X(\filter_0/n9527 ) );
  nand_x1_sg U46001 ( .A(n26669), .B(n26670), .X(\filter_0/n9593 ) );
  nand_x1_sg U46002 ( .A(n26663), .B(n26664), .X(\filter_0/n9596 ) );
  nand_x1_sg U46003 ( .A(n26657), .B(n26658), .X(\filter_0/n9599 ) );
  nand_x1_sg U46004 ( .A(n26651), .B(n26652), .X(\filter_0/n9602 ) );
  nand_x1_sg U46005 ( .A(n26645), .B(n26646), .X(\filter_0/n9605 ) );
  nand_x1_sg U46006 ( .A(n26639), .B(n26640), .X(\filter_0/n9608 ) );
  nand_x1_sg U46007 ( .A(n27933), .B(n27934), .X(\filter_0/n8961 ) );
  nand_x1_sg U46008 ( .A(n27931), .B(n27932), .X(\filter_0/n8962 ) );
  nand_x1_sg U46009 ( .A(n27927), .B(n27928), .X(\filter_0/n8964 ) );
  nand_x1_sg U46010 ( .A(n27925), .B(n27926), .X(\filter_0/n8965 ) );
  nand_x1_sg U46011 ( .A(n27921), .B(n27922), .X(\filter_0/n8967 ) );
  nand_x1_sg U46012 ( .A(n27919), .B(n27920), .X(\filter_0/n8968 ) );
  nand_x1_sg U46013 ( .A(n27915), .B(n27916), .X(\filter_0/n8970 ) );
  nand_x1_sg U46014 ( .A(n27913), .B(n27914), .X(\filter_0/n8971 ) );
  nand_x1_sg U46015 ( .A(n27909), .B(n27910), .X(\filter_0/n8973 ) );
  nand_x1_sg U46016 ( .A(n27907), .B(n27908), .X(\filter_0/n8974 ) );
  nand_x1_sg U46017 ( .A(n27903), .B(n27904), .X(\filter_0/n8976 ) );
  nand_x1_sg U46018 ( .A(n27901), .B(n27902), .X(\filter_0/n8977 ) );
  nand_x1_sg U46019 ( .A(n27843), .B(n27844), .X(\filter_0/n9006 ) );
  nand_x1_sg U46020 ( .A(n27841), .B(n27842), .X(\filter_0/n9007 ) );
  nand_x1_sg U46021 ( .A(n27837), .B(n27838), .X(\filter_0/n9009 ) );
  nand_x1_sg U46022 ( .A(n27835), .B(n27836), .X(\filter_0/n9010 ) );
  nand_x1_sg U46023 ( .A(n27831), .B(n27832), .X(\filter_0/n9012 ) );
  nand_x1_sg U46024 ( .A(n27829), .B(n27830), .X(\filter_0/n9013 ) );
  nand_x1_sg U46025 ( .A(n27825), .B(n27826), .X(\filter_0/n9015 ) );
  nand_x1_sg U46026 ( .A(n27823), .B(n27824), .X(\filter_0/n9016 ) );
  nand_x1_sg U46027 ( .A(n27819), .B(n27820), .X(\filter_0/n9018 ) );
  nand_x1_sg U46028 ( .A(n27817), .B(n27818), .X(\filter_0/n9019 ) );
  nand_x1_sg U46029 ( .A(n27813), .B(n27814), .X(\filter_0/n9021 ) );
  nand_x1_sg U46030 ( .A(n27811), .B(n27812), .X(\filter_0/n9022 ) );
  nand_x1_sg U46031 ( .A(n27771), .B(n27772), .X(\filter_0/n9042 ) );
  nand_x1_sg U46032 ( .A(n27769), .B(n27770), .X(\filter_0/n9043 ) );
  nand_x1_sg U46033 ( .A(n27765), .B(n27766), .X(\filter_0/n9045 ) );
  nand_x1_sg U46034 ( .A(n27763), .B(n27764), .X(\filter_0/n9046 ) );
  nand_x1_sg U46035 ( .A(n27759), .B(n27760), .X(\filter_0/n9048 ) );
  nand_x1_sg U46036 ( .A(n27757), .B(n27758), .X(\filter_0/n9049 ) );
  nand_x1_sg U46037 ( .A(n27753), .B(n27754), .X(\filter_0/n9051 ) );
  nand_x1_sg U46038 ( .A(n27751), .B(n27752), .X(\filter_0/n9052 ) );
  nand_x1_sg U46039 ( .A(n27747), .B(n27748), .X(\filter_0/n9054 ) );
  nand_x1_sg U46040 ( .A(n27745), .B(n27746), .X(\filter_0/n9055 ) );
  nand_x1_sg U46041 ( .A(n27741), .B(n27742), .X(\filter_0/n9057 ) );
  nand_x1_sg U46042 ( .A(n27739), .B(n27740), .X(\filter_0/n9058 ) );
  nand_x1_sg U46043 ( .A(n27735), .B(n27736), .X(\filter_0/n9060 ) );
  nand_x1_sg U46044 ( .A(n27721), .B(n27722), .X(\filter_0/n9067 ) );
  nand_x1_sg U46045 ( .A(n27607), .B(n27608), .X(\filter_0/n9124 ) );
  nand_x1_sg U46046 ( .A(n27603), .B(n27604), .X(\filter_0/n9126 ) );
  nand_x1_sg U46047 ( .A(n27601), .B(n27602), .X(\filter_0/n9127 ) );
  nand_x1_sg U46048 ( .A(n27597), .B(n27598), .X(\filter_0/n9129 ) );
  nand_x1_sg U46049 ( .A(n27555), .B(n27556), .X(\filter_0/n9150 ) );
  nand_x1_sg U46050 ( .A(n27553), .B(n27554), .X(\filter_0/n9151 ) );
  nand_x1_sg U46051 ( .A(n27549), .B(n27550), .X(\filter_0/n9153 ) );
  nand_x1_sg U46052 ( .A(n27547), .B(n27548), .X(\filter_0/n9154 ) );
  nand_x1_sg U46053 ( .A(n27543), .B(n27544), .X(\filter_0/n9156 ) );
  nand_x1_sg U46054 ( .A(n27541), .B(n27542), .X(\filter_0/n9157 ) );
  nand_x1_sg U46055 ( .A(n27537), .B(n27538), .X(\filter_0/n9159 ) );
  nand_x1_sg U46056 ( .A(n27535), .B(n27536), .X(\filter_0/n9160 ) );
  nand_x1_sg U46057 ( .A(n27453), .B(n27454), .X(\filter_0/n9201 ) );
  nand_x1_sg U46058 ( .A(n27451), .B(n27452), .X(\filter_0/n9202 ) );
  nand_x1_sg U46059 ( .A(n27447), .B(n27448), .X(\filter_0/n9204 ) );
  nand_x1_sg U46060 ( .A(n27445), .B(n27446), .X(\filter_0/n9205 ) );
  nand_x1_sg U46061 ( .A(n27441), .B(n27442), .X(\filter_0/n9207 ) );
  nand_x1_sg U46062 ( .A(n27439), .B(n27440), .X(\filter_0/n9208 ) );
  nand_x1_sg U46063 ( .A(n27435), .B(n27436), .X(\filter_0/n9210 ) );
  nand_x1_sg U46064 ( .A(n27433), .B(n27434), .X(\filter_0/n9211 ) );
  nand_x1_sg U46065 ( .A(n27405), .B(n27406), .X(\filter_0/n9225 ) );
  nand_x1_sg U46066 ( .A(n27403), .B(n27404), .X(\filter_0/n9226 ) );
  nand_x1_sg U46067 ( .A(n27399), .B(n27400), .X(\filter_0/n9228 ) );
  nand_x1_sg U46068 ( .A(n27397), .B(n27398), .X(\filter_0/n9229 ) );
  nand_x1_sg U46069 ( .A(n27393), .B(n27394), .X(\filter_0/n9231 ) );
  nand_x1_sg U46070 ( .A(n27391), .B(n27392), .X(\filter_0/n9232 ) );
  nand_x1_sg U46071 ( .A(n27387), .B(n27388), .X(\filter_0/n9234 ) );
  nand_x1_sg U46072 ( .A(n27385), .B(n27386), .X(\filter_0/n9235 ) );
  nand_x1_sg U46073 ( .A(n27381), .B(n27382), .X(\filter_0/n9237 ) );
  nand_x1_sg U46074 ( .A(n27379), .B(n27380), .X(\filter_0/n9238 ) );
  nand_x1_sg U46075 ( .A(n27375), .B(n27376), .X(\filter_0/n9240 ) );
  nand_x1_sg U46076 ( .A(n27373), .B(n27374), .X(\filter_0/n9241 ) );
  nand_x1_sg U46077 ( .A(n27369), .B(n27370), .X(\filter_0/n9243 ) );
  nand_x1_sg U46078 ( .A(n27343), .B(n27344), .X(\filter_0/n9256 ) );
  nand_x1_sg U46079 ( .A(n27339), .B(n27340), .X(\filter_0/n9258 ) );
  nand_x1_sg U46080 ( .A(n27337), .B(n27338), .X(\filter_0/n9259 ) );
  nand_x1_sg U46081 ( .A(n27333), .B(n27334), .X(\filter_0/n9261 ) );
  nand_x1_sg U46082 ( .A(n27331), .B(n27332), .X(\filter_0/n9262 ) );
  nand_x1_sg U46083 ( .A(n27241), .B(n27242), .X(\filter_0/n9307 ) );
  nand_x1_sg U46084 ( .A(n27237), .B(n27238), .X(\filter_0/n9309 ) );
  nand_x1_sg U46085 ( .A(n27235), .B(n27236), .X(\filter_0/n9310 ) );
  nand_x1_sg U46086 ( .A(n27231), .B(n27232), .X(\filter_0/n9312 ) );
  nand_x1_sg U46087 ( .A(n27229), .B(n27230), .X(\filter_0/n9313 ) );
  nand_x1_sg U46088 ( .A(n27225), .B(n27226), .X(\filter_0/n9315 ) );
  nand_x1_sg U46089 ( .A(n27223), .B(n27224), .X(\filter_0/n9316 ) );
  nand_x1_sg U46090 ( .A(n27219), .B(n27220), .X(\filter_0/n9318 ) );
  nand_x1_sg U46091 ( .A(n27177), .B(n27178), .X(\filter_0/n9339 ) );
  nand_x1_sg U46092 ( .A(n27175), .B(n27176), .X(\filter_0/n9340 ) );
  nand_x1_sg U46093 ( .A(n27171), .B(n27172), .X(\filter_0/n9342 ) );
  nand_x1_sg U46094 ( .A(n27169), .B(n27170), .X(\filter_0/n9343 ) );
  nand_x1_sg U46095 ( .A(n27063), .B(n27064), .X(\filter_0/n9396 ) );
  nand_x1_sg U46096 ( .A(n27061), .B(n27062), .X(\filter_0/n9397 ) );
  nand_x1_sg U46097 ( .A(n27057), .B(n27058), .X(\filter_0/n9399 ) );
  nand_x1_sg U46098 ( .A(n27055), .B(n27056), .X(\filter_0/n9400 ) );
  nand_x1_sg U46099 ( .A(n27039), .B(n27040), .X(\filter_0/n9408 ) );
  nand_x1_sg U46100 ( .A(n27037), .B(n27038), .X(\filter_0/n9409 ) );
  nand_x1_sg U46101 ( .A(n27033), .B(n27034), .X(\filter_0/n9411 ) );
  nand_x1_sg U46102 ( .A(n27031), .B(n27032), .X(\filter_0/n9412 ) );
  nand_x1_sg U46103 ( .A(n27027), .B(n27028), .X(\filter_0/n9414 ) );
  nand_x1_sg U46104 ( .A(n27025), .B(n27026), .X(\filter_0/n9415 ) );
  nand_x1_sg U46105 ( .A(n27021), .B(n27022), .X(\filter_0/n9417 ) );
  nand_x1_sg U46106 ( .A(n27019), .B(n27020), .X(\filter_0/n9418 ) );
  nand_x1_sg U46107 ( .A(n27015), .B(n27016), .X(\filter_0/n9420 ) );
  nand_x1_sg U46108 ( .A(n27013), .B(n27014), .X(\filter_0/n9421 ) );
  nand_x1_sg U46109 ( .A(n27009), .B(n27010), .X(\filter_0/n9423 ) );
  nand_x1_sg U46110 ( .A(n27007), .B(n27008), .X(\filter_0/n9424 ) );
  nand_x1_sg U46111 ( .A(n27003), .B(n27004), .X(\filter_0/n9426 ) );
  nand_x1_sg U46112 ( .A(n26965), .B(n26966), .X(\filter_0/n9445 ) );
  nand_x1_sg U46113 ( .A(n26961), .B(n26962), .X(\filter_0/n9447 ) );
  nand_x1_sg U46114 ( .A(n26959), .B(n26960), .X(\filter_0/n9448 ) );
  nand_x1_sg U46115 ( .A(n26955), .B(n26956), .X(\filter_0/n9450 ) );
  nand_x1_sg U46116 ( .A(n26953), .B(n26954), .X(\filter_0/n9451 ) );
  nand_x1_sg U46117 ( .A(n26949), .B(n26950), .X(\filter_0/n9453 ) );
  nand_x1_sg U46118 ( .A(n26947), .B(n26948), .X(\filter_0/n9454 ) );
  nand_x1_sg U46119 ( .A(n26943), .B(n26944), .X(\filter_0/n9456 ) );
  nand_x1_sg U46120 ( .A(n26941), .B(n26942), .X(\filter_0/n9457 ) );
  nand_x1_sg U46121 ( .A(n26875), .B(n26876), .X(\filter_0/n9490 ) );
  nand_x1_sg U46122 ( .A(n26871), .B(n26872), .X(\filter_0/n9492 ) );
  nand_x1_sg U46123 ( .A(n26869), .B(n26870), .X(\filter_0/n9493 ) );
  nand_x1_sg U46124 ( .A(n26865), .B(n26866), .X(\filter_0/n9495 ) );
  nand_x1_sg U46125 ( .A(n26863), .B(n26864), .X(\filter_0/n9496 ) );
  nand_x1_sg U46126 ( .A(n26859), .B(n26860), .X(\filter_0/n9498 ) );
  nand_x1_sg U46127 ( .A(n26857), .B(n26858), .X(\filter_0/n9499 ) );
  nand_x1_sg U46128 ( .A(n26853), .B(n26854), .X(\filter_0/n9501 ) );
  nand_x1_sg U46129 ( .A(n26851), .B(n26852), .X(\filter_0/n9502 ) );
  nand_x1_sg U46130 ( .A(n26847), .B(n26848), .X(\filter_0/n9504 ) );
  nand_x1_sg U46131 ( .A(n26845), .B(n26846), .X(\filter_0/n9505 ) );
  nand_x1_sg U46132 ( .A(n26841), .B(n26842), .X(\filter_0/n9507 ) );
  nand_x1_sg U46133 ( .A(n26673), .B(n26674), .X(\filter_0/n9591 ) );
  nand_x1_sg U46134 ( .A(n26671), .B(n26672), .X(\filter_0/n9592 ) );
  nand_x1_sg U46135 ( .A(n26667), .B(n26668), .X(\filter_0/n9594 ) );
  nand_x1_sg U46136 ( .A(n26665), .B(n26666), .X(\filter_0/n9595 ) );
  nand_x1_sg U46137 ( .A(n26661), .B(n26662), .X(\filter_0/n9597 ) );
  nand_x1_sg U46138 ( .A(n26659), .B(n26660), .X(\filter_0/n9598 ) );
  nand_x1_sg U46139 ( .A(n26655), .B(n26656), .X(\filter_0/n9600 ) );
  nand_x1_sg U46140 ( .A(n26653), .B(n26654), .X(\filter_0/n9601 ) );
  nand_x1_sg U46141 ( .A(n26649), .B(n26650), .X(\filter_0/n9603 ) );
  nand_x1_sg U46142 ( .A(n26647), .B(n26648), .X(\filter_0/n9604 ) );
  nand_x1_sg U46143 ( .A(n26643), .B(n26644), .X(\filter_0/n9606 ) );
  nand_x1_sg U46144 ( .A(n26641), .B(n26642), .X(\filter_0/n9607 ) );
  nand_x1_sg U46145 ( .A(n26637), .B(n26638), .X(\filter_0/n9609 ) );
  nand_x1_sg U46146 ( .A(n22225), .B(n22226), .X(n5978) );
  nand_x1_sg U46147 ( .A(n22231), .B(n22232), .X(n5975) );
  nand_x1_sg U46148 ( .A(n22237), .B(n22238), .X(n5972) );
  nand_x1_sg U46149 ( .A(n22243), .B(n22244), .X(n5969) );
  nand_x1_sg U46150 ( .A(n22249), .B(n22250), .X(n5966) );
  nand_x1_sg U46151 ( .A(n22255), .B(n22256), .X(n5963) );
  nand_x1_sg U46152 ( .A(n22261), .B(n22262), .X(n5960) );
  nand_x1_sg U46153 ( .A(n22267), .B(n22268), .X(n5957) );
  nand_x1_sg U46154 ( .A(n22273), .B(n22274), .X(n5954) );
  nand_x1_sg U46155 ( .A(n22279), .B(n22280), .X(n5951) );
  nand_x1_sg U46156 ( .A(n22285), .B(n22286), .X(n5948) );
  nand_x1_sg U46157 ( .A(n22291), .B(n22292), .X(n5945) );
  nand_x1_sg U46158 ( .A(n22297), .B(n22298), .X(n5942) );
  nand_x1_sg U46159 ( .A(n22303), .B(n22304), .X(n5939) );
  nand_x1_sg U46160 ( .A(n22309), .B(n22310), .X(n5936) );
  nand_x1_sg U46161 ( .A(n22315), .B(n22316), .X(n5933) );
  nand_x1_sg U46162 ( .A(n22321), .B(n22322), .X(n5930) );
  nand_x1_sg U46163 ( .A(n22327), .B(n22328), .X(n5927) );
  nand_x1_sg U46164 ( .A(n22333), .B(n22334), .X(n5924) );
  nand_x1_sg U46165 ( .A(n22339), .B(n22340), .X(n5921) );
  nand_x1_sg U46166 ( .A(n22345), .B(n22346), .X(n5918) );
  nand_x1_sg U46167 ( .A(n22351), .B(n22352), .X(n5915) );
  nand_x1_sg U46168 ( .A(n22357), .B(n22358), .X(n5912) );
  nand_x1_sg U46169 ( .A(n22363), .B(n22364), .X(n5909) );
  nand_x1_sg U46170 ( .A(n22369), .B(n22370), .X(n5906) );
  nand_x1_sg U46171 ( .A(n22375), .B(n22376), .X(n5903) );
  nand_x1_sg U46172 ( .A(n22381), .B(n22382), .X(n5900) );
  nand_x1_sg U46173 ( .A(n22387), .B(n22388), .X(n5897) );
  nand_x1_sg U46174 ( .A(n22393), .B(n22394), .X(n5894) );
  nand_x1_sg U46175 ( .A(n22399), .B(n22400), .X(n5891) );
  nand_x1_sg U46176 ( .A(n22405), .B(n22406), .X(n5888) );
  nand_x1_sg U46177 ( .A(n22411), .B(n22412), .X(n5885) );
  nand_x1_sg U46178 ( .A(n22417), .B(n22418), .X(n5882) );
  nand_x1_sg U46179 ( .A(n22423), .B(n22424), .X(n5879) );
  nand_x1_sg U46180 ( .A(n22429), .B(n22430), .X(n5876) );
  nand_x1_sg U46181 ( .A(n22435), .B(n22436), .X(n5873) );
  nand_x1_sg U46182 ( .A(n22441), .B(n22442), .X(n5870) );
  nand_x1_sg U46183 ( .A(n22447), .B(n22448), .X(n5867) );
  nand_x1_sg U46184 ( .A(n22453), .B(n22454), .X(n5864) );
  nand_x1_sg U46185 ( .A(n22459), .B(n22460), .X(n5861) );
  nand_x1_sg U46186 ( .A(n22465), .B(n22466), .X(n5858) );
  nand_x1_sg U46187 ( .A(n22471), .B(n22472), .X(n5855) );
  nand_x1_sg U46188 ( .A(n22477), .B(n22478), .X(n5852) );
  nand_x1_sg U46189 ( .A(n22483), .B(n22484), .X(n5849) );
  nand_x1_sg U46190 ( .A(n22489), .B(n22490), .X(n5846) );
  nand_x1_sg U46191 ( .A(n22495), .B(n22496), .X(n5843) );
  nand_x1_sg U46192 ( .A(n22501), .B(n22502), .X(n5840) );
  nand_x1_sg U46193 ( .A(n22507), .B(n22508), .X(n5837) );
  nand_x1_sg U46194 ( .A(n22513), .B(n22514), .X(n5834) );
  nand_x1_sg U46195 ( .A(n22519), .B(n22520), .X(n5831) );
  nand_x1_sg U46196 ( .A(n22525), .B(n22526), .X(n5828) );
  nand_x1_sg U46197 ( .A(n22531), .B(n22532), .X(n5825) );
  nand_x1_sg U46198 ( .A(n22537), .B(n22538), .X(n5822) );
  nand_x1_sg U46199 ( .A(n22543), .B(n22544), .X(n5819) );
  nand_x1_sg U46200 ( .A(n22549), .B(n22550), .X(n5816) );
  nand_x1_sg U46201 ( .A(n22555), .B(n22556), .X(n5813) );
  nand_x1_sg U46202 ( .A(n22561), .B(n22562), .X(n5810) );
  nand_x1_sg U46203 ( .A(n22567), .B(n22568), .X(n5807) );
  nand_x1_sg U46204 ( .A(n22573), .B(n22574), .X(n5804) );
  nand_x1_sg U46205 ( .A(n22579), .B(n22580), .X(n5801) );
  nand_x1_sg U46206 ( .A(n22585), .B(n22586), .X(n5798) );
  nand_x1_sg U46207 ( .A(n22591), .B(n22592), .X(n5795) );
  nand_x1_sg U46208 ( .A(n22597), .B(n22598), .X(n5792) );
  nand_x1_sg U46209 ( .A(n22603), .B(n22604), .X(n5789) );
  nand_x1_sg U46210 ( .A(n22609), .B(n22610), .X(n5786) );
  nand_x1_sg U46211 ( .A(n22615), .B(n22616), .X(n5783) );
  nand_x1_sg U46212 ( .A(n22621), .B(n22622), .X(n5780) );
  nand_x1_sg U46213 ( .A(n22627), .B(n22628), .X(n5777) );
  nand_x1_sg U46214 ( .A(n22633), .B(n22634), .X(n5774) );
  nand_x1_sg U46215 ( .A(n22639), .B(n22640), .X(n5771) );
  nand_x1_sg U46216 ( .A(n22645), .B(n22646), .X(n5768) );
  nand_x1_sg U46217 ( .A(n22651), .B(n22652), .X(n5765) );
  nand_x1_sg U46218 ( .A(n22657), .B(n22658), .X(n5762) );
  nand_x1_sg U46219 ( .A(n22663), .B(n22664), .X(n5759) );
  nand_x1_sg U46220 ( .A(n22669), .B(n22670), .X(n5756) );
  nand_x1_sg U46221 ( .A(n22675), .B(n22676), .X(n5753) );
  nand_x1_sg U46222 ( .A(n22681), .B(n22682), .X(n5750) );
  nand_x1_sg U46223 ( .A(n22687), .B(n22688), .X(n5747) );
  nand_x1_sg U46224 ( .A(n22693), .B(n22694), .X(n5744) );
  nand_x1_sg U46225 ( .A(n22699), .B(n22700), .X(n5741) );
  nand_x1_sg U46226 ( .A(n22705), .B(n22706), .X(n5738) );
  nand_x1_sg U46227 ( .A(n22711), .B(n22712), .X(n5735) );
  nand_x1_sg U46228 ( .A(n22717), .B(n22718), .X(n5732) );
  nand_x1_sg U46229 ( .A(n22723), .B(n22724), .X(n5729) );
  nand_x1_sg U46230 ( .A(n22729), .B(n22730), .X(n5726) );
  nand_x1_sg U46231 ( .A(n22735), .B(n22736), .X(n5723) );
  nand_x1_sg U46232 ( .A(n22741), .B(n22742), .X(n5720) );
  nand_x1_sg U46233 ( .A(n22747), .B(n22748), .X(n5717) );
  nand_x1_sg U46234 ( .A(n22753), .B(n22754), .X(n5714) );
  nand_x1_sg U46235 ( .A(n22759), .B(n22760), .X(n5711) );
  nand_x1_sg U46236 ( .A(n22765), .B(n22766), .X(n5708) );
  nand_x1_sg U46237 ( .A(n22771), .B(n22772), .X(n5705) );
  nand_x1_sg U46238 ( .A(n22777), .B(n22778), .X(n5702) );
  nand_x1_sg U46239 ( .A(n22783), .B(n22784), .X(n5699) );
  nand_x1_sg U46240 ( .A(n22789), .B(n22790), .X(n5696) );
  nand_x1_sg U46241 ( .A(n22795), .B(n22796), .X(n5693) );
  nand_x1_sg U46242 ( .A(n22801), .B(n22802), .X(n5690) );
  nand_x1_sg U46243 ( .A(n22807), .B(n22808), .X(n5687) );
  nand_x1_sg U46244 ( .A(n22813), .B(n22814), .X(n5684) );
  nand_x1_sg U46245 ( .A(n22819), .B(n22820), .X(n5681) );
  nand_x1_sg U46246 ( .A(n22825), .B(n22826), .X(n5678) );
  nand_x1_sg U46247 ( .A(n22831), .B(n22832), .X(n5675) );
  nand_x1_sg U46248 ( .A(n22837), .B(n22838), .X(n5672) );
  nand_x1_sg U46249 ( .A(n22843), .B(n22844), .X(n5669) );
  nand_x1_sg U46250 ( .A(n22849), .B(n22850), .X(n5666) );
  nand_x1_sg U46251 ( .A(n22855), .B(n22856), .X(n5663) );
  nand_x1_sg U46252 ( .A(n22861), .B(n22862), .X(n5660) );
  nand_x1_sg U46253 ( .A(n22867), .B(n22868), .X(n5657) );
  nand_x1_sg U46254 ( .A(n22873), .B(n22874), .X(n5654) );
  nand_x1_sg U46255 ( .A(n22879), .B(n22880), .X(n5651) );
  nand_x1_sg U46256 ( .A(n22885), .B(n22886), .X(n5648) );
  nand_x1_sg U46257 ( .A(n22891), .B(n22892), .X(n5645) );
  nand_x1_sg U46258 ( .A(n22897), .B(n22898), .X(n5642) );
  nand_x1_sg U46259 ( .A(n22903), .B(n22904), .X(n5639) );
  nand_x1_sg U46260 ( .A(n22909), .B(n22910), .X(n5636) );
  nand_x1_sg U46261 ( .A(n22915), .B(n22916), .X(n5633) );
  nand_x1_sg U46262 ( .A(n22921), .B(n22922), .X(n5630) );
  nand_x1_sg U46263 ( .A(n22927), .B(n22928), .X(n5627) );
  nand_x1_sg U46264 ( .A(n22933), .B(n22934), .X(n5624) );
  nand_x1_sg U46265 ( .A(n22939), .B(n22940), .X(n5621) );
  nand_x1_sg U46266 ( .A(n22945), .B(n22946), .X(n5618) );
  nand_x1_sg U46267 ( .A(n22951), .B(n22952), .X(n5615) );
  nand_x1_sg U46268 ( .A(n22957), .B(n22958), .X(n5612) );
  nand_x1_sg U46269 ( .A(n22963), .B(n22964), .X(n5609) );
  nand_x1_sg U46270 ( .A(n22969), .B(n22970), .X(n5606) );
  nand_x1_sg U46271 ( .A(n22975), .B(n22976), .X(n5603) );
  nand_x1_sg U46272 ( .A(n22981), .B(n22982), .X(n5600) );
  nand_x1_sg U46273 ( .A(n22987), .B(n22988), .X(n5597) );
  nand_x1_sg U46274 ( .A(n22993), .B(n22994), .X(n5594) );
  nand_x1_sg U46275 ( .A(n22999), .B(n23000), .X(n5591) );
  nand_x1_sg U46276 ( .A(n23005), .B(n23006), .X(n5588) );
  nand_x1_sg U46277 ( .A(n23011), .B(n23012), .X(n5585) );
  nand_x1_sg U46278 ( .A(n23017), .B(n23018), .X(n5582) );
  nand_x1_sg U46279 ( .A(n23023), .B(n23024), .X(n5579) );
  nand_x1_sg U46280 ( .A(n23029), .B(n23030), .X(n5576) );
  nand_x1_sg U46281 ( .A(n23035), .B(n23036), .X(n5573) );
  nand_x1_sg U46282 ( .A(n23041), .B(n23042), .X(n5570) );
  nand_x1_sg U46283 ( .A(n23047), .B(n23048), .X(n5567) );
  nand_x1_sg U46284 ( .A(n23053), .B(n23054), .X(n5564) );
  nand_x1_sg U46285 ( .A(n23059), .B(n23060), .X(n5561) );
  nand_x1_sg U46286 ( .A(n23065), .B(n23066), .X(n5558) );
  nand_x1_sg U46287 ( .A(n23071), .B(n23072), .X(n5555) );
  nand_x1_sg U46288 ( .A(n23077), .B(n23078), .X(n5552) );
  nand_x1_sg U46289 ( .A(n23083), .B(n23084), .X(n5549) );
  nand_x1_sg U46290 ( .A(n23089), .B(n23090), .X(n5546) );
  nand_x1_sg U46291 ( .A(n23095), .B(n23096), .X(n5543) );
  nand_x1_sg U46292 ( .A(n23101), .B(n23102), .X(n5540) );
  nand_x1_sg U46293 ( .A(n23107), .B(n23108), .X(n5537) );
  nand_x1_sg U46294 ( .A(n23113), .B(n23114), .X(n5534) );
  nand_x1_sg U46295 ( .A(n23119), .B(n23120), .X(n5531) );
  nand_x1_sg U46296 ( .A(n23125), .B(n23126), .X(n5528) );
  nand_x1_sg U46297 ( .A(n23131), .B(n23132), .X(n5525) );
  nand_x1_sg U46298 ( .A(n23137), .B(n23138), .X(n5522) );
  nand_x1_sg U46299 ( .A(n23143), .B(n23144), .X(n5519) );
  nand_x1_sg U46300 ( .A(n23149), .B(n23150), .X(n5516) );
  nand_x1_sg U46301 ( .A(n23155), .B(n23156), .X(n5513) );
  nand_x1_sg U46302 ( .A(n23161), .B(n23162), .X(n5510) );
  nand_x1_sg U46303 ( .A(n23167), .B(n23168), .X(n5507) );
  nand_x1_sg U46304 ( .A(n23173), .B(n23174), .X(n5504) );
  nand_x1_sg U46305 ( .A(n23179), .B(n23180), .X(n5501) );
  nand_x1_sg U46306 ( .A(n23185), .B(n23186), .X(n5498) );
  nand_x1_sg U46307 ( .A(n23191), .B(n23192), .X(n5495) );
  nand_x1_sg U46308 ( .A(n23197), .B(n23198), .X(n5492) );
  nand_x1_sg U46309 ( .A(n23203), .B(n23204), .X(n5489) );
  nand_x1_sg U46310 ( .A(n23209), .B(n23210), .X(n5486) );
  nand_x1_sg U46311 ( .A(n23215), .B(n23216), .X(n5483) );
  nand_x1_sg U46312 ( .A(n23221), .B(n23222), .X(n5480) );
  nand_x1_sg U46313 ( .A(n23227), .B(n23228), .X(n5477) );
  nand_x1_sg U46314 ( .A(n23233), .B(n23234), .X(n5474) );
  nand_x1_sg U46315 ( .A(n23239), .B(n23240), .X(n5471) );
  nand_x1_sg U46316 ( .A(n23245), .B(n23246), .X(n5468) );
  nand_x1_sg U46317 ( .A(n23251), .B(n23252), .X(n5465) );
  nand_x1_sg U46318 ( .A(n23257), .B(n23258), .X(n5462) );
  nand_x1_sg U46319 ( .A(n23263), .B(n23264), .X(n5459) );
  nand_x1_sg U46320 ( .A(n23269), .B(n23270), .X(n5456) );
  nand_x1_sg U46321 ( .A(n23275), .B(n23276), .X(n5453) );
  nand_x1_sg U46322 ( .A(n23281), .B(n23282), .X(n5450) );
  nand_x1_sg U46323 ( .A(n23287), .B(n23288), .X(n5447) );
  nand_x1_sg U46324 ( .A(n23293), .B(n23294), .X(n5444) );
  nand_x1_sg U46325 ( .A(n23299), .B(n23300), .X(n5441) );
  nand_x1_sg U46326 ( .A(n23305), .B(n23306), .X(n5438) );
  nand_x1_sg U46327 ( .A(n23311), .B(n23312), .X(n5435) );
  nand_x1_sg U46328 ( .A(n23317), .B(n23318), .X(n5432) );
  nand_x1_sg U46329 ( .A(n23323), .B(n23324), .X(n5429) );
  nand_x1_sg U46330 ( .A(n23329), .B(n23330), .X(n5426) );
  nand_x1_sg U46331 ( .A(n23335), .B(n23336), .X(n5423) );
  nand_x1_sg U46332 ( .A(n23341), .B(n23342), .X(n5420) );
  nand_x1_sg U46333 ( .A(n23347), .B(n23348), .X(n5417) );
  nand_x1_sg U46334 ( .A(n23353), .B(n23354), .X(n5414) );
  nand_x1_sg U46335 ( .A(n23359), .B(n23360), .X(n5411) );
  nand_x1_sg U46336 ( .A(n23365), .B(n23366), .X(n5408) );
  nand_x1_sg U46337 ( .A(n23371), .B(n23372), .X(n5405) );
  nand_x1_sg U46338 ( .A(n23377), .B(n23378), .X(n5402) );
  nand_x1_sg U46339 ( .A(n23383), .B(n23384), .X(n5399) );
  nand_x1_sg U46340 ( .A(n23389), .B(n23390), .X(n5396) );
  nand_x1_sg U46341 ( .A(n23395), .B(n23396), .X(n5393) );
  nand_x1_sg U46342 ( .A(n23401), .B(n23402), .X(n5390) );
  nand_x1_sg U46343 ( .A(n23407), .B(n23408), .X(n5387) );
  nand_x1_sg U46344 ( .A(n23413), .B(n23414), .X(n5384) );
  nand_x1_sg U46345 ( .A(n23419), .B(n23420), .X(n5381) );
  nand_x1_sg U46346 ( .A(n23425), .B(n23426), .X(n5378) );
  nand_x1_sg U46347 ( .A(n23431), .B(n23432), .X(n5375) );
  nand_x1_sg U46348 ( .A(n23437), .B(n23438), .X(n5372) );
  nand_x1_sg U46349 ( .A(n23443), .B(n23444), .X(n5369) );
  nand_x1_sg U46350 ( .A(n23449), .B(n23450), .X(n5366) );
  nand_x1_sg U46351 ( .A(n23455), .B(n23456), .X(n5363) );
  nand_x1_sg U46352 ( .A(n23461), .B(n23462), .X(n5360) );
  nand_x1_sg U46353 ( .A(n23467), .B(n23468), .X(n5357) );
  nand_x1_sg U46354 ( .A(n23473), .B(n23474), .X(n5354) );
  nand_x1_sg U46355 ( .A(n23479), .B(n23480), .X(n5351) );
  nand_x1_sg U46356 ( .A(n23485), .B(n23486), .X(n5348) );
  nand_x1_sg U46357 ( .A(n23491), .B(n23492), .X(n5345) );
  nand_x1_sg U46358 ( .A(n23497), .B(n23498), .X(n5342) );
  nand_x1_sg U46359 ( .A(n23503), .B(n23504), .X(n5339) );
  nand_x1_sg U46360 ( .A(n23509), .B(n23510), .X(n5336) );
  nand_x1_sg U46361 ( .A(n23515), .B(n23516), .X(n5333) );
  nand_x1_sg U46362 ( .A(n23521), .B(n23522), .X(n5330) );
  nand_x1_sg U46363 ( .A(n23527), .B(n23528), .X(n5327) );
  nand_x1_sg U46364 ( .A(n23533), .B(n23534), .X(n5324) );
  nand_x1_sg U46365 ( .A(n23539), .B(n23540), .X(n5321) );
  nand_x1_sg U46366 ( .A(n23545), .B(n23546), .X(n5318) );
  nand_x1_sg U46367 ( .A(n23551), .B(n23552), .X(n5315) );
  nand_x1_sg U46368 ( .A(n23557), .B(n23558), .X(n5312) );
  nand_x1_sg U46369 ( .A(n23563), .B(n23564), .X(n5309) );
  nand_x1_sg U46370 ( .A(n23569), .B(n23570), .X(n5306) );
  nand_x1_sg U46371 ( .A(n23575), .B(n23576), .X(n5303) );
  nand_x1_sg U46372 ( .A(n23581), .B(n23582), .X(n5300) );
  nand_x1_sg U46373 ( .A(n23587), .B(n23588), .X(n5297) );
  nand_x1_sg U46374 ( .A(n23593), .B(n23594), .X(n5294) );
  nand_x1_sg U46375 ( .A(n23599), .B(n23600), .X(n5291) );
  nand_x1_sg U46376 ( .A(n23605), .B(n23606), .X(n5288) );
  nand_x1_sg U46377 ( .A(n23611), .B(n23612), .X(n5285) );
  nand_x1_sg U46378 ( .A(n23617), .B(n23618), .X(n5282) );
  nand_x1_sg U46379 ( .A(n23623), .B(n23624), .X(n5279) );
  nand_x1_sg U46380 ( .A(n22221), .B(n22222), .X(n5980) );
  nand_x1_sg U46381 ( .A(n22223), .B(n22224), .X(n5979) );
  nand_x1_sg U46382 ( .A(n22227), .B(n22228), .X(n5977) );
  nand_x1_sg U46383 ( .A(n22229), .B(n22230), .X(n5976) );
  nand_x1_sg U46384 ( .A(n22233), .B(n22234), .X(n5974) );
  nand_x1_sg U46385 ( .A(n22235), .B(n22236), .X(n5973) );
  nand_x1_sg U46386 ( .A(n22239), .B(n22240), .X(n5971) );
  nand_x1_sg U46387 ( .A(n22241), .B(n22242), .X(n5970) );
  nand_x1_sg U46388 ( .A(n22245), .B(n22246), .X(n5968) );
  nand_x1_sg U46389 ( .A(n22247), .B(n22248), .X(n5967) );
  nand_x1_sg U46390 ( .A(n22251), .B(n22252), .X(n5965) );
  nand_x1_sg U46391 ( .A(n22253), .B(n22254), .X(n5964) );
  nand_x1_sg U46392 ( .A(n22257), .B(n22258), .X(n5962) );
  nand_x1_sg U46393 ( .A(n22259), .B(n22260), .X(n5961) );
  nand_x1_sg U46394 ( .A(n22263), .B(n22264), .X(n5959) );
  nand_x1_sg U46395 ( .A(n22265), .B(n22266), .X(n5958) );
  nand_x1_sg U46396 ( .A(n22269), .B(n22270), .X(n5956) );
  nand_x1_sg U46397 ( .A(n22271), .B(n22272), .X(n5955) );
  nand_x1_sg U46398 ( .A(n22275), .B(n22276), .X(n5953) );
  nand_x1_sg U46399 ( .A(n22277), .B(n22278), .X(n5952) );
  nand_x1_sg U46400 ( .A(n22281), .B(n22282), .X(n5950) );
  nand_x1_sg U46401 ( .A(n22283), .B(n22284), .X(n5949) );
  nand_x1_sg U46402 ( .A(n22287), .B(n22288), .X(n5947) );
  nand_x1_sg U46403 ( .A(n22289), .B(n22290), .X(n5946) );
  nand_x1_sg U46404 ( .A(n22293), .B(n22294), .X(n5944) );
  nand_x1_sg U46405 ( .A(n22295), .B(n22296), .X(n5943) );
  nand_x1_sg U46406 ( .A(n22299), .B(n22300), .X(n5941) );
  nand_x1_sg U46407 ( .A(n22301), .B(n22302), .X(n5940) );
  nand_x1_sg U46408 ( .A(n22305), .B(n22306), .X(n5938) );
  nand_x1_sg U46409 ( .A(n22307), .B(n22308), .X(n5937) );
  nand_x1_sg U46410 ( .A(n22311), .B(n22312), .X(n5935) );
  nand_x1_sg U46411 ( .A(n22313), .B(n22314), .X(n5934) );
  nand_x1_sg U46412 ( .A(n22317), .B(n22318), .X(n5932) );
  nand_x1_sg U46413 ( .A(n22319), .B(n22320), .X(n5931) );
  nand_x1_sg U46414 ( .A(n22323), .B(n22324), .X(n5929) );
  nand_x1_sg U46415 ( .A(n22325), .B(n22326), .X(n5928) );
  nand_x1_sg U46416 ( .A(n22329), .B(n22330), .X(n5926) );
  nand_x1_sg U46417 ( .A(n22331), .B(n22332), .X(n5925) );
  nand_x1_sg U46418 ( .A(n22335), .B(n22336), .X(n5923) );
  nand_x1_sg U46419 ( .A(n22337), .B(n22338), .X(n5922) );
  nand_x1_sg U46420 ( .A(n22341), .B(n22342), .X(n5920) );
  nand_x1_sg U46421 ( .A(n22343), .B(n22344), .X(n5919) );
  nand_x1_sg U46422 ( .A(n22347), .B(n22348), .X(n5917) );
  nand_x1_sg U46423 ( .A(n22349), .B(n22350), .X(n5916) );
  nand_x1_sg U46424 ( .A(n22353), .B(n22354), .X(n5914) );
  nand_x1_sg U46425 ( .A(n22355), .B(n22356), .X(n5913) );
  nand_x1_sg U46426 ( .A(n22359), .B(n22360), .X(n5911) );
  nand_x1_sg U46427 ( .A(n22361), .B(n22362), .X(n5910) );
  nand_x1_sg U46428 ( .A(n22365), .B(n22366), .X(n5908) );
  nand_x1_sg U46429 ( .A(n22367), .B(n22368), .X(n5907) );
  nand_x1_sg U46430 ( .A(n22371), .B(n22372), .X(n5905) );
  nand_x1_sg U46431 ( .A(n22373), .B(n22374), .X(n5904) );
  nand_x1_sg U46432 ( .A(n22377), .B(n22378), .X(n5902) );
  nand_x1_sg U46433 ( .A(n22379), .B(n22380), .X(n5901) );
  nand_x1_sg U46434 ( .A(n22383), .B(n22384), .X(n5899) );
  nand_x1_sg U46435 ( .A(n22385), .B(n22386), .X(n5898) );
  nand_x1_sg U46436 ( .A(n22389), .B(n22390), .X(n5896) );
  nand_x1_sg U46437 ( .A(n22391), .B(n22392), .X(n5895) );
  nand_x1_sg U46438 ( .A(n22395), .B(n22396), .X(n5893) );
  nand_x1_sg U46439 ( .A(n22397), .B(n22398), .X(n5892) );
  nand_x1_sg U46440 ( .A(n22401), .B(n22402), .X(n5890) );
  nand_x1_sg U46441 ( .A(n22403), .B(n22404), .X(n5889) );
  nand_x1_sg U46442 ( .A(n22407), .B(n22408), .X(n5887) );
  nand_x1_sg U46443 ( .A(n22409), .B(n22410), .X(n5886) );
  nand_x1_sg U46444 ( .A(n22413), .B(n22414), .X(n5884) );
  nand_x1_sg U46445 ( .A(n22415), .B(n22416), .X(n5883) );
  nand_x1_sg U46446 ( .A(n22419), .B(n22420), .X(n5881) );
  nand_x1_sg U46447 ( .A(n22421), .B(n22422), .X(n5880) );
  nand_x1_sg U46448 ( .A(n22425), .B(n22426), .X(n5878) );
  nand_x1_sg U46449 ( .A(n22427), .B(n22428), .X(n5877) );
  nand_x1_sg U46450 ( .A(n22431), .B(n22432), .X(n5875) );
  nand_x1_sg U46451 ( .A(n22433), .B(n22434), .X(n5874) );
  nand_x1_sg U46452 ( .A(n22437), .B(n22438), .X(n5872) );
  nand_x1_sg U46453 ( .A(n22439), .B(n22440), .X(n5871) );
  nand_x1_sg U46454 ( .A(n22443), .B(n22444), .X(n5869) );
  nand_x1_sg U46455 ( .A(n22445), .B(n22446), .X(n5868) );
  nand_x1_sg U46456 ( .A(n22449), .B(n22450), .X(n5866) );
  nand_x1_sg U46457 ( .A(n22451), .B(n22452), .X(n5865) );
  nand_x1_sg U46458 ( .A(n22455), .B(n22456), .X(n5863) );
  nand_x1_sg U46459 ( .A(n22457), .B(n22458), .X(n5862) );
  nand_x1_sg U46460 ( .A(n22461), .B(n22462), .X(n5860) );
  nand_x1_sg U46461 ( .A(n22463), .B(n22464), .X(n5859) );
  nand_x1_sg U46462 ( .A(n22467), .B(n22468), .X(n5857) );
  nand_x1_sg U46463 ( .A(n22469), .B(n22470), .X(n5856) );
  nand_x1_sg U46464 ( .A(n22473), .B(n22474), .X(n5854) );
  nand_x1_sg U46465 ( .A(n22475), .B(n22476), .X(n5853) );
  nand_x1_sg U46466 ( .A(n22479), .B(n22480), .X(n5851) );
  nand_x1_sg U46467 ( .A(n22481), .B(n22482), .X(n5850) );
  nand_x1_sg U46468 ( .A(n22485), .B(n22486), .X(n5848) );
  nand_x1_sg U46469 ( .A(n22487), .B(n22488), .X(n5847) );
  nand_x1_sg U46470 ( .A(n22491), .B(n22492), .X(n5845) );
  nand_x1_sg U46471 ( .A(n22493), .B(n22494), .X(n5844) );
  nand_x1_sg U46472 ( .A(n22497), .B(n22498), .X(n5842) );
  nand_x1_sg U46473 ( .A(n22499), .B(n22500), .X(n5841) );
  nand_x1_sg U46474 ( .A(n22503), .B(n22504), .X(n5839) );
  nand_x1_sg U46475 ( .A(n22505), .B(n22506), .X(n5838) );
  nand_x1_sg U46476 ( .A(n22509), .B(n22510), .X(n5836) );
  nand_x1_sg U46477 ( .A(n22511), .B(n22512), .X(n5835) );
  nand_x1_sg U46478 ( .A(n22515), .B(n22516), .X(n5833) );
  nand_x1_sg U46479 ( .A(n22517), .B(n22518), .X(n5832) );
  nand_x1_sg U46480 ( .A(n22521), .B(n22522), .X(n5830) );
  nand_x1_sg U46481 ( .A(n22523), .B(n22524), .X(n5829) );
  nand_x1_sg U46482 ( .A(n22527), .B(n22528), .X(n5827) );
  nand_x1_sg U46483 ( .A(n22529), .B(n22530), .X(n5826) );
  nand_x1_sg U46484 ( .A(n22533), .B(n22534), .X(n5824) );
  nand_x1_sg U46485 ( .A(n22535), .B(n22536), .X(n5823) );
  nand_x1_sg U46486 ( .A(n22539), .B(n22540), .X(n5821) );
  nand_x1_sg U46487 ( .A(n22541), .B(n22542), .X(n5820) );
  nand_x1_sg U46488 ( .A(n22545), .B(n22546), .X(n5818) );
  nand_x1_sg U46489 ( .A(n22547), .B(n22548), .X(n5817) );
  nand_x1_sg U46490 ( .A(n22551), .B(n22552), .X(n5815) );
  nand_x1_sg U46491 ( .A(n22553), .B(n22554), .X(n5814) );
  nand_x1_sg U46492 ( .A(n22557), .B(n22558), .X(n5812) );
  nand_x1_sg U46493 ( .A(n22559), .B(n22560), .X(n5811) );
  nand_x1_sg U46494 ( .A(n22563), .B(n22564), .X(n5809) );
  nand_x1_sg U46495 ( .A(n22565), .B(n22566), .X(n5808) );
  nand_x1_sg U46496 ( .A(n22569), .B(n22570), .X(n5806) );
  nand_x1_sg U46497 ( .A(n22571), .B(n22572), .X(n5805) );
  nand_x1_sg U46498 ( .A(n22575), .B(n22576), .X(n5803) );
  nand_x1_sg U46499 ( .A(n22577), .B(n22578), .X(n5802) );
  nand_x1_sg U46500 ( .A(n22581), .B(n22582), .X(n5800) );
  nand_x1_sg U46501 ( .A(n22583), .B(n22584), .X(n5799) );
  nand_x1_sg U46502 ( .A(n22587), .B(n22588), .X(n5797) );
  nand_x1_sg U46503 ( .A(n22589), .B(n22590), .X(n5796) );
  nand_x1_sg U46504 ( .A(n22593), .B(n22594), .X(n5794) );
  nand_x1_sg U46505 ( .A(n22595), .B(n22596), .X(n5793) );
  nand_x1_sg U46506 ( .A(n22599), .B(n22600), .X(n5791) );
  nand_x1_sg U46507 ( .A(n22601), .B(n22602), .X(n5790) );
  nand_x1_sg U46508 ( .A(n22605), .B(n22606), .X(n5788) );
  nand_x1_sg U46509 ( .A(n22607), .B(n22608), .X(n5787) );
  nand_x1_sg U46510 ( .A(n22611), .B(n22612), .X(n5785) );
  nand_x1_sg U46511 ( .A(n22613), .B(n22614), .X(n5784) );
  nand_x1_sg U46512 ( .A(n22617), .B(n22618), .X(n5782) );
  nand_x1_sg U46513 ( .A(n22619), .B(n22620), .X(n5781) );
  nand_x1_sg U46514 ( .A(n22623), .B(n22624), .X(n5779) );
  nand_x1_sg U46515 ( .A(n22625), .B(n22626), .X(n5778) );
  nand_x1_sg U46516 ( .A(n22629), .B(n22630), .X(n5776) );
  nand_x1_sg U46517 ( .A(n22631), .B(n22632), .X(n5775) );
  nand_x1_sg U46518 ( .A(n22635), .B(n22636), .X(n5773) );
  nand_x1_sg U46519 ( .A(n22637), .B(n22638), .X(n5772) );
  nand_x1_sg U46520 ( .A(n22641), .B(n22642), .X(n5770) );
  nand_x1_sg U46521 ( .A(n22643), .B(n22644), .X(n5769) );
  nand_x1_sg U46522 ( .A(n22647), .B(n22648), .X(n5767) );
  nand_x1_sg U46523 ( .A(n22649), .B(n22650), .X(n5766) );
  nand_x1_sg U46524 ( .A(n22653), .B(n22654), .X(n5764) );
  nand_x1_sg U46525 ( .A(n22655), .B(n22656), .X(n5763) );
  nand_x1_sg U46526 ( .A(n22659), .B(n22660), .X(n5761) );
  nand_x1_sg U46527 ( .A(n22661), .B(n22662), .X(n5760) );
  nand_x1_sg U46528 ( .A(n22665), .B(n22666), .X(n5758) );
  nand_x1_sg U46529 ( .A(n22667), .B(n22668), .X(n5757) );
  nand_x1_sg U46530 ( .A(n22671), .B(n22672), .X(n5755) );
  nand_x1_sg U46531 ( .A(n22673), .B(n22674), .X(n5754) );
  nand_x1_sg U46532 ( .A(n22677), .B(n22678), .X(n5752) );
  nand_x1_sg U46533 ( .A(n22679), .B(n22680), .X(n5751) );
  nand_x1_sg U46534 ( .A(n22683), .B(n22684), .X(n5749) );
  nand_x1_sg U46535 ( .A(n22685), .B(n22686), .X(n5748) );
  nand_x1_sg U46536 ( .A(n22689), .B(n22690), .X(n5746) );
  nand_x1_sg U46537 ( .A(n22691), .B(n22692), .X(n5745) );
  nand_x1_sg U46538 ( .A(n22695), .B(n22696), .X(n5743) );
  nand_x1_sg U46539 ( .A(n22697), .B(n22698), .X(n5742) );
  nand_x1_sg U46540 ( .A(n22701), .B(n22702), .X(n5740) );
  nand_x1_sg U46541 ( .A(n22703), .B(n22704), .X(n5739) );
  nand_x1_sg U46542 ( .A(n22707), .B(n22708), .X(n5737) );
  nand_x1_sg U46543 ( .A(n22709), .B(n22710), .X(n5736) );
  nand_x1_sg U46544 ( .A(n22713), .B(n22714), .X(n5734) );
  nand_x1_sg U46545 ( .A(n22715), .B(n22716), .X(n5733) );
  nand_x1_sg U46546 ( .A(n22719), .B(n22720), .X(n5731) );
  nand_x1_sg U46547 ( .A(n22721), .B(n22722), .X(n5730) );
  nand_x1_sg U46548 ( .A(n22725), .B(n22726), .X(n5728) );
  nand_x1_sg U46549 ( .A(n22727), .B(n22728), .X(n5727) );
  nand_x1_sg U46550 ( .A(n22731), .B(n22732), .X(n5725) );
  nand_x1_sg U46551 ( .A(n22733), .B(n22734), .X(n5724) );
  nand_x1_sg U46552 ( .A(n22737), .B(n22738), .X(n5722) );
  nand_x1_sg U46553 ( .A(n22739), .B(n22740), .X(n5721) );
  nand_x1_sg U46554 ( .A(n22743), .B(n22744), .X(n5719) );
  nand_x1_sg U46555 ( .A(n22745), .B(n22746), .X(n5718) );
  nand_x1_sg U46556 ( .A(n22749), .B(n22750), .X(n5716) );
  nand_x1_sg U46557 ( .A(n22751), .B(n22752), .X(n5715) );
  nand_x1_sg U46558 ( .A(n22755), .B(n22756), .X(n5713) );
  nand_x1_sg U46559 ( .A(n22757), .B(n22758), .X(n5712) );
  nand_x1_sg U46560 ( .A(n22761), .B(n22762), .X(n5710) );
  nand_x1_sg U46561 ( .A(n22763), .B(n22764), .X(n5709) );
  nand_x1_sg U46562 ( .A(n22767), .B(n22768), .X(n5707) );
  nand_x1_sg U46563 ( .A(n22769), .B(n22770), .X(n5706) );
  nand_x1_sg U46564 ( .A(n22773), .B(n22774), .X(n5704) );
  nand_x1_sg U46565 ( .A(n22775), .B(n22776), .X(n5703) );
  nand_x1_sg U46566 ( .A(n22779), .B(n22780), .X(n5701) );
  nand_x1_sg U46567 ( .A(n22781), .B(n22782), .X(n5700) );
  nand_x1_sg U46568 ( .A(n22785), .B(n22786), .X(n5698) );
  nand_x1_sg U46569 ( .A(n22787), .B(n22788), .X(n5697) );
  nand_x1_sg U46570 ( .A(n22791), .B(n22792), .X(n5695) );
  nand_x1_sg U46571 ( .A(n22793), .B(n22794), .X(n5694) );
  nand_x1_sg U46572 ( .A(n22797), .B(n22798), .X(n5692) );
  nand_x1_sg U46573 ( .A(n22799), .B(n22800), .X(n5691) );
  nand_x1_sg U46574 ( .A(n22803), .B(n22804), .X(n5689) );
  nand_x1_sg U46575 ( .A(n22805), .B(n22806), .X(n5688) );
  nand_x1_sg U46576 ( .A(n22809), .B(n22810), .X(n5686) );
  nand_x1_sg U46577 ( .A(n22811), .B(n22812), .X(n5685) );
  nand_x1_sg U46578 ( .A(n22815), .B(n22816), .X(n5683) );
  nand_x1_sg U46579 ( .A(n22817), .B(n22818), .X(n5682) );
  nand_x1_sg U46580 ( .A(n22821), .B(n22822), .X(n5680) );
  nand_x1_sg U46581 ( .A(n22823), .B(n22824), .X(n5679) );
  nand_x1_sg U46582 ( .A(n22827), .B(n22828), .X(n5677) );
  nand_x1_sg U46583 ( .A(n22829), .B(n22830), .X(n5676) );
  nand_x1_sg U46584 ( .A(n22833), .B(n22834), .X(n5674) );
  nand_x1_sg U46585 ( .A(n22835), .B(n22836), .X(n5673) );
  nand_x1_sg U46586 ( .A(n22839), .B(n22840), .X(n5671) );
  nand_x1_sg U46587 ( .A(n22841), .B(n22842), .X(n5670) );
  nand_x1_sg U46588 ( .A(n22845), .B(n22846), .X(n5668) );
  nand_x1_sg U46589 ( .A(n22847), .B(n22848), .X(n5667) );
  nand_x1_sg U46590 ( .A(n22851), .B(n22852), .X(n5665) );
  nand_x1_sg U46591 ( .A(n22853), .B(n22854), .X(n5664) );
  nand_x1_sg U46592 ( .A(n22857), .B(n22858), .X(n5662) );
  nand_x1_sg U46593 ( .A(n22859), .B(n22860), .X(n5661) );
  nand_x1_sg U46594 ( .A(n22863), .B(n22864), .X(n5659) );
  nand_x1_sg U46595 ( .A(n22865), .B(n22866), .X(n5658) );
  nand_x1_sg U46596 ( .A(n22869), .B(n22870), .X(n5656) );
  nand_x1_sg U46597 ( .A(n22871), .B(n22872), .X(n5655) );
  nand_x1_sg U46598 ( .A(n22875), .B(n22876), .X(n5653) );
  nand_x1_sg U46599 ( .A(n22877), .B(n22878), .X(n5652) );
  nand_x1_sg U46600 ( .A(n22881), .B(n22882), .X(n5650) );
  nand_x1_sg U46601 ( .A(n22883), .B(n22884), .X(n5649) );
  nand_x1_sg U46602 ( .A(n22887), .B(n22888), .X(n5647) );
  nand_x1_sg U46603 ( .A(n22889), .B(n22890), .X(n5646) );
  nand_x1_sg U46604 ( .A(n22893), .B(n22894), .X(n5644) );
  nand_x1_sg U46605 ( .A(n22895), .B(n22896), .X(n5643) );
  nand_x1_sg U46606 ( .A(n22899), .B(n22900), .X(n5641) );
  nand_x1_sg U46607 ( .A(n22901), .B(n22902), .X(n5640) );
  nand_x1_sg U46608 ( .A(n22905), .B(n22906), .X(n5638) );
  nand_x1_sg U46609 ( .A(n22907), .B(n22908), .X(n5637) );
  nand_x1_sg U46610 ( .A(n22911), .B(n22912), .X(n5635) );
  nand_x1_sg U46611 ( .A(n22913), .B(n22914), .X(n5634) );
  nand_x1_sg U46612 ( .A(n22917), .B(n22918), .X(n5632) );
  nand_x1_sg U46613 ( .A(n22919), .B(n22920), .X(n5631) );
  nand_x1_sg U46614 ( .A(n22923), .B(n22924), .X(n5629) );
  nand_x1_sg U46615 ( .A(n22925), .B(n22926), .X(n5628) );
  nand_x1_sg U46616 ( .A(n22929), .B(n22930), .X(n5626) );
  nand_x1_sg U46617 ( .A(n22931), .B(n22932), .X(n5625) );
  nand_x1_sg U46618 ( .A(n22935), .B(n22936), .X(n5623) );
  nand_x1_sg U46619 ( .A(n22937), .B(n22938), .X(n5622) );
  nand_x1_sg U46620 ( .A(n22941), .B(n22942), .X(n5620) );
  nand_x1_sg U46621 ( .A(n22943), .B(n22944), .X(n5619) );
  nand_x1_sg U46622 ( .A(n22947), .B(n22948), .X(n5617) );
  nand_x1_sg U46623 ( .A(n22949), .B(n22950), .X(n5616) );
  nand_x1_sg U46624 ( .A(n22953), .B(n22954), .X(n5614) );
  nand_x1_sg U46625 ( .A(n22955), .B(n22956), .X(n5613) );
  nand_x1_sg U46626 ( .A(n22959), .B(n22960), .X(n5611) );
  nand_x1_sg U46627 ( .A(n22961), .B(n22962), .X(n5610) );
  nand_x1_sg U46628 ( .A(n22965), .B(n22966), .X(n5608) );
  nand_x1_sg U46629 ( .A(n22967), .B(n22968), .X(n5607) );
  nand_x1_sg U46630 ( .A(n22971), .B(n22972), .X(n5605) );
  nand_x1_sg U46631 ( .A(n22973), .B(n22974), .X(n5604) );
  nand_x1_sg U46632 ( .A(n22977), .B(n22978), .X(n5602) );
  nand_x1_sg U46633 ( .A(n22979), .B(n22980), .X(n5601) );
  nand_x1_sg U46634 ( .A(n22983), .B(n22984), .X(n5599) );
  nand_x1_sg U46635 ( .A(n22985), .B(n22986), .X(n5598) );
  nand_x1_sg U46636 ( .A(n22989), .B(n22990), .X(n5596) );
  nand_x1_sg U46637 ( .A(n22991), .B(n22992), .X(n5595) );
  nand_x1_sg U46638 ( .A(n22995), .B(n22996), .X(n5593) );
  nand_x1_sg U46639 ( .A(n22997), .B(n22998), .X(n5592) );
  nand_x1_sg U46640 ( .A(n23001), .B(n23002), .X(n5590) );
  nand_x1_sg U46641 ( .A(n23003), .B(n23004), .X(n5589) );
  nand_x1_sg U46642 ( .A(n23007), .B(n23008), .X(n5587) );
  nand_x1_sg U46643 ( .A(n23009), .B(n23010), .X(n5586) );
  nand_x1_sg U46644 ( .A(n23013), .B(n23014), .X(n5584) );
  nand_x1_sg U46645 ( .A(n23015), .B(n23016), .X(n5583) );
  nand_x1_sg U46646 ( .A(n23019), .B(n23020), .X(n5581) );
  nand_x1_sg U46647 ( .A(n23021), .B(n23022), .X(n5580) );
  nand_x1_sg U46648 ( .A(n23025), .B(n23026), .X(n5578) );
  nand_x1_sg U46649 ( .A(n23027), .B(n23028), .X(n5577) );
  nand_x1_sg U46650 ( .A(n23031), .B(n23032), .X(n5575) );
  nand_x1_sg U46651 ( .A(n23033), .B(n23034), .X(n5574) );
  nand_x1_sg U46652 ( .A(n23037), .B(n23038), .X(n5572) );
  nand_x1_sg U46653 ( .A(n23039), .B(n23040), .X(n5571) );
  nand_x1_sg U46654 ( .A(n23043), .B(n23044), .X(n5569) );
  nand_x1_sg U46655 ( .A(n23045), .B(n23046), .X(n5568) );
  nand_x1_sg U46656 ( .A(n23049), .B(n23050), .X(n5566) );
  nand_x1_sg U46657 ( .A(n23051), .B(n23052), .X(n5565) );
  nand_x1_sg U46658 ( .A(n23055), .B(n23056), .X(n5563) );
  nand_x1_sg U46659 ( .A(n23057), .B(n23058), .X(n5562) );
  nand_x1_sg U46660 ( .A(n23061), .B(n23062), .X(n5560) );
  nand_x1_sg U46661 ( .A(n23063), .B(n23064), .X(n5559) );
  nand_x1_sg U46662 ( .A(n23067), .B(n23068), .X(n5557) );
  nand_x1_sg U46663 ( .A(n23069), .B(n23070), .X(n5556) );
  nand_x1_sg U46664 ( .A(n23073), .B(n23074), .X(n5554) );
  nand_x1_sg U46665 ( .A(n23075), .B(n23076), .X(n5553) );
  nand_x1_sg U46666 ( .A(n23079), .B(n23080), .X(n5551) );
  nand_x1_sg U46667 ( .A(n23081), .B(n23082), .X(n5550) );
  nand_x1_sg U46668 ( .A(n23085), .B(n23086), .X(n5548) );
  nand_x1_sg U46669 ( .A(n23087), .B(n23088), .X(n5547) );
  nand_x1_sg U46670 ( .A(n23091), .B(n23092), .X(n5545) );
  nand_x1_sg U46671 ( .A(n23093), .B(n23094), .X(n5544) );
  nand_x1_sg U46672 ( .A(n23097), .B(n23098), .X(n5542) );
  nand_x1_sg U46673 ( .A(n23099), .B(n23100), .X(n5541) );
  nand_x1_sg U46674 ( .A(n23103), .B(n23104), .X(n5539) );
  nand_x1_sg U46675 ( .A(n23105), .B(n23106), .X(n5538) );
  nand_x1_sg U46676 ( .A(n23109), .B(n23110), .X(n5536) );
  nand_x1_sg U46677 ( .A(n23111), .B(n23112), .X(n5535) );
  nand_x1_sg U46678 ( .A(n23115), .B(n23116), .X(n5533) );
  nand_x1_sg U46679 ( .A(n23117), .B(n23118), .X(n5532) );
  nand_x1_sg U46680 ( .A(n23121), .B(n23122), .X(n5530) );
  nand_x1_sg U46681 ( .A(n23123), .B(n23124), .X(n5529) );
  nand_x1_sg U46682 ( .A(n23127), .B(n23128), .X(n5527) );
  nand_x1_sg U46683 ( .A(n23129), .B(n23130), .X(n5526) );
  nand_x1_sg U46684 ( .A(n23133), .B(n23134), .X(n5524) );
  nand_x1_sg U46685 ( .A(n23135), .B(n23136), .X(n5523) );
  nand_x1_sg U46686 ( .A(n23139), .B(n23140), .X(n5521) );
  nand_x1_sg U46687 ( .A(n23141), .B(n23142), .X(n5520) );
  nand_x1_sg U46688 ( .A(n23145), .B(n23146), .X(n5518) );
  nand_x1_sg U46689 ( .A(n23147), .B(n23148), .X(n5517) );
  nand_x1_sg U46690 ( .A(n23151), .B(n23152), .X(n5515) );
  nand_x1_sg U46691 ( .A(n23153), .B(n23154), .X(n5514) );
  nand_x1_sg U46692 ( .A(n23157), .B(n23158), .X(n5512) );
  nand_x1_sg U46693 ( .A(n23159), .B(n23160), .X(n5511) );
  nand_x1_sg U46694 ( .A(n23163), .B(n23164), .X(n5509) );
  nand_x1_sg U46695 ( .A(n23165), .B(n23166), .X(n5508) );
  nand_x1_sg U46696 ( .A(n23169), .B(n23170), .X(n5506) );
  nand_x1_sg U46697 ( .A(n23171), .B(n23172), .X(n5505) );
  nand_x1_sg U46698 ( .A(n23175), .B(n23176), .X(n5503) );
  nand_x1_sg U46699 ( .A(n23177), .B(n23178), .X(n5502) );
  nand_x1_sg U46700 ( .A(n23181), .B(n23182), .X(n5500) );
  nand_x1_sg U46701 ( .A(n23183), .B(n23184), .X(n5499) );
  nand_x1_sg U46702 ( .A(n23187), .B(n23188), .X(n5497) );
  nand_x1_sg U46703 ( .A(n23189), .B(n23190), .X(n5496) );
  nand_x1_sg U46704 ( .A(n23193), .B(n23194), .X(n5494) );
  nand_x1_sg U46705 ( .A(n23195), .B(n23196), .X(n5493) );
  nand_x1_sg U46706 ( .A(n23199), .B(n23200), .X(n5491) );
  nand_x1_sg U46707 ( .A(n23201), .B(n23202), .X(n5490) );
  nand_x1_sg U46708 ( .A(n23205), .B(n23206), .X(n5488) );
  nand_x1_sg U46709 ( .A(n23207), .B(n23208), .X(n5487) );
  nand_x1_sg U46710 ( .A(n23211), .B(n23212), .X(n5485) );
  nand_x1_sg U46711 ( .A(n23213), .B(n23214), .X(n5484) );
  nand_x1_sg U46712 ( .A(n23217), .B(n23218), .X(n5482) );
  nand_x1_sg U46713 ( .A(n23219), .B(n23220), .X(n5481) );
  nand_x1_sg U46714 ( .A(n23223), .B(n23224), .X(n5479) );
  nand_x1_sg U46715 ( .A(n23225), .B(n23226), .X(n5478) );
  nand_x1_sg U46716 ( .A(n23229), .B(n23230), .X(n5476) );
  nand_x1_sg U46717 ( .A(n23231), .B(n23232), .X(n5475) );
  nand_x1_sg U46718 ( .A(n23235), .B(n23236), .X(n5473) );
  nand_x1_sg U46719 ( .A(n23237), .B(n23238), .X(n5472) );
  nand_x1_sg U46720 ( .A(n23241), .B(n23242), .X(n5470) );
  nand_x1_sg U46721 ( .A(n23243), .B(n23244), .X(n5469) );
  nand_x1_sg U46722 ( .A(n23247), .B(n23248), .X(n5467) );
  nand_x1_sg U46723 ( .A(n23249), .B(n23250), .X(n5466) );
  nand_x1_sg U46724 ( .A(n23253), .B(n23254), .X(n5464) );
  nand_x1_sg U46725 ( .A(n23255), .B(n23256), .X(n5463) );
  nand_x1_sg U46726 ( .A(n23259), .B(n23260), .X(n5461) );
  nand_x1_sg U46727 ( .A(n23261), .B(n23262), .X(n5460) );
  nand_x1_sg U46728 ( .A(n23265), .B(n23266), .X(n5458) );
  nand_x1_sg U46729 ( .A(n23267), .B(n23268), .X(n5457) );
  nand_x1_sg U46730 ( .A(n23271), .B(n23272), .X(n5455) );
  nand_x1_sg U46731 ( .A(n23273), .B(n23274), .X(n5454) );
  nand_x1_sg U46732 ( .A(n23277), .B(n23278), .X(n5452) );
  nand_x1_sg U46733 ( .A(n23279), .B(n23280), .X(n5451) );
  nand_x1_sg U46734 ( .A(n23283), .B(n23284), .X(n5449) );
  nand_x1_sg U46735 ( .A(n23285), .B(n23286), .X(n5448) );
  nand_x1_sg U46736 ( .A(n23289), .B(n23290), .X(n5446) );
  nand_x1_sg U46737 ( .A(n23291), .B(n23292), .X(n5445) );
  nand_x1_sg U46738 ( .A(n23295), .B(n23296), .X(n5443) );
  nand_x1_sg U46739 ( .A(n23297), .B(n23298), .X(n5442) );
  nand_x1_sg U46740 ( .A(n23301), .B(n23302), .X(n5440) );
  nand_x1_sg U46741 ( .A(n23303), .B(n23304), .X(n5439) );
  nand_x1_sg U46742 ( .A(n23307), .B(n23308), .X(n5437) );
  nand_x1_sg U46743 ( .A(n23309), .B(n23310), .X(n5436) );
  nand_x1_sg U46744 ( .A(n23313), .B(n23314), .X(n5434) );
  nand_x1_sg U46745 ( .A(n23315), .B(n23316), .X(n5433) );
  nand_x1_sg U46746 ( .A(n23319), .B(n23320), .X(n5431) );
  nand_x1_sg U46747 ( .A(n23321), .B(n23322), .X(n5430) );
  nand_x1_sg U46748 ( .A(n23325), .B(n23326), .X(n5428) );
  nand_x1_sg U46749 ( .A(n23327), .B(n23328), .X(n5427) );
  nand_x1_sg U46750 ( .A(n23331), .B(n23332), .X(n5425) );
  nand_x1_sg U46751 ( .A(n23333), .B(n23334), .X(n5424) );
  nand_x1_sg U46752 ( .A(n23337), .B(n23338), .X(n5422) );
  nand_x1_sg U46753 ( .A(n23339), .B(n23340), .X(n5421) );
  nand_x1_sg U46754 ( .A(n23343), .B(n23344), .X(n5419) );
  nand_x1_sg U46755 ( .A(n23345), .B(n23346), .X(n5418) );
  nand_x1_sg U46756 ( .A(n23349), .B(n23350), .X(n5416) );
  nand_x1_sg U46757 ( .A(n23351), .B(n23352), .X(n5415) );
  nand_x1_sg U46758 ( .A(n23355), .B(n23356), .X(n5413) );
  nand_x1_sg U46759 ( .A(n23357), .B(n23358), .X(n5412) );
  nand_x1_sg U46760 ( .A(n23361), .B(n23362), .X(n5410) );
  nand_x1_sg U46761 ( .A(n23363), .B(n23364), .X(n5409) );
  nand_x1_sg U46762 ( .A(n23367), .B(n23368), .X(n5407) );
  nand_x1_sg U46763 ( .A(n23369), .B(n23370), .X(n5406) );
  nand_x1_sg U46764 ( .A(n23373), .B(n23374), .X(n5404) );
  nand_x1_sg U46765 ( .A(n23375), .B(n23376), .X(n5403) );
  nand_x1_sg U46766 ( .A(n23379), .B(n23380), .X(n5401) );
  nand_x1_sg U46767 ( .A(n23381), .B(n23382), .X(n5400) );
  nand_x1_sg U46768 ( .A(n23385), .B(n23386), .X(n5398) );
  nand_x1_sg U46769 ( .A(n23387), .B(n23388), .X(n5397) );
  nand_x1_sg U46770 ( .A(n23391), .B(n23392), .X(n5395) );
  nand_x1_sg U46771 ( .A(n23393), .B(n23394), .X(n5394) );
  nand_x1_sg U46772 ( .A(n23397), .B(n23398), .X(n5392) );
  nand_x1_sg U46773 ( .A(n23399), .B(n23400), .X(n5391) );
  nand_x1_sg U46774 ( .A(n23403), .B(n23404), .X(n5389) );
  nand_x1_sg U46775 ( .A(n23405), .B(n23406), .X(n5388) );
  nand_x1_sg U46776 ( .A(n23409), .B(n23410), .X(n5386) );
  nand_x1_sg U46777 ( .A(n23411), .B(n23412), .X(n5385) );
  nand_x1_sg U46778 ( .A(n23415), .B(n23416), .X(n5383) );
  nand_x1_sg U46779 ( .A(n23417), .B(n23418), .X(n5382) );
  nand_x1_sg U46780 ( .A(n23421), .B(n23422), .X(n5380) );
  nand_x1_sg U46781 ( .A(n23423), .B(n23424), .X(n5379) );
  nand_x1_sg U46782 ( .A(n23427), .B(n23428), .X(n5377) );
  nand_x1_sg U46783 ( .A(n23429), .B(n23430), .X(n5376) );
  nand_x1_sg U46784 ( .A(n23433), .B(n23434), .X(n5374) );
  nand_x1_sg U46785 ( .A(n23435), .B(n23436), .X(n5373) );
  nand_x1_sg U46786 ( .A(n23439), .B(n23440), .X(n5371) );
  nand_x1_sg U46787 ( .A(n23441), .B(n23442), .X(n5370) );
  nand_x1_sg U46788 ( .A(n23445), .B(n23446), .X(n5368) );
  nand_x1_sg U46789 ( .A(n23447), .B(n23448), .X(n5367) );
  nand_x1_sg U46790 ( .A(n23451), .B(n23452), .X(n5365) );
  nand_x1_sg U46791 ( .A(n23453), .B(n23454), .X(n5364) );
  nand_x1_sg U46792 ( .A(n23457), .B(n23458), .X(n5362) );
  nand_x1_sg U46793 ( .A(n23459), .B(n23460), .X(n5361) );
  nand_x1_sg U46794 ( .A(n23463), .B(n23464), .X(n5359) );
  nand_x1_sg U46795 ( .A(n23465), .B(n23466), .X(n5358) );
  nand_x1_sg U46796 ( .A(n23469), .B(n23470), .X(n5356) );
  nand_x1_sg U46797 ( .A(n23471), .B(n23472), .X(n5355) );
  nand_x1_sg U46798 ( .A(n23475), .B(n23476), .X(n5353) );
  nand_x1_sg U46799 ( .A(n23477), .B(n23478), .X(n5352) );
  nand_x1_sg U46800 ( .A(n23481), .B(n23482), .X(n5350) );
  nand_x1_sg U46801 ( .A(n23483), .B(n23484), .X(n5349) );
  nand_x1_sg U46802 ( .A(n23487), .B(n23488), .X(n5347) );
  nand_x1_sg U46803 ( .A(n23489), .B(n23490), .X(n5346) );
  nand_x1_sg U46804 ( .A(n23493), .B(n23494), .X(n5344) );
  nand_x1_sg U46805 ( .A(n23495), .B(n23496), .X(n5343) );
  nand_x1_sg U46806 ( .A(n23499), .B(n23500), .X(n5341) );
  nand_x1_sg U46807 ( .A(n23501), .B(n23502), .X(n5340) );
  nand_x1_sg U46808 ( .A(n23505), .B(n23506), .X(n5338) );
  nand_x1_sg U46809 ( .A(n23507), .B(n23508), .X(n5337) );
  nand_x1_sg U46810 ( .A(n23511), .B(n23512), .X(n5335) );
  nand_x1_sg U46811 ( .A(n23513), .B(n23514), .X(n5334) );
  nand_x1_sg U46812 ( .A(n23517), .B(n23518), .X(n5332) );
  nand_x1_sg U46813 ( .A(n23519), .B(n23520), .X(n5331) );
  nand_x1_sg U46814 ( .A(n23523), .B(n23524), .X(n5329) );
  nand_x1_sg U46815 ( .A(n23525), .B(n23526), .X(n5328) );
  nand_x1_sg U46816 ( .A(n23529), .B(n23530), .X(n5326) );
  nand_x1_sg U46817 ( .A(n23531), .B(n23532), .X(n5325) );
  nand_x1_sg U46818 ( .A(n23535), .B(n23536), .X(n5323) );
  nand_x1_sg U46819 ( .A(n23537), .B(n23538), .X(n5322) );
  nand_x1_sg U46820 ( .A(n23541), .B(n23542), .X(n5320) );
  nand_x1_sg U46821 ( .A(n23543), .B(n23544), .X(n5319) );
  nand_x1_sg U46822 ( .A(n23547), .B(n23548), .X(n5317) );
  nand_x1_sg U46823 ( .A(n23549), .B(n23550), .X(n5316) );
  nand_x1_sg U46824 ( .A(n23553), .B(n23554), .X(n5314) );
  nand_x1_sg U46825 ( .A(n23555), .B(n23556), .X(n5313) );
  nand_x1_sg U46826 ( .A(n23559), .B(n23560), .X(n5311) );
  nand_x1_sg U46827 ( .A(n23561), .B(n23562), .X(n5310) );
  nand_x1_sg U46828 ( .A(n23565), .B(n23566), .X(n5308) );
  nand_x1_sg U46829 ( .A(n23567), .B(n23568), .X(n5307) );
  nand_x1_sg U46830 ( .A(n23571), .B(n23572), .X(n5305) );
  nand_x1_sg U46831 ( .A(n23573), .B(n23574), .X(n5304) );
  nand_x1_sg U46832 ( .A(n23577), .B(n23578), .X(n5302) );
  nand_x1_sg U46833 ( .A(n23579), .B(n23580), .X(n5301) );
  nand_x1_sg U46834 ( .A(n23583), .B(n23584), .X(n5299) );
  nand_x1_sg U46835 ( .A(n23585), .B(n23586), .X(n5298) );
  nand_x1_sg U46836 ( .A(n23589), .B(n23590), .X(n5296) );
  nand_x1_sg U46837 ( .A(n23591), .B(n23592), .X(n5295) );
  nand_x1_sg U46838 ( .A(n23595), .B(n23596), .X(n5293) );
  nand_x1_sg U46839 ( .A(n23597), .B(n23598), .X(n5292) );
  nand_x1_sg U46840 ( .A(n23601), .B(n23602), .X(n5290) );
  nand_x1_sg U46841 ( .A(n23603), .B(n23604), .X(n5289) );
  nand_x1_sg U46842 ( .A(n23607), .B(n23608), .X(n5287) );
  nand_x1_sg U46843 ( .A(n23609), .B(n23610), .X(n5286) );
  nand_x1_sg U46844 ( .A(n23613), .B(n23614), .X(n5284) );
  nand_x1_sg U46845 ( .A(n23615), .B(n23616), .X(n5283) );
  nand_x1_sg U46846 ( .A(n23619), .B(n23620), .X(n5281) );
  nand_x1_sg U46847 ( .A(n23621), .B(n23622), .X(n5280) );
  nand_x1_sg U46848 ( .A(n23625), .B(n23626), .X(n5278) );
  nand_x1_sg U46849 ( .A(n23627), .B(n23628), .X(n5277) );
  nand_x1_sg U46850 ( .A(n22212), .B(n22213), .X(n5982) );
  nand_x1_sg U46851 ( .A(n23629), .B(n23630), .X(n5276) );
  nand_x1_sg U46852 ( .A(n20895), .B(n20896), .X(\shifter_0/n10241 ) );
  nand_x1_sg U46853 ( .A(n20571), .B(n20572), .X(\shifter_0/n10402 ) );
  nand_x1_sg U46854 ( .A(n20569), .B(n20570), .X(\shifter_0/n10403 ) );
  nand_x1_sg U46855 ( .A(n20567), .B(n20568), .X(\shifter_0/n10404 ) );
  nand_x1_sg U46856 ( .A(n20565), .B(n20566), .X(\shifter_0/n10405 ) );
  nand_x1_sg U46857 ( .A(n20563), .B(n20564), .X(\shifter_0/n10406 ) );
  nand_x1_sg U46858 ( .A(n20561), .B(n20562), .X(\shifter_0/n10407 ) );
  nand_x1_sg U46859 ( .A(n20559), .B(n20560), .X(\shifter_0/n10408 ) );
  nand_x1_sg U46860 ( .A(n20557), .B(n20558), .X(\shifter_0/n10409 ) );
  nand_x1_sg U46861 ( .A(n20537), .B(n20538), .X(\shifter_0/n10419 ) );
  nand_x1_sg U46862 ( .A(n20535), .B(n20536), .X(\shifter_0/n10420 ) );
  nand_x1_sg U46863 ( .A(n20533), .B(n20534), .X(\shifter_0/n10421 ) );
  nand_x1_sg U46864 ( .A(n19925), .B(n19926), .X(\shifter_0/n10725 ) );
  nand_x1_sg U46865 ( .A(n19923), .B(n19924), .X(\shifter_0/n10726 ) );
  nand_x1_sg U46866 ( .A(n19921), .B(n19922), .X(\shifter_0/n10727 ) );
  nand_x1_sg U46867 ( .A(n19919), .B(n19920), .X(\shifter_0/n10728 ) );
  nand_x1_sg U46868 ( .A(n19917), .B(n19918), .X(\shifter_0/n10729 ) );
  nand_x1_sg U46869 ( .A(n19915), .B(n19916), .X(\shifter_0/n10730 ) );
  nand_x1_sg U46870 ( .A(n19913), .B(n19914), .X(\shifter_0/n10731 ) );
  nand_x1_sg U46871 ( .A(n19911), .B(n19912), .X(\shifter_0/n10732 ) );
  nand_x1_sg U46872 ( .A(n19909), .B(n19910), .X(\shifter_0/n10733 ) );
  nand_x1_sg U46873 ( .A(n19907), .B(n19908), .X(\shifter_0/n10734 ) );
  nand_x1_sg U46874 ( .A(n19905), .B(n19906), .X(\shifter_0/n10735 ) );
  nand_x1_sg U46875 ( .A(n19903), .B(n19904), .X(\shifter_0/n10736 ) );
  nand_x1_sg U46876 ( .A(n19899), .B(n19900), .X(\shifter_0/n10738 ) );
  nand_x1_sg U46877 ( .A(n19895), .B(n19896), .X(\shifter_0/n10740 ) );
  nand_x1_sg U46878 ( .A(n19893), .B(n19894), .X(\shifter_0/n10741 ) );
  nand_x1_sg U46879 ( .A(n20891), .B(n20892), .X(\shifter_0/n10242 ) );
  nand_x1_sg U46880 ( .A(n20889), .B(n20890), .X(\shifter_0/n10243 ) );
  nand_x1_sg U46881 ( .A(n20887), .B(n20888), .X(\shifter_0/n10244 ) );
  nand_x1_sg U46882 ( .A(n20885), .B(n20886), .X(\shifter_0/n10245 ) );
  nand_x1_sg U46883 ( .A(n20883), .B(n20884), .X(\shifter_0/n10246 ) );
  nand_x1_sg U46884 ( .A(n20881), .B(n20882), .X(\shifter_0/n10247 ) );
  nand_x1_sg U46885 ( .A(n20879), .B(n20880), .X(\shifter_0/n10248 ) );
  nand_x1_sg U46886 ( .A(n20877), .B(n20878), .X(\shifter_0/n10249 ) );
  nand_x1_sg U46887 ( .A(n20875), .B(n20876), .X(\shifter_0/n10250 ) );
  nand_x1_sg U46888 ( .A(n20873), .B(n20874), .X(\shifter_0/n10251 ) );
  nand_x1_sg U46889 ( .A(n20871), .B(n20872), .X(\shifter_0/n10252 ) );
  nand_x1_sg U46890 ( .A(n20869), .B(n20870), .X(\shifter_0/n10253 ) );
  nand_x1_sg U46891 ( .A(n20867), .B(n20868), .X(\shifter_0/n10254 ) );
  nand_x1_sg U46892 ( .A(n20865), .B(n20866), .X(\shifter_0/n10255 ) );
  nand_x1_sg U46893 ( .A(n20863), .B(n20864), .X(\shifter_0/n10256 ) );
  nand_x1_sg U46894 ( .A(n20861), .B(n20862), .X(\shifter_0/n10257 ) );
  nand_x1_sg U46895 ( .A(n20859), .B(n20860), .X(\shifter_0/n10258 ) );
  nand_x1_sg U46896 ( .A(n20857), .B(n20858), .X(\shifter_0/n10259 ) );
  nand_x1_sg U46897 ( .A(n20855), .B(n20856), .X(\shifter_0/n10260 ) );
  nand_x1_sg U46898 ( .A(n20853), .B(n20854), .X(\shifter_0/n10261 ) );
  nand_x1_sg U46899 ( .A(n20851), .B(n20852), .X(\shifter_0/n10262 ) );
  nand_x1_sg U46900 ( .A(n20849), .B(n20850), .X(\shifter_0/n10263 ) );
  nand_x1_sg U46901 ( .A(n20847), .B(n20848), .X(\shifter_0/n10264 ) );
  nand_x1_sg U46902 ( .A(n20845), .B(n20846), .X(\shifter_0/n10265 ) );
  nand_x1_sg U46903 ( .A(n20843), .B(n20844), .X(\shifter_0/n10266 ) );
  nand_x1_sg U46904 ( .A(n20841), .B(n20842), .X(\shifter_0/n10267 ) );
  nand_x1_sg U46905 ( .A(n20839), .B(n20840), .X(\shifter_0/n10268 ) );
  nand_x1_sg U46906 ( .A(n20837), .B(n20838), .X(\shifter_0/n10269 ) );
  nand_x1_sg U46907 ( .A(n20835), .B(n20836), .X(\shifter_0/n10270 ) );
  nand_x1_sg U46908 ( .A(n20833), .B(n20834), .X(\shifter_0/n10271 ) );
  nand_x1_sg U46909 ( .A(n20831), .B(n20832), .X(\shifter_0/n10272 ) );
  nand_x1_sg U46910 ( .A(n20829), .B(n20830), .X(\shifter_0/n10273 ) );
  nand_x1_sg U46911 ( .A(n20827), .B(n20828), .X(\shifter_0/n10274 ) );
  nand_x1_sg U46912 ( .A(n20825), .B(n20826), .X(\shifter_0/n10275 ) );
  nand_x1_sg U46913 ( .A(n20823), .B(n20824), .X(\shifter_0/n10276 ) );
  nand_x1_sg U46914 ( .A(n20821), .B(n20822), .X(\shifter_0/n10277 ) );
  nand_x1_sg U46915 ( .A(n20819), .B(n20820), .X(\shifter_0/n10278 ) );
  nand_x1_sg U46916 ( .A(n20817), .B(n20818), .X(\shifter_0/n10279 ) );
  nand_x1_sg U46917 ( .A(n20815), .B(n20816), .X(\shifter_0/n10280 ) );
  nand_x1_sg U46918 ( .A(n20813), .B(n20814), .X(\shifter_0/n10281 ) );
  nand_x1_sg U46919 ( .A(n20811), .B(n20812), .X(\shifter_0/n10282 ) );
  nand_x1_sg U46920 ( .A(n20809), .B(n20810), .X(\shifter_0/n10283 ) );
  nand_x1_sg U46921 ( .A(n20807), .B(n20808), .X(\shifter_0/n10284 ) );
  nand_x1_sg U46922 ( .A(n20805), .B(n20806), .X(\shifter_0/n10285 ) );
  nand_x1_sg U46923 ( .A(n20803), .B(n20804), .X(\shifter_0/n10286 ) );
  nand_x1_sg U46924 ( .A(n20801), .B(n20802), .X(\shifter_0/n10287 ) );
  nand_x1_sg U46925 ( .A(n20799), .B(n20800), .X(\shifter_0/n10288 ) );
  nand_x1_sg U46926 ( .A(n20797), .B(n20798), .X(\shifter_0/n10289 ) );
  nand_x1_sg U46927 ( .A(n20795), .B(n20796), .X(\shifter_0/n10290 ) );
  nand_x1_sg U46928 ( .A(n20773), .B(n20774), .X(\shifter_0/n10301 ) );
  nand_x1_sg U46929 ( .A(n20771), .B(n20772), .X(\shifter_0/n10302 ) );
  nand_x1_sg U46930 ( .A(n20769), .B(n20770), .X(\shifter_0/n10303 ) );
  nand_x1_sg U46931 ( .A(n20767), .B(n20768), .X(\shifter_0/n10304 ) );
  nand_x1_sg U46932 ( .A(n20765), .B(n20766), .X(\shifter_0/n10305 ) );
  nand_x1_sg U46933 ( .A(n20763), .B(n20764), .X(\shifter_0/n10306 ) );
  nand_x1_sg U46934 ( .A(n20761), .B(n20762), .X(\shifter_0/n10307 ) );
  nand_x1_sg U46935 ( .A(n20759), .B(n20760), .X(\shifter_0/n10308 ) );
  nand_x1_sg U46936 ( .A(n20757), .B(n20758), .X(\shifter_0/n10309 ) );
  nand_x1_sg U46937 ( .A(n20755), .B(n20756), .X(\shifter_0/n10310 ) );
  nand_x1_sg U46938 ( .A(n20753), .B(n20754), .X(\shifter_0/n10311 ) );
  nand_x1_sg U46939 ( .A(n20751), .B(n20752), .X(\shifter_0/n10312 ) );
  nand_x1_sg U46940 ( .A(n20749), .B(n20750), .X(\shifter_0/n10313 ) );
  nand_x1_sg U46941 ( .A(n20747), .B(n20748), .X(\shifter_0/n10314 ) );
  nand_x1_sg U46942 ( .A(n20745), .B(n20746), .X(\shifter_0/n10315 ) );
  nand_x1_sg U46943 ( .A(n20743), .B(n20744), .X(\shifter_0/n10316 ) );
  nand_x1_sg U46944 ( .A(n20741), .B(n20742), .X(\shifter_0/n10317 ) );
  nand_x1_sg U46945 ( .A(n20739), .B(n20740), .X(\shifter_0/n10318 ) );
  nand_x1_sg U46946 ( .A(n20737), .B(n20738), .X(\shifter_0/n10319 ) );
  nand_x1_sg U46947 ( .A(n20735), .B(n20736), .X(\shifter_0/n10320 ) );
  nand_x1_sg U46948 ( .A(n20733), .B(n20734), .X(\shifter_0/n10321 ) );
  nand_x1_sg U46949 ( .A(n20731), .B(n20732), .X(\shifter_0/n10322 ) );
  nand_x1_sg U46950 ( .A(n20729), .B(n20730), .X(\shifter_0/n10323 ) );
  nand_x1_sg U46951 ( .A(n20727), .B(n20728), .X(\shifter_0/n10324 ) );
  nand_x1_sg U46952 ( .A(n20725), .B(n20726), .X(\shifter_0/n10325 ) );
  nand_x1_sg U46953 ( .A(n20723), .B(n20724), .X(\shifter_0/n10326 ) );
  nand_x1_sg U46954 ( .A(n20721), .B(n20722), .X(\shifter_0/n10327 ) );
  nand_x1_sg U46955 ( .A(n20719), .B(n20720), .X(\shifter_0/n10328 ) );
  nand_x1_sg U46956 ( .A(n20717), .B(n20718), .X(\shifter_0/n10329 ) );
  nand_x1_sg U46957 ( .A(n20715), .B(n20716), .X(\shifter_0/n10330 ) );
  nand_x1_sg U46958 ( .A(n20713), .B(n20714), .X(\shifter_0/n10331 ) );
  nand_x1_sg U46959 ( .A(n20711), .B(n20712), .X(\shifter_0/n10332 ) );
  nand_x1_sg U46960 ( .A(n20693), .B(n20694), .X(\shifter_0/n10341 ) );
  nand_x1_sg U46961 ( .A(n20691), .B(n20692), .X(\shifter_0/n10342 ) );
  nand_x1_sg U46962 ( .A(n20689), .B(n20690), .X(\shifter_0/n10343 ) );
  nand_x1_sg U46963 ( .A(n20687), .B(n20688), .X(\shifter_0/n10344 ) );
  nand_x1_sg U46964 ( .A(n20685), .B(n20686), .X(\shifter_0/n10345 ) );
  nand_x1_sg U46965 ( .A(n20683), .B(n20684), .X(\shifter_0/n10346 ) );
  nand_x1_sg U46966 ( .A(n20681), .B(n20682), .X(\shifter_0/n10347 ) );
  nand_x1_sg U46967 ( .A(n20679), .B(n20680), .X(\shifter_0/n10348 ) );
  nand_x1_sg U46968 ( .A(n20677), .B(n20678), .X(\shifter_0/n10349 ) );
  nand_x1_sg U46969 ( .A(n20675), .B(n20676), .X(\shifter_0/n10350 ) );
  nand_x1_sg U46970 ( .A(n20655), .B(n20656), .X(\shifter_0/n10360 ) );
  nand_x1_sg U46971 ( .A(n20653), .B(n20654), .X(\shifter_0/n10361 ) );
  nand_x1_sg U46972 ( .A(n20651), .B(n20652), .X(\shifter_0/n10362 ) );
  nand_x1_sg U46973 ( .A(n20649), .B(n20650), .X(\shifter_0/n10363 ) );
  nand_x1_sg U46974 ( .A(n20647), .B(n20648), .X(\shifter_0/n10364 ) );
  nand_x1_sg U46975 ( .A(n20645), .B(n20646), .X(\shifter_0/n10365 ) );
  nand_x1_sg U46976 ( .A(n20643), .B(n20644), .X(\shifter_0/n10366 ) );
  nand_x1_sg U46977 ( .A(n20641), .B(n20642), .X(\shifter_0/n10367 ) );
  nand_x1_sg U46978 ( .A(n20639), .B(n20640), .X(\shifter_0/n10368 ) );
  nand_x1_sg U46979 ( .A(n20637), .B(n20638), .X(\shifter_0/n10369 ) );
  nand_x1_sg U46980 ( .A(n20635), .B(n20636), .X(\shifter_0/n10370 ) );
  nand_x1_sg U46981 ( .A(n20633), .B(n20634), .X(\shifter_0/n10371 ) );
  nand_x1_sg U46982 ( .A(n20631), .B(n20632), .X(\shifter_0/n10372 ) );
  nand_x1_sg U46983 ( .A(n20629), .B(n20630), .X(\shifter_0/n10373 ) );
  nand_x1_sg U46984 ( .A(n20627), .B(n20628), .X(\shifter_0/n10374 ) );
  nand_x1_sg U46985 ( .A(n20625), .B(n20626), .X(\shifter_0/n10375 ) );
  nand_x1_sg U46986 ( .A(n20623), .B(n20624), .X(\shifter_0/n10376 ) );
  nand_x1_sg U46987 ( .A(n20621), .B(n20622), .X(\shifter_0/n10377 ) );
  nand_x1_sg U46988 ( .A(n20619), .B(n20620), .X(\shifter_0/n10378 ) );
  nand_x1_sg U46989 ( .A(n20617), .B(n20618), .X(\shifter_0/n10379 ) );
  nand_x1_sg U46990 ( .A(n20615), .B(n20616), .X(\shifter_0/n10380 ) );
  nand_x1_sg U46991 ( .A(n20613), .B(n20614), .X(\shifter_0/n10381 ) );
  nand_x1_sg U46992 ( .A(n20529), .B(n20530), .X(\shifter_0/n10423 ) );
  nand_x1_sg U46993 ( .A(n20527), .B(n20528), .X(\shifter_0/n10424 ) );
  nand_x1_sg U46994 ( .A(n20519), .B(n20520), .X(\shifter_0/n10428 ) );
  nand_x1_sg U46995 ( .A(n20517), .B(n20518), .X(\shifter_0/n10429 ) );
  nand_x1_sg U46996 ( .A(n20511), .B(n20512), .X(\shifter_0/n10432 ) );
  nand_x1_sg U46997 ( .A(n20509), .B(n20510), .X(\shifter_0/n10433 ) );
  nand_x1_sg U46998 ( .A(n20501), .B(n20502), .X(\shifter_0/n10437 ) );
  nand_x1_sg U46999 ( .A(n20499), .B(n20500), .X(\shifter_0/n10438 ) );
  nand_x1_sg U47000 ( .A(n20491), .B(n20492), .X(\shifter_0/n10442 ) );
  nand_x1_sg U47001 ( .A(n20489), .B(n20490), .X(\shifter_0/n10443 ) );
  nand_x1_sg U47002 ( .A(n20487), .B(n20488), .X(\shifter_0/n10444 ) );
  nand_x1_sg U47003 ( .A(n20485), .B(n20486), .X(\shifter_0/n10445 ) );
  nand_x1_sg U47004 ( .A(n20483), .B(n20484), .X(\shifter_0/n10446 ) );
  nand_x1_sg U47005 ( .A(n20481), .B(n20482), .X(\shifter_0/n10447 ) );
  nand_x1_sg U47006 ( .A(n20479), .B(n20480), .X(\shifter_0/n10448 ) );
  nand_x1_sg U47007 ( .A(n20477), .B(n20478), .X(\shifter_0/n10449 ) );
  nand_x1_sg U47008 ( .A(n20475), .B(n20476), .X(\shifter_0/n10450 ) );
  nand_x1_sg U47009 ( .A(n20473), .B(n20474), .X(\shifter_0/n10451 ) );
  nand_x1_sg U47010 ( .A(n20471), .B(n20472), .X(\shifter_0/n10452 ) );
  nand_x1_sg U47011 ( .A(n20469), .B(n20470), .X(\shifter_0/n10453 ) );
  nand_x1_sg U47012 ( .A(n20467), .B(n20468), .X(\shifter_0/n10454 ) );
  nand_x1_sg U47013 ( .A(n20465), .B(n20466), .X(\shifter_0/n10455 ) );
  nand_x1_sg U47014 ( .A(n20463), .B(n20464), .X(\shifter_0/n10456 ) );
  nand_x1_sg U47015 ( .A(n20461), .B(n20462), .X(\shifter_0/n10457 ) );
  nand_x1_sg U47016 ( .A(n20459), .B(n20460), .X(\shifter_0/n10458 ) );
  nand_x1_sg U47017 ( .A(n20457), .B(n20458), .X(\shifter_0/n10459 ) );
  nand_x1_sg U47018 ( .A(n20455), .B(n20456), .X(\shifter_0/n10460 ) );
  nand_x1_sg U47019 ( .A(n20453), .B(n20454), .X(\shifter_0/n10461 ) );
  nand_x1_sg U47020 ( .A(n20451), .B(n20452), .X(\shifter_0/n10462 ) );
  nand_x1_sg U47021 ( .A(n20449), .B(n20450), .X(\shifter_0/n10463 ) );
  nand_x1_sg U47022 ( .A(n20447), .B(n20448), .X(\shifter_0/n10464 ) );
  nand_x1_sg U47023 ( .A(n20445), .B(n20446), .X(\shifter_0/n10465 ) );
  nand_x1_sg U47024 ( .A(n20443), .B(n20444), .X(\shifter_0/n10466 ) );
  nand_x1_sg U47025 ( .A(n20441), .B(n20442), .X(\shifter_0/n10467 ) );
  nand_x1_sg U47026 ( .A(n20439), .B(n20440), .X(\shifter_0/n10468 ) );
  nand_x1_sg U47027 ( .A(n20419), .B(n20420), .X(\shifter_0/n10478 ) );
  nand_x1_sg U47028 ( .A(n20417), .B(n20418), .X(\shifter_0/n10479 ) );
  nand_x1_sg U47029 ( .A(n20415), .B(n20416), .X(\shifter_0/n10480 ) );
  nand_x1_sg U47030 ( .A(n20413), .B(n20414), .X(\shifter_0/n10481 ) );
  nand_x1_sg U47031 ( .A(n20411), .B(n20412), .X(\shifter_0/n10482 ) );
  nand_x1_sg U47032 ( .A(n20409), .B(n20410), .X(\shifter_0/n10483 ) );
  nand_x1_sg U47033 ( .A(n20407), .B(n20408), .X(\shifter_0/n10484 ) );
  nand_x1_sg U47034 ( .A(n20405), .B(n20406), .X(\shifter_0/n10485 ) );
  nand_x1_sg U47035 ( .A(n20403), .B(n20404), .X(\shifter_0/n10486 ) );
  nand_x1_sg U47036 ( .A(n20401), .B(n20402), .X(\shifter_0/n10487 ) );
  nand_x1_sg U47037 ( .A(n20399), .B(n20400), .X(\shifter_0/n10488 ) );
  nand_x1_sg U47038 ( .A(n20397), .B(n20398), .X(\shifter_0/n10489 ) );
  nand_x1_sg U47039 ( .A(n20395), .B(n20396), .X(\shifter_0/n10490 ) );
  nand_x1_sg U47040 ( .A(n20393), .B(n20394), .X(\shifter_0/n10491 ) );
  nand_x1_sg U47041 ( .A(n20391), .B(n20392), .X(\shifter_0/n10492 ) );
  nand_x1_sg U47042 ( .A(n20389), .B(n20390), .X(\shifter_0/n10493 ) );
  nand_x1_sg U47043 ( .A(n20387), .B(n20388), .X(\shifter_0/n10494 ) );
  nand_x1_sg U47044 ( .A(n20385), .B(n20386), .X(\shifter_0/n10495 ) );
  nand_x1_sg U47045 ( .A(n20383), .B(n20384), .X(\shifter_0/n10496 ) );
  nand_x1_sg U47046 ( .A(n20381), .B(n20382), .X(\shifter_0/n10497 ) );
  nand_x1_sg U47047 ( .A(n20379), .B(n20380), .X(\shifter_0/n10498 ) );
  nand_x1_sg U47048 ( .A(n20377), .B(n20378), .X(\shifter_0/n10499 ) );
  nand_x1_sg U47049 ( .A(n20375), .B(n20376), .X(\shifter_0/n10500 ) );
  nand_x1_sg U47050 ( .A(n20373), .B(n20374), .X(\shifter_0/n10501 ) );
  nand_x1_sg U47051 ( .A(n20369), .B(n20370), .X(\shifter_0/n10503 ) );
  nand_x1_sg U47052 ( .A(n20367), .B(n20368), .X(\shifter_0/n10504 ) );
  nand_x1_sg U47053 ( .A(n20359), .B(n20360), .X(\shifter_0/n10508 ) );
  nand_x1_sg U47054 ( .A(n20357), .B(n20358), .X(\shifter_0/n10509 ) );
  nand_x1_sg U47055 ( .A(n20351), .B(n20352), .X(\shifter_0/n10512 ) );
  nand_x1_sg U47056 ( .A(n20349), .B(n20350), .X(\shifter_0/n10513 ) );
  nand_x1_sg U47057 ( .A(n20341), .B(n20342), .X(\shifter_0/n10517 ) );
  nand_x1_sg U47058 ( .A(n20339), .B(n20340), .X(\shifter_0/n10518 ) );
  nand_x1_sg U47059 ( .A(n20331), .B(n20332), .X(\shifter_0/n10522 ) );
  nand_x1_sg U47060 ( .A(n20329), .B(n20330), .X(\shifter_0/n10523 ) );
  nand_x1_sg U47061 ( .A(n20327), .B(n20328), .X(\shifter_0/n10524 ) );
  nand_x1_sg U47062 ( .A(n20325), .B(n20326), .X(\shifter_0/n10525 ) );
  nand_x1_sg U47063 ( .A(n20323), .B(n20324), .X(\shifter_0/n10526 ) );
  nand_x1_sg U47064 ( .A(n20321), .B(n20322), .X(\shifter_0/n10527 ) );
  nand_x1_sg U47065 ( .A(n20309), .B(n20310), .X(\shifter_0/n10533 ) );
  nand_x1_sg U47066 ( .A(n20307), .B(n20308), .X(\shifter_0/n10534 ) );
  nand_x1_sg U47067 ( .A(n20305), .B(n20306), .X(\shifter_0/n10535 ) );
  nand_x1_sg U47068 ( .A(n20303), .B(n20304), .X(\shifter_0/n10536 ) );
  nand_x1_sg U47069 ( .A(n20301), .B(n20302), .X(\shifter_0/n10537 ) );
  nand_x1_sg U47070 ( .A(n20299), .B(n20300), .X(\shifter_0/n10538 ) );
  nand_x1_sg U47071 ( .A(n20297), .B(n20298), .X(\shifter_0/n10539 ) );
  nand_x1_sg U47072 ( .A(n20295), .B(n20296), .X(\shifter_0/n10540 ) );
  nand_x1_sg U47073 ( .A(n20293), .B(n20294), .X(\shifter_0/n10541 ) );
  nand_x1_sg U47074 ( .A(n20283), .B(n20284), .X(\shifter_0/n10546 ) );
  nand_x1_sg U47075 ( .A(n20281), .B(n20282), .X(\shifter_0/n10547 ) );
  nand_x1_sg U47076 ( .A(n20279), .B(n20280), .X(\shifter_0/n10548 ) );
  nand_x1_sg U47077 ( .A(n20277), .B(n20278), .X(\shifter_0/n10549 ) );
  nand_x1_sg U47078 ( .A(n20275), .B(n20276), .X(\shifter_0/n10550 ) );
  nand_x1_sg U47079 ( .A(n20273), .B(n20274), .X(\shifter_0/n10551 ) );
  nand_x1_sg U47080 ( .A(n20271), .B(n20272), .X(\shifter_0/n10552 ) );
  nand_x1_sg U47081 ( .A(n20269), .B(n20270), .X(\shifter_0/n10553 ) );
  nand_x1_sg U47082 ( .A(n20267), .B(n20268), .X(\shifter_0/n10554 ) );
  nand_x1_sg U47083 ( .A(n20265), .B(n20266), .X(\shifter_0/n10555 ) );
  nand_x1_sg U47084 ( .A(n20263), .B(n20264), .X(\shifter_0/n10556 ) );
  nand_x1_sg U47085 ( .A(n20261), .B(n20262), .X(\shifter_0/n10557 ) );
  nand_x1_sg U47086 ( .A(n20259), .B(n20260), .X(\shifter_0/n10558 ) );
  nand_x1_sg U47087 ( .A(n20257), .B(n20258), .X(\shifter_0/n10559 ) );
  nand_x1_sg U47088 ( .A(n20255), .B(n20256), .X(\shifter_0/n10560 ) );
  nand_x1_sg U47089 ( .A(n20253), .B(n20254), .X(\shifter_0/n10561 ) );
  nand_x1_sg U47090 ( .A(n20251), .B(n20252), .X(\shifter_0/n10562 ) );
  nand_x1_sg U47091 ( .A(n20249), .B(n20250), .X(\shifter_0/n10563 ) );
  nand_x1_sg U47092 ( .A(n20245), .B(n20246), .X(\shifter_0/n10565 ) );
  nand_x1_sg U47093 ( .A(n20243), .B(n20244), .X(\shifter_0/n10566 ) );
  nand_x1_sg U47094 ( .A(n20241), .B(n20242), .X(\shifter_0/n10567 ) );
  nand_x1_sg U47095 ( .A(n20239), .B(n20240), .X(\shifter_0/n10568 ) );
  nand_x1_sg U47096 ( .A(n20237), .B(n20238), .X(\shifter_0/n10569 ) );
  nand_x1_sg U47097 ( .A(n20235), .B(n20236), .X(\shifter_0/n10570 ) );
  nand_x1_sg U47098 ( .A(n20233), .B(n20234), .X(\shifter_0/n10571 ) );
  nand_x1_sg U47099 ( .A(n20231), .B(n20232), .X(\shifter_0/n10572 ) );
  nand_x1_sg U47100 ( .A(n20229), .B(n20230), .X(\shifter_0/n10573 ) );
  nand_x1_sg U47101 ( .A(n20227), .B(n20228), .X(\shifter_0/n10574 ) );
  nand_x1_sg U47102 ( .A(n20225), .B(n20226), .X(\shifter_0/n10575 ) );
  nand_x1_sg U47103 ( .A(n20223), .B(n20224), .X(\shifter_0/n10576 ) );
  nand_x1_sg U47104 ( .A(n20221), .B(n20222), .X(\shifter_0/n10577 ) );
  nand_x1_sg U47105 ( .A(n20219), .B(n20220), .X(\shifter_0/n10578 ) );
  nand_x1_sg U47106 ( .A(n20215), .B(n20216), .X(\shifter_0/n10580 ) );
  nand_x1_sg U47107 ( .A(n20213), .B(n20214), .X(\shifter_0/n10581 ) );
  nand_x1_sg U47108 ( .A(n20211), .B(n20212), .X(\shifter_0/n10582 ) );
  nand_x1_sg U47109 ( .A(n20209), .B(n20210), .X(\shifter_0/n10583 ) );
  nand_x1_sg U47110 ( .A(n20207), .B(n20208), .X(\shifter_0/n10584 ) );
  nand_x1_sg U47111 ( .A(n20205), .B(n20206), .X(\shifter_0/n10585 ) );
  nand_x1_sg U47112 ( .A(n20203), .B(n20204), .X(\shifter_0/n10586 ) );
  nand_x1_sg U47113 ( .A(n20191), .B(n20192), .X(\shifter_0/n10592 ) );
  nand_x1_sg U47114 ( .A(n20189), .B(n20190), .X(\shifter_0/n10593 ) );
  nand_x1_sg U47115 ( .A(n20187), .B(n20188), .X(\shifter_0/n10594 ) );
  nand_x1_sg U47116 ( .A(n20185), .B(n20186), .X(\shifter_0/n10595 ) );
  nand_x1_sg U47117 ( .A(n20165), .B(n20166), .X(\shifter_0/n10605 ) );
  nand_x1_sg U47118 ( .A(n20163), .B(n20164), .X(\shifter_0/n10606 ) );
  nand_x1_sg U47119 ( .A(n20161), .B(n20162), .X(\shifter_0/n10607 ) );
  nand_x1_sg U47120 ( .A(n20159), .B(n20160), .X(\shifter_0/n10608 ) );
  nand_x1_sg U47121 ( .A(n20157), .B(n20158), .X(\shifter_0/n10609 ) );
  nand_x1_sg U47122 ( .A(n20155), .B(n20156), .X(\shifter_0/n10610 ) );
  nand_x1_sg U47123 ( .A(n20153), .B(n20154), .X(\shifter_0/n10611 ) );
  nand_x1_sg U47124 ( .A(n20151), .B(n20152), .X(\shifter_0/n10612 ) );
  nand_x1_sg U47125 ( .A(n20149), .B(n20150), .X(\shifter_0/n10613 ) );
  nand_x1_sg U47126 ( .A(n20147), .B(n20148), .X(\shifter_0/n10614 ) );
  nand_x1_sg U47127 ( .A(n20145), .B(n20146), .X(\shifter_0/n10615 ) );
  nand_x1_sg U47128 ( .A(n20143), .B(n20144), .X(\shifter_0/n10616 ) );
  nand_x1_sg U47129 ( .A(n20141), .B(n20142), .X(\shifter_0/n10617 ) );
  nand_x1_sg U47130 ( .A(n20139), .B(n20140), .X(\shifter_0/n10618 ) );
  nand_x1_sg U47131 ( .A(n20137), .B(n20138), .X(\shifter_0/n10619 ) );
  nand_x1_sg U47132 ( .A(n20135), .B(n20136), .X(\shifter_0/n10620 ) );
  nand_x1_sg U47133 ( .A(n20133), .B(n20134), .X(\shifter_0/n10621 ) );
  nand_x1_sg U47134 ( .A(n20131), .B(n20132), .X(\shifter_0/n10622 ) );
  nand_x1_sg U47135 ( .A(n20129), .B(n20130), .X(\shifter_0/n10623 ) );
  nand_x1_sg U47136 ( .A(n20127), .B(n20128), .X(\shifter_0/n10624 ) );
  nand_x1_sg U47137 ( .A(n20125), .B(n20126), .X(\shifter_0/n10625 ) );
  nand_x1_sg U47138 ( .A(n20123), .B(n20124), .X(\shifter_0/n10626 ) );
  nand_x1_sg U47139 ( .A(n20121), .B(n20122), .X(\shifter_0/n10627 ) );
  nand_x1_sg U47140 ( .A(n20119), .B(n20120), .X(\shifter_0/n10628 ) );
  nand_x1_sg U47141 ( .A(n20117), .B(n20118), .X(\shifter_0/n10629 ) );
  nand_x1_sg U47142 ( .A(n20115), .B(n20116), .X(\shifter_0/n10630 ) );
  nand_x1_sg U47143 ( .A(n20113), .B(n20114), .X(\shifter_0/n10631 ) );
  nand_x1_sg U47144 ( .A(n20111), .B(n20112), .X(\shifter_0/n10632 ) );
  nand_x1_sg U47145 ( .A(n20101), .B(n20102), .X(\shifter_0/n10637 ) );
  nand_x1_sg U47146 ( .A(n20099), .B(n20100), .X(\shifter_0/n10638 ) );
  nand_x1_sg U47147 ( .A(n20097), .B(n20098), .X(\shifter_0/n10639 ) );
  nand_x1_sg U47148 ( .A(n20095), .B(n20096), .X(\shifter_0/n10640 ) );
  nand_x1_sg U47149 ( .A(n20093), .B(n20094), .X(\shifter_0/n10641 ) );
  nand_x1_sg U47150 ( .A(n20091), .B(n20092), .X(\shifter_0/n10642 ) );
  nand_x1_sg U47151 ( .A(n20089), .B(n20090), .X(\shifter_0/n10643 ) );
  nand_x1_sg U47152 ( .A(n20087), .B(n20088), .X(\shifter_0/n10644 ) );
  nand_x1_sg U47153 ( .A(n20085), .B(n20086), .X(\shifter_0/n10645 ) );
  nand_x1_sg U47154 ( .A(n20083), .B(n20084), .X(\shifter_0/n10646 ) );
  nand_x1_sg U47155 ( .A(n20081), .B(n20082), .X(\shifter_0/n10647 ) );
  nand_x1_sg U47156 ( .A(n20079), .B(n20080), .X(\shifter_0/n10648 ) );
  nand_x1_sg U47157 ( .A(n20077), .B(n20078), .X(\shifter_0/n10649 ) );
  nand_x1_sg U47158 ( .A(n20075), .B(n20076), .X(\shifter_0/n10650 ) );
  nand_x1_sg U47159 ( .A(n20073), .B(n20074), .X(\shifter_0/n10651 ) );
  nand_x1_sg U47160 ( .A(n20071), .B(n20072), .X(\shifter_0/n10652 ) );
  nand_x1_sg U47161 ( .A(n20069), .B(n20070), .X(\shifter_0/n10653 ) );
  nand_x1_sg U47162 ( .A(n20067), .B(n20068), .X(\shifter_0/n10654 ) );
  nand_x1_sg U47163 ( .A(n20047), .B(n20048), .X(\shifter_0/n10664 ) );
  nand_x1_sg U47164 ( .A(n20045), .B(n20046), .X(\shifter_0/n10665 ) );
  nand_x1_sg U47165 ( .A(n20043), .B(n20044), .X(\shifter_0/n10666 ) );
  nand_x1_sg U47166 ( .A(n20041), .B(n20042), .X(\shifter_0/n10667 ) );
  nand_x1_sg U47167 ( .A(n20039), .B(n20040), .X(\shifter_0/n10668 ) );
  nand_x1_sg U47168 ( .A(n20037), .B(n20038), .X(\shifter_0/n10669 ) );
  nand_x1_sg U47169 ( .A(n20035), .B(n20036), .X(\shifter_0/n10670 ) );
  nand_x1_sg U47170 ( .A(n20033), .B(n20034), .X(\shifter_0/n10671 ) );
  nand_x1_sg U47171 ( .A(n20031), .B(n20032), .X(\shifter_0/n10672 ) );
  nand_x1_sg U47172 ( .A(n20029), .B(n20030), .X(\shifter_0/n10673 ) );
  nand_x1_sg U47173 ( .A(n20027), .B(n20028), .X(\shifter_0/n10674 ) );
  nand_x1_sg U47174 ( .A(n20025), .B(n20026), .X(\shifter_0/n10675 ) );
  nand_x1_sg U47175 ( .A(n20023), .B(n20024), .X(\shifter_0/n10676 ) );
  nand_x1_sg U47176 ( .A(n20021), .B(n20022), .X(\shifter_0/n10677 ) );
  nand_x1_sg U47177 ( .A(n20019), .B(n20020), .X(\shifter_0/n10678 ) );
  nand_x1_sg U47178 ( .A(n20017), .B(n20018), .X(\shifter_0/n10679 ) );
  nand_x1_sg U47179 ( .A(n20015), .B(n20016), .X(\shifter_0/n10680 ) );
  nand_x1_sg U47180 ( .A(n20013), .B(n20014), .X(\shifter_0/n10681 ) );
  nand_x1_sg U47181 ( .A(n20011), .B(n20012), .X(\shifter_0/n10682 ) );
  nand_x1_sg U47182 ( .A(n20009), .B(n20010), .X(\shifter_0/n10683 ) );
  nand_x1_sg U47183 ( .A(n20007), .B(n20008), .X(\shifter_0/n10684 ) );
  nand_x1_sg U47184 ( .A(n20005), .B(n20006), .X(\shifter_0/n10685 ) );
  nand_x1_sg U47185 ( .A(n20003), .B(n20004), .X(\shifter_0/n10686 ) );
  nand_x1_sg U47186 ( .A(n20001), .B(n20002), .X(\shifter_0/n10687 ) );
  nand_x1_sg U47187 ( .A(n19999), .B(n20000), .X(\shifter_0/n10688 ) );
  nand_x1_sg U47188 ( .A(n19997), .B(n19998), .X(\shifter_0/n10689 ) );
  nand_x1_sg U47189 ( .A(n19995), .B(n19996), .X(\shifter_0/n10690 ) );
  nand_x1_sg U47190 ( .A(n19993), .B(n19994), .X(\shifter_0/n10691 ) );
  nand_x1_sg U47191 ( .A(n19991), .B(n19992), .X(\shifter_0/n10692 ) );
  nand_x1_sg U47192 ( .A(n19989), .B(n19990), .X(\shifter_0/n10693 ) );
  nand_x1_sg U47193 ( .A(n19987), .B(n19988), .X(\shifter_0/n10694 ) );
  nand_x1_sg U47194 ( .A(n19985), .B(n19986), .X(\shifter_0/n10695 ) );
  nand_x1_sg U47195 ( .A(n19983), .B(n19984), .X(\shifter_0/n10696 ) );
  nand_x1_sg U47196 ( .A(n19981), .B(n19982), .X(\shifter_0/n10697 ) );
  nand_x1_sg U47197 ( .A(n19979), .B(n19980), .X(\shifter_0/n10698 ) );
  nand_x1_sg U47198 ( .A(n19977), .B(n19978), .X(\shifter_0/n10699 ) );
  nand_x1_sg U47199 ( .A(n19975), .B(n19976), .X(\shifter_0/n10700 ) );
  nand_x1_sg U47200 ( .A(n19973), .B(n19974), .X(\shifter_0/n10701 ) );
  nand_x1_sg U47201 ( .A(n19901), .B(n19902), .X(\shifter_0/n10737 ) );
  nand_x1_sg U47202 ( .A(n19889), .B(n19890), .X(\shifter_0/n10743 ) );
  nand_x1_sg U47203 ( .A(n19887), .B(n19888), .X(\shifter_0/n10744 ) );
  nand_x1_sg U47204 ( .A(n19879), .B(n19880), .X(\shifter_0/n10748 ) );
  nand_x1_sg U47205 ( .A(n19877), .B(n19878), .X(\shifter_0/n10749 ) );
  nand_x1_sg U47206 ( .A(n19871), .B(n19872), .X(\shifter_0/n10752 ) );
  nand_x1_sg U47207 ( .A(n19869), .B(n19870), .X(\shifter_0/n10753 ) );
  nand_x1_sg U47208 ( .A(n19861), .B(n19862), .X(\shifter_0/n10757 ) );
  nand_x1_sg U47209 ( .A(n19859), .B(n19860), .X(\shifter_0/n10758 ) );
  nand_x1_sg U47210 ( .A(n19851), .B(n19852), .X(\shifter_0/n10762 ) );
  nand_x1_sg U47211 ( .A(n19849), .B(n19850), .X(\shifter_0/n10763 ) );
  nand_x1_sg U47212 ( .A(n19847), .B(n19848), .X(\shifter_0/n10764 ) );
  nand_x1_sg U47213 ( .A(n19845), .B(n19846), .X(\shifter_0/n10765 ) );
  nand_x1_sg U47214 ( .A(n19843), .B(n19844), .X(\shifter_0/n10766 ) );
  nand_x1_sg U47215 ( .A(n19841), .B(n19842), .X(\shifter_0/n10767 ) );
  nand_x1_sg U47216 ( .A(n19839), .B(n19840), .X(\shifter_0/n10768 ) );
  nand_x1_sg U47217 ( .A(n19837), .B(n19838), .X(\shifter_0/n10769 ) );
  nand_x1_sg U47218 ( .A(n19835), .B(n19836), .X(\shifter_0/n10770 ) );
  nand_x1_sg U47219 ( .A(n19833), .B(n19834), .X(\shifter_0/n10771 ) );
  nand_x1_sg U47220 ( .A(n19831), .B(n19832), .X(\shifter_0/n10772 ) );
  nand_x1_sg U47221 ( .A(n19811), .B(n19812), .X(\shifter_0/n10782 ) );
  nand_x1_sg U47222 ( .A(n19809), .B(n19810), .X(\shifter_0/n10783 ) );
  nand_x1_sg U47223 ( .A(n19807), .B(n19808), .X(\shifter_0/n10784 ) );
  nand_x1_sg U47224 ( .A(n19805), .B(n19806), .X(\shifter_0/n10785 ) );
  nand_x1_sg U47225 ( .A(n19803), .B(n19804), .X(\shifter_0/n10786 ) );
  nand_x1_sg U47226 ( .A(n19801), .B(n19802), .X(\shifter_0/n10787 ) );
  nand_x1_sg U47227 ( .A(n19799), .B(n19800), .X(\shifter_0/n10788 ) );
  nand_x1_sg U47228 ( .A(n19797), .B(n19798), .X(\shifter_0/n10789 ) );
  nand_x1_sg U47229 ( .A(n19795), .B(n19796), .X(\shifter_0/n10790 ) );
  nand_x1_sg U47230 ( .A(n19793), .B(n19794), .X(\shifter_0/n10791 ) );
  nand_x1_sg U47231 ( .A(n19791), .B(n19792), .X(\shifter_0/n10792 ) );
  nand_x1_sg U47232 ( .A(n19789), .B(n19790), .X(\shifter_0/n10793 ) );
  nand_x1_sg U47233 ( .A(n19787), .B(n19788), .X(\shifter_0/n10794 ) );
  nand_x1_sg U47234 ( .A(n19785), .B(n19786), .X(\shifter_0/n10795 ) );
  nand_x1_sg U47235 ( .A(n19783), .B(n19784), .X(\shifter_0/n10796 ) );
  nand_x1_sg U47236 ( .A(n19781), .B(n19782), .X(\shifter_0/n10797 ) );
  nand_x1_sg U47237 ( .A(n19779), .B(n19780), .X(\shifter_0/n10798 ) );
  nand_x1_sg U47238 ( .A(n19777), .B(n19778), .X(\shifter_0/n10799 ) );
  nand_x1_sg U47239 ( .A(n19775), .B(n19776), .X(\shifter_0/n10800 ) );
  nand_x1_sg U47240 ( .A(n19773), .B(n19774), .X(\shifter_0/n10801 ) );
  nand_x1_sg U47241 ( .A(n19771), .B(n19772), .X(\shifter_0/n10802 ) );
  nand_x1_sg U47242 ( .A(n19769), .B(n19770), .X(\shifter_0/n10803 ) );
  nand_x1_sg U47243 ( .A(n19767), .B(n19768), .X(\shifter_0/n10804 ) );
  nand_x1_sg U47244 ( .A(n19765), .B(n19766), .X(\shifter_0/n10805 ) );
  nand_x1_sg U47245 ( .A(n19763), .B(n19764), .X(\shifter_0/n10806 ) );
  nand_x1_sg U47246 ( .A(n19761), .B(n19762), .X(\shifter_0/n10807 ) );
  nand_x1_sg U47247 ( .A(n19759), .B(n19760), .X(\shifter_0/n10808 ) );
  nand_x1_sg U47248 ( .A(n19757), .B(n19758), .X(\shifter_0/n10809 ) );
  nand_x1_sg U47249 ( .A(n19755), .B(n19756), .X(\shifter_0/n10810 ) );
  nand_x1_sg U47250 ( .A(n19753), .B(n19754), .X(\shifter_0/n10811 ) );
  nand_x1_sg U47251 ( .A(n19751), .B(n19752), .X(\shifter_0/n10812 ) );
  nand_x1_sg U47252 ( .A(n19749), .B(n19750), .X(\shifter_0/n10813 ) );
  nand_x1_sg U47253 ( .A(n19747), .B(n19748), .X(\shifter_0/n10814 ) );
  nand_x1_sg U47254 ( .A(n19745), .B(n19746), .X(\shifter_0/n10815 ) );
  nand_x1_sg U47255 ( .A(n19743), .B(n19744), .X(\shifter_0/n10816 ) );
  nand_x1_sg U47256 ( .A(n19741), .B(n19742), .X(\shifter_0/n10817 ) );
  nand_x1_sg U47257 ( .A(n19739), .B(n19740), .X(\shifter_0/n10818 ) );
  nand_x1_sg U47258 ( .A(n19737), .B(n19738), .X(\shifter_0/n10819 ) );
  nand_x1_sg U47259 ( .A(n19735), .B(n19736), .X(\shifter_0/n10820 ) );
  nand_x1_sg U47260 ( .A(n19733), .B(n19734), .X(\shifter_0/n10821 ) );
  nand_x1_sg U47261 ( .A(n19729), .B(n19730), .X(\shifter_0/n10823 ) );
  nand_x1_sg U47262 ( .A(n19727), .B(n19728), .X(\shifter_0/n10824 ) );
  nand_x1_sg U47263 ( .A(n19719), .B(n19720), .X(\shifter_0/n10828 ) );
  nand_x1_sg U47264 ( .A(n19717), .B(n19718), .X(\shifter_0/n10829 ) );
  nand_x1_sg U47265 ( .A(n19709), .B(n19710), .X(\shifter_0/n10833 ) );
  nand_x1_sg U47266 ( .A(n19701), .B(n19702), .X(\shifter_0/n10837 ) );
  nand_x1_sg U47267 ( .A(n19699), .B(n19700), .X(\shifter_0/n10838 ) );
  nand_x1_sg U47268 ( .A(n19675), .B(n19676), .X(\shifter_0/n10850 ) );
  nand_x1_sg U47269 ( .A(n19673), .B(n19674), .X(\shifter_0/n10851 ) );
  nand_x1_sg U47270 ( .A(n19671), .B(n19672), .X(\shifter_0/n10852 ) );
  nand_x1_sg U47271 ( .A(n19669), .B(n19670), .X(\shifter_0/n10853 ) );
  nand_x1_sg U47272 ( .A(n19667), .B(n19668), .X(\shifter_0/n10854 ) );
  nand_x1_sg U47273 ( .A(n19665), .B(n19666), .X(\shifter_0/n10855 ) );
  nand_x1_sg U47274 ( .A(n19663), .B(n19664), .X(\shifter_0/n10856 ) );
  nand_x1_sg U47275 ( .A(n19661), .B(n19662), .X(\shifter_0/n10857 ) );
  nand_x1_sg U47276 ( .A(n19659), .B(n19660), .X(\shifter_0/n10858 ) );
  nand_x1_sg U47277 ( .A(n19657), .B(n19658), .X(\shifter_0/n10859 ) );
  nand_x1_sg U47278 ( .A(n19655), .B(n19656), .X(\shifter_0/n10860 ) );
  nand_x1_sg U47279 ( .A(n19653), .B(n19654), .X(\shifter_0/n10861 ) );
  nand_x1_sg U47280 ( .A(n19651), .B(n19652), .X(\shifter_0/n10862 ) );
  nand_x1_sg U47281 ( .A(n19649), .B(n19650), .X(\shifter_0/n10863 ) );
  nand_x1_sg U47282 ( .A(n19647), .B(n19648), .X(\shifter_0/n10864 ) );
  nand_x1_sg U47283 ( .A(n19645), .B(n19646), .X(\shifter_0/n10865 ) );
  nand_x1_sg U47284 ( .A(n19643), .B(n19644), .X(\shifter_0/n10866 ) );
  nand_x1_sg U47285 ( .A(n19641), .B(n19642), .X(\shifter_0/n10867 ) );
  nand_x1_sg U47286 ( .A(n19639), .B(n19640), .X(\shifter_0/n10868 ) );
  nand_x1_sg U47287 ( .A(n19637), .B(n19638), .X(\shifter_0/n10869 ) );
  nand_x1_sg U47288 ( .A(n19635), .B(n19636), .X(\shifter_0/n10870 ) );
  nand_x1_sg U47289 ( .A(n19633), .B(n19634), .X(\shifter_0/n10871 ) );
  nand_x1_sg U47290 ( .A(n19631), .B(n19632), .X(\shifter_0/n10872 ) );
  nand_x1_sg U47291 ( .A(n19629), .B(n19630), .X(\shifter_0/n10873 ) );
  nand_x1_sg U47292 ( .A(n19627), .B(n19628), .X(\shifter_0/n10874 ) );
  nand_x1_sg U47293 ( .A(n19625), .B(n19626), .X(\shifter_0/n10875 ) );
  nand_x1_sg U47294 ( .A(n19623), .B(n19624), .X(\shifter_0/n10876 ) );
  nand_x1_sg U47295 ( .A(n19621), .B(n19622), .X(\shifter_0/n10877 ) );
  nand_x1_sg U47296 ( .A(n19619), .B(n19620), .X(\shifter_0/n10878 ) );
  nand_x1_sg U47297 ( .A(n19617), .B(n19618), .X(\shifter_0/n10879 ) );
  nand_x1_sg U47298 ( .A(n19615), .B(n19616), .X(\shifter_0/n10880 ) );
  nand_x1_sg U47299 ( .A(n19613), .B(n19614), .X(\shifter_0/n10881 ) );
  nand_x1_sg U47300 ( .A(n20525), .B(n20526), .X(\shifter_0/n10425 ) );
  nand_x1_sg U47301 ( .A(n20611), .B(n20612), .X(\shifter_0/n10382 ) );
  nand_x1_sg U47302 ( .A(n20609), .B(n20610), .X(\shifter_0/n10383 ) );
  nand_x1_sg U47303 ( .A(n20607), .B(n20608), .X(\shifter_0/n10384 ) );
  nand_x1_sg U47304 ( .A(n20605), .B(n20606), .X(\shifter_0/n10385 ) );
  nand_x1_sg U47305 ( .A(n20603), .B(n20604), .X(\shifter_0/n10386 ) );
  nand_x1_sg U47306 ( .A(n20601), .B(n20602), .X(\shifter_0/n10387 ) );
  nand_x1_sg U47307 ( .A(n20599), .B(n20600), .X(\shifter_0/n10388 ) );
  nand_x1_sg U47308 ( .A(n20597), .B(n20598), .X(\shifter_0/n10389 ) );
  nand_x1_sg U47309 ( .A(n20595), .B(n20596), .X(\shifter_0/n10390 ) );
  nand_x1_sg U47310 ( .A(n20593), .B(n20594), .X(\shifter_0/n10391 ) );
  nand_x1_sg U47311 ( .A(n20591), .B(n20592), .X(\shifter_0/n10392 ) );
  nand_x1_sg U47312 ( .A(n20589), .B(n20590), .X(\shifter_0/n10393 ) );
  nand_x1_sg U47313 ( .A(n20587), .B(n20588), .X(\shifter_0/n10394 ) );
  nand_x1_sg U47314 ( .A(n20585), .B(n20586), .X(\shifter_0/n10395 ) );
  nand_x1_sg U47315 ( .A(n20583), .B(n20584), .X(\shifter_0/n10396 ) );
  nand_x1_sg U47316 ( .A(n20581), .B(n20582), .X(\shifter_0/n10397 ) );
  nand_x1_sg U47317 ( .A(n20579), .B(n20580), .X(\shifter_0/n10398 ) );
  nand_x1_sg U47318 ( .A(n20577), .B(n20578), .X(\shifter_0/n10399 ) );
  nand_x1_sg U47319 ( .A(n20575), .B(n20576), .X(\shifter_0/n10400 ) );
  nand_x1_sg U47320 ( .A(n20573), .B(n20574), .X(\shifter_0/n10401 ) );
  nand_x1_sg U47321 ( .A(n20531), .B(n20532), .X(\shifter_0/n10422 ) );
  nand_x1_sg U47322 ( .A(n20507), .B(n20508), .X(\shifter_0/n10434 ) );
  nand_x1_sg U47323 ( .A(n20505), .B(n20506), .X(\shifter_0/n10435 ) );
  nand_x1_sg U47324 ( .A(n20503), .B(n20504), .X(\shifter_0/n10436 ) );
  nand_x1_sg U47325 ( .A(n20497), .B(n20498), .X(\shifter_0/n10439 ) );
  nand_x1_sg U47326 ( .A(n20495), .B(n20496), .X(\shifter_0/n10440 ) );
  nand_x1_sg U47327 ( .A(n20493), .B(n20494), .X(\shifter_0/n10441 ) );
  nand_x1_sg U47328 ( .A(n20247), .B(n20248), .X(\shifter_0/n10564 ) );
  nand_x1_sg U47329 ( .A(n20217), .B(n20218), .X(\shifter_0/n10579 ) );
  nand_x1_sg U47330 ( .A(n19971), .B(n19972), .X(\shifter_0/n10702 ) );
  nand_x1_sg U47331 ( .A(n19969), .B(n19970), .X(\shifter_0/n10703 ) );
  nand_x1_sg U47332 ( .A(n19967), .B(n19968), .X(\shifter_0/n10704 ) );
  nand_x1_sg U47333 ( .A(n19965), .B(n19966), .X(\shifter_0/n10705 ) );
  nand_x1_sg U47334 ( .A(n19963), .B(n19964), .X(\shifter_0/n10706 ) );
  nand_x1_sg U47335 ( .A(n19961), .B(n19962), .X(\shifter_0/n10707 ) );
  nand_x1_sg U47336 ( .A(n19959), .B(n19960), .X(\shifter_0/n10708 ) );
  nand_x1_sg U47337 ( .A(n19957), .B(n19958), .X(\shifter_0/n10709 ) );
  nand_x1_sg U47338 ( .A(n19955), .B(n19956), .X(\shifter_0/n10710 ) );
  nand_x1_sg U47339 ( .A(n19953), .B(n19954), .X(\shifter_0/n10711 ) );
  nand_x1_sg U47340 ( .A(n19951), .B(n19952), .X(\shifter_0/n10712 ) );
  nand_x1_sg U47341 ( .A(n19949), .B(n19950), .X(\shifter_0/n10713 ) );
  nand_x1_sg U47342 ( .A(n19929), .B(n19930), .X(\shifter_0/n10723 ) );
  nand_x1_sg U47343 ( .A(n19927), .B(n19928), .X(\shifter_0/n10724 ) );
  nand_x1_sg U47344 ( .A(n19897), .B(n19898), .X(\shifter_0/n10739 ) );
  nand_x1_sg U47345 ( .A(n19891), .B(n19892), .X(\shifter_0/n10742 ) );
  nand_x1_sg U47346 ( .A(n19885), .B(n19886), .X(\shifter_0/n10745 ) );
  nand_x1_sg U47347 ( .A(n19883), .B(n19884), .X(\shifter_0/n10746 ) );
  nand_x1_sg U47348 ( .A(n19881), .B(n19882), .X(\shifter_0/n10747 ) );
  nand_x1_sg U47349 ( .A(n19875), .B(n19876), .X(\shifter_0/n10750 ) );
  nand_x1_sg U47350 ( .A(n19873), .B(n19874), .X(\shifter_0/n10751 ) );
  nand_x1_sg U47351 ( .A(n19731), .B(n19732), .X(\shifter_0/n10822 ) );
  nand_x1_sg U47352 ( .A(n19725), .B(n19726), .X(\shifter_0/n10825 ) );
  nand_x1_sg U47353 ( .A(n19723), .B(n19724), .X(\shifter_0/n10826 ) );
  nand_x1_sg U47354 ( .A(n19721), .B(n19722), .X(\shifter_0/n10827 ) );
  nand_x1_sg U47355 ( .A(n19715), .B(n19716), .X(\shifter_0/n10830 ) );
  nand_x1_sg U47356 ( .A(n19713), .B(n19714), .X(\shifter_0/n10831 ) );
  nand_x1_sg U47357 ( .A(n19707), .B(n19708), .X(\shifter_0/n10834 ) );
  nand_x1_sg U47358 ( .A(n19705), .B(n19706), .X(\shifter_0/n10835 ) );
  nand_x1_sg U47359 ( .A(n19703), .B(n19704), .X(\shifter_0/n10836 ) );
  nand_x1_sg U47360 ( .A(n19697), .B(n19698), .X(\shifter_0/n10839 ) );
  nand_x1_sg U47361 ( .A(n19695), .B(n19696), .X(\shifter_0/n10840 ) );
  nand_x1_sg U47362 ( .A(n19693), .B(n19694), .X(\shifter_0/n10841 ) );
  nand_x1_sg U47363 ( .A(n20523), .B(n20524), .X(\shifter_0/n10426 ) );
  nand_x1_sg U47364 ( .A(n20521), .B(n20522), .X(\shifter_0/n10427 ) );
  nand_x1_sg U47365 ( .A(n20515), .B(n20516), .X(\shifter_0/n10430 ) );
  nand_x1_sg U47366 ( .A(n20513), .B(n20514), .X(\shifter_0/n10431 ) );
  nand_x1_sg U47367 ( .A(n20371), .B(n20372), .X(\shifter_0/n10502 ) );
  nand_x1_sg U47368 ( .A(n20365), .B(n20366), .X(\shifter_0/n10505 ) );
  nand_x1_sg U47369 ( .A(n20363), .B(n20364), .X(\shifter_0/n10506 ) );
  nand_x1_sg U47370 ( .A(n20361), .B(n20362), .X(\shifter_0/n10507 ) );
  nand_x1_sg U47371 ( .A(n20355), .B(n20356), .X(\shifter_0/n10510 ) );
  nand_x1_sg U47372 ( .A(n20353), .B(n20354), .X(\shifter_0/n10511 ) );
  nand_x1_sg U47373 ( .A(n20347), .B(n20348), .X(\shifter_0/n10514 ) );
  nand_x1_sg U47374 ( .A(n20345), .B(n20346), .X(\shifter_0/n10515 ) );
  nand_x1_sg U47375 ( .A(n20343), .B(n20344), .X(\shifter_0/n10516 ) );
  nand_x1_sg U47376 ( .A(n20337), .B(n20338), .X(\shifter_0/n10519 ) );
  nand_x1_sg U47377 ( .A(n20335), .B(n20336), .X(\shifter_0/n10520 ) );
  nand_x1_sg U47378 ( .A(n20333), .B(n20334), .X(\shifter_0/n10521 ) );
  nand_x1_sg U47379 ( .A(n19867), .B(n19868), .X(\shifter_0/n10754 ) );
  nand_x1_sg U47380 ( .A(n19865), .B(n19866), .X(\shifter_0/n10755 ) );
  nand_x1_sg U47381 ( .A(n19863), .B(n19864), .X(\shifter_0/n10756 ) );
  nand_x1_sg U47382 ( .A(n19857), .B(n19858), .X(\shifter_0/n10759 ) );
  nand_x1_sg U47383 ( .A(n19855), .B(n19856), .X(\shifter_0/n10760 ) );
  nand_x1_sg U47384 ( .A(n19853), .B(n19854), .X(\shifter_0/n10761 ) );
  nand_x1_sg U47385 ( .A(n20555), .B(n20556), .X(\shifter_0/n10410 ) );
  nand_x1_sg U47386 ( .A(n20553), .B(n20554), .X(\shifter_0/n10411 ) );
  nand_x1_sg U47387 ( .A(n20551), .B(n20552), .X(\shifter_0/n10412 ) );
  nand_x1_sg U47388 ( .A(n20549), .B(n20550), .X(\shifter_0/n10413 ) );
  nand_x1_sg U47389 ( .A(n20547), .B(n20548), .X(\shifter_0/n10414 ) );
  nand_x1_sg U47390 ( .A(n20545), .B(n20546), .X(\shifter_0/n10415 ) );
  nand_x1_sg U47391 ( .A(n20543), .B(n20544), .X(\shifter_0/n10416 ) );
  nand_x1_sg U47392 ( .A(n20541), .B(n20542), .X(\shifter_0/n10417 ) );
  nand_x1_sg U47393 ( .A(n20539), .B(n20540), .X(\shifter_0/n10418 ) );
  nand_x1_sg U47394 ( .A(n19931), .B(n19932), .X(\shifter_0/n10722 ) );
  nand_x1_sg U47395 ( .A(n20793), .B(n20794), .X(\shifter_0/n10291 ) );
  nand_x1_sg U47396 ( .A(n20787), .B(n20788), .X(\shifter_0/n10294 ) );
  nand_x1_sg U47397 ( .A(n20785), .B(n20786), .X(\shifter_0/n10295 ) );
  nand_x1_sg U47398 ( .A(n20783), .B(n20784), .X(\shifter_0/n10296 ) );
  nand_x1_sg U47399 ( .A(n20777), .B(n20778), .X(\shifter_0/n10299 ) );
  nand_x1_sg U47400 ( .A(n20775), .B(n20776), .X(\shifter_0/n10300 ) );
  nand_x1_sg U47401 ( .A(n20707), .B(n20708), .X(\shifter_0/n10334 ) );
  nand_x1_sg U47402 ( .A(n20705), .B(n20706), .X(\shifter_0/n10335 ) );
  nand_x1_sg U47403 ( .A(n20703), .B(n20704), .X(\shifter_0/n10336 ) );
  nand_x1_sg U47404 ( .A(n20697), .B(n20698), .X(\shifter_0/n10339 ) );
  nand_x1_sg U47405 ( .A(n20695), .B(n20696), .X(\shifter_0/n10340 ) );
  nand_x1_sg U47406 ( .A(n20673), .B(n20674), .X(\shifter_0/n10351 ) );
  nand_x1_sg U47407 ( .A(n20671), .B(n20672), .X(\shifter_0/n10352 ) );
  nand_x1_sg U47408 ( .A(n20669), .B(n20670), .X(\shifter_0/n10353 ) );
  nand_x1_sg U47409 ( .A(n20667), .B(n20668), .X(\shifter_0/n10354 ) );
  nand_x1_sg U47410 ( .A(n20665), .B(n20666), .X(\shifter_0/n10355 ) );
  nand_x1_sg U47411 ( .A(n20663), .B(n20664), .X(\shifter_0/n10356 ) );
  nand_x1_sg U47412 ( .A(n20661), .B(n20662), .X(\shifter_0/n10357 ) );
  nand_x1_sg U47413 ( .A(n20659), .B(n20660), .X(\shifter_0/n10358 ) );
  nand_x1_sg U47414 ( .A(n20657), .B(n20658), .X(\shifter_0/n10359 ) );
  nand_x1_sg U47415 ( .A(n20201), .B(n20202), .X(\shifter_0/n10587 ) );
  nand_x1_sg U47416 ( .A(n20195), .B(n20196), .X(\shifter_0/n10590 ) );
  nand_x1_sg U47417 ( .A(n20193), .B(n20194), .X(\shifter_0/n10591 ) );
  nand_x1_sg U47418 ( .A(n20183), .B(n20184), .X(\shifter_0/n10596 ) );
  nand_x1_sg U47419 ( .A(n20179), .B(n20180), .X(\shifter_0/n10598 ) );
  nand_x1_sg U47420 ( .A(n20175), .B(n20176), .X(\shifter_0/n10600 ) );
  nand_x1_sg U47421 ( .A(n20173), .B(n20174), .X(\shifter_0/n10601 ) );
  nand_x1_sg U47422 ( .A(n20171), .B(n20172), .X(\shifter_0/n10602 ) );
  nand_x1_sg U47423 ( .A(n20107), .B(n20108), .X(\shifter_0/n10634 ) );
  nand_x1_sg U47424 ( .A(n20105), .B(n20106), .X(\shifter_0/n10635 ) );
  nand_x1_sg U47425 ( .A(n20103), .B(n20104), .X(\shifter_0/n10636 ) );
  nand_x1_sg U47426 ( .A(n20065), .B(n20066), .X(\shifter_0/n10655 ) );
  nand_x1_sg U47427 ( .A(n20063), .B(n20064), .X(\shifter_0/n10656 ) );
  nand_x1_sg U47428 ( .A(n20059), .B(n20060), .X(\shifter_0/n10658 ) );
  nand_x1_sg U47429 ( .A(n20055), .B(n20056), .X(\shifter_0/n10660 ) );
  nand_x1_sg U47430 ( .A(n20053), .B(n20054), .X(\shifter_0/n10661 ) );
  nand_x1_sg U47431 ( .A(n20051), .B(n20052), .X(\shifter_0/n10662 ) );
  nand_x1_sg U47432 ( .A(n19827), .B(n19828), .X(\shifter_0/n10774 ) );
  nand_x1_sg U47433 ( .A(n19825), .B(n19826), .X(\shifter_0/n10775 ) );
  nand_x1_sg U47434 ( .A(n19823), .B(n19824), .X(\shifter_0/n10776 ) );
  nand_x1_sg U47435 ( .A(n19817), .B(n19818), .X(\shifter_0/n10779 ) );
  nand_x1_sg U47436 ( .A(n19815), .B(n19816), .X(\shifter_0/n10780 ) );
  nand_x1_sg U47437 ( .A(n19813), .B(n19814), .X(\shifter_0/n10781 ) );
  nand_x1_sg U47438 ( .A(n19939), .B(n19940), .X(\shifter_0/n10718 ) );
  nand_x1_sg U47439 ( .A(n19937), .B(n19938), .X(\shifter_0/n10719 ) );
  nand_x1_sg U47440 ( .A(n19947), .B(n19948), .X(\shifter_0/n10714 ) );
  nand_x1_sg U47441 ( .A(n19945), .B(n19946), .X(\shifter_0/n10715 ) );
  nand_x1_sg U47442 ( .A(n19943), .B(n19944), .X(\shifter_0/n10716 ) );
  nand_x1_sg U47443 ( .A(n19941), .B(n19942), .X(\shifter_0/n10717 ) );
  nand_x1_sg U47444 ( .A(n19935), .B(n19936), .X(\shifter_0/n10720 ) );
  nand_x1_sg U47445 ( .A(n19933), .B(n19934), .X(\shifter_0/n10721 ) );
  nand_x1_sg U47446 ( .A(n20061), .B(n20062), .X(\shifter_0/n10657 ) );
  nand_x1_sg U47447 ( .A(n20791), .B(n20792), .X(\shifter_0/n10292 ) );
  nand_x1_sg U47448 ( .A(n20789), .B(n20790), .X(\shifter_0/n10293 ) );
  nand_x1_sg U47449 ( .A(n20781), .B(n20782), .X(\shifter_0/n10297 ) );
  nand_x1_sg U47450 ( .A(n20779), .B(n20780), .X(\shifter_0/n10298 ) );
  nand_x1_sg U47451 ( .A(n20709), .B(n20710), .X(\shifter_0/n10333 ) );
  nand_x1_sg U47452 ( .A(n20701), .B(n20702), .X(\shifter_0/n10337 ) );
  nand_x1_sg U47453 ( .A(n20319), .B(n20320), .X(\shifter_0/n10528 ) );
  nand_x1_sg U47454 ( .A(n20317), .B(n20318), .X(\shifter_0/n10529 ) );
  nand_x1_sg U47455 ( .A(n20315), .B(n20316), .X(\shifter_0/n10530 ) );
  nand_x1_sg U47456 ( .A(n20313), .B(n20314), .X(\shifter_0/n10531 ) );
  nand_x1_sg U47457 ( .A(n20311), .B(n20312), .X(\shifter_0/n10532 ) );
  nand_x1_sg U47458 ( .A(n20291), .B(n20292), .X(\shifter_0/n10542 ) );
  nand_x1_sg U47459 ( .A(n20289), .B(n20290), .X(\shifter_0/n10543 ) );
  nand_x1_sg U47460 ( .A(n20287), .B(n20288), .X(\shifter_0/n10544 ) );
  nand_x1_sg U47461 ( .A(n20285), .B(n20286), .X(\shifter_0/n10545 ) );
  nand_x1_sg U47462 ( .A(n20199), .B(n20200), .X(\shifter_0/n10588 ) );
  nand_x1_sg U47463 ( .A(n20197), .B(n20198), .X(\shifter_0/n10589 ) );
  nand_x1_sg U47464 ( .A(n20181), .B(n20182), .X(\shifter_0/n10597 ) );
  nand_x1_sg U47465 ( .A(n20177), .B(n20178), .X(\shifter_0/n10599 ) );
  nand_x1_sg U47466 ( .A(n20169), .B(n20170), .X(\shifter_0/n10603 ) );
  nand_x1_sg U47467 ( .A(n20167), .B(n20168), .X(\shifter_0/n10604 ) );
  nand_x1_sg U47468 ( .A(n20057), .B(n20058), .X(\shifter_0/n10659 ) );
  nand_x1_sg U47469 ( .A(n20049), .B(n20050), .X(\shifter_0/n10663 ) );
  nand_x1_sg U47470 ( .A(n19711), .B(n19712), .X(\shifter_0/n10832 ) );
  nand_x1_sg U47471 ( .A(n19691), .B(n19692), .X(\shifter_0/n10842 ) );
  nand_x1_sg U47472 ( .A(n19689), .B(n19690), .X(\shifter_0/n10843 ) );
  nand_x1_sg U47473 ( .A(n19687), .B(n19688), .X(\shifter_0/n10844 ) );
  nand_x1_sg U47474 ( .A(n19685), .B(n19686), .X(\shifter_0/n10845 ) );
  nand_x1_sg U47475 ( .A(n19683), .B(n19684), .X(\shifter_0/n10846 ) );
  nand_x1_sg U47476 ( .A(n19681), .B(n19682), .X(\shifter_0/n10847 ) );
  nand_x1_sg U47477 ( .A(n19679), .B(n19680), .X(\shifter_0/n10848 ) );
  nand_x1_sg U47478 ( .A(n19677), .B(n19678), .X(\shifter_0/n10849 ) );
  nand_x1_sg U47479 ( .A(n20699), .B(n20700), .X(\shifter_0/n10338 ) );
  nand_x1_sg U47480 ( .A(n20437), .B(n20438), .X(\shifter_0/n10469 ) );
  nand_x1_sg U47481 ( .A(n20435), .B(n20436), .X(\shifter_0/n10470 ) );
  nand_x1_sg U47482 ( .A(n20433), .B(n20434), .X(\shifter_0/n10471 ) );
  nand_x1_sg U47483 ( .A(n20431), .B(n20432), .X(\shifter_0/n10472 ) );
  nand_x1_sg U47484 ( .A(n20429), .B(n20430), .X(\shifter_0/n10473 ) );
  nand_x1_sg U47485 ( .A(n20427), .B(n20428), .X(\shifter_0/n10474 ) );
  nand_x1_sg U47486 ( .A(n20425), .B(n20426), .X(\shifter_0/n10475 ) );
  nand_x1_sg U47487 ( .A(n20423), .B(n20424), .X(\shifter_0/n10476 ) );
  nand_x1_sg U47488 ( .A(n20421), .B(n20422), .X(\shifter_0/n10477 ) );
  nand_x1_sg U47489 ( .A(n20109), .B(n20110), .X(\shifter_0/n10633 ) );
  nand_x1_sg U47490 ( .A(n19829), .B(n19830), .X(\shifter_0/n10773 ) );
  nand_x1_sg U47491 ( .A(n19821), .B(n19822), .X(\shifter_0/n10777 ) );
  nand_x1_sg U47492 ( .A(n19819), .B(n19820), .X(\shifter_0/n10778 ) );
  nand_x1_sg U47493 ( .A(n31112), .B(n19610), .X(\shifter_0/n10882 ) );
  nand_x1_sg U47494 ( .A(n26348), .B(n26349), .X(\mask_0/n706 ) );
  nand_x1_sg U47495 ( .A(n26353), .B(n26354), .X(\mask_0/n705 ) );
  nand_x1_sg U47496 ( .A(n26356), .B(n26357), .X(\mask_0/n704 ) );
  nand_x1_sg U47497 ( .A(n26359), .B(n26360), .X(\mask_0/n703 ) );
  nand_x1_sg U47498 ( .A(n26362), .B(n26363), .X(\mask_0/n702 ) );
  nand_x1_sg U47499 ( .A(n26365), .B(n26366), .X(\mask_0/n701 ) );
  nand_x1_sg U47500 ( .A(n26368), .B(n26369), .X(\mask_0/n700 ) );
  nand_x1_sg U47501 ( .A(n26371), .B(n26372), .X(\mask_0/n699 ) );
  nand_x1_sg U47502 ( .A(n26374), .B(n26375), .X(\mask_0/n698 ) );
  nand_x1_sg U47503 ( .A(n26377), .B(n26378), .X(\mask_0/n697 ) );
  nand_x1_sg U47504 ( .A(n26380), .B(n26381), .X(\mask_0/n696 ) );
  nand_x1_sg U47505 ( .A(n26383), .B(n26384), .X(\mask_0/n695 ) );
  nand_x1_sg U47506 ( .A(n26386), .B(n26387), .X(\mask_0/n694 ) );
  nand_x1_sg U47507 ( .A(n26389), .B(n26390), .X(\mask_0/n693 ) );
  nand_x1_sg U47508 ( .A(n26392), .B(n26393), .X(\mask_0/n692 ) );
  nand_x1_sg U47509 ( .A(n26395), .B(n26396), .X(\mask_0/n691 ) );
  nand_x1_sg U47510 ( .A(n26398), .B(n26399), .X(\mask_0/n690 ) );
  nand_x1_sg U47511 ( .A(n26401), .B(n26402), .X(\mask_0/n689 ) );
  nand_x1_sg U47512 ( .A(n26404), .B(n26405), .X(\mask_0/n688 ) );
  nand_x1_sg U47513 ( .A(n26407), .B(n26408), .X(\mask_0/n687 ) );
  nand_x1_sg U47514 ( .A(n26410), .B(n26411), .X(\mask_0/n686 ) );
  nand_x1_sg U47515 ( .A(n26413), .B(n26414), .X(\mask_0/n685 ) );
  nand_x1_sg U47516 ( .A(n26416), .B(n26417), .X(\mask_0/n684 ) );
  nand_x1_sg U47517 ( .A(n26419), .B(n26420), .X(\mask_0/n683 ) );
  nand_x1_sg U47518 ( .A(n26422), .B(n26423), .X(\mask_0/n682 ) );
  nand_x1_sg U47519 ( .A(n26425), .B(n26426), .X(\mask_0/n681 ) );
  nand_x1_sg U47520 ( .A(n26428), .B(n26429), .X(\mask_0/n680 ) );
  nand_x1_sg U47521 ( .A(n26431), .B(n26432), .X(\mask_0/n679 ) );
  nand_x1_sg U47522 ( .A(n26434), .B(n26435), .X(\mask_0/n678 ) );
  nand_x1_sg U47523 ( .A(n26437), .B(n26438), .X(\mask_0/n677 ) );
  nand_x1_sg U47524 ( .A(n26440), .B(n26441), .X(\mask_0/n676 ) );
  nand_x1_sg U47525 ( .A(n26443), .B(n26444), .X(\mask_0/n675 ) );
  nand_x1_sg U47526 ( .A(n26470), .B(n26471), .X(\mask_0/n662 ) );
  nand_x1_sg U47527 ( .A(n26472), .B(n26473), .X(\mask_0/n661 ) );
  nand_x1_sg U47528 ( .A(n26482), .B(n26483), .X(\mask_0/n656 ) );
  nand_x1_sg U47529 ( .A(n26446), .B(n26447), .X(\mask_0/n674 ) );
  nand_x1_sg U47530 ( .A(n26448), .B(n26449), .X(\mask_0/n673 ) );
  nand_x1_sg U47531 ( .A(n26450), .B(n26451), .X(\mask_0/n672 ) );
  nand_x1_sg U47532 ( .A(n26452), .B(n26453), .X(\mask_0/n671 ) );
  nand_x1_sg U47533 ( .A(n26454), .B(n26455), .X(\mask_0/n670 ) );
  nand_x1_sg U47534 ( .A(n26456), .B(n26457), .X(\mask_0/n669 ) );
  nand_x1_sg U47535 ( .A(n26458), .B(n26459), .X(\mask_0/n668 ) );
  nand_x1_sg U47536 ( .A(n26460), .B(n26461), .X(\mask_0/n667 ) );
  nand_x1_sg U47537 ( .A(n26462), .B(n26463), .X(\mask_0/n666 ) );
  nand_x1_sg U47538 ( .A(n26464), .B(n26465), .X(\mask_0/n665 ) );
  nand_x1_sg U47539 ( .A(n26466), .B(n26467), .X(\mask_0/n664 ) );
  nand_x1_sg U47540 ( .A(n26468), .B(n26469), .X(\mask_0/n663 ) );
  nand_x1_sg U47541 ( .A(n26474), .B(n26475), .X(\mask_0/n660 ) );
  nand_x1_sg U47542 ( .A(n26476), .B(n26477), .X(\mask_0/n659 ) );
  nand_x1_sg U47543 ( .A(n26478), .B(n26479), .X(\mask_0/n658 ) );
  nand_x1_sg U47544 ( .A(n26480), .B(n26481), .X(\mask_0/n657 ) );
  nand_x1_sg U47545 ( .A(n26484), .B(n26485), .X(\mask_0/n655 ) );
  nand_x1_sg U47546 ( .A(n26486), .B(n26487), .X(\mask_0/n654 ) );
  nand_x1_sg U47547 ( .A(n26488), .B(n26489), .X(\mask_0/n653 ) );
  nand_x1_sg U47548 ( .A(n26490), .B(n26491), .X(\mask_0/n652 ) );
  nand_x1_sg U47549 ( .A(n26492), .B(n26493), .X(\mask_0/n651 ) );
  nand_x1_sg U47550 ( .A(n26494), .B(n26495), .X(\mask_0/n650 ) );
  nand_x1_sg U47551 ( .A(n26496), .B(n26497), .X(\mask_0/n649 ) );
  nand_x1_sg U47552 ( .A(n26498), .B(n26499), .X(\mask_0/n648 ) );
  nand_x1_sg U47553 ( .A(n26500), .B(n26501), .X(\mask_0/n647 ) );
  nand_x1_sg U47554 ( .A(n26502), .B(n26503), .X(\mask_0/n646 ) );
  nand_x1_sg U47555 ( .A(n26504), .B(n26505), .X(\mask_0/n645 ) );
  nand_x1_sg U47556 ( .A(n26506), .B(n26507), .X(\mask_0/n644 ) );
  nand_x1_sg U47557 ( .A(n26508), .B(n26509), .X(\mask_0/n643 ) );
  nand_x1_sg U47558 ( .A(n26510), .B(n26511), .X(\mask_0/n642 ) );
  nand_x1_sg U47559 ( .A(n26512), .B(n26513), .X(\mask_0/n641 ) );
  nand_x1_sg U47560 ( .A(n26514), .B(n26515), .X(\mask_0/n640 ) );
  nand_x1_sg U47561 ( .A(n26516), .B(n26517), .X(\mask_0/n639 ) );
  nand_x1_sg U47562 ( .A(n26518), .B(n26519), .X(\mask_0/n638 ) );
  nand_x1_sg U47563 ( .A(n26520), .B(n26521), .X(\mask_0/n637 ) );
  nand_x1_sg U47564 ( .A(n26522), .B(n26523), .X(\mask_0/n636 ) );
  nand_x1_sg U47565 ( .A(n26524), .B(n26525), .X(\mask_0/n635 ) );
  nand_x1_sg U47566 ( .A(n26526), .B(n26527), .X(\mask_0/n634 ) );
  nand_x1_sg U47567 ( .A(n26528), .B(n26529), .X(\mask_0/n633 ) );
  nand_x1_sg U47568 ( .A(n26530), .B(n26531), .X(\mask_0/n632 ) );
  nand_x1_sg U47569 ( .A(n26532), .B(n26533), .X(\mask_0/n631 ) );
  nand_x1_sg U47570 ( .A(n26534), .B(n26535), .X(\mask_0/n630 ) );
  nand_x1_sg U47571 ( .A(n26536), .B(n26537), .X(\mask_0/n629 ) );
  nand_x1_sg U47572 ( .A(n26538), .B(n26539), .X(\mask_0/n628 ) );
  nand_x1_sg U47573 ( .A(n26540), .B(n26541), .X(\mask_0/n627 ) );
  nand_x1_sg U47574 ( .A(n26542), .B(n26543), .X(\mask_0/n626 ) );
  nand_x1_sg U47575 ( .A(n26544), .B(n26545), .X(\mask_0/n625 ) );
  nand_x1_sg U47576 ( .A(n26546), .B(n26547), .X(\mask_0/n624 ) );
  nand_x1_sg U47577 ( .A(n26548), .B(n26549), .X(\mask_0/n623 ) );
  nand_x1_sg U47578 ( .A(n26550), .B(n26551), .X(\mask_0/n622 ) );
  nand_x1_sg U47579 ( .A(n26552), .B(n26553), .X(\mask_0/n621 ) );
  nand_x1_sg U47580 ( .A(n26554), .B(n26555), .X(\mask_0/n620 ) );
  nand_x1_sg U47581 ( .A(n26556), .B(n26557), .X(\mask_0/n619 ) );
  nand_x1_sg U47582 ( .A(n26558), .B(n26559), .X(\mask_0/n618 ) );
  nand_x1_sg U47583 ( .A(n26560), .B(n26561), .X(\mask_0/n617 ) );
  nand_x1_sg U47584 ( .A(n26562), .B(n26563), .X(\mask_0/n616 ) );
  nand_x1_sg U47585 ( .A(n26564), .B(n26565), .X(\mask_0/n615 ) );
  nand_x1_sg U47586 ( .A(n26566), .B(n26567), .X(\mask_0/n614 ) );
  nand_x1_sg U47587 ( .A(n26568), .B(n26569), .X(\mask_0/n613 ) );
  nand_x1_sg U47588 ( .A(n26570), .B(n26571), .X(\mask_0/n612 ) );
  nand_x1_sg U47589 ( .A(n26572), .B(n26573), .X(\mask_0/n611 ) );
  nand_x1_sg U47590 ( .A(n28968), .B(n28969), .X(\filter_0/n8567 ) );
  nand_x1_sg U47591 ( .A(n28974), .B(n28975), .X(\filter_0/n8564 ) );
  nand_x1_sg U47592 ( .A(n32886), .B(\filter_0/n8240 ), .X(n28974) );
  nand_x1_sg U47593 ( .A(n28274), .B(n28275), .X(\filter_0/n8888 ) );
  nand_x1_sg U47594 ( .A(n32887), .B(\filter_0/n7911 ), .X(n28274) );
  nand_x1_sg U47595 ( .A(n28970), .B(n28971), .X(\filter_0/n8566 ) );
  nand_x1_sg U47596 ( .A(n28972), .B(n28973), .X(\filter_0/n8565 ) );
  nand_x1_sg U47597 ( .A(n32887), .B(\filter_0/n8241 ), .X(n28972) );
  nand_x1_sg U47598 ( .A(n28257), .B(n28258), .X(\filter_0/n8896 ) );
  nand_x1_sg U47599 ( .A(n28262), .B(n28263), .X(\filter_0/n8894 ) );
  nand_x1_sg U47600 ( .A(n28268), .B(n28269), .X(\filter_0/n8891 ) );
  nand_x1_sg U47601 ( .A(n28272), .B(n28273), .X(\filter_0/n8889 ) );
  nand_x1_sg U47602 ( .A(n28260), .B(n28261), .X(\filter_0/n8895 ) );
  nand_x1_sg U47603 ( .A(n26291), .B(n26292), .X(\mask_0/n734 ) );
  nand_x1_sg U47604 ( .A(n26273), .B(n26274), .X(\mask_0/n743 ) );
  nand_x1_sg U47605 ( .A(n26271), .B(n26272), .X(\mask_0/n744 ) );
  nand_x1_sg U47606 ( .A(n26269), .B(n26270), .X(\mask_0/n745 ) );
  nand_x1_sg U47607 ( .A(n26267), .B(n26268), .X(\mask_0/n746 ) );
  nand_x1_sg U47608 ( .A(n26265), .B(n26266), .X(\mask_0/n747 ) );
  nand_x1_sg U47609 ( .A(n26263), .B(n26264), .X(\mask_0/n748 ) );
  nand_x1_sg U47610 ( .A(n26345), .B(n26346), .X(\mask_0/n707 ) );
  nand_x1_sg U47611 ( .A(n26343), .B(n26344), .X(\mask_0/n708 ) );
  nand_x1_sg U47612 ( .A(n26341), .B(n26342), .X(\mask_0/n709 ) );
  nand_x1_sg U47613 ( .A(n26339), .B(n26340), .X(\mask_0/n710 ) );
  nand_x1_sg U47614 ( .A(n26337), .B(n26338), .X(\mask_0/n711 ) );
  nand_x1_sg U47615 ( .A(n26335), .B(n26336), .X(\mask_0/n712 ) );
  nand_x1_sg U47616 ( .A(n26333), .B(n26334), .X(\mask_0/n713 ) );
  nand_x1_sg U47617 ( .A(n26331), .B(n26332), .X(\mask_0/n714 ) );
  nand_x1_sg U47618 ( .A(n26329), .B(n26330), .X(\mask_0/n715 ) );
  nand_x1_sg U47619 ( .A(n26327), .B(n26328), .X(\mask_0/n716 ) );
  nand_x1_sg U47620 ( .A(n26325), .B(n26326), .X(\mask_0/n717 ) );
  nand_x1_sg U47621 ( .A(n26323), .B(n26324), .X(\mask_0/n718 ) );
  nand_x1_sg U47622 ( .A(n26321), .B(n26322), .X(\mask_0/n719 ) );
  nand_x1_sg U47623 ( .A(n26319), .B(n26320), .X(\mask_0/n720 ) );
  nand_x1_sg U47624 ( .A(n26317), .B(n26318), .X(\mask_0/n721 ) );
  nand_x1_sg U47625 ( .A(n26315), .B(n26316), .X(\mask_0/n722 ) );
  nand_x1_sg U47626 ( .A(n26313), .B(n26314), .X(\mask_0/n723 ) );
  nand_x1_sg U47627 ( .A(n26311), .B(n26312), .X(\mask_0/n724 ) );
  nand_x1_sg U47628 ( .A(n26309), .B(n26310), .X(\mask_0/n725 ) );
  nand_x1_sg U47629 ( .A(n26307), .B(n26308), .X(\mask_0/n726 ) );
  nand_x1_sg U47630 ( .A(n26305), .B(n26306), .X(\mask_0/n727 ) );
  nand_x1_sg U47631 ( .A(n26303), .B(n26304), .X(\mask_0/n728 ) );
  nand_x1_sg U47632 ( .A(n26301), .B(n26302), .X(\mask_0/n729 ) );
  nand_x1_sg U47633 ( .A(n26299), .B(n26300), .X(\mask_0/n730 ) );
  nand_x1_sg U47634 ( .A(n26297), .B(n26298), .X(\mask_0/n731 ) );
  nand_x1_sg U47635 ( .A(n26295), .B(n26296), .X(\mask_0/n732 ) );
  nand_x1_sg U47636 ( .A(n26293), .B(n26294), .X(\mask_0/n733 ) );
  nand_x1_sg U47637 ( .A(n26289), .B(n26290), .X(\mask_0/n735 ) );
  nand_x1_sg U47638 ( .A(n26287), .B(n26288), .X(\mask_0/n736 ) );
  nand_x1_sg U47639 ( .A(n26285), .B(n26286), .X(\mask_0/n737 ) );
  nand_x1_sg U47640 ( .A(n26283), .B(n26284), .X(\mask_0/n738 ) );
  nand_x1_sg U47641 ( .A(n26281), .B(n26282), .X(\mask_0/n739 ) );
  nand_x1_sg U47642 ( .A(n26279), .B(n26280), .X(\mask_0/n740 ) );
  nand_x1_sg U47643 ( .A(n26277), .B(n26278), .X(\mask_0/n741 ) );
  nand_x1_sg U47644 ( .A(n26275), .B(n26276), .X(\mask_0/n742 ) );
  nand_x1_sg U47645 ( .A(n26261), .B(n26262), .X(\mask_0/n749 ) );
  nand_x1_sg U47646 ( .A(n26259), .B(n26260), .X(\mask_0/n750 ) );
  nand_x1_sg U47647 ( .A(n26257), .B(n26258), .X(\mask_0/n751 ) );
  nand_x1_sg U47648 ( .A(n26255), .B(n26256), .X(\mask_0/n752 ) );
  nand_x1_sg U47649 ( .A(n26253), .B(n26254), .X(\mask_0/n753 ) );
  nand_x1_sg U47650 ( .A(n26251), .B(n26252), .X(\mask_0/n754 ) );
  nand_x1_sg U47651 ( .A(n26249), .B(n26250), .X(\mask_0/n755 ) );
  nand_x1_sg U47652 ( .A(n26247), .B(n26248), .X(\mask_0/n756 ) );
  nand_x1_sg U47653 ( .A(n26245), .B(n26246), .X(\mask_0/n757 ) );
  nand_x1_sg U47654 ( .A(n26243), .B(n26244), .X(\mask_0/n758 ) );
  nand_x1_sg U47655 ( .A(n26241), .B(n26242), .X(\mask_0/n759 ) );
  nand_x1_sg U47656 ( .A(n26239), .B(n26240), .X(\mask_0/n760 ) );
  nand_x1_sg U47657 ( .A(n26237), .B(n26238), .X(\mask_0/n761 ) );
  nand_x1_sg U47658 ( .A(n26235), .B(n26236), .X(\mask_0/n762 ) );
  nand_x1_sg U47659 ( .A(n26233), .B(n26234), .X(\mask_0/n763 ) );
  nand_x1_sg U47660 ( .A(n26231), .B(n26232), .X(\mask_0/n764 ) );
  nand_x1_sg U47661 ( .A(n26229), .B(n26230), .X(\mask_0/n765 ) );
  nand_x1_sg U47662 ( .A(n26227), .B(n26228), .X(\mask_0/n766 ) );
  nand_x1_sg U47663 ( .A(n26225), .B(n26226), .X(\mask_0/n767 ) );
  nand_x1_sg U47664 ( .A(n26223), .B(n26224), .X(\mask_0/n768 ) );
  nand_x1_sg U47665 ( .A(n26221), .B(n26222), .X(\mask_0/n769 ) );
  nand_x1_sg U47666 ( .A(n26217), .B(n26218), .X(\mask_0/n770 ) );
  nand_x1_sg U47667 ( .A(n28270), .B(n28271), .X(\filter_0/n8890 ) );
  nand_x1_sg U47668 ( .A(n28266), .B(n28267), .X(\filter_0/n8892 ) );
  nand_x1_sg U47669 ( .A(n28264), .B(n28265), .X(\filter_0/n8893 ) );
  inv_x1_sg U47670 ( .A(n21146), .X(n42717) );
  inv_x1_sg U47671 ( .A(n21138), .X(n42715) );
  inv_x1_sg U47672 ( .A(n21135), .X(n42714) );
  inv_x1_sg U47673 ( .A(n21143), .X(n42716) );
  inv_x1_sg U47674 ( .A(n26585), .X(n42412) );
  inv_x1_sg U47675 ( .A(n21238), .X(n42719) );
  inv_x1_sg U47676 ( .A(n21235), .X(n42718) );
  inv_x1_sg U47677 ( .A(n21246), .X(n42721) );
  nand_x1_sg U47678 ( .A(n26580), .B(n26581), .X(\filter_0/n9634 ) );
  inv_x1_sg U47679 ( .A(n21534), .X(n42605) );
  inv_x1_sg U47680 ( .A(n21539), .X(n42606) );
  inv_x1_sg U47681 ( .A(n21243), .X(n42720) );
  nand_x1_sg U47682 ( .A(n26576), .B(n26577), .X(\filter_0/n9635 ) );
  inv_x1_sg U47683 ( .A(n21591), .X(n42608) );
  inv_x1_sg U47684 ( .A(n21256), .X(n42731) );
  inv_x1_sg U47685 ( .A(n21253), .X(n42730) );
  inv_x1_sg U47686 ( .A(n21264), .X(n42733) );
  inv_x1_sg U47687 ( .A(n21695), .X(n42629) );
  inv_x1_sg U47688 ( .A(n21596), .X(n42609) );
  inv_x1_sg U47689 ( .A(n21261), .X(n42732) );
  inv_x1_sg U47690 ( .A(n21588), .X(n42607) );
  inv_x1_sg U47691 ( .A(n21713), .X(n42643) );
  inv_x1_sg U47692 ( .A(n21674), .X(n42636) );
  inv_x1_sg U47693 ( .A(n21599), .X(n42610) );
  inv_x1_sg U47694 ( .A(n21609), .X(n42619) );
  inv_x1_sg U47695 ( .A(n21614), .X(n42620) );
  inv_x1_sg U47696 ( .A(n21606), .X(n42618) );
  inv_x1_sg U47697 ( .A(n21617), .X(n42621) );
  inv_x1_sg U47698 ( .A(n21644), .X(n42611) );
  inv_x1_sg U47699 ( .A(n21626), .X(n42622) );
  nand_x1_sg U47700 ( .A(n26210), .B(n26211), .X(\mask_0/n771 ) );
  nand_x1_sg U47701 ( .A(n26212), .B(n35418), .X(n26211) );
  nand_x1_sg U47702 ( .A(n26207), .B(n26208), .X(\mask_0/n772 ) );
  nand_x1_sg U47703 ( .A(n26201), .B(n26202), .X(\mask_0/n773 ) );
  inv_x1_sg U47704 ( .A(n28254), .X(n42478) );
  inv_x1_sg U47705 ( .A(n28249), .X(n42477) );
  inv_x1_sg U47706 ( .A(n28244), .X(n42476) );
  inv_x1_sg U47707 ( .A(n28239), .X(n42475) );
  inv_x1_sg U47708 ( .A(n28234), .X(n42474) );
  inv_x1_sg U47709 ( .A(n28229), .X(n42473) );
  inv_x1_sg U47710 ( .A(n28224), .X(n42472) );
  inv_x1_sg U47711 ( .A(n28219), .X(n42471) );
  inv_x1_sg U47712 ( .A(n28214), .X(n42470) );
  inv_x1_sg U47713 ( .A(n28209), .X(n42469) );
  inv_x1_sg U47714 ( .A(n28204), .X(n42468) );
  inv_x1_sg U47715 ( .A(n28199), .X(n42467) );
  inv_x1_sg U47716 ( .A(n28194), .X(n42466) );
  inv_x1_sg U47717 ( .A(n28189), .X(n42465) );
  inv_x1_sg U47718 ( .A(n28184), .X(n42464) );
  inv_x1_sg U47719 ( .A(n28179), .X(n42463) );
  inv_x1_sg U47720 ( .A(n28174), .X(n42462) );
  inv_x1_sg U47721 ( .A(n28169), .X(n42461) );
  inv_x1_sg U47722 ( .A(n28164), .X(n42460) );
  inv_x1_sg U47723 ( .A(n28159), .X(n42459) );
  inv_x1_sg U47724 ( .A(n28154), .X(n42458) );
  inv_x1_sg U47725 ( .A(n28149), .X(n42457) );
  inv_x1_sg U47726 ( .A(n28144), .X(n42456) );
  inv_x1_sg U47727 ( .A(n28139), .X(n42455) );
  inv_x1_sg U47728 ( .A(n28134), .X(n42454) );
  inv_x1_sg U47729 ( .A(n28129), .X(n42453) );
  inv_x1_sg U47730 ( .A(n28124), .X(n42452) );
  inv_x1_sg U47731 ( .A(n28119), .X(n42451) );
  inv_x1_sg U47732 ( .A(n28114), .X(n42450) );
  inv_x1_sg U47733 ( .A(n28109), .X(n42449) );
  inv_x1_sg U47734 ( .A(n28104), .X(n42448) );
  inv_x1_sg U47735 ( .A(n28099), .X(n42447) );
  inv_x1_sg U47736 ( .A(n28094), .X(n42446) );
  inv_x1_sg U47737 ( .A(n28089), .X(n42445) );
  inv_x1_sg U47738 ( .A(n28084), .X(n42444) );
  inv_x1_sg U47739 ( .A(n28079), .X(n42443) );
  inv_x1_sg U47740 ( .A(n28074), .X(n42442) );
  inv_x1_sg U47741 ( .A(n28069), .X(n42441) );
  inv_x1_sg U47742 ( .A(n28064), .X(n42440) );
  inv_x1_sg U47743 ( .A(n28059), .X(n42439) );
  inv_x1_sg U47744 ( .A(n28054), .X(n42438) );
  inv_x1_sg U47745 ( .A(n28049), .X(n42437) );
  inv_x1_sg U47746 ( .A(n28044), .X(n42436) );
  inv_x1_sg U47747 ( .A(n28039), .X(n42435) );
  inv_x1_sg U47748 ( .A(n28034), .X(n42434) );
  inv_x1_sg U47749 ( .A(n28029), .X(n42433) );
  inv_x1_sg U47750 ( .A(n28024), .X(n42432) );
  inv_x1_sg U47751 ( .A(n28019), .X(n42431) );
  inv_x1_sg U47752 ( .A(n28014), .X(n42430) );
  inv_x1_sg U47753 ( .A(n28009), .X(n42429) );
  inv_x1_sg U47754 ( .A(n28004), .X(n42428) );
  inv_x1_sg U47755 ( .A(n27999), .X(n42427) );
  inv_x1_sg U47756 ( .A(n27994), .X(n42426) );
  inv_x1_sg U47757 ( .A(n27989), .X(n42425) );
  inv_x1_sg U47758 ( .A(n27984), .X(n42424) );
  inv_x1_sg U47759 ( .A(n27979), .X(n42423) );
  inv_x1_sg U47760 ( .A(n27974), .X(n42422) );
  inv_x1_sg U47761 ( .A(n27969), .X(n42421) );
  inv_x1_sg U47762 ( .A(n27964), .X(n42420) );
  inv_x1_sg U47763 ( .A(n27959), .X(n42419) );
  inv_x1_sg U47764 ( .A(n27954), .X(n42418) );
  inv_x1_sg U47765 ( .A(n27949), .X(n42417) );
  inv_x1_sg U47766 ( .A(n27944), .X(n42416) );
  inv_x1_sg U47767 ( .A(n27939), .X(n42415) );
  inv_x1_sg U47768 ( .A(n14266), .X(n40924) );
  inv_x1_sg U47769 ( .A(n14390), .X(n40918) );
  inv_x1_sg U47770 ( .A(n14453), .X(n41069) );
  inv_x1_sg U47771 ( .A(n14579), .X(n41063) );
  inv_x1_sg U47772 ( .A(n14641), .X(n41059) );
  inv_x1_sg U47773 ( .A(n14765), .X(n41053) );
  inv_x1_sg U47774 ( .A(n14889), .X(n41047) );
  inv_x1_sg U47775 ( .A(n14952), .X(n41044) );
  inv_x1_sg U47776 ( .A(n14204), .X(n40928) );
  inv_x1_sg U47777 ( .A(n14328), .X(n40921) );
  inv_x1_sg U47778 ( .A(n14517), .X(n41066) );
  inv_x1_sg U47779 ( .A(n14703), .X(n41057) );
  inv_x1_sg U47780 ( .A(n14827), .X(n41051) );
  inv_x1_sg U47781 ( .A(n13987), .X(n40938) );
  inv_x1_sg U47782 ( .A(n14018), .X(n40936) );
  inv_x1_sg U47783 ( .A(n14111), .X(n40932) );
  inv_x1_sg U47784 ( .A(n14142), .X(n40930) );
  inv_x1_sg U47785 ( .A(n14235), .X(n40926) );
  inv_x1_sg U47786 ( .A(n14297), .X(n40922) );
  inv_x1_sg U47787 ( .A(n14422), .X(n41071) );
  inv_x1_sg U47788 ( .A(n14610), .X(n41061) );
  inv_x1_sg U47789 ( .A(n14734), .X(n41055) );
  inv_x1_sg U47790 ( .A(n14858), .X(n41049) );
  inv_x1_sg U47791 ( .A(n14920), .X(n41045) );
  inv_x1_sg U47792 ( .A(n15013), .X(n41041) );
  inv_x1_sg U47793 ( .A(n13795), .X(n40948) );
  inv_x1_sg U47794 ( .A(n13832), .X(n40946) );
  inv_x1_sg U47795 ( .A(n13863), .X(n40944) );
  inv_x1_sg U47796 ( .A(n13956), .X(n40940) );
  inv_x1_sg U47797 ( .A(n14485), .X(n41067) );
  inv_x1_sg U47798 ( .A(n14549), .X(n41065) );
  inv_x1_sg U47799 ( .A(n14983), .X(n41043) );
  inv_x1_sg U47800 ( .A(n14049), .X(n40935) );
  inv_x1_sg U47801 ( .A(n14080), .X(n40934) );
  inv_x1_sg U47802 ( .A(n14173), .X(n40929) );
  inv_x1_sg U47803 ( .A(n14359), .X(n40920) );
  inv_x1_sg U47804 ( .A(n14672), .X(n41058) );
  inv_x1_sg U47805 ( .A(n14796), .X(n41052) );
  inv_x1_sg U47806 ( .A(n13894), .X(n40943) );
  inv_x1_sg U47807 ( .A(n13925), .X(n40942) );
  inv_x1_sg U47808 ( .A(n15150), .X(n42373) );
  inv_x1_sg U47809 ( .A(n15279), .X(n42375) );
  inv_x1_sg U47810 ( .A(n15117), .X(n42372) );
  inv_x1_sg U47811 ( .A(n15246), .X(n42374) );
  inv_x1_sg U47812 ( .A(n15064), .X(n42404) );
  inv_x1_sg U47813 ( .A(n15200), .X(n42397) );
  nand_x1_sg U47814 ( .A(n31413), .B(n40911), .X(n14121) );
  nand_x1_sg U47815 ( .A(n30076), .B(n40910), .X(n14152) );
  nand_x1_sg U47816 ( .A(n34204), .B(n40909), .X(n14245) );
  nand_x1_sg U47817 ( .A(n34206), .B(n40908), .X(n14276) );
  inv_x1_sg U47818 ( .A(n15092), .X(n42367) );
  inv_x1_sg U47819 ( .A(n15226), .X(n42368) );
  nand_x1_sg U47820 ( .A(n12458), .B(n12459), .X(\shifter_0/n7657 ) );
  inv_x1_sg U47821 ( .A(n15222), .X(n42384) );
  inv_x1_sg U47822 ( .A(n15086), .X(n42383) );
  inv_x1_sg U47823 ( .A(n15136), .X(n42392) );
  inv_x1_sg U47824 ( .A(n15265), .X(n42389) );
  nand_x1_sg U47825 ( .A(n12446), .B(n12447), .X(\shifter_0/n7666 ) );
  nand_x1_sg U47826 ( .A(n12455), .B(n12456), .X(\shifter_0/n7658 ) );
  nand_x1_sg U47827 ( .A(n12508), .B(n12509), .X(\shifter_0/n7606 ) );
  nand_x1_sg U47828 ( .A(n12513), .B(n12514), .X(\shifter_0/n7602 ) );
  nand_x1_sg U47829 ( .A(n12347), .B(n12348), .X(\shifter_0/n7754 ) );
  nand_x1_sg U47830 ( .A(n12354), .B(n12355), .X(\shifter_0/n7750 ) );
  nand_x1_sg U47831 ( .A(n12358), .B(n12359), .X(\shifter_0/n7746 ) );
  nand_x1_sg U47832 ( .A(n12362), .B(n12363), .X(\shifter_0/n7742 ) );
  nand_x1_sg U47833 ( .A(n12366), .B(n12367), .X(\shifter_0/n7738 ) );
  nand_x1_sg U47834 ( .A(n12370), .B(n12371), .X(\shifter_0/n7734 ) );
  nand_x1_sg U47835 ( .A(n12374), .B(n12375), .X(\shifter_0/n7730 ) );
  nand_x1_sg U47836 ( .A(n12378), .B(n12379), .X(\shifter_0/n7726 ) );
  nand_x1_sg U47837 ( .A(n12382), .B(n12383), .X(\shifter_0/n7722 ) );
  nand_x1_sg U47838 ( .A(n12386), .B(n12387), .X(\shifter_0/n7718 ) );
  nand_x1_sg U47839 ( .A(n12390), .B(n12391), .X(\shifter_0/n7714 ) );
  nand_x1_sg U47840 ( .A(n12394), .B(n12395), .X(\shifter_0/n7710 ) );
  nand_x1_sg U47841 ( .A(n12398), .B(n12399), .X(\shifter_0/n7706 ) );
  nand_x1_sg U47842 ( .A(n12402), .B(n12403), .X(\shifter_0/n7702 ) );
  nand_x1_sg U47843 ( .A(n12406), .B(n12407), .X(\shifter_0/n7698 ) );
  nand_x1_sg U47844 ( .A(n12410), .B(n12411), .X(\shifter_0/n7694 ) );
  nand_x1_sg U47845 ( .A(n12414), .B(n12415), .X(\shifter_0/n7690 ) );
  nand_x1_sg U47846 ( .A(n12418), .B(n12419), .X(\shifter_0/n7686 ) );
  nand_x1_sg U47847 ( .A(n12422), .B(n12423), .X(\shifter_0/n7682 ) );
  nand_x1_sg U47848 ( .A(n12426), .B(n12427), .X(\shifter_0/n7678 ) );
  nand_x1_sg U47849 ( .A(n12435), .B(n12436), .X(\shifter_0/n7674 ) );
  nand_x1_sg U47850 ( .A(n12442), .B(n12443), .X(\shifter_0/n7670 ) );
  nand_x1_sg U47851 ( .A(n12451), .B(n12452), .X(\shifter_0/n7662 ) );
  nand_x1_sg U47852 ( .A(n12460), .B(n12461), .X(\shifter_0/n7654 ) );
  nand_x1_sg U47853 ( .A(n12464), .B(n12465), .X(\shifter_0/n7650 ) );
  nand_x1_sg U47854 ( .A(n12468), .B(n12469), .X(\shifter_0/n7646 ) );
  nand_x1_sg U47855 ( .A(n12472), .B(n12473), .X(\shifter_0/n7642 ) );
  nand_x1_sg U47856 ( .A(n12476), .B(n12477), .X(\shifter_0/n7638 ) );
  nand_x1_sg U47857 ( .A(n12480), .B(n12481), .X(\shifter_0/n7634 ) );
  nand_x1_sg U47858 ( .A(n12484), .B(n12485), .X(\shifter_0/n7630 ) );
  nand_x1_sg U47859 ( .A(n12488), .B(n12489), .X(\shifter_0/n7626 ) );
  nand_x1_sg U47860 ( .A(n12492), .B(n12493), .X(\shifter_0/n7622 ) );
  nand_x1_sg U47861 ( .A(n12496), .B(n12497), .X(\shifter_0/n7618 ) );
  nand_x1_sg U47862 ( .A(n12500), .B(n12501), .X(\shifter_0/n7614 ) );
  nand_x1_sg U47863 ( .A(n12504), .B(n12505), .X(\shifter_0/n7610 ) );
  nand_x1_sg U47864 ( .A(n12518), .B(n12519), .X(\shifter_0/n7598 ) );
  nand_x1_sg U47865 ( .A(n11907), .B(n11908), .X(\shifter_0/n7910 ) );
  nand_x1_sg U47866 ( .A(n11929), .B(n11930), .X(\shifter_0/n7902 ) );
  nand_x1_sg U47867 ( .A(n11951), .B(n11952), .X(\shifter_0/n7894 ) );
  nand_x1_sg U47868 ( .A(n11973), .B(n11974), .X(\shifter_0/n7886 ) );
  nand_x1_sg U47869 ( .A(n11995), .B(n11996), .X(\shifter_0/n7878 ) );
  nand_x1_sg U47870 ( .A(n12017), .B(n12018), .X(\shifter_0/n7870 ) );
  nand_x1_sg U47871 ( .A(n12039), .B(n12040), .X(\shifter_0/n7862 ) );
  nand_x1_sg U47872 ( .A(n12135), .B(n12136), .X(\shifter_0/n7830 ) );
  nand_x1_sg U47873 ( .A(n12157), .B(n12158), .X(\shifter_0/n7822 ) );
  nand_x1_sg U47874 ( .A(n12179), .B(n12180), .X(\shifter_0/n7814 ) );
  nand_x1_sg U47875 ( .A(n12201), .B(n12202), .X(\shifter_0/n7806 ) );
  nand_x1_sg U47876 ( .A(n12223), .B(n12224), .X(\shifter_0/n7798 ) );
  nand_x1_sg U47877 ( .A(n12245), .B(n12246), .X(\shifter_0/n7790 ) );
  nand_x1_sg U47878 ( .A(n12267), .B(n12268), .X(\shifter_0/n7782 ) );
  nand_x1_sg U47879 ( .A(n11893), .B(n11894), .X(\shifter_0/n7914 ) );
  nand_x1_sg U47880 ( .A(n11918), .B(n11919), .X(\shifter_0/n7906 ) );
  nand_x1_sg U47881 ( .A(n11940), .B(n11941), .X(\shifter_0/n7898 ) );
  nand_x1_sg U47882 ( .A(n11962), .B(n11963), .X(\shifter_0/n7890 ) );
  nand_x1_sg U47883 ( .A(n11984), .B(n11985), .X(\shifter_0/n7882 ) );
  nand_x1_sg U47884 ( .A(n12006), .B(n12007), .X(\shifter_0/n7874 ) );
  nand_x1_sg U47885 ( .A(n12028), .B(n12029), .X(\shifter_0/n7866 ) );
  nand_x1_sg U47886 ( .A(n12050), .B(n12051), .X(\shifter_0/n7858 ) );
  nand_x1_sg U47887 ( .A(n12061), .B(n12062), .X(\shifter_0/n7854 ) );
  nand_x1_sg U47888 ( .A(n12072), .B(n12073), .X(\shifter_0/n7850 ) );
  nand_x1_sg U47889 ( .A(n12083), .B(n12084), .X(\shifter_0/n7846 ) );
  nand_x1_sg U47890 ( .A(n12094), .B(n12095), .X(\shifter_0/n7842 ) );
  nand_x1_sg U47891 ( .A(n12105), .B(n12106), .X(\shifter_0/n7838 ) );
  nand_x1_sg U47892 ( .A(n12121), .B(n12122), .X(\shifter_0/n7834 ) );
  nand_x1_sg U47893 ( .A(n12146), .B(n12147), .X(\shifter_0/n7826 ) );
  nand_x1_sg U47894 ( .A(n12168), .B(n12169), .X(\shifter_0/n7818 ) );
  nand_x1_sg U47895 ( .A(n12190), .B(n12191), .X(\shifter_0/n7810 ) );
  nand_x1_sg U47896 ( .A(n12212), .B(n12213), .X(\shifter_0/n7802 ) );
  nand_x1_sg U47897 ( .A(n12234), .B(n12235), .X(\shifter_0/n7794 ) );
  nand_x1_sg U47898 ( .A(n12256), .B(n12257), .X(\shifter_0/n7786 ) );
  nand_x1_sg U47899 ( .A(n12278), .B(n12279), .X(\shifter_0/n7778 ) );
  nand_x1_sg U47900 ( .A(n12289), .B(n12290), .X(\shifter_0/n7774 ) );
  nand_x1_sg U47901 ( .A(n12300), .B(n12301), .X(\shifter_0/n7770 ) );
  nand_x1_sg U47902 ( .A(n12311), .B(n12312), .X(\shifter_0/n7766 ) );
  nand_x1_sg U47903 ( .A(n12322), .B(n12323), .X(\shifter_0/n7762 ) );
  nand_x1_sg U47904 ( .A(n12333), .B(n12334), .X(\shifter_0/n7758 ) );
  nand_x1_sg U47905 ( .A(n20975), .B(n20976), .X(n20974) );
  nand_x1_sg U47906 ( .A(n20964), .B(n20965), .X(n20963) );
  nand_x1_sg U47907 ( .A(n21474), .B(n21475), .X(n21473) );
  nand_x1_sg U47908 ( .A(n20995), .B(n20996), .X(n20994) );
  nand_x1_sg U47909 ( .A(n21381), .B(n21382), .X(n21380) );
  nand_x1_sg U47910 ( .A(n21568), .B(n21569), .X(n21567) );
  nor_x1_sg U47911 ( .A(n11640), .B(n34435), .X(n11664) );
  nor_x1_sg U47912 ( .A(n11798), .B(n35655), .X(n11843) );
  nor_x1_sg U47913 ( .A(n41499), .B(n32186), .X(n12120) );
  inv_x1_sg U47914 ( .A(n11843), .X(n41499) );
  inv_x1_sg U47915 ( .A(n11798), .X(n41418) );
  inv_x1_sg U47916 ( .A(n11640), .X(n41183) );
  nand_x1_sg U47917 ( .A(n30539), .B(n35656), .X(n11798) );
  nand_x1_sg U47918 ( .A(n11559), .B(n35456), .X(n11640) );
  nor_x1_sg U47919 ( .A(n33763), .B(n34067), .X(n35676) );
  nor_x1_sg U47920 ( .A(n42544), .B(n31704), .X(n21006) );
  nor_x1_sg U47921 ( .A(n42543), .B(n32024), .X(n21005) );
  nor_x1_sg U47922 ( .A(n42539), .B(n35278), .X(n21365) );
  nor_x1_sg U47923 ( .A(n42541), .B(n31704), .X(n21364) );
  nor_x1_sg U47924 ( .A(n42540), .B(n32022), .X(n21363) );
  nor_x1_sg U47925 ( .A(n32023), .B(n32509), .X(n19585) );
  nor_x1_sg U47926 ( .A(n31601), .B(n33962), .X(n12116) );
  nor_x1_sg U47927 ( .A(n31601), .B(n32510), .X(n11716) );
  nor_x1_sg U47928 ( .A(n35098), .B(n33805), .X(n35651) );
  nor_x1_sg U47929 ( .A(n35098), .B(n33814), .X(n11895) );
  nor_x1_sg U47930 ( .A(n34444), .B(n31980), .X(n11559) );
  nor_x1_sg U47931 ( .A(n31705), .B(n32508), .X(n13291) );
  nor_x1_sg U47932 ( .A(n30977), .B(n30535), .X(n11906) );
  nor_x1_sg U47933 ( .A(n33804), .B(n12116), .X(n12134) );
  nor_x1_sg U47934 ( .A(n19584), .B(n32507), .X(n19582) );
  nor_x1_sg U47935 ( .A(n33622), .B(n34070), .X(n35663) );
  nor_x1_sg U47936 ( .A(n33598), .B(n34070), .X(n29447) );
  nor_x1_sg U47937 ( .A(n33606), .B(n34066), .X(n35664) );
  nor_x1_sg U47938 ( .A(n33702), .B(n34065), .X(n29623) );
  nor_x1_sg U47939 ( .A(n33771), .B(n34066), .X(n35678) );
  nor_x1_sg U47940 ( .A(n33566), .B(n34068), .X(n35675) );
  nor_x1_sg U47941 ( .A(n33574), .B(n34070), .X(n35673) );
  nor_x1_sg U47942 ( .A(n33678), .B(n34069), .X(n28705) );
  nor_x1_sg U47943 ( .A(n33638), .B(n34064), .X(n35680) );
  nor_x1_sg U47944 ( .A(n33646), .B(n34064), .X(n28621) );
  nor_x1_sg U47945 ( .A(n33662), .B(n34063), .X(n35672) );
  nor_x1_sg U47946 ( .A(n33686), .B(n34062), .X(n35681) );
  nor_x1_sg U47947 ( .A(n33787), .B(n34065), .X(n28452) );
  nor_x1_sg U47948 ( .A(n33542), .B(n34069), .X(n35674) );
  nor_x1_sg U47949 ( .A(n33550), .B(n34069), .X(n35671) );
  nor_x1_sg U47950 ( .A(n33534), .B(n34066), .X(n35660) );
  nor_x1_sg U47951 ( .A(n33694), .B(n34068), .X(n35658) );
  nor_x1_sg U47952 ( .A(n33526), .B(n34068), .X(n35670) );
  nor_x1_sg U47953 ( .A(n21089), .B(n21090), .X(n21088) );
  nor_x1_sg U47954 ( .A(n21127), .B(n21128), .X(n21087) );
  nand_x4_sg U47955 ( .A(n21003), .B(n21004), .X(n20940) );
  nor_x1_sg U47956 ( .A(n21165), .B(n21166), .X(n21003) );
  nor_x1_sg U47957 ( .A(n21005), .B(n21006), .X(n21004) );
  nor_x1_sg U47958 ( .A(n20916), .B(n31663), .X(n21166) );
  nor_x1_sg U47959 ( .A(n21010), .B(n21011), .X(n21009) );
  nor_x1_sg U47960 ( .A(n21048), .B(n21049), .X(n21008) );
  nand_x4_sg U47961 ( .A(n21361), .B(n21362), .X(n21336) );
  nor_x1_sg U47962 ( .A(n21365), .B(n21366), .X(n21361) );
  nor_x1_sg U47963 ( .A(n21363), .B(n21364), .X(n21362) );
  nor_x1_sg U47964 ( .A(n21367), .B(n31663), .X(n21366) );
  nor_x1_sg U47965 ( .A(n21485), .B(n21486), .X(n21484) );
  nor_x1_sg U47966 ( .A(n21523), .B(n21524), .X(n21483) );
  nor_x1_sg U47967 ( .A(n21393), .B(n21394), .X(n21392) );
  nor_x1_sg U47968 ( .A(n21431), .B(n21432), .X(n21391) );
  nor_x1_sg U47969 ( .A(n21580), .B(n21581), .X(n21579) );
  nor_x1_sg U47970 ( .A(n21618), .B(n21619), .X(n21578) );
  nor_x1_sg U47971 ( .A(n42542), .B(n35278), .X(n21165) );
  nor_x1_sg U47972 ( .A(n19585), .B(n19600), .X(n19598) );
  nor_x1_sg U47973 ( .A(n35100), .B(n42536), .X(n21335) );
  nor_x1_sg U47974 ( .A(n35101), .B(n35563), .X(n20957) );
  nor_x1_sg U47975 ( .A(n31706), .B(n32517), .X(n13699) );
  nor_x1_sg U47976 ( .A(n32519), .B(n19584), .X(n11611) );
  nor_x1_sg U47977 ( .A(n32219), .B(n35158), .X(n13804) );
  nor_x1_sg U47978 ( .A(n33960), .B(n32932), .X(n13805) );
  nor_x1_sg U47979 ( .A(n32518), .B(n32933), .X(n13816) );
  nor_x1_sg U47980 ( .A(n31666), .B(n31705), .X(n13290) );
  nor_x1_sg U47981 ( .A(n31652), .B(n31663), .X(n35657) );
  nor_x1_sg U47982 ( .A(n32509), .B(n32934), .X(n35650) );
  nor_x1_sg U47983 ( .A(n32024), .B(n32520), .X(n12834) );
  inv_x1_sg U47984 ( .A(n11663), .X(n41110) );
  nor_x1_sg U47985 ( .A(n13097), .B(n32519), .X(n13096) );
  nand_x1_sg U47986 ( .A(n34516), .B(n11663), .X(n11711) );
  nand_x1_sg U47987 ( .A(n32420), .B(n11635), .X(n11738) );
  nand_x1_sg U47988 ( .A(n32410), .B(n11635), .X(n11792) );
  nor_x1_sg U47989 ( .A(n32056), .B(n34859), .X(n19588) );
  nor_x1_sg U47990 ( .A(n42537), .B(n31604), .X(n35684) );
  inv_x1_sg U47991 ( .A(n19607), .X(n42537) );
  nor_x1_sg U47992 ( .A(n31603), .B(n33825), .X(n18763) );
  nor_x1_sg U47993 ( .A(n29755), .B(n42407), .X(n35683) );
  nor_x1_sg U47994 ( .A(n19608), .B(n31604), .X(n19602) );
  nand_x1_sg U47995 ( .A(n42537), .B(n19609), .X(n19608) );
  nor_x1_sg U47996 ( .A(n33514), .B(n34065), .X(n35668) );
  nor_x1_sg U47997 ( .A(n33670), .B(n34070), .X(n35662) );
  nor_x1_sg U47998 ( .A(n33490), .B(n34062), .X(n28978) );
  nor_x1_sg U47999 ( .A(n33482), .B(n34063), .X(n29492) );
  nor_x1_sg U48000 ( .A(n33474), .B(n34066), .X(n35659) );
  nand_x1_sg U48001 ( .A(n32169), .B(n32935), .X(n19584) );
  nand_x1_sg U48002 ( .A(n28790), .B(n35270), .X(n28789) );
  nor_x1_sg U48003 ( .A(n32508), .B(n20981), .X(n21128) );
  nor_x1_sg U48004 ( .A(n32508), .B(n20971), .X(n21049) );
  nor_x1_sg U48005 ( .A(n32507), .B(n21001), .X(n21266) );
  nor_x1_sg U48006 ( .A(n32507), .B(n21480), .X(n21524) );
  nor_x1_sg U48007 ( .A(n32509), .B(n21387), .X(n21432) );
  nor_x1_sg U48008 ( .A(n32510), .B(n21574), .X(n21619) );
  nor_x1_sg U48009 ( .A(n21227), .B(n21228), .X(n21226) );
  nor_x1_sg U48010 ( .A(n21265), .B(n21266), .X(n21225) );
  nor_x1_sg U48011 ( .A(n33959), .B(n20997), .X(n21228) );
  nand_x1_sg U48012 ( .A(n20919), .B(n31708), .X(n20918) );
  nor_x1_sg U48013 ( .A(n30136), .B(n32896), .X(n20968) );
  nor_x1_sg U48014 ( .A(n42546), .B(n21167), .X(n20916) );
  nor_x1_sg U48015 ( .A(n20991), .B(n32517), .X(n21167) );
  nor_x1_sg U48016 ( .A(n21187), .B(n21188), .X(n21186) );
  nor_x1_sg U48017 ( .A(n32219), .B(n20992), .X(n21187) );
  nor_x1_sg U48018 ( .A(n42545), .B(n21667), .X(n21367) );
  nor_x1_sg U48019 ( .A(n21665), .B(n32520), .X(n21667) );
  nor_x1_sg U48020 ( .A(n21687), .B(n21688), .X(n21686) );
  nor_x1_sg U48021 ( .A(n32221), .B(n21666), .X(n21687) );
  nor_x1_sg U48022 ( .A(n20960), .B(n20961), .X(n20959) );
  nor_x1_sg U48023 ( .A(n20983), .B(n20984), .X(n20958) );
  nor_x1_sg U48024 ( .A(n20928), .B(n32022), .X(n20960) );
  nor_x1_sg U48025 ( .A(n21353), .B(n21354), .X(n21352) );
  nor_x1_sg U48026 ( .A(n21357), .B(n21358), .X(n21351) );
  nor_x1_sg U48027 ( .A(n21356), .B(n32023), .X(n21353) );
  nor_x1_sg U48028 ( .A(n32220), .B(n20978), .X(n21089) );
  nor_x1_sg U48029 ( .A(n32220), .B(n20967), .X(n21010) );
  nor_x1_sg U48030 ( .A(n32222), .B(n20998), .X(n21227) );
  nor_x1_sg U48031 ( .A(n32222), .B(n21477), .X(n21485) );
  nor_x1_sg U48032 ( .A(n32221), .B(n21384), .X(n21393) );
  nor_x1_sg U48033 ( .A(n32219), .B(n21571), .X(n21580) );
  nand_x1_sg U48034 ( .A(n19594), .B(n32167), .X(n19595) );
  nand_x1_sg U48035 ( .A(n35266), .B(n19597), .X(n19596) );
  nand_x1_sg U48036 ( .A(n19598), .B(n19599), .X(n19597) );
  nand_x1_sg U48037 ( .A(n32940), .B(n20900), .X(n20899) );
  nand_x1_sg U48038 ( .A(n30585), .B(n31992), .X(n20898) );
  nand_x1_sg U48039 ( .A(n35463), .B(n20901), .X(n20900) );
  nor_x1_sg U48040 ( .A(n20931), .B(n32937), .X(n20930) );
  nor_x1_sg U48041 ( .A(n31708), .B(n20932), .X(n20931) );
  nand_x1_sg U48042 ( .A(n20967), .B(n20968), .X(n20964) );
  nor_x1_sg U48043 ( .A(n33959), .B(n20988), .X(n21188) );
  nor_x1_sg U48044 ( .A(n32517), .B(n20982), .X(n21127) );
  nor_x1_sg U48045 ( .A(n32938), .B(n20920), .X(n20917) );
  nor_x1_sg U48046 ( .A(n20921), .B(n35303), .X(n20920) );
  nand_x1_sg U48047 ( .A(n20998), .B(n20968), .X(n20995) );
  nand_x1_sg U48048 ( .A(n20978), .B(n20968), .X(n20975) );
  nand_x1_sg U48049 ( .A(n20971), .B(n31665), .X(n20970) );
  nor_x1_sg U48050 ( .A(n32519), .B(n21002), .X(n21265) );
  nor_x1_sg U48051 ( .A(n32518), .B(n21481), .X(n21523) );
  nand_x1_sg U48052 ( .A(n21001), .B(n31666), .X(n21000) );
  nor_x1_sg U48053 ( .A(n20921), .B(n35278), .X(n20983) );
  nor_x1_sg U48054 ( .A(n20932), .B(n31705), .X(n20961) );
  nor_x1_sg U48055 ( .A(n21355), .B(n31706), .X(n21354) );
  nand_x1_sg U48056 ( .A(n20981), .B(n31666), .X(n20980) );
  nand_x1_sg U48057 ( .A(n21384), .B(n31600), .X(n21381) );
  nand_x1_sg U48058 ( .A(n21477), .B(n31600), .X(n21474) );
  nor_x1_sg U48059 ( .A(n21360), .B(n35278), .X(n21357) );
  nor_x1_sg U48060 ( .A(n32520), .B(n20972), .X(n21048) );
  nand_x1_sg U48061 ( .A(n21571), .B(n31600), .X(n21568) );
  nor_x1_sg U48062 ( .A(n32518), .B(n21388), .X(n21431) );
  nor_x1_sg U48063 ( .A(n32519), .B(n21575), .X(n21618) );
  nor_x1_sg U48064 ( .A(n33961), .B(n21662), .X(n21688) );
  nand_x1_sg U48065 ( .A(n35266), .B(n32507), .X(n20901) );
  nand_x1_sg U48066 ( .A(n30784), .B(n32510), .X(n19599) );
  nor_x1_sg U48067 ( .A(n33960), .B(n20977), .X(n21090) );
  nor_x1_sg U48068 ( .A(n31670), .B(n21360), .X(n21565) );
  nand_x1_sg U48069 ( .A(n21574), .B(n31665), .X(n21573) );
  nand_x1_sg U48070 ( .A(n21387), .B(n31665), .X(n21386) );
  nand_x1_sg U48071 ( .A(n21480), .B(n31666), .X(n21479) );
  nor_x1_sg U48072 ( .A(n31668), .B(n21355), .X(n21378) );
  nand_x1_sg U48073 ( .A(n32426), .B(n35104), .X(n29148) );
  nor_x1_sg U48074 ( .A(n33962), .B(n21570), .X(n21581) );
  nor_x1_sg U48075 ( .A(n30016), .B(n20966), .X(n21011) );
  nor_x1_sg U48076 ( .A(n31652), .B(n21476), .X(n21486) );
  nor_x1_sg U48077 ( .A(n31653), .B(n21383), .X(n21394) );
  nor_x1_sg U48078 ( .A(n35158), .B(n34549), .X(n13221) );
  nor_x1_sg U48079 ( .A(n31604), .B(n33819), .X(n35685) );
  nor_x1_sg U48080 ( .A(n31603), .B(n35266), .X(n19594) );
  nand_x1_sg U48081 ( .A(n20966), .B(n33985), .X(n20965) );
  nand_x1_sg U48082 ( .A(n20977), .B(n33986), .X(n20976) );
  nand_x1_sg U48083 ( .A(n20997), .B(n33987), .X(n20996) );
  nand_x1_sg U48084 ( .A(n21570), .B(n30908), .X(n21569) );
  nand_x1_sg U48085 ( .A(n21662), .B(n31696), .X(n21661) );
  nand_x1_sg U48086 ( .A(n21476), .B(n30909), .X(n21475) );
  nor_x1_sg U48087 ( .A(n32395), .B(n32936), .X(n19600) );
  nand_x1_sg U48088 ( .A(n21383), .B(n33984), .X(n21382) );
  nor_x1_sg U48089 ( .A(n32936), .B(n34550), .X(n13224) );
  nand_x1_sg U48090 ( .A(n30585), .B(n34806), .X(n19592) );
  nand_x1_sg U48091 ( .A(n19594), .B(n34858), .X(n19593) );
  nand_x1_sg U48092 ( .A(n20991), .B(n29771), .X(n20990) );
  nand_x1_sg U48093 ( .A(n21665), .B(n32889), .X(n21664) );
  inv_x1_sg U48094 ( .A(n12968), .X(n42536) );
  nor_x1_sg U48095 ( .A(n33964), .B(n35582), .X(n15052) );
  nor_x1_sg U48096 ( .A(n35304), .B(n35280), .X(n11635) );
  nand_x1_sg U48097 ( .A(n28790), .B(n31662), .X(n15056) );
  nor_x1_sg U48098 ( .A(n32220), .B(n32940), .X(n14496) );
  nor_x1_sg U48099 ( .A(n29688), .B(n32937), .X(n14497) );
  nor_x1_sg U48100 ( .A(n35302), .B(n35279), .X(n11663) );
  nand_x1_sg U48101 ( .A(n35529), .B(n42402), .X(n35632) );
  nand_x1_sg U48102 ( .A(n35552), .B(n35553), .X(n35630) );
  nand_x1_sg U48103 ( .A(n35552), .B(n35504), .X(n35629) );
  nand_x1_sg U48104 ( .A(n32925), .B(n32390), .X(n12533) );
  nor_x1_sg U48105 ( .A(n32387), .B(n41139), .X(n12630) );
  nor_x1_sg U48106 ( .A(n32392), .B(n41140), .X(n12639) );
  nor_x1_sg U48107 ( .A(n32388), .B(n41141), .X(n12692) );
  nor_x1_sg U48108 ( .A(n32391), .B(n41142), .X(n12697) );
  nand_x1_sg U48109 ( .A(n35529), .B(n35516), .X(n35633) );
  nor_x1_sg U48110 ( .A(n34560), .B(n32922), .X(n35647) );
  nor_x1_sg U48111 ( .A(n34561), .B(n32917), .X(n35641) );
  nand_x1_sg U48112 ( .A(n32054), .B(n30143), .X(n12717) );
  nor_x1_sg U48113 ( .A(n32917), .B(n32171), .X(n35640) );
  nor_x1_sg U48114 ( .A(n33836), .B(n34548), .X(n12531) );
  nor_x1_sg U48115 ( .A(n32396), .B(n33809), .X(n12353) );
  nor_x1_sg U48116 ( .A(n32397), .B(n30985), .X(n12976) );
  nor_x1_sg U48117 ( .A(n32922), .B(n31299), .X(n35646) );
  nand_x1_sg U48118 ( .A(n13220), .B(n31867), .X(n13219) );
  nand_x1_sg U48119 ( .A(n13223), .B(n12968), .X(n13218) );
  nor_x1_sg U48120 ( .A(n30525), .B(n33962), .X(n13220) );
  nor_x1_sg U48121 ( .A(n30979), .B(n34559), .X(n35648) );
  nor_x1_sg U48122 ( .A(n29750), .B(n31704), .X(n13787) );
  nor_x1_sg U48123 ( .A(n30011), .B(n34551), .X(n35642) );
  nand_x1_sg U48124 ( .A(n13781), .B(n31983), .X(n14411) );
  nor_x1_sg U48125 ( .A(n35563), .B(n35105), .X(n13097) );
  nor_x1_sg U48126 ( .A(n12630), .B(n14481), .X(n13301) );
  nor_x1_sg U48127 ( .A(n32023), .B(n41135), .X(n14481) );
  nor_x1_sg U48128 ( .A(n12639), .B(n14545), .X(n13308) );
  nor_x1_sg U48129 ( .A(n32022), .B(n41136), .X(n14545) );
  nor_x1_sg U48130 ( .A(n12692), .B(n14948), .X(n13348) );
  nor_x1_sg U48131 ( .A(n32024), .B(n41137), .X(n14948) );
  nor_x1_sg U48132 ( .A(n12697), .B(n14979), .X(n13352) );
  nor_x1_sg U48133 ( .A(n32024), .B(n41138), .X(n14979) );
  nor_x1_sg U48134 ( .A(n35158), .B(n34545), .X(n12839) );
  nand_x1_sg U48135 ( .A(n31507), .B(n13781), .X(n13778) );
  nand_x1_sg U48136 ( .A(n33957), .B(n13700), .X(n13696) );
  nor_x1_sg U48137 ( .A(n12610), .B(n35419), .X(n35645) );
  nor_x1_sg U48138 ( .A(n12703), .B(n41705), .X(n35644) );
  nand_x1_sg U48139 ( .A(n12840), .B(n34559), .X(n12433) );
  nor_x1_sg U48140 ( .A(n32022), .B(n30137), .X(n12613) );
  nor_x1_sg U48141 ( .A(n13290), .B(n35101), .X(n13289) );
  nor_x1_sg U48142 ( .A(n34429), .B(n42547), .X(n13698) );
  nand_x1_sg U48143 ( .A(n13097), .B(n30784), .X(n13091) );
  nand_x1_sg U48144 ( .A(n11713), .B(n30527), .X(n11712) );
  nand_x1_sg U48145 ( .A(n11740), .B(n30529), .X(n11739) );
  nor_x1_sg U48146 ( .A(n32520), .B(n32938), .X(n13808) );
  nor_x1_sg U48147 ( .A(n13290), .B(n35100), .X(n13359) );
  nor_x1_sg U48148 ( .A(n34430), .B(n42533), .X(n13780) );
  nor_x1_sg U48149 ( .A(n13608), .B(n33828), .X(n13613) );
  nand_x1_sg U48150 ( .A(n34537), .B(n31696), .X(n35634) );
  nand_x1_sg U48151 ( .A(n13608), .B(n31704), .X(n13607) );
  nand_x1_sg U48152 ( .A(n42402), .B(n35250), .X(n15037) );
  nand_x1_sg U48153 ( .A(n35510), .B(n35250), .X(n15038) );
  nand_x1_sg U48154 ( .A(n35516), .B(n35250), .X(n15039) );
  nand_x1_sg U48155 ( .A(n35530), .B(n35249), .X(n15170) );
  nand_x1_sg U48156 ( .A(n35553), .B(n35249), .X(n15172) );
  nand_x1_sg U48157 ( .A(n12968), .B(n32170), .X(n12525) );
  nor_x1_sg U48158 ( .A(n30134), .B(n35106), .X(n13223) );
  nor_x1_sg U48159 ( .A(n11843), .B(n42533), .X(n11890) );
  nor_x1_sg U48160 ( .A(n13095), .B(n13096), .X(n13094) );
  nor_x1_sg U48161 ( .A(n13098), .B(n32023), .X(n13093) );
  nor_x1_sg U48162 ( .A(n13097), .B(n31303), .X(n13095) );
  nor_x1_sg U48163 ( .A(n35262), .B(n35099), .X(n15035) );
  nor_x1_sg U48164 ( .A(n35262), .B(n41110), .X(n15034) );
  nor_x1_sg U48165 ( .A(n34445), .B(n31709), .X(n11560) );
  nor_x1_sg U48166 ( .A(n32192), .B(n31669), .X(n11585) );
  nor_x1_sg U48167 ( .A(n14062), .B(n14063), .X(n14052) );
  nand_x1_sg U48168 ( .A(n14065), .B(n14066), .X(n14062) );
  nor_x1_sg U48169 ( .A(n14093), .B(n14094), .X(n14083) );
  nand_x1_sg U48170 ( .A(n14096), .B(n14097), .X(n14093) );
  nor_x1_sg U48171 ( .A(n14186), .B(n14187), .X(n14176) );
  nand_x1_sg U48172 ( .A(n14189), .B(n14190), .X(n14186) );
  nor_x1_sg U48173 ( .A(n14217), .B(n14218), .X(n14207) );
  nand_x1_sg U48174 ( .A(n14220), .B(n14221), .X(n14217) );
  inv_x1_sg U48175 ( .A(n19583), .X(n41109) );
  nand_x1_sg U48176 ( .A(n35303), .B(n35279), .X(n11770) );
  nor_x1_sg U48177 ( .A(n29988), .B(n35537), .X(\shifter_0/n6553 ) );
  nor_x1_sg U48178 ( .A(n33004), .B(n35520), .X(\shifter_0/n6549 ) );
  nor_x1_sg U48179 ( .A(n33003), .B(n35550), .X(\shifter_0/n6545 ) );
  nor_x1_sg U48180 ( .A(n33005), .B(n14507), .X(\shifter_0/n6541 ) );
  nor_x1_sg U48181 ( .A(n33006), .B(n35471), .X(\shifter_0/n6537 ) );
  nor_x1_sg U48182 ( .A(n33004), .B(n35536), .X(\shifter_0/n6533 ) );
  nor_x1_sg U48183 ( .A(n33005), .B(n35535), .X(\shifter_0/n6529 ) );
  nor_x1_sg U48184 ( .A(n35405), .B(n35534), .X(\shifter_0/n6525 ) );
  nor_x1_sg U48185 ( .A(n33003), .B(n35496), .X(\shifter_0/n6521 ) );
  nor_x1_sg U48186 ( .A(n33003), .B(n35470), .X(\shifter_0/n6517 ) );
  nor_x1_sg U48187 ( .A(n33004), .B(n35519), .X(\shifter_0/n6513 ) );
  nor_x1_sg U48188 ( .A(n33005), .B(n35518), .X(\shifter_0/n6509 ) );
  nor_x1_sg U48189 ( .A(n29988), .B(n35468), .X(\shifter_0/n6505 ) );
  nor_x1_sg U48190 ( .A(n33005), .B(n35495), .X(\shifter_0/n6501 ) );
  nor_x1_sg U48191 ( .A(n33006), .B(n35533), .X(\shifter_0/n6497 ) );
  nor_x1_sg U48192 ( .A(n33006), .B(n35532), .X(\shifter_0/n6493 ) );
  nor_x1_sg U48193 ( .A(n33004), .B(n35531), .X(\shifter_0/n6489 ) );
  nor_x1_sg U48194 ( .A(n35405), .B(n35469), .X(\shifter_0/n6485 ) );
  nor_x1_sg U48195 ( .A(n33003), .B(n35467), .X(\shifter_0/n6481 ) );
  nor_x1_sg U48196 ( .A(n33006), .B(n35517), .X(\shifter_0/n6477 ) );
  inv_x1_sg U48197 ( .A(n13372), .X(n41410) );
  inv_x1_sg U48198 ( .A(n13378), .X(n41406) );
  inv_x1_sg U48199 ( .A(n13402), .X(n41390) );
  inv_x1_sg U48200 ( .A(n13426), .X(n41374) );
  inv_x1_sg U48201 ( .A(n13432), .X(n41370) );
  inv_x1_sg U48202 ( .A(n13456), .X(n41354) );
  inv_x1_sg U48203 ( .A(n13480), .X(n41338) );
  inv_x1_sg U48204 ( .A(n13493), .X(n41337) );
  inv_x1_sg U48205 ( .A(n13527), .X(n41333) );
  inv_x1_sg U48206 ( .A(n13551), .X(n41329) );
  inv_x1_sg U48207 ( .A(n13557), .X(n41328) );
  inv_x1_sg U48208 ( .A(n13581), .X(n41324) );
  inv_x1_sg U48209 ( .A(n13364), .X(n41414) );
  inv_x1_sg U48210 ( .A(n13384), .X(n41402) );
  inv_x1_sg U48211 ( .A(n13390), .X(n41398) );
  inv_x1_sg U48212 ( .A(n13396), .X(n41394) );
  inv_x1_sg U48213 ( .A(n13408), .X(n41386) );
  inv_x1_sg U48214 ( .A(n13414), .X(n41382) );
  inv_x1_sg U48215 ( .A(n13420), .X(n41378) );
  inv_x1_sg U48216 ( .A(n13438), .X(n41366) );
  inv_x1_sg U48217 ( .A(n13444), .X(n41362) );
  inv_x1_sg U48218 ( .A(n13450), .X(n41358) );
  inv_x1_sg U48219 ( .A(n13462), .X(n41350) );
  inv_x1_sg U48220 ( .A(n13468), .X(n41346) );
  inv_x1_sg U48221 ( .A(n13474), .X(n41342) );
  inv_x1_sg U48222 ( .A(n13499), .X(n41336) );
  inv_x1_sg U48223 ( .A(n13510), .X(n41335) );
  inv_x1_sg U48224 ( .A(n13521), .X(n41334) );
  inv_x1_sg U48225 ( .A(n13533), .X(n41332) );
  inv_x1_sg U48226 ( .A(n13539), .X(n41331) );
  inv_x1_sg U48227 ( .A(n13545), .X(n41330) );
  inv_x1_sg U48228 ( .A(n13563), .X(n41327) );
  inv_x1_sg U48229 ( .A(n13569), .X(n41326) );
  inv_x1_sg U48230 ( .A(n13575), .X(n41325) );
  inv_x1_sg U48231 ( .A(n13587), .X(n41323) );
  inv_x1_sg U48232 ( .A(n13603), .X(n41322) );
  nor_x1_sg U48233 ( .A(n32984), .B(n35523), .X(\shifter_0/n6633 ) );
  nor_x1_sg U48234 ( .A(n32986), .B(n35546), .X(\shifter_0/n6629 ) );
  nor_x1_sg U48235 ( .A(n32983), .B(n35545), .X(\shifter_0/n6625 ) );
  nor_x1_sg U48236 ( .A(n32984), .B(n35502), .X(\shifter_0/n6621 ) );
  nor_x1_sg U48237 ( .A(n32984), .B(n35501), .X(\shifter_0/n6617 ) );
  nor_x1_sg U48238 ( .A(n32985), .B(n35544), .X(\shifter_0/n6613 ) );
  nor_x1_sg U48239 ( .A(n29990), .B(n35543), .X(\shifter_0/n6609 ) );
  nor_x1_sg U48240 ( .A(n32983), .B(n35542), .X(\shifter_0/n6605 ) );
  nor_x1_sg U48241 ( .A(n32985), .B(n35500), .X(\shifter_0/n6601 ) );
  nor_x1_sg U48242 ( .A(n32983), .B(n35473), .X(\shifter_0/n6597 ) );
  nor_x1_sg U48243 ( .A(n32986), .B(n35541), .X(\shifter_0/n6593 ) );
  nor_x1_sg U48244 ( .A(n32986), .B(n35522), .X(\shifter_0/n6589 ) );
  nor_x1_sg U48245 ( .A(n32985), .B(n35499), .X(\shifter_0/n6585 ) );
  nor_x1_sg U48246 ( .A(n29990), .B(n35498), .X(\shifter_0/n6581 ) );
  nor_x1_sg U48247 ( .A(n32984), .B(n35540), .X(\shifter_0/n6577 ) );
  nor_x1_sg U48248 ( .A(n41321), .B(n35539), .X(\shifter_0/n6573 ) );
  nor_x1_sg U48249 ( .A(n32985), .B(n35538), .X(\shifter_0/n6569 ) );
  nor_x1_sg U48250 ( .A(n41321), .B(n35472), .X(\shifter_0/n6565 ) );
  nor_x1_sg U48251 ( .A(n32983), .B(n35497), .X(\shifter_0/n6561 ) );
  nor_x1_sg U48252 ( .A(n32986), .B(n35521), .X(\shifter_0/n6557 ) );
  nor_x1_sg U48253 ( .A(n33018), .B(n35549), .X(\shifter_0/n6953 ) );
  nor_x1_sg U48254 ( .A(n30004), .B(n35557), .X(\shifter_0/n6949 ) );
  nor_x1_sg U48255 ( .A(n35244), .B(n35548), .X(\shifter_0/n6945 ) );
  nor_x1_sg U48256 ( .A(n30004), .B(n35559), .X(\shifter_0/n6941 ) );
  nor_x1_sg U48257 ( .A(n33019), .B(n35556), .X(\shifter_0/n6937 ) );
  nor_x1_sg U48258 ( .A(n33021), .B(n35555), .X(\shifter_0/n6933 ) );
  nor_x1_sg U48259 ( .A(n33021), .B(n35554), .X(\shifter_0/n6929 ) );
  nor_x1_sg U48260 ( .A(n33019), .B(n35547), .X(\shifter_0/n6925 ) );
  nor_x1_sg U48261 ( .A(n33020), .B(n35526), .X(\shifter_0/n6921 ) );
  nor_x1_sg U48262 ( .A(n33019), .B(n35525), .X(\shifter_0/n6917 ) );
  nor_x1_sg U48263 ( .A(n33019), .B(n35524), .X(\shifter_0/n6913 ) );
  nor_x1_sg U48264 ( .A(n33020), .B(n35494), .X(\shifter_0/n6909 ) );
  nor_x1_sg U48265 ( .A(n33018), .B(n35493), .X(\shifter_0/n6905 ) );
  nor_x1_sg U48266 ( .A(n33018), .B(n35492), .X(\shifter_0/n6901 ) );
  nor_x1_sg U48267 ( .A(n35244), .B(n35491), .X(\shifter_0/n6897 ) );
  nor_x1_sg U48268 ( .A(n33021), .B(n35490), .X(\shifter_0/n6893 ) );
  nor_x1_sg U48269 ( .A(n33021), .B(n35482), .X(\shifter_0/n6889 ) );
  nor_x1_sg U48270 ( .A(n33018), .B(n35489), .X(\shifter_0/n6885 ) );
  nor_x1_sg U48271 ( .A(n33020), .B(n35488), .X(\shifter_0/n6881 ) );
  nor_x1_sg U48272 ( .A(n33020), .B(n35487), .X(\shifter_0/n6877 ) );
  nor_x1_sg U48273 ( .A(n29994), .B(n35449), .X(\shifter_0/n7433 ) );
  nor_x1_sg U48274 ( .A(n32996), .B(n12719), .X(\shifter_0/n7429 ) );
  nor_x1_sg U48275 ( .A(n32993), .B(n35450), .X(\shifter_0/n7425 ) );
  nor_x1_sg U48276 ( .A(n32993), .B(n12731), .X(\shifter_0/n7421 ) );
  nor_x1_sg U48277 ( .A(n32996), .B(n12737), .X(\shifter_0/n7417 ) );
  nor_x1_sg U48278 ( .A(n32996), .B(n35451), .X(\shifter_0/n7413 ) );
  nor_x1_sg U48279 ( .A(n35407), .B(n35452), .X(\shifter_0/n7409 ) );
  nor_x1_sg U48280 ( .A(n32993), .B(n12755), .X(\shifter_0/n7405 ) );
  nor_x1_sg U48281 ( .A(n32994), .B(n35445), .X(\shifter_0/n7401 ) );
  nor_x1_sg U48282 ( .A(n32995), .B(n35446), .X(\shifter_0/n7397 ) );
  nor_x1_sg U48283 ( .A(n32994), .B(n35447), .X(\shifter_0/n7393 ) );
  nor_x1_sg U48284 ( .A(n29994), .B(n35448), .X(\shifter_0/n7389 ) );
  nor_x1_sg U48285 ( .A(n32994), .B(n12785), .X(\shifter_0/n7385 ) );
  nor_x1_sg U48286 ( .A(n32995), .B(n35441), .X(\shifter_0/n7381 ) );
  nor_x1_sg U48287 ( .A(n35407), .B(n12797), .X(\shifter_0/n7377 ) );
  nor_x1_sg U48288 ( .A(n32995), .B(n35442), .X(\shifter_0/n7373 ) );
  nor_x1_sg U48289 ( .A(n32996), .B(n35443), .X(\shifter_0/n7369 ) );
  nor_x1_sg U48290 ( .A(n32995), .B(n35444), .X(\shifter_0/n7365 ) );
  nor_x1_sg U48291 ( .A(n32994), .B(n35437), .X(\shifter_0/n7361 ) );
  nor_x1_sg U48292 ( .A(n32993), .B(n35438), .X(\shifter_0/n7357 ) );
  nor_x1_sg U48293 ( .A(n32989), .B(n35439), .X(\shifter_0/n7353 ) );
  nor_x1_sg U48294 ( .A(n32991), .B(n35440), .X(\shifter_0/n7349 ) );
  nor_x1_sg U48295 ( .A(n35408), .B(n35433), .X(\shifter_0/n7345 ) );
  nor_x1_sg U48296 ( .A(n32988), .B(n12861), .X(\shifter_0/n7341 ) );
  nor_x1_sg U48297 ( .A(n32988), .B(n35434), .X(\shifter_0/n7337 ) );
  nor_x1_sg U48298 ( .A(n30012), .B(n35435), .X(\shifter_0/n7333 ) );
  nor_x1_sg U48299 ( .A(n32988), .B(n35436), .X(\shifter_0/n7329 ) );
  nor_x1_sg U48300 ( .A(n32989), .B(n35429), .X(\shifter_0/n7325 ) );
  nor_x1_sg U48301 ( .A(n32990), .B(n35430), .X(\shifter_0/n7321 ) );
  nor_x1_sg U48302 ( .A(n32991), .B(n35431), .X(\shifter_0/n7317 ) );
  nor_x1_sg U48303 ( .A(n32990), .B(n35432), .X(\shifter_0/n7313 ) );
  nor_x1_sg U48304 ( .A(n32991), .B(n35425), .X(\shifter_0/n7309 ) );
  nor_x1_sg U48305 ( .A(n35408), .B(n35426), .X(\shifter_0/n7305 ) );
  nor_x1_sg U48306 ( .A(n32990), .B(n35427), .X(\shifter_0/n7301 ) );
  nor_x1_sg U48307 ( .A(n32989), .B(n35428), .X(\shifter_0/n7297 ) );
  nor_x1_sg U48308 ( .A(n32991), .B(n35421), .X(\shifter_0/n7293 ) );
  nor_x1_sg U48309 ( .A(n32989), .B(n35422), .X(\shifter_0/n7289 ) );
  nor_x1_sg U48310 ( .A(n32988), .B(n35423), .X(\shifter_0/n7285 ) );
  nor_x1_sg U48311 ( .A(n32990), .B(n35424), .X(\shifter_0/n7281 ) );
  nor_x1_sg U48312 ( .A(n30012), .B(n35420), .X(\shifter_0/n7277 ) );
  nor_x1_sg U48313 ( .A(n33031), .B(n35481), .X(\shifter_0/n6873 ) );
  nor_x1_sg U48314 ( .A(n29996), .B(n13497), .X(\shifter_0/n6869 ) );
  nor_x1_sg U48315 ( .A(n33028), .B(n13503), .X(\shifter_0/n6865 ) );
  nor_x1_sg U48316 ( .A(n33030), .B(n35558), .X(\shifter_0/n6861 ) );
  nor_x1_sg U48317 ( .A(n33029), .B(n13514), .X(\shifter_0/n6857 ) );
  nor_x1_sg U48318 ( .A(n33031), .B(n35480), .X(\shifter_0/n6853 ) );
  nor_x1_sg U48319 ( .A(n33029), .B(n35479), .X(\shifter_0/n6849 ) );
  nor_x1_sg U48320 ( .A(n33028), .B(n35478), .X(\shifter_0/n6845 ) );
  nor_x1_sg U48321 ( .A(n33029), .B(n35486), .X(\shifter_0/n6841 ) );
  nor_x1_sg U48322 ( .A(n33030), .B(n13543), .X(\shifter_0/n6837 ) );
  nor_x1_sg U48323 ( .A(n33029), .B(n35477), .X(\shifter_0/n6833 ) );
  nor_x1_sg U48324 ( .A(n29996), .B(n35476), .X(\shifter_0/n6829 ) );
  nor_x1_sg U48325 ( .A(n33030), .B(n35475), .X(\shifter_0/n6825 ) );
  nor_x1_sg U48326 ( .A(n33028), .B(n35474), .X(\shifter_0/n6821 ) );
  nor_x1_sg U48327 ( .A(n35242), .B(n13573), .X(\shifter_0/n6817 ) );
  nor_x1_sg U48328 ( .A(n33028), .B(n13579), .X(\shifter_0/n6813 ) );
  nor_x1_sg U48329 ( .A(n35242), .B(n13585), .X(\shifter_0/n6809 ) );
  nor_x1_sg U48330 ( .A(n33031), .B(n13591), .X(\shifter_0/n6805 ) );
  nor_x1_sg U48331 ( .A(n33031), .B(n13596), .X(\shifter_0/n6801 ) );
  nor_x1_sg U48332 ( .A(n33030), .B(n13601), .X(\shifter_0/n6797 ) );
  nor_x1_sg U48333 ( .A(n31461), .B(n41420), .X(\shifter_0/n8390 ) );
  nor_x1_sg U48334 ( .A(n34127), .B(n41421), .X(\shifter_0/n8386 ) );
  nor_x1_sg U48335 ( .A(n34124), .B(n41422), .X(\shifter_0/n8382 ) );
  nor_x1_sg U48336 ( .A(n31461), .B(n41423), .X(\shifter_0/n8378 ) );
  nor_x1_sg U48337 ( .A(n31851), .B(n41424), .X(\shifter_0/n8374 ) );
  nor_x1_sg U48338 ( .A(n31462), .B(n41425), .X(\shifter_0/n8370 ) );
  nor_x1_sg U48339 ( .A(n30058), .B(n41426), .X(\shifter_0/n8366 ) );
  nor_x1_sg U48340 ( .A(n34124), .B(n41427), .X(\shifter_0/n8362 ) );
  nor_x1_sg U48341 ( .A(n34127), .B(n41428), .X(\shifter_0/n8358 ) );
  nor_x1_sg U48342 ( .A(n34126), .B(n41429), .X(\shifter_0/n8354 ) );
  nor_x1_sg U48343 ( .A(n31462), .B(n41430), .X(\shifter_0/n8350 ) );
  nor_x1_sg U48344 ( .A(n31462), .B(n41431), .X(\shifter_0/n8346 ) );
  nor_x1_sg U48345 ( .A(n34125), .B(n41432), .X(\shifter_0/n8342 ) );
  nor_x1_sg U48346 ( .A(n31850), .B(n41433), .X(\shifter_0/n8338 ) );
  nor_x1_sg U48347 ( .A(n34126), .B(n41434), .X(\shifter_0/n8334 ) );
  nor_x1_sg U48348 ( .A(n30057), .B(n41435), .X(\shifter_0/n8330 ) );
  nor_x1_sg U48349 ( .A(n30057), .B(n41436), .X(\shifter_0/n8326 ) );
  nor_x1_sg U48350 ( .A(n34127), .B(n41437), .X(\shifter_0/n8322 ) );
  nor_x1_sg U48351 ( .A(n31850), .B(n41438), .X(\shifter_0/n8318 ) );
  nor_x1_sg U48352 ( .A(n31467), .B(n41440), .X(\shifter_0/n8310 ) );
  nor_x1_sg U48353 ( .A(n34119), .B(n41441), .X(\shifter_0/n8306 ) );
  nor_x1_sg U48354 ( .A(n31468), .B(n41442), .X(\shifter_0/n8302 ) );
  nor_x1_sg U48355 ( .A(n31468), .B(n41443), .X(\shifter_0/n8298 ) );
  nor_x1_sg U48356 ( .A(n30052), .B(n41444), .X(\shifter_0/n8294 ) );
  nor_x1_sg U48357 ( .A(n31467), .B(n41445), .X(\shifter_0/n8290 ) );
  nor_x1_sg U48358 ( .A(n34116), .B(n41446), .X(\shifter_0/n8286 ) );
  nor_x1_sg U48359 ( .A(n34118), .B(n41447), .X(\shifter_0/n8282 ) );
  nor_x1_sg U48360 ( .A(n31855), .B(n41448), .X(\shifter_0/n8278 ) );
  nor_x1_sg U48361 ( .A(n34117), .B(n41449), .X(\shifter_0/n8274 ) );
  nor_x1_sg U48362 ( .A(n31854), .B(n41450), .X(\shifter_0/n8270 ) );
  nor_x1_sg U48363 ( .A(n34116), .B(n41451), .X(\shifter_0/n8266 ) );
  nor_x1_sg U48364 ( .A(n31854), .B(n41452), .X(\shifter_0/n8262 ) );
  nor_x1_sg U48365 ( .A(n30052), .B(n41453), .X(\shifter_0/n8258 ) );
  nor_x1_sg U48366 ( .A(n34117), .B(n41454), .X(\shifter_0/n8254 ) );
  nor_x1_sg U48367 ( .A(n30052), .B(n41455), .X(\shifter_0/n8250 ) );
  nor_x1_sg U48368 ( .A(n30051), .B(n41456), .X(\shifter_0/n8246 ) );
  nor_x1_sg U48369 ( .A(n31855), .B(n41457), .X(\shifter_0/n8242 ) );
  nor_x1_sg U48370 ( .A(n34118), .B(n41458), .X(\shifter_0/n8238 ) );
  nor_x1_sg U48371 ( .A(n34112), .B(n41460), .X(\shifter_0/n8230 ) );
  nor_x1_sg U48372 ( .A(n31856), .B(n41461), .X(\shifter_0/n8226 ) );
  nor_x1_sg U48373 ( .A(n31471), .B(n41462), .X(\shifter_0/n8222 ) );
  nor_x1_sg U48374 ( .A(n31471), .B(n41463), .X(\shifter_0/n8218 ) );
  nor_x1_sg U48375 ( .A(n31470), .B(n41464), .X(\shifter_0/n8214 ) );
  nor_x1_sg U48376 ( .A(n31470), .B(n41465), .X(\shifter_0/n8210 ) );
  nor_x1_sg U48377 ( .A(n30049), .B(n41466), .X(\shifter_0/n8206 ) );
  nor_x1_sg U48378 ( .A(n34113), .B(n41467), .X(\shifter_0/n8202 ) );
  nor_x1_sg U48379 ( .A(n30048), .B(n41468), .X(\shifter_0/n8198 ) );
  nor_x1_sg U48380 ( .A(n30048), .B(n41469), .X(\shifter_0/n8194 ) );
  nor_x1_sg U48381 ( .A(n34115), .B(n41470), .X(\shifter_0/n8190 ) );
  nor_x1_sg U48382 ( .A(n34113), .B(n41471), .X(\shifter_0/n8186 ) );
  nor_x1_sg U48383 ( .A(n34114), .B(n41472), .X(\shifter_0/n8182 ) );
  nor_x1_sg U48384 ( .A(n31857), .B(n41473), .X(\shifter_0/n8178 ) );
  nor_x1_sg U48385 ( .A(n34114), .B(n41474), .X(\shifter_0/n8174 ) );
  nor_x1_sg U48386 ( .A(n31856), .B(n41475), .X(\shifter_0/n8170 ) );
  nor_x1_sg U48387 ( .A(n30048), .B(n41476), .X(\shifter_0/n8166 ) );
  nor_x1_sg U48388 ( .A(n34115), .B(n41477), .X(\shifter_0/n8162 ) );
  nor_x1_sg U48389 ( .A(n31471), .B(n41478), .X(\shifter_0/n8158 ) );
  nor_x1_sg U48390 ( .A(n34123), .B(n41480), .X(\shifter_0/n8150 ) );
  nor_x1_sg U48391 ( .A(n34122), .B(n41481), .X(\shifter_0/n8146 ) );
  nor_x1_sg U48392 ( .A(n34121), .B(n41482), .X(\shifter_0/n8142 ) );
  nor_x1_sg U48393 ( .A(n31464), .B(n41483), .X(\shifter_0/n8138 ) );
  nor_x1_sg U48394 ( .A(n31464), .B(n41484), .X(\shifter_0/n8134 ) );
  nor_x1_sg U48395 ( .A(n31465), .B(n41485), .X(\shifter_0/n8130 ) );
  nor_x1_sg U48396 ( .A(n34120), .B(n41486), .X(\shifter_0/n8126 ) );
  nor_x1_sg U48397 ( .A(n31464), .B(n41487), .X(\shifter_0/n8122 ) );
  nor_x1_sg U48398 ( .A(n31852), .B(n41488), .X(\shifter_0/n8118 ) );
  nor_x1_sg U48399 ( .A(n31464), .B(n41489), .X(\shifter_0/n8114 ) );
  nor_x1_sg U48400 ( .A(n31853), .B(n41490), .X(\shifter_0/n8110 ) );
  nor_x1_sg U48401 ( .A(n34122), .B(n41491), .X(\shifter_0/n8106 ) );
  nor_x1_sg U48402 ( .A(n34120), .B(n41492), .X(\shifter_0/n8102 ) );
  nor_x1_sg U48403 ( .A(n34121), .B(n41493), .X(\shifter_0/n8098 ) );
  nor_x1_sg U48404 ( .A(n31852), .B(n41494), .X(\shifter_0/n8094 ) );
  nor_x1_sg U48405 ( .A(n34123), .B(n41495), .X(\shifter_0/n8090 ) );
  nor_x1_sg U48406 ( .A(n30054), .B(n41496), .X(\shifter_0/n8086 ) );
  nor_x1_sg U48407 ( .A(n31465), .B(n41497), .X(\shifter_0/n8082 ) );
  nor_x1_sg U48408 ( .A(n30054), .B(n41498), .X(\shifter_0/n8078 ) );
  nor_x1_sg U48409 ( .A(n33965), .B(n15155), .X(\filter_0/n6296 ) );
  nor_x1_sg U48410 ( .A(n33966), .B(n15165), .X(\filter_0/n6280 ) );
  nor_x1_sg U48411 ( .A(n15202), .B(n30017), .X(\filter_0/n4989 ) );
  nor_x1_sg U48412 ( .A(n42399), .B(n15203), .X(n15202) );
  inv_x1_sg U48413 ( .A(n15205), .X(n42399) );
  nor_x1_sg U48414 ( .A(n35305), .B(n15204), .X(n15203) );
  nor_x1_sg U48415 ( .A(n41233), .B(n31315), .X(\shifter_0/n8518 ) );
  nor_x1_sg U48416 ( .A(n41213), .B(n34375), .X(\shifter_0/n8598 ) );
  nor_x1_sg U48417 ( .A(n41253), .B(n31368), .X(\shifter_0/n8438 ) );
  nor_x1_sg U48418 ( .A(n41224), .B(n31314), .X(\shifter_0/n8554 ) );
  nor_x1_sg U48419 ( .A(n41225), .B(n31314), .X(\shifter_0/n8550 ) );
  nor_x1_sg U48420 ( .A(n41226), .B(n34370), .X(\shifter_0/n8546 ) );
  nor_x1_sg U48421 ( .A(n41227), .B(n34371), .X(\shifter_0/n8542 ) );
  nor_x1_sg U48422 ( .A(n41228), .B(n30358), .X(\shifter_0/n8538 ) );
  nor_x1_sg U48423 ( .A(n41229), .B(n31759), .X(\shifter_0/n8534 ) );
  nor_x1_sg U48424 ( .A(n41230), .B(n31760), .X(\shifter_0/n8530 ) );
  nor_x1_sg U48425 ( .A(n41231), .B(n11641), .X(\shifter_0/n8526 ) );
  nor_x1_sg U48426 ( .A(n41232), .B(n30358), .X(\shifter_0/n8522 ) );
  nor_x1_sg U48427 ( .A(n41234), .B(n34369), .X(\shifter_0/n8514 ) );
  nor_x1_sg U48428 ( .A(n41235), .B(n29708), .X(\shifter_0/n8510 ) );
  nor_x1_sg U48429 ( .A(n41236), .B(n31315), .X(\shifter_0/n8506 ) );
  nor_x1_sg U48430 ( .A(n41237), .B(n34370), .X(\shifter_0/n8502 ) );
  nor_x1_sg U48431 ( .A(n41238), .B(n30109), .X(\shifter_0/n8498 ) );
  nor_x1_sg U48432 ( .A(n41239), .B(n34370), .X(\shifter_0/n8494 ) );
  nor_x1_sg U48433 ( .A(n41240), .B(n31759), .X(\shifter_0/n8490 ) );
  nor_x1_sg U48434 ( .A(n41241), .B(n31759), .X(\shifter_0/n8486 ) );
  nor_x1_sg U48435 ( .A(n41242), .B(n31760), .X(\shifter_0/n8482 ) );
  nor_x1_sg U48436 ( .A(n41243), .B(n31315), .X(\shifter_0/n8478 ) );
  nor_x1_sg U48437 ( .A(n41204), .B(n34374), .X(\shifter_0/n8634 ) );
  nor_x1_sg U48438 ( .A(n41205), .B(n30110), .X(\shifter_0/n8630 ) );
  nor_x1_sg U48439 ( .A(n41206), .B(n34377), .X(\shifter_0/n8626 ) );
  nor_x1_sg U48440 ( .A(n41207), .B(n30360), .X(\shifter_0/n8622 ) );
  nor_x1_sg U48441 ( .A(n41208), .B(n34377), .X(\shifter_0/n8618 ) );
  nor_x1_sg U48442 ( .A(n41209), .B(n30360), .X(\shifter_0/n8614 ) );
  nor_x1_sg U48443 ( .A(n41210), .B(n34374), .X(\shifter_0/n8610 ) );
  nor_x1_sg U48444 ( .A(n41211), .B(n31758), .X(\shifter_0/n8606 ) );
  nor_x1_sg U48445 ( .A(n41212), .B(n35458), .X(\shifter_0/n8602 ) );
  nor_x1_sg U48446 ( .A(n41214), .B(n31312), .X(\shifter_0/n8594 ) );
  nor_x1_sg U48447 ( .A(n41215), .B(n34376), .X(\shifter_0/n8590 ) );
  nor_x1_sg U48448 ( .A(n41216), .B(n31311), .X(\shifter_0/n8586 ) );
  nor_x1_sg U48449 ( .A(n41217), .B(n31757), .X(\shifter_0/n8582 ) );
  nor_x1_sg U48450 ( .A(n41218), .B(n31757), .X(\shifter_0/n8578 ) );
  nor_x1_sg U48451 ( .A(n41219), .B(n31312), .X(\shifter_0/n8574 ) );
  nor_x1_sg U48452 ( .A(n41220), .B(n30360), .X(\shifter_0/n8570 ) );
  nor_x1_sg U48453 ( .A(n41221), .B(n31311), .X(\shifter_0/n8566 ) );
  nor_x1_sg U48454 ( .A(n41222), .B(n31758), .X(\shifter_0/n8562 ) );
  nor_x1_sg U48455 ( .A(n41223), .B(n31757), .X(\shifter_0/n8558 ) );
  nor_x1_sg U48456 ( .A(n41244), .B(n11667), .X(\shifter_0/n8474 ) );
  nor_x1_sg U48457 ( .A(n41245), .B(n30322), .X(\shifter_0/n8470 ) );
  nor_x1_sg U48458 ( .A(n41246), .B(n29726), .X(\shifter_0/n8466 ) );
  nor_x1_sg U48459 ( .A(n41247), .B(n34282), .X(\shifter_0/n8462 ) );
  nor_x1_sg U48460 ( .A(n41248), .B(n31796), .X(\shifter_0/n8458 ) );
  nor_x1_sg U48461 ( .A(n41249), .B(n30322), .X(\shifter_0/n8454 ) );
  nor_x1_sg U48462 ( .A(n41250), .B(n31795), .X(\shifter_0/n8450 ) );
  nor_x1_sg U48463 ( .A(n41251), .B(n31368), .X(\shifter_0/n8446 ) );
  nor_x1_sg U48464 ( .A(n41252), .B(n31796), .X(\shifter_0/n8442 ) );
  nor_x1_sg U48465 ( .A(n41254), .B(n31796), .X(\shifter_0/n8434 ) );
  nor_x1_sg U48466 ( .A(n41255), .B(n31796), .X(\shifter_0/n8430 ) );
  nor_x1_sg U48467 ( .A(n41256), .B(n34282), .X(\shifter_0/n8426 ) );
  nor_x1_sg U48468 ( .A(n41257), .B(n34280), .X(\shifter_0/n8422 ) );
  nor_x1_sg U48469 ( .A(n41258), .B(n31795), .X(\shifter_0/n8418 ) );
  nor_x1_sg U48470 ( .A(n41259), .B(n30091), .X(\shifter_0/n8414 ) );
  nor_x1_sg U48471 ( .A(n41260), .B(n30091), .X(\shifter_0/n8410 ) );
  nor_x1_sg U48472 ( .A(n41261), .B(n31795), .X(\shifter_0/n8406 ) );
  nor_x1_sg U48473 ( .A(n41262), .B(n34281), .X(\shifter_0/n8402 ) );
  nor_x1_sg U48474 ( .A(n41263), .B(n34281), .X(\shifter_0/n8398 ) );
  nor_x1_sg U48475 ( .A(n42393), .B(n31651), .X(\filter_0/n6297 ) );
  inv_x1_sg U48476 ( .A(n15155), .X(n42393) );
  nor_x1_sg U48477 ( .A(n42391), .B(n33964), .X(\filter_0/n6281 ) );
  inv_x1_sg U48478 ( .A(n15165), .X(n42391) );
  nor_x1_sg U48479 ( .A(n41143), .B(n30108), .X(\shifter_0/n8874 ) );
  nor_x1_sg U48480 ( .A(n41144), .B(n31317), .X(\shifter_0/n8870 ) );
  nor_x1_sg U48481 ( .A(n41145), .B(n34367), .X(\shifter_0/n8866 ) );
  nor_x1_sg U48482 ( .A(n41146), .B(n30356), .X(\shifter_0/n8862 ) );
  nor_x1_sg U48483 ( .A(n41147), .B(n34365), .X(\shifter_0/n8858 ) );
  nor_x1_sg U48484 ( .A(n41148), .B(n31761), .X(\shifter_0/n8854 ) );
  nor_x1_sg U48485 ( .A(n41149), .B(n34367), .X(\shifter_0/n8850 ) );
  nor_x1_sg U48486 ( .A(n41150), .B(n31761), .X(\shifter_0/n8846 ) );
  nor_x1_sg U48487 ( .A(n41151), .B(n30356), .X(\shifter_0/n8842 ) );
  nor_x1_sg U48488 ( .A(n41152), .B(n34365), .X(\shifter_0/n8838 ) );
  nor_x1_sg U48489 ( .A(n41153), .B(n34364), .X(\shifter_0/n8834 ) );
  nor_x1_sg U48490 ( .A(n41154), .B(n34366), .X(\shifter_0/n8830 ) );
  nor_x1_sg U48491 ( .A(n41155), .B(n34366), .X(\shifter_0/n8826 ) );
  nor_x1_sg U48492 ( .A(n41156), .B(n31762), .X(\shifter_0/n8822 ) );
  nor_x1_sg U48493 ( .A(n41157), .B(n31318), .X(\shifter_0/n8818 ) );
  nor_x1_sg U48494 ( .A(n41158), .B(n31317), .X(\shifter_0/n8814 ) );
  nor_x1_sg U48495 ( .A(n41159), .B(n34365), .X(\shifter_0/n8810 ) );
  nor_x1_sg U48496 ( .A(n41160), .B(n34365), .X(\shifter_0/n8806 ) );
  nor_x1_sg U48497 ( .A(n41161), .B(n31761), .X(\shifter_0/n8802 ) );
  nor_x1_sg U48498 ( .A(n41162), .B(n31762), .X(\shifter_0/n8798 ) );
  nor_x1_sg U48499 ( .A(n41163), .B(n34354), .X(\shifter_0/n8794 ) );
  nor_x1_sg U48500 ( .A(n41164), .B(n29711), .X(\shifter_0/n8790 ) );
  nor_x1_sg U48501 ( .A(n41165), .B(n30352), .X(\shifter_0/n8786 ) );
  nor_x1_sg U48502 ( .A(n41166), .B(n34356), .X(\shifter_0/n8782 ) );
  nor_x1_sg U48503 ( .A(n41167), .B(n29711), .X(\shifter_0/n8778 ) );
  nor_x1_sg U48504 ( .A(n41168), .B(n30352), .X(\shifter_0/n8774 ) );
  nor_x1_sg U48505 ( .A(n41169), .B(n31324), .X(\shifter_0/n8770 ) );
  nor_x1_sg U48506 ( .A(n41170), .B(n31766), .X(\shifter_0/n8766 ) );
  nor_x1_sg U48507 ( .A(n41171), .B(n30106), .X(\shifter_0/n8762 ) );
  nor_x1_sg U48508 ( .A(n41172), .B(n31765), .X(\shifter_0/n8758 ) );
  nor_x1_sg U48509 ( .A(n41173), .B(n31324), .X(\shifter_0/n8754 ) );
  nor_x1_sg U48510 ( .A(n41174), .B(n34355), .X(\shifter_0/n8750 ) );
  nor_x1_sg U48511 ( .A(n41175), .B(n30106), .X(\shifter_0/n8746 ) );
  nor_x1_sg U48512 ( .A(n41176), .B(n34355), .X(\shifter_0/n8742 ) );
  nor_x1_sg U48513 ( .A(n41177), .B(n34357), .X(\shifter_0/n8738 ) );
  nor_x1_sg U48514 ( .A(n41178), .B(n34354), .X(\shifter_0/n8734 ) );
  nor_x1_sg U48515 ( .A(n41179), .B(n34357), .X(\shifter_0/n8730 ) );
  nor_x1_sg U48516 ( .A(n41180), .B(n34355), .X(\shifter_0/n8726 ) );
  nor_x1_sg U48517 ( .A(n41181), .B(n31323), .X(\shifter_0/n8722 ) );
  nor_x1_sg U48518 ( .A(n41182), .B(n34356), .X(\shifter_0/n8718 ) );
  nor_x1_sg U48519 ( .A(n41184), .B(n34359), .X(\shifter_0/n8714 ) );
  nor_x1_sg U48520 ( .A(n41185), .B(n34362), .X(\shifter_0/n8710 ) );
  nor_x1_sg U48521 ( .A(n41186), .B(n29710), .X(\shifter_0/n8706 ) );
  nor_x1_sg U48522 ( .A(n41187), .B(n34361), .X(\shifter_0/n8702 ) );
  nor_x1_sg U48523 ( .A(n41188), .B(n34361), .X(\shifter_0/n8698 ) );
  nor_x1_sg U48524 ( .A(n41189), .B(n31764), .X(\shifter_0/n8694 ) );
  nor_x1_sg U48525 ( .A(n41190), .B(n34359), .X(\shifter_0/n8690 ) );
  nor_x1_sg U48526 ( .A(n41191), .B(n30107), .X(\shifter_0/n8686 ) );
  nor_x1_sg U48527 ( .A(n41192), .B(n30107), .X(\shifter_0/n8682 ) );
  nor_x1_sg U48528 ( .A(n41193), .B(n34362), .X(\shifter_0/n8678 ) );
  nor_x1_sg U48529 ( .A(n41194), .B(n29710), .X(\shifter_0/n8674 ) );
  nor_x1_sg U48530 ( .A(n41195), .B(n31764), .X(\shifter_0/n8670 ) );
  nor_x1_sg U48531 ( .A(n41196), .B(n31764), .X(\shifter_0/n8666 ) );
  nor_x1_sg U48532 ( .A(n41197), .B(n31320), .X(\shifter_0/n8662 ) );
  nor_x1_sg U48533 ( .A(n41198), .B(n30107), .X(\shifter_0/n8658 ) );
  nor_x1_sg U48534 ( .A(n41199), .B(n31321), .X(\shifter_0/n8654 ) );
  nor_x1_sg U48535 ( .A(n41200), .B(n31763), .X(\shifter_0/n8650 ) );
  nor_x1_sg U48536 ( .A(n41201), .B(n34360), .X(\shifter_0/n8646 ) );
  nor_x1_sg U48537 ( .A(n41202), .B(n31320), .X(\shifter_0/n8642 ) );
  nor_x1_sg U48538 ( .A(n41203), .B(n34359), .X(\shifter_0/n8638 ) );
  nor_x1_sg U48539 ( .A(n41419), .B(n31850), .X(\shifter_0/n8394 ) );
  nor_x1_sg U48540 ( .A(n41439), .B(n31468), .X(\shifter_0/n8314 ) );
  nor_x1_sg U48541 ( .A(n41459), .B(n34113), .X(\shifter_0/n8234 ) );
  nor_x1_sg U48542 ( .A(n41479), .B(n34123), .X(\shifter_0/n8154 ) );
  nand_x1_sg U48543 ( .A(n41135), .B(n33868), .X(n13119) );
  nand_x1_sg U48544 ( .A(n33871), .B(n41139), .X(n13118) );
  nand_x1_sg U48545 ( .A(n41136), .B(n33866), .X(n13130) );
  nand_x1_sg U48546 ( .A(n30944), .B(n41140), .X(n13129) );
  nand_x1_sg U48547 ( .A(n41137), .B(n33865), .X(n13207) );
  nand_x1_sg U48548 ( .A(n30943), .B(n41141), .X(n13206) );
  nand_x1_sg U48549 ( .A(n41138), .B(n33866), .X(n13212) );
  nand_x1_sg U48550 ( .A(n30943), .B(n41142), .X(n13211) );
  nand_x1_sg U48551 ( .A(n35638), .B(n13497), .X(n13496) );
  nand_x1_sg U48552 ( .A(n33721), .B(n13519), .X(n13518) );
  nand_x1_sg U48553 ( .A(n29997), .B(n13531), .X(n13530) );
  nand_x1_sg U48554 ( .A(n29997), .B(n13543), .X(n13542) );
  nand_x1_sg U48555 ( .A(n33720), .B(n13491), .X(n13489) );
  nand_x1_sg U48556 ( .A(n33720), .B(n13503), .X(n13502) );
  nand_x1_sg U48557 ( .A(n30997), .B(n13514), .X(n13513) );
  nand_x1_sg U48558 ( .A(n33722), .B(n13525), .X(n13524) );
  nand_x1_sg U48559 ( .A(n35638), .B(n13537), .X(n13536) );
  nand_x1_sg U48560 ( .A(n33721), .B(n13549), .X(n13548) );
  nand_x1_sg U48561 ( .A(n33722), .B(n13561), .X(n13560) );
  nand_x1_sg U48562 ( .A(n29997), .B(n13573), .X(n13572) );
  nand_x1_sg U48563 ( .A(n30997), .B(n13579), .X(n13578) );
  nand_x1_sg U48564 ( .A(n33722), .B(n13585), .X(n13584) );
  nand_x1_sg U48565 ( .A(n30997), .B(n13591), .X(n13590) );
  nand_x1_sg U48566 ( .A(n33721), .B(n13596), .X(n13595) );
  nand_x1_sg U48567 ( .A(n30013), .B(n35440), .X(n12848) );
  nand_x1_sg U48568 ( .A(n12842), .B(n35435), .X(n12872) );
  nand_x1_sg U48569 ( .A(n12842), .B(n35429), .X(n12884) );
  nand_x1_sg U48570 ( .A(n30987), .B(n35431), .X(n12896) );
  nand_x1_sg U48571 ( .A(n33718), .B(n12719), .X(n12718) );
  nand_x1_sg U48572 ( .A(n29995), .B(n35451), .X(n12742) );
  nand_x1_sg U48573 ( .A(n30998), .B(n12755), .X(n12754) );
  nand_x1_sg U48574 ( .A(n33718), .B(n35446), .X(n12766) );
  nand_x1_sg U48575 ( .A(n30987), .B(n35439), .X(n12841) );
  nand_x1_sg U48576 ( .A(n33796), .B(n35433), .X(n12854) );
  nand_x1_sg U48577 ( .A(n33797), .B(n35434), .X(n12866) );
  nand_x1_sg U48578 ( .A(n33796), .B(n35436), .X(n12878) );
  nand_x1_sg U48579 ( .A(n30987), .B(n35430), .X(n12890) );
  nand_x1_sg U48580 ( .A(n33798), .B(n35432), .X(n12902) );
  nand_x1_sg U48581 ( .A(n33798), .B(n35426), .X(n12914) );
  nand_x1_sg U48582 ( .A(n33797), .B(n35428), .X(n12926) );
  nand_x1_sg U48583 ( .A(n30013), .B(n35421), .X(n12932) );
  nand_x1_sg U48584 ( .A(n30013), .B(n35422), .X(n12938) );
  nand_x1_sg U48585 ( .A(n30987), .B(n35423), .X(n12944) );
  nand_x1_sg U48586 ( .A(n33797), .B(n35424), .X(n12950) );
  nand_x1_sg U48587 ( .A(n35620), .B(n13370), .X(n13369) );
  nand_x1_sg U48588 ( .A(n30992), .B(n13394), .X(n13393) );
  nand_x1_sg U48589 ( .A(n30005), .B(n13406), .X(n13405) );
  nand_x1_sg U48590 ( .A(n33741), .B(n13418), .X(n13417) );
  nand_x1_sg U48591 ( .A(n29995), .B(n35449), .X(n12710) );
  nand_x1_sg U48592 ( .A(n33717), .B(n35450), .X(n12724) );
  nand_x1_sg U48593 ( .A(n33717), .B(n12737), .X(n12736) );
  nand_x1_sg U48594 ( .A(n33717), .B(n35452), .X(n12748) );
  nand_x1_sg U48595 ( .A(n30998), .B(n35445), .X(n12760) );
  nand_x1_sg U48596 ( .A(n30998), .B(n35447), .X(n12772) );
  nand_x1_sg U48597 ( .A(n35622), .B(n12785), .X(n12784) );
  nand_x1_sg U48598 ( .A(n29995), .B(n12797), .X(n12796) );
  nand_x1_sg U48599 ( .A(n33716), .B(n35442), .X(n12802) );
  nand_x1_sg U48600 ( .A(n30998), .B(n35443), .X(n12808) );
  nand_x1_sg U48601 ( .A(n33716), .B(n35444), .X(n12814) );
  nand_x1_sg U48602 ( .A(n29995), .B(n35437), .X(n12820) );
  nand_x1_sg U48603 ( .A(n35620), .B(n13362), .X(n13360) );
  nand_x1_sg U48604 ( .A(n33741), .B(n13376), .X(n13375) );
  nand_x1_sg U48605 ( .A(n33743), .B(n13388), .X(n13387) );
  nand_x1_sg U48606 ( .A(n33742), .B(n13400), .X(n13399) );
  nand_x1_sg U48607 ( .A(n33743), .B(n13412), .X(n13411) );
  nand_x1_sg U48608 ( .A(n33742), .B(n13424), .X(n13423) );
  nand_x1_sg U48609 ( .A(n30992), .B(n13436), .X(n13435) );
  nand_x1_sg U48610 ( .A(n30005), .B(n13448), .X(n13447) );
  nand_x1_sg U48611 ( .A(n30992), .B(n13454), .X(n13453) );
  nand_x1_sg U48612 ( .A(n30992), .B(n13460), .X(n13459) );
  nand_x1_sg U48613 ( .A(n30005), .B(n13466), .X(n13465) );
  nand_x1_sg U48614 ( .A(n30005), .B(n13472), .X(n13471) );
  nand_x1_sg U48615 ( .A(n31001), .B(n13822), .X(n13821) );
  nand_x1_sg U48616 ( .A(n35635), .B(n13884), .X(n13883) );
  nand_x1_sg U48617 ( .A(n33633), .B(n13946), .X(n13945) );
  nand_x1_sg U48618 ( .A(n33631), .B(n14008), .X(n14007) );
  nand_x1_sg U48619 ( .A(n35635), .B(n14070), .X(n14069) );
  nand_x1_sg U48620 ( .A(n29991), .B(n13784), .X(n13782) );
  nand_x1_sg U48621 ( .A(n33631), .B(n13853), .X(n13852) );
  nand_x1_sg U48622 ( .A(n31001), .B(n13915), .X(n13914) );
  nand_x1_sg U48623 ( .A(n29991), .B(n13977), .X(n13976) );
  nand_x1_sg U48624 ( .A(n33633), .B(n14039), .X(n14038) );
  nand_x1_sg U48625 ( .A(n31001), .B(n14101), .X(n14100) );
  nand_x1_sg U48626 ( .A(n33632), .B(n14163), .X(n14162) );
  nand_x1_sg U48627 ( .A(n29991), .B(n14225), .X(n14224) );
  nand_x1_sg U48628 ( .A(n33632), .B(n14256), .X(n14255) );
  nand_x1_sg U48629 ( .A(n33633), .B(n14287), .X(n14286) );
  nand_x1_sg U48630 ( .A(n29991), .B(n14318), .X(n14317) );
  nand_x1_sg U48631 ( .A(n33632), .B(n14349), .X(n14348) );
  nand_x1_sg U48632 ( .A(n14411), .B(n14569), .X(n14568) );
  nand_x1_sg U48633 ( .A(n31002), .B(n14662), .X(n14661) );
  nand_x1_sg U48634 ( .A(n29989), .B(n14724), .X(n14723) );
  nand_x1_sg U48635 ( .A(n31002), .B(n14786), .X(n14785) );
  nand_x1_sg U48636 ( .A(n33524), .B(n14848), .X(n14847) );
  nand_x1_sg U48637 ( .A(n14411), .B(n14910), .X(n14909) );
  nand_x1_sg U48638 ( .A(n31002), .B(n14972), .X(n14971) );
  nand_x1_sg U48639 ( .A(n31002), .B(n14443), .X(n14442) );
  nand_x1_sg U48640 ( .A(n29989), .B(n14538), .X(n14537) );
  nand_x1_sg U48641 ( .A(n33525), .B(n14631), .X(n14630) );
  nand_x1_sg U48642 ( .A(n33523), .B(n14412), .X(n14410) );
  nand_x1_sg U48643 ( .A(n33525), .B(n35095), .X(n14506) );
  nand_x1_sg U48644 ( .A(n33524), .B(n14600), .X(n14599) );
  nand_x1_sg U48645 ( .A(n33524), .B(n14693), .X(n14692) );
  nand_x1_sg U48646 ( .A(n29989), .B(n14755), .X(n14754) );
  nand_x1_sg U48647 ( .A(n33523), .B(n14817), .X(n14816) );
  nand_x1_sg U48648 ( .A(n29989), .B(n14879), .X(n14878) );
  nand_x1_sg U48649 ( .A(n33524), .B(n14941), .X(n14940) );
  nand_x1_sg U48650 ( .A(n33525), .B(n15003), .X(n15002) );
  nor_x1_sg U48651 ( .A(n22209), .B(n35251), .X(n19607) );
  nand_x1_sg U48652 ( .A(n31978), .B(n35551), .X(n22209) );
  nand_x1_sg U48653 ( .A(n22220), .B(n30541), .X(n26194) );
  nor_x1_sg U48654 ( .A(n35605), .B(n21303), .X(n20906) );
  nand_x1_sg U48655 ( .A(n31883), .B(n30540), .X(n20949) );
  nand_x1_sg U48656 ( .A(n31701), .B(n30540), .X(n20941) );
  nand_x1_sg U48657 ( .A(n20906), .B(n20943), .X(n20942) );
  nand_x1_sg U48658 ( .A(n20944), .B(n20945), .X(n20943) );
  nor_x1_sg U48659 ( .A(n21303), .B(n42408), .X(n21327) );
  inv_x1_sg U48660 ( .A(n21370), .X(n42408) );
  nand_x4_sg U48661 ( .A(n21732), .B(n21733), .X(n21727) );
  nand_x1_sg U48662 ( .A(n32005), .B(n21326), .X(n21325) );
  nand_x1_sg U48663 ( .A(n21329), .B(n21330), .X(n21328) );
  nand_x1_sg U48664 ( .A(n31698), .B(n21326), .X(n21338) );
  nand_x1_sg U48665 ( .A(n21327), .B(n21339), .X(n21337) );
  nand_x1_sg U48666 ( .A(n21340), .B(n21341), .X(n21339) );
  nor_x1_sg U48667 ( .A(n31886), .B(n35265), .X(n26590) );
  nand_x1_sg U48668 ( .A(n29489), .B(n31880), .X(n29488) );
  nor_x1_sg U48669 ( .A(n34062), .B(n35272), .X(n29489) );
  nor_x1_sg U48670 ( .A(n15306), .B(n42380), .X(n15305) );
  nand_x4_sg U48671 ( .A(n15310), .B(n42386), .X(n15306) );
  nor_x1_sg U48672 ( .A(n15308), .B(n15309), .X(n15307) );
  nand_x1_sg U48673 ( .A(\filter_0/N16 ), .B(n15320), .X(n15285) );
  nor_x1_sg U48674 ( .A(n15339), .B(n42382), .X(n15338) );
  nor_x1_sg U48675 ( .A(n15291), .B(n42385), .X(n15290) );
  nand_x4_sg U48676 ( .A(n15295), .B(n42369), .X(n15291) );
  nor_x1_sg U48677 ( .A(n15293), .B(n15294), .X(n15292) );
  nor_x1_sg U48678 ( .A(n15324), .B(n42387), .X(n15323) );
  nor_x1_sg U48679 ( .A(n15318), .B(n15319), .X(n15315) );
  nor_x1_sg U48680 ( .A(n35306), .B(n15317), .X(n15316) );
  nand_x1_sg U48681 ( .A(n28967), .B(n35270), .X(n28966) );
  nand_x1_sg U48682 ( .A(n29666), .B(n35270), .X(n29665) );
  nand_x1_sg U48683 ( .A(n28878), .B(n35270), .X(n28877) );
  nand_x1_sg U48684 ( .A(n28834), .B(n34061), .X(n28833) );
  nor_x1_sg U48685 ( .A(n20922), .B(n20923), .X(n20907) );
  nor_x1_sg U48686 ( .A(n20929), .B(n42538), .X(n20922) );
  nand_x1_sg U48687 ( .A(n20924), .B(n32390), .X(n20923) );
  nand_x1_sg U48688 ( .A(n32172), .B(n21561), .X(n21372) );
  nand_x1_sg U48689 ( .A(n21656), .B(n32936), .X(n21562) );
  nand_x1_sg U48690 ( .A(n32004), .B(n21336), .X(n21329) );
  nand_x1_sg U48691 ( .A(n31882), .B(n20940), .X(n20952) );
  nand_x1_sg U48692 ( .A(n31702), .B(n20940), .X(n20944) );
  nand_x1_sg U48693 ( .A(n31699), .B(n21336), .X(n21340) );
  nand_x1_sg U48694 ( .A(n21374), .B(n34563), .X(n21373) );
  nand_x1_sg U48695 ( .A(n21469), .B(n32940), .X(n21375) );
  nor_x1_sg U48696 ( .A(n26584), .B(n26587), .X(n26579) );
  nor_x1_sg U48697 ( .A(n34562), .B(n20909), .X(n20908) );
  nand_x1_sg U48698 ( .A(n20912), .B(n32939), .X(n20911) );
  nor_x1_sg U48699 ( .A(n20915), .B(n19584), .X(n20984) );
  nor_x1_sg U48700 ( .A(n21359), .B(n19584), .X(n21358) );
  nand_x1_sg U48701 ( .A(n31884), .B(n35101), .X(n20956) );
  nor_x1_sg U48702 ( .A(n19583), .B(n20957), .X(n20955) );
  nand_x1_sg U48703 ( .A(n20938), .B(n20939), .X(n20937) );
  nand_x1_sg U48704 ( .A(n42547), .B(n19586), .X(n20939) );
  nand_x1_sg U48705 ( .A(n42533), .B(n19587), .X(n21350) );
  nand_x1_sg U48706 ( .A(n32006), .B(n35100), .X(n21334) );
  nor_x1_sg U48707 ( .A(n19581), .B(n21335), .X(n21333) );
  nand_x1_sg U48708 ( .A(n19579), .B(n35279), .X(n20947) );
  nand_x1_sg U48709 ( .A(n31701), .B(n35101), .X(n20948) );
  nand_x1_sg U48710 ( .A(n19580), .B(n35280), .X(n21343) );
  nand_x1_sg U48711 ( .A(n31698), .B(n35100), .X(n21344) );
  nand_x1_sg U48712 ( .A(n22215), .B(n35455), .X(n23629) );
  nor_x1_sg U48713 ( .A(n22214), .B(n22216), .X(n5981) );
  nor_x1_sg U48714 ( .A(n22217), .B(n34503), .X(n22216) );
  nor_x1_sg U48715 ( .A(n35455), .B(n42414), .X(n22217) );
  nand_x1_sg U48716 ( .A(n20972), .B(n30135), .X(n20969) );
  nand_x1_sg U48717 ( .A(n21002), .B(n34540), .X(n20999) );
  nand_x1_sg U48718 ( .A(n20982), .B(n34541), .X(n20979) );
  nand_x1_sg U48719 ( .A(n21388), .B(n32060), .X(n21385) );
  nand_x1_sg U48720 ( .A(n21575), .B(n32059), .X(n21572) );
  nand_x1_sg U48721 ( .A(n32424), .B(n29620), .X(n29487) );
  nand_x1_sg U48722 ( .A(n32427), .B(n29444), .X(n29317) );
  nand_x1_sg U48723 ( .A(n32424), .B(n28921), .X(n28788) );
  nand_x1_sg U48724 ( .A(n32425), .B(n28745), .X(n28618) );
  nor_x1_sg U48725 ( .A(n31885), .B(n29664), .X(n29663) );
  nor_x1_sg U48726 ( .A(n31886), .B(n28965), .X(n28964) );
  nand_x1_sg U48727 ( .A(n35251), .B(n19606), .X(n20893) );
  nor_x1_sg U48728 ( .A(n31120), .B(n35269), .X(n28790) );
  inv_x1_sg U48729 ( .A(n22215), .X(n42407) );
  nor_x1_sg U48730 ( .A(n31886), .B(n32885), .X(n28259) );
  nor_x1_sg U48731 ( .A(n35267), .B(n31668), .X(n19580) );
  nor_x1_sg U48732 ( .A(n35459), .B(n26350), .X(n26352) );
  nor_x1_sg U48733 ( .A(n35271), .B(n35303), .X(n19579) );
  nand_x4_sg U48734 ( .A(n21141), .B(n21142), .X(n21140) );
  nand_x4_sg U48735 ( .A(n21540), .B(n21541), .X(n21535) );
  nor_x1_sg U48736 ( .A(n35628), .B(n34388), .X(n26219) );
  nor_x1_sg U48737 ( .A(n35454), .B(n31201), .X(n35682) );
  nor_x1_sg U48738 ( .A(n29669), .B(n29670), .X(\filter_0/N1845 ) );
  nand_x1_sg U48739 ( .A(n31876), .B(n32000), .X(n29670) );
  inv_x1_sg U48740 ( .A(n11637), .X(n42533) );
  nand_x4_sg U48741 ( .A(n21241), .B(n21242), .X(n21240) );
  nand_x4_sg U48742 ( .A(n21597), .B(n21598), .X(n21592) );
  nand_x4_sg U48743 ( .A(n21719), .B(n21720), .X(n21718) );
  nand_x4_sg U48744 ( .A(n21701), .B(n21702), .X(n21700) );
  nand_x4_sg U48745 ( .A(n21219), .B(n21220), .X(n21218) );
  nand_x4_sg U48746 ( .A(n21062), .B(n21063), .X(n21061) );
  nand_x4_sg U48747 ( .A(n21201), .B(n21202), .X(n21200) );
  nand_x4_sg U48748 ( .A(n21650), .B(n21651), .X(n21649) );
  inv_x1_sg U48749 ( .A(n11612), .X(n42547) );
  nand_x4_sg U48750 ( .A(n21615), .B(n21616), .X(n21610) );
  nand_x4_sg U48751 ( .A(n21632), .B(n21633), .X(n21631) );
  nand_x4_sg U48752 ( .A(n21445), .B(n21446), .X(n21444) );
  nand_x4_sg U48753 ( .A(n21259), .B(n21260), .X(n21258) );
  nand_x4_sg U48754 ( .A(n21121), .B(n21122), .X(n21120) );
  nand_x4_sg U48755 ( .A(n21159), .B(n21160), .X(n21158) );
  nand_x4_sg U48756 ( .A(n21680), .B(n21681), .X(n21679) );
  nand_x4_sg U48757 ( .A(n21042), .B(n21043), .X(n21041) );
  nand_x4_sg U48758 ( .A(n21517), .B(n21518), .X(n21516) );
  nor_x1_sg U48759 ( .A(n31697), .B(n32005), .X(n12968) );
  nand_x4_sg U48760 ( .A(n21555), .B(n21556), .X(n21554) );
  nand_x4_sg U48761 ( .A(n21297), .B(n21298), .X(n21296) );
  nor_x1_sg U48762 ( .A(n31700), .B(n31883), .X(n12840) );
  nand_x4_sg U48763 ( .A(n21180), .B(n21181), .X(n21179) );
  nand_x4_sg U48764 ( .A(n21279), .B(n21280), .X(n21278) );
  nand_x4_sg U48765 ( .A(n21425), .B(n21426), .X(n21424) );
  nand_x4_sg U48766 ( .A(n21080), .B(n21081), .X(n21079) );
  nand_x4_sg U48767 ( .A(n21463), .B(n21464), .X(n21462) );
  nor_x1_sg U48768 ( .A(n35459), .B(n26206), .X(n26350) );
  nand_x4_sg U48769 ( .A(n21024), .B(n21025), .X(n21023) );
  nand_x4_sg U48770 ( .A(n21103), .B(n21104), .X(n21102) );
  nand_x1_sg U48771 ( .A(n42770), .B(n42771), .X(n21314) );
  nor_x1_sg U48772 ( .A(n35304), .B(n31699), .X(n19581) );
  nand_x4_sg U48773 ( .A(n21407), .B(n21408), .X(n21406) );
  nand_x4_sg U48774 ( .A(n21499), .B(n21500), .X(n21498) );
  nor_x1_sg U48775 ( .A(n31881), .B(n31702), .X(n19583) );
  nor_x1_sg U48776 ( .A(n26215), .B(n31201), .X(n26209) );
  nand_x1_sg U48777 ( .A(n26214), .B(n35454), .X(n26215) );
  inv_x1_sg U48778 ( .A(n26206), .X(n42528) );
  inv_x1_sg U48779 ( .A(n26214), .X(n42527) );
  nand_x1_sg U48780 ( .A(n42528), .B(n42530), .X(n26197) );
  nand_x1_sg U48781 ( .A(n26200), .B(n26206), .X(n26205) );
  nor_x1_sg U48782 ( .A(n31884), .B(n31701), .X(n13098) );
  nor_x1_sg U48783 ( .A(n31698), .B(n32006), .X(n13222) );
  nand_x1_sg U48784 ( .A(n28878), .B(n31661), .X(n15051) );
  nand_x1_sg U48785 ( .A(n28834), .B(n31662), .X(n15054) );
  nor_x1_sg U48786 ( .A(n31880), .B(n35272), .X(n15186) );
  nor_x1_sg U48787 ( .A(n35272), .B(n35305), .X(n15192) );
  nand_x1_sg U48788 ( .A(n30537), .B(n32004), .X(n12522) );
  nand_x1_sg U48789 ( .A(n30529), .B(n12524), .X(n12523) );
  nand_x1_sg U48790 ( .A(n12525), .B(n12526), .X(n12524) );
  nand_x1_sg U48791 ( .A(n31200), .B(n11609), .X(n13700) );
  nor_x1_sg U48792 ( .A(n12433), .B(n19586), .X(n12610) );
  nor_x1_sg U48793 ( .A(n12525), .B(n19587), .X(n12703) );
  nand_x1_sg U48794 ( .A(n15122), .B(n31876), .X(n15080) );
  nand_x1_sg U48795 ( .A(n15251), .B(n31876), .X(n15216) );
  nand_x1_sg U48796 ( .A(n13222), .B(n11639), .X(n13781) );
  nor_x1_sg U48797 ( .A(n12120), .B(n41604), .X(n12346) );
  inv_x1_sg U48798 ( .A(n19581), .X(n41604) );
  nand_x1_sg U48799 ( .A(n12433), .B(n12434), .X(n12432) );
  nand_x1_sg U48800 ( .A(n19585), .B(n31701), .X(n12434) );
  nand_x1_sg U48801 ( .A(n30522), .B(n35508), .X(n15049) );
  nand_x1_sg U48802 ( .A(n28965), .B(n35516), .X(n15055) );
  nand_x1_sg U48803 ( .A(n30520), .B(n35504), .X(n15182) );
  nand_x1_sg U48804 ( .A(n29664), .B(n35553), .X(n15190) );
  nand_x1_sg U48805 ( .A(n12116), .B(n31884), .X(n12117) );
  nand_x1_sg U48806 ( .A(n12116), .B(n32005), .X(n12344) );
  nand_x1_sg U48807 ( .A(n11612), .B(n12837), .X(n12832) );
  nand_x1_sg U48808 ( .A(n12433), .B(n12838), .X(n12837) );
  nand_x1_sg U48809 ( .A(n12839), .B(n12840), .X(n12838) );
  nor_x1_sg U48810 ( .A(n12120), .B(n41109), .X(n12119) );
  nor_x1_sg U48811 ( .A(n35102), .B(n19587), .X(n13608) );
  nand_x1_sg U48812 ( .A(n15045), .B(n35508), .X(n15044) );
  nand_x1_sg U48813 ( .A(n15045), .B(n35516), .X(n15048) );
  nand_x1_sg U48814 ( .A(n30523), .B(n35504), .X(n15177) );
  nand_x1_sg U48815 ( .A(n15178), .B(n35515), .X(n15180) );
  nand_x1_sg U48816 ( .A(n15178), .B(n35553), .X(n15181) );
  nor_x1_sg U48817 ( .A(n11843), .B(n41109), .X(n11842) );
  nand_x1_sg U48818 ( .A(n19585), .B(n31883), .X(n12430) );
  nand_x1_sg U48819 ( .A(n12525), .B(n12967), .X(n12966) );
  nand_x1_sg U48820 ( .A(n12839), .B(n12968), .X(n12967) );
  nor_x1_sg U48821 ( .A(n13488), .B(n19586), .X(n13487) );
  nor_x1_sg U48822 ( .A(n32939), .B(n31752), .X(n13488) );
  nand_x1_sg U48823 ( .A(n32175), .B(n11663), .X(n11764) );
  nand_x1_sg U48824 ( .A(n11794), .B(n32006), .X(n11793) );
  nor_x1_sg U48825 ( .A(n13364), .B(n35627), .X(n13617) );
  nor_x1_sg U48826 ( .A(n13789), .B(n13790), .X(n13788) );
  nor_x1_sg U48827 ( .A(n13372), .B(n35626), .X(n13622) );
  nor_x1_sg U48828 ( .A(n13826), .B(n13827), .X(n13825) );
  nor_x1_sg U48829 ( .A(n13378), .B(n35625), .X(n13626) );
  nor_x1_sg U48830 ( .A(n13857), .B(n13858), .X(n13856) );
  nor_x1_sg U48831 ( .A(n13384), .B(n41288), .X(n13630) );
  nor_x1_sg U48832 ( .A(n13888), .B(n13889), .X(n13887) );
  nor_x1_sg U48833 ( .A(n13390), .B(n41289), .X(n13634) );
  nor_x1_sg U48834 ( .A(n13919), .B(n13920), .X(n13918) );
  nor_x1_sg U48835 ( .A(n13396), .B(n41290), .X(n13638) );
  nor_x1_sg U48836 ( .A(n13950), .B(n13951), .X(n13949) );
  nor_x1_sg U48837 ( .A(n13402), .B(n41291), .X(n13642) );
  nand_x1_sg U48838 ( .A(n34220), .B(n13980), .X(n13979) );
  nor_x1_sg U48839 ( .A(n13981), .B(n13982), .X(n13980) );
  nor_x1_sg U48840 ( .A(n13408), .B(n41292), .X(n13646) );
  nand_x1_sg U48841 ( .A(n34222), .B(n14011), .X(n14010) );
  nor_x1_sg U48842 ( .A(n14012), .B(n14013), .X(n14011) );
  nor_x1_sg U48843 ( .A(n13414), .B(n41293), .X(n13650) );
  nand_x1_sg U48844 ( .A(n31404), .B(n14042), .X(n14041) );
  nor_x1_sg U48845 ( .A(n14043), .B(n14044), .X(n14042) );
  nor_x1_sg U48846 ( .A(n13420), .B(n41294), .X(n13654) );
  nand_x1_sg U48847 ( .A(n30294), .B(n14073), .X(n14072) );
  nor_x1_sg U48848 ( .A(n14074), .B(n14075), .X(n14073) );
  nor_x1_sg U48849 ( .A(n13426), .B(n41295), .X(n13658) );
  nand_x1_sg U48850 ( .A(n34222), .B(n14104), .X(n14103) );
  nor_x1_sg U48851 ( .A(n14105), .B(n14106), .X(n14104) );
  nor_x1_sg U48852 ( .A(n13432), .B(n41296), .X(n13662) );
  nand_x1_sg U48853 ( .A(n31404), .B(n14135), .X(n14134) );
  nor_x1_sg U48854 ( .A(n14136), .B(n14137), .X(n14135) );
  nor_x1_sg U48855 ( .A(n13438), .B(n41297), .X(n13666) );
  nand_x1_sg U48856 ( .A(n30294), .B(n14166), .X(n14165) );
  nor_x1_sg U48857 ( .A(n14167), .B(n14168), .X(n14166) );
  nor_x1_sg U48858 ( .A(n13444), .B(n41298), .X(n13670) );
  nand_x1_sg U48859 ( .A(n30079), .B(n14197), .X(n14196) );
  nor_x1_sg U48860 ( .A(n14198), .B(n14199), .X(n14197) );
  nor_x1_sg U48861 ( .A(n13450), .B(n41299), .X(n13674) );
  nand_x1_sg U48862 ( .A(n31814), .B(n14228), .X(n14227) );
  nor_x1_sg U48863 ( .A(n14229), .B(n14230), .X(n14228) );
  nor_x1_sg U48864 ( .A(n13456), .B(n41300), .X(n13678) );
  nand_x1_sg U48865 ( .A(n30294), .B(n14259), .X(n14258) );
  nor_x1_sg U48866 ( .A(n14260), .B(n14261), .X(n14259) );
  nor_x1_sg U48867 ( .A(n13462), .B(n41301), .X(n13682) );
  nand_x1_sg U48868 ( .A(n30079), .B(n14290), .X(n14289) );
  nor_x1_sg U48869 ( .A(n14291), .B(n14292), .X(n14290) );
  nor_x1_sg U48870 ( .A(n13468), .B(n41302), .X(n13686) );
  nand_x1_sg U48871 ( .A(n34220), .B(n14321), .X(n14320) );
  nor_x1_sg U48872 ( .A(n14322), .B(n14323), .X(n14321) );
  nor_x1_sg U48873 ( .A(n13474), .B(n41303), .X(n13690) );
  nand_x1_sg U48874 ( .A(n30294), .B(n14352), .X(n14351) );
  nor_x1_sg U48875 ( .A(n14353), .B(n14354), .X(n14352) );
  nor_x1_sg U48876 ( .A(n13480), .B(n41304), .X(n13694) );
  nand_x1_sg U48877 ( .A(n34221), .B(n14383), .X(n14382) );
  nor_x1_sg U48878 ( .A(n14384), .B(n14385), .X(n14383) );
  nor_x1_sg U48879 ( .A(n13493), .B(n41305), .X(n13704) );
  nand_x1_sg U48880 ( .A(n31404), .B(n14415), .X(n14414) );
  nor_x1_sg U48881 ( .A(n14416), .B(n14417), .X(n14415) );
  nor_x1_sg U48882 ( .A(n13499), .B(n41306), .X(n13708) );
  nand_x1_sg U48883 ( .A(n30079), .B(n14446), .X(n14445) );
  nor_x1_sg U48884 ( .A(n14447), .B(n14448), .X(n14446) );
  nor_x1_sg U48885 ( .A(n13510), .B(n41307), .X(n13715) );
  nand_x1_sg U48886 ( .A(n34219), .B(n14510), .X(n14509) );
  nor_x1_sg U48887 ( .A(n14511), .B(n14512), .X(n14510) );
  nor_x1_sg U48888 ( .A(n13521), .B(n41308), .X(n13722) );
  nand_x1_sg U48889 ( .A(n34220), .B(n14572), .X(n14571) );
  nor_x1_sg U48890 ( .A(n14573), .B(n14574), .X(n14572) );
  nor_x1_sg U48891 ( .A(n13527), .B(n41309), .X(n13726) );
  nand_x1_sg U48892 ( .A(n31405), .B(n14603), .X(n14602) );
  nor_x1_sg U48893 ( .A(n14604), .B(n14605), .X(n14603) );
  nor_x1_sg U48894 ( .A(n13533), .B(n41310), .X(n13730) );
  nand_x1_sg U48895 ( .A(n31814), .B(n14634), .X(n14633) );
  nor_x1_sg U48896 ( .A(n14635), .B(n14636), .X(n14634) );
  nor_x1_sg U48897 ( .A(n13539), .B(n41311), .X(n13734) );
  nand_x1_sg U48898 ( .A(n31405), .B(n14665), .X(n14664) );
  nor_x1_sg U48899 ( .A(n14666), .B(n14667), .X(n14665) );
  nor_x1_sg U48900 ( .A(n13545), .B(n41312), .X(n13738) );
  nand_x1_sg U48901 ( .A(n34220), .B(n14696), .X(n14695) );
  nor_x1_sg U48902 ( .A(n14697), .B(n14698), .X(n14696) );
  nor_x1_sg U48903 ( .A(n13551), .B(n41313), .X(n13742) );
  nand_x1_sg U48904 ( .A(n30292), .B(n14727), .X(n14726) );
  nor_x1_sg U48905 ( .A(n14728), .B(n14729), .X(n14727) );
  nor_x1_sg U48906 ( .A(n13557), .B(n41314), .X(n13746) );
  nand_x1_sg U48907 ( .A(n30292), .B(n14758), .X(n14757) );
  nor_x1_sg U48908 ( .A(n14759), .B(n14760), .X(n14758) );
  nor_x1_sg U48909 ( .A(n13563), .B(n41315), .X(n13750) );
  nand_x1_sg U48910 ( .A(n31405), .B(n14789), .X(n14788) );
  nor_x1_sg U48911 ( .A(n14790), .B(n14791), .X(n14789) );
  nor_x1_sg U48912 ( .A(n13569), .B(n41316), .X(n13754) );
  nand_x1_sg U48913 ( .A(n31814), .B(n14820), .X(n14819) );
  nor_x1_sg U48914 ( .A(n14821), .B(n14822), .X(n14820) );
  nor_x1_sg U48915 ( .A(n13575), .B(n41317), .X(n13758) );
  nand_x1_sg U48916 ( .A(n34219), .B(n14851), .X(n14850) );
  nor_x1_sg U48917 ( .A(n14852), .B(n14853), .X(n14851) );
  nor_x1_sg U48918 ( .A(n13581), .B(n41318), .X(n13762) );
  nand_x1_sg U48919 ( .A(n30079), .B(n14882), .X(n14881) );
  nor_x1_sg U48920 ( .A(n14883), .B(n14884), .X(n14882) );
  nor_x1_sg U48921 ( .A(n13587), .B(n41319), .X(n13766) );
  nand_x1_sg U48922 ( .A(n34221), .B(n14913), .X(n14912) );
  nor_x1_sg U48923 ( .A(n14914), .B(n14915), .X(n14913) );
  nor_x1_sg U48924 ( .A(n13603), .B(n41320), .X(n13776) );
  nand_x1_sg U48925 ( .A(n31814), .B(n15006), .X(n15005) );
  nor_x1_sg U48926 ( .A(n15007), .B(n15008), .X(n15006) );
  nand_x1_sg U48927 ( .A(n35515), .B(n35249), .X(n15171) );
  nor_x1_sg U48928 ( .A(n34424), .B(n11612), .X(n11610) );
  nor_x1_sg U48929 ( .A(n35096), .B(n35272), .X(n15201) );
  nor_x1_sg U48930 ( .A(n12617), .B(n33833), .X(n12614) );
  nor_x1_sg U48931 ( .A(n35563), .B(n19586), .X(n12617) );
  nor_x1_sg U48932 ( .A(n12709), .B(n33839), .X(n12706) );
  nor_x1_sg U48933 ( .A(n42536), .B(n19587), .X(n12709) );
  nand_x1_sg U48934 ( .A(n35302), .B(n12836), .X(n12835) );
  nand_x1_sg U48935 ( .A(n31702), .B(n35105), .X(n12836) );
  nand_x1_sg U48936 ( .A(n35304), .B(n12965), .X(n12964) );
  nand_x1_sg U48937 ( .A(n31698), .B(n35106), .X(n12965) );
  nor_x1_sg U48938 ( .A(n35267), .B(n35280), .X(n12708) );
  nor_x1_sg U48939 ( .A(n41183), .B(n11636), .X(n11634) );
  nor_x1_sg U48940 ( .A(n11637), .B(n11638), .X(n11636) );
  nor_x1_sg U48941 ( .A(n11639), .B(n35456), .X(n11638) );
  nor_x1_sg U48942 ( .A(n30539), .B(n11689), .X(n11688) );
  nor_x1_sg U48943 ( .A(n30517), .B(n32198), .X(n11689) );
  nand_x1_sg U48944 ( .A(n41110), .B(n11846), .X(n11845) );
  nand_x1_sg U48945 ( .A(n31882), .B(n35105), .X(n11846) );
  nand_x1_sg U48946 ( .A(n35099), .B(n11892), .X(n11891) );
  nand_x1_sg U48947 ( .A(n32005), .B(n35106), .X(n11892) );
  nor_x1_sg U48948 ( .A(n13611), .B(n13612), .X(n13610) );
  nor_x1_sg U48949 ( .A(n13613), .B(n32058), .X(n13609) );
  nand_x1_sg U48950 ( .A(n32934), .B(n32396), .X(n13612) );
  nor_x1_sg U48951 ( .A(n11664), .B(n11665), .X(n11662) );
  nor_x1_sg U48952 ( .A(n11609), .B(n34434), .X(n11665) );
  nand_x1_sg U48953 ( .A(n30138), .B(n13940), .X(n13939) );
  nand_x1_sg U48954 ( .A(n31751), .B(n42735), .X(n13940) );
  nand_x1_sg U48955 ( .A(n32171), .B(n14095), .X(n14094) );
  nand_x1_sg U48956 ( .A(n34411), .B(n42737), .X(n14095) );
  nand_x1_sg U48957 ( .A(n31299), .B(n14219), .X(n14218) );
  nand_x1_sg U48958 ( .A(n34409), .B(n42739), .X(n14219) );
  nand_x1_sg U48959 ( .A(n32170), .B(n14374), .X(n14373) );
  nand_x1_sg U48960 ( .A(n31750), .B(n42741), .X(n14374) );
  nand_x1_sg U48961 ( .A(n32167), .B(n14718), .X(n14717) );
  nand_x1_sg U48962 ( .A(n30114), .B(n42624), .X(n14718) );
  nand_x1_sg U48963 ( .A(n30138), .B(n14842), .X(n14841) );
  nand_x1_sg U48964 ( .A(n34410), .B(n42626), .X(n14842) );
  nor_x1_sg U48965 ( .A(n35279), .B(n35271), .X(n12616) );
  nand_x1_sg U48966 ( .A(n14502), .B(n14503), .X(n14498) );
  nand_x1_sg U48967 ( .A(n14564), .B(n14565), .X(n14560) );
  nand_x1_sg U48968 ( .A(n14967), .B(n14968), .X(n14963) );
  nand_x1_sg U48969 ( .A(n14998), .B(n14999), .X(n14994) );
  nor_x1_sg U48970 ( .A(n11795), .B(n35267), .X(n11794) );
  nor_x1_sg U48971 ( .A(n11796), .B(n34519), .X(n11795) );
  nor_x1_sg U48972 ( .A(n41418), .B(n11797), .X(n11796) );
  nand_x1_sg U48973 ( .A(n31670), .B(n35280), .X(n11797) );
  nand_x1_sg U48974 ( .A(n34559), .B(n13909), .X(n13908) );
  nand_x1_sg U48975 ( .A(n34411), .B(n42734), .X(n13909) );
  nand_x1_sg U48976 ( .A(n32172), .B(n14064), .X(n14063) );
  nand_x1_sg U48977 ( .A(n31750), .B(n42736), .X(n14064) );
  nand_x1_sg U48978 ( .A(n32168), .B(n14188), .X(n14187) );
  nand_x1_sg U48979 ( .A(n31750), .B(n42738), .X(n14188) );
  nand_x1_sg U48980 ( .A(n32167), .B(n14343), .X(n14342) );
  nand_x1_sg U48981 ( .A(n34410), .B(n42740), .X(n14343) );
  nand_x1_sg U48982 ( .A(n32171), .B(n14687), .X(n14686) );
  nand_x1_sg U48983 ( .A(n34408), .B(n42623), .X(n14687) );
  nand_x1_sg U48984 ( .A(n34551), .B(n14811), .X(n14810) );
  nand_x1_sg U48985 ( .A(n31750), .B(n42625), .X(n14811) );
  nand_x1_sg U48986 ( .A(n32168), .B(n14935), .X(n14934) );
  nand_x1_sg U48987 ( .A(n34408), .B(n42628), .X(n14935) );
  nor_x1_sg U48988 ( .A(n13505), .B(n13506), .X(n13504) );
  nor_x1_sg U48989 ( .A(n35151), .B(n30090), .X(n13506) );
  nor_x1_sg U48990 ( .A(n34344), .B(n41094), .X(n13505) );
  nor_x1_sg U48991 ( .A(n13516), .B(n13517), .X(n13515) );
  nor_x1_sg U48992 ( .A(n42573), .B(n31371), .X(n13517) );
  nor_x1_sg U48993 ( .A(n31770), .B(n42565), .X(n13516) );
  nor_x1_sg U48994 ( .A(n13593), .B(n13594), .X(n13592) );
  nor_x1_sg U48995 ( .A(n42578), .B(n34274), .X(n13594) );
  nor_x1_sg U48996 ( .A(n34344), .B(n42570), .X(n13593) );
  nor_x1_sg U48997 ( .A(n13598), .B(n13599), .X(n13597) );
  nor_x1_sg U48998 ( .A(n42579), .B(n30320), .X(n13599) );
  nor_x1_sg U48999 ( .A(n31770), .B(n42571), .X(n13598) );
  nor_x1_sg U49000 ( .A(n11714), .B(n35302), .X(n11713) );
  nor_x1_sg U49001 ( .A(n11715), .B(n34516), .X(n11714) );
  nor_x1_sg U49002 ( .A(n31702), .B(n11664), .X(n11715) );
  nor_x1_sg U49003 ( .A(n11741), .B(n35304), .X(n11740) );
  nor_x1_sg U49004 ( .A(n11742), .B(n34515), .X(n11741) );
  nor_x1_sg U49005 ( .A(n31699), .B(n11664), .X(n11742) );
  nor_x1_sg U49006 ( .A(n11559), .B(n11585), .X(n11584) );
  nor_x1_sg U49007 ( .A(n35267), .B(n35099), .X(n11583) );
  nor_x1_sg U49008 ( .A(n41110), .B(n35271), .X(n11557) );
  nor_x1_sg U49009 ( .A(n11559), .B(n11560), .X(n11558) );
  nor_x1_sg U49010 ( .A(n11610), .B(n41110), .X(n11607) );
  nor_x1_sg U49011 ( .A(n41183), .B(n30518), .X(n11608) );
  nor_x1_sg U49012 ( .A(n15123), .B(n15124), .X(n15122) );
  nand_x4_sg U49013 ( .A(n15147), .B(n15148), .X(n15140) );
  nor_x1_sg U49014 ( .A(n15252), .B(n15253), .X(n15251) );
  nand_x4_sg U49015 ( .A(n15276), .B(n15277), .X(n15269) );
  nand_x1_sg U49016 ( .A(n34088), .B(n12980), .X(n13828) );
  nand_x1_sg U49017 ( .A(n34089), .B(n12986), .X(n13859) );
  nand_x1_sg U49018 ( .A(n31866), .B(n13010), .X(n13983) );
  nand_x1_sg U49019 ( .A(n30040), .B(n13034), .X(n14107) );
  nand_x1_sg U49020 ( .A(n34089), .B(n13040), .X(n14138) );
  nand_x1_sg U49021 ( .A(n30039), .B(n13064), .X(n14262) );
  nand_x1_sg U49022 ( .A(n31495), .B(n13088), .X(n14386) );
  nand_x1_sg U49023 ( .A(n31867), .B(n13103), .X(n14418) );
  nand_x1_sg U49024 ( .A(n34087), .B(n13139), .X(n14606) );
  nand_x1_sg U49025 ( .A(n31866), .B(n13163), .X(n14730) );
  nand_x1_sg U49026 ( .A(n34087), .B(n13169), .X(n14761) );
  nand_x1_sg U49027 ( .A(n30040), .B(n13193), .X(n14885) );
  nand_x1_sg U49028 ( .A(n31495), .B(n12972), .X(n13791) );
  nand_x1_sg U49029 ( .A(n31866), .B(n12998), .X(n13921) );
  nand_x1_sg U49030 ( .A(n30039), .B(n13004), .X(n13952) );
  nand_x1_sg U49031 ( .A(n31867), .B(n13028), .X(n14076) );
  nand_x1_sg U49032 ( .A(n34086), .B(n13052), .X(n14200) );
  nand_x1_sg U49033 ( .A(n31866), .B(n13058), .X(n14231) );
  nand_x1_sg U49034 ( .A(n34087), .B(n13082), .X(n14355) );
  nand_x1_sg U49035 ( .A(n30040), .B(n13122), .X(n14513) );
  nand_x1_sg U49036 ( .A(n34086), .B(n13133), .X(n14575) );
  nand_x1_sg U49037 ( .A(n34088), .B(n13157), .X(n14699) );
  nand_x1_sg U49038 ( .A(n31867), .B(n13181), .X(n14823) );
  nand_x1_sg U49039 ( .A(n31495), .B(n13187), .X(n14854) );
  nand_x1_sg U49040 ( .A(n31494), .B(n12992), .X(n13890) );
  nand_x1_sg U49041 ( .A(n34087), .B(n13016), .X(n14014) );
  nand_x1_sg U49042 ( .A(n34089), .B(n13022), .X(n14045) );
  nand_x1_sg U49043 ( .A(n30039), .B(n13046), .X(n14169) );
  nand_x1_sg U49044 ( .A(n34086), .B(n13070), .X(n14293) );
  nand_x1_sg U49045 ( .A(n31495), .B(n13076), .X(n14324) );
  nand_x1_sg U49046 ( .A(n31494), .B(n13111), .X(n14449) );
  nand_x1_sg U49047 ( .A(n34088), .B(n13145), .X(n14637) );
  nand_x1_sg U49048 ( .A(n31494), .B(n13151), .X(n14668) );
  nand_x1_sg U49049 ( .A(n31494), .B(n13175), .X(n14792) );
  nand_x1_sg U49050 ( .A(n34088), .B(n13199), .X(n14916) );
  nand_x1_sg U49051 ( .A(n34089), .B(n13215), .X(n15009) );
  nor_x1_sg U49052 ( .A(n31875), .B(n15106), .X(n15082) );
  nand_x4_sg U49053 ( .A(n15114), .B(n15115), .X(n15107) );
  nand_x4_sg U49054 ( .A(n15109), .B(n15110), .X(n15108) );
  nor_x1_sg U49055 ( .A(n31875), .B(n15235), .X(n15218) );
  nand_x4_sg U49056 ( .A(n15243), .B(n15244), .X(n15236) );
  nand_x4_sg U49057 ( .A(n15238), .B(n15239), .X(n15237) );
  nand_x1_sg U49058 ( .A(n30537), .B(n31699), .X(n12526) );
  nand_x1_sg U49059 ( .A(n32000), .B(n32504), .X(n15157) );
  nand_x1_sg U49060 ( .A(n35460), .B(n31203), .X(n15156) );
  nand_x1_sg U49061 ( .A(n31875), .B(n15167), .X(n15166) );
  nor_x1_sg U49062 ( .A(n15167), .B(n31876), .X(n15168) );
  nor_x1_sg U49063 ( .A(n13811), .B(n13812), .X(n13798) );
  nand_x1_sg U49064 ( .A(n13814), .B(n13815), .X(n13811) );
  nor_x1_sg U49065 ( .A(n13845), .B(n13846), .X(n13835) );
  nand_x1_sg U49066 ( .A(n13848), .B(n13849), .X(n13845) );
  nor_x1_sg U49067 ( .A(n13876), .B(n13877), .X(n13866) );
  nand_x1_sg U49068 ( .A(n13879), .B(n13880), .X(n13876) );
  nand_x1_sg U49069 ( .A(n13910), .B(n13911), .X(n13907) );
  nand_x1_sg U49070 ( .A(n13941), .B(n13942), .X(n13938) );
  nor_x1_sg U49071 ( .A(n13969), .B(n13970), .X(n13959) );
  nand_x1_sg U49072 ( .A(n13972), .B(n13973), .X(n13969) );
  nor_x1_sg U49073 ( .A(n14000), .B(n14001), .X(n13990) );
  nand_x1_sg U49074 ( .A(n14003), .B(n14004), .X(n14000) );
  nor_x1_sg U49075 ( .A(n14031), .B(n14032), .X(n14021) );
  nand_x1_sg U49076 ( .A(n14034), .B(n14035), .X(n14031) );
  nor_x1_sg U49077 ( .A(n14124), .B(n14125), .X(n14114) );
  nand_x1_sg U49078 ( .A(n14127), .B(n14128), .X(n14124) );
  nor_x1_sg U49079 ( .A(n14155), .B(n14156), .X(n14145) );
  nand_x1_sg U49080 ( .A(n14158), .B(n14159), .X(n14155) );
  nor_x1_sg U49081 ( .A(n14248), .B(n14249), .X(n14238) );
  nand_x1_sg U49082 ( .A(n14251), .B(n14252), .X(n14248) );
  nor_x1_sg U49083 ( .A(n14279), .B(n14280), .X(n14269) );
  nand_x1_sg U49084 ( .A(n14282), .B(n14283), .X(n14279) );
  nor_x1_sg U49085 ( .A(n14310), .B(n14311), .X(n14300) );
  nand_x1_sg U49086 ( .A(n14313), .B(n14314), .X(n14310) );
  nand_x1_sg U49087 ( .A(n14344), .B(n14345), .X(n14341) );
  nand_x1_sg U49088 ( .A(n14375), .B(n14376), .X(n14372) );
  nor_x1_sg U49089 ( .A(n14403), .B(n14404), .X(n14393) );
  nand_x1_sg U49090 ( .A(n14406), .B(n14407), .X(n14403) );
  nor_x1_sg U49091 ( .A(n14435), .B(n14436), .X(n14425) );
  nand_x1_sg U49092 ( .A(n14438), .B(n14439), .X(n14435) );
  nor_x1_sg U49093 ( .A(n14466), .B(n14467), .X(n14456) );
  nand_x1_sg U49094 ( .A(n14469), .B(n14470), .X(n14466) );
  nor_x1_sg U49095 ( .A(n14530), .B(n14531), .X(n14520) );
  nand_x1_sg U49096 ( .A(n14533), .B(n14534), .X(n14530) );
  nor_x1_sg U49097 ( .A(n14592), .B(n14593), .X(n14582) );
  nand_x1_sg U49098 ( .A(n14595), .B(n14596), .X(n14592) );
  nor_x1_sg U49099 ( .A(n14623), .B(n14624), .X(n14613) );
  nand_x1_sg U49100 ( .A(n14626), .B(n14627), .X(n14623) );
  nor_x1_sg U49101 ( .A(n14654), .B(n14655), .X(n14644) );
  nand_x1_sg U49102 ( .A(n14657), .B(n14658), .X(n14654) );
  nand_x1_sg U49103 ( .A(n14688), .B(n14689), .X(n14685) );
  nand_x1_sg U49104 ( .A(n14719), .B(n14720), .X(n14716) );
  nor_x1_sg U49105 ( .A(n14747), .B(n14748), .X(n14737) );
  nand_x1_sg U49106 ( .A(n14750), .B(n14751), .X(n14747) );
  nor_x1_sg U49107 ( .A(n14778), .B(n14779), .X(n14768) );
  nand_x1_sg U49108 ( .A(n14781), .B(n14782), .X(n14778) );
  nand_x1_sg U49109 ( .A(n14812), .B(n14813), .X(n14809) );
  nand_x1_sg U49110 ( .A(n14843), .B(n14844), .X(n14840) );
  nor_x1_sg U49111 ( .A(n14871), .B(n14872), .X(n14861) );
  nand_x1_sg U49112 ( .A(n14874), .B(n14875), .X(n14871) );
  nor_x1_sg U49113 ( .A(n14902), .B(n14903), .X(n14892) );
  nand_x1_sg U49114 ( .A(n14905), .B(n14906), .X(n14902) );
  nand_x1_sg U49115 ( .A(n14936), .B(n14937), .X(n14933) );
  nor_x1_sg U49116 ( .A(n15026), .B(n15027), .X(n15016) );
  nand_x1_sg U49117 ( .A(n15029), .B(n15030), .X(n15026) );
  nand_x1_sg U49118 ( .A(n12858), .B(n34562), .X(n12857) );
  nor_x1_sg U49119 ( .A(n12630), .B(n12859), .X(n12856) );
  nor_x1_sg U49120 ( .A(n34406), .B(n41082), .X(n12859) );
  nand_x1_sg U49121 ( .A(n12870), .B(n32393), .X(n12869) );
  nor_x1_sg U49122 ( .A(n12639), .B(n12871), .X(n12868) );
  nor_x1_sg U49123 ( .A(n34405), .B(n42589), .X(n12871) );
  nand_x1_sg U49124 ( .A(n12948), .B(n34561), .X(n12947) );
  nor_x1_sg U49125 ( .A(n12692), .B(n12949), .X(n12946) );
  nor_x1_sg U49126 ( .A(n31996), .B(n42594), .X(n12949) );
  nand_x1_sg U49127 ( .A(n12954), .B(n32391), .X(n12953) );
  nor_x1_sg U49128 ( .A(n12697), .B(n12955), .X(n12952) );
  nor_x1_sg U49129 ( .A(n30113), .B(n42595), .X(n12955) );
  nor_x1_sg U49130 ( .A(n35614), .B(n12716), .X(n12713) );
  nand_x1_sg U49131 ( .A(n12715), .B(n32398), .X(n12714) );
  nor_x1_sg U49132 ( .A(n31998), .B(n40961), .X(n12716) );
  nor_x1_sg U49133 ( .A(n35561), .B(n12723), .X(n12720) );
  nand_x1_sg U49134 ( .A(n12722), .B(n32393), .X(n12721) );
  nor_x1_sg U49135 ( .A(n31996), .B(n40960), .X(n12723) );
  nor_x1_sg U49136 ( .A(n35613), .B(n12729), .X(n12726) );
  nand_x1_sg U49137 ( .A(n12728), .B(n34560), .X(n12727) );
  nor_x1_sg U49138 ( .A(n34403), .B(n40959), .X(n12729) );
  nor_x1_sg U49139 ( .A(n35509), .B(n12735), .X(n12732) );
  nand_x1_sg U49140 ( .A(n12734), .B(n30142), .X(n12733) );
  nor_x1_sg U49141 ( .A(n34403), .B(n42698), .X(n12735) );
  nor_x1_sg U49142 ( .A(n35604), .B(n12741), .X(n12738) );
  nand_x1_sg U49143 ( .A(n12740), .B(n32388), .X(n12739) );
  nor_x1_sg U49144 ( .A(n12717), .B(n42699), .X(n12741) );
  nor_x1_sg U49145 ( .A(n35619), .B(n12747), .X(n12744) );
  nand_x1_sg U49146 ( .A(n12746), .B(n32397), .X(n12745) );
  nor_x1_sg U49147 ( .A(n30857), .B(n40958), .X(n12747) );
  nand_x1_sg U49148 ( .A(n12752), .B(n30143), .X(n12751) );
  nor_x1_sg U49149 ( .A(n35514), .B(n12753), .X(n12750) );
  nor_x1_sg U49150 ( .A(n12717), .B(n40957), .X(n12753) );
  nand_x1_sg U49151 ( .A(n12758), .B(n34563), .X(n12757) );
  nor_x1_sg U49152 ( .A(n35618), .B(n12759), .X(n12756) );
  nor_x1_sg U49153 ( .A(n34404), .B(n40956), .X(n12759) );
  nand_x1_sg U49154 ( .A(n12764), .B(n32392), .X(n12763) );
  nor_x1_sg U49155 ( .A(n35612), .B(n12765), .X(n12762) );
  nor_x1_sg U49156 ( .A(n34406), .B(n42700), .X(n12765) );
  nand_x1_sg U49157 ( .A(n12770), .B(n34560), .X(n12769) );
  nor_x1_sg U49158 ( .A(n35617), .B(n12771), .X(n12768) );
  nor_x1_sg U49159 ( .A(n31998), .B(n42701), .X(n12771) );
  nand_x1_sg U49160 ( .A(n12776), .B(n32388), .X(n12775) );
  nor_x1_sg U49161 ( .A(n35602), .B(n12777), .X(n12774) );
  nor_x1_sg U49162 ( .A(n34405), .B(n40955), .X(n12777) );
  nand_x1_sg U49163 ( .A(n12782), .B(n32392), .X(n12781) );
  nor_x1_sg U49164 ( .A(n35616), .B(n12783), .X(n12780) );
  nor_x1_sg U49165 ( .A(n31997), .B(n40954), .X(n12783) );
  nand_x1_sg U49166 ( .A(n12788), .B(n32387), .X(n12787) );
  nor_x1_sg U49167 ( .A(n35611), .B(n12789), .X(n12786) );
  nor_x1_sg U49168 ( .A(n31997), .B(n42702), .X(n12789) );
  nand_x1_sg U49169 ( .A(n12794), .B(n32396), .X(n12793) );
  nor_x1_sg U49170 ( .A(n35615), .B(n12795), .X(n12792) );
  nor_x1_sg U49171 ( .A(n34406), .B(n42703), .X(n12795) );
  nand_x1_sg U49172 ( .A(n12800), .B(n34563), .X(n12799) );
  nor_x1_sg U49173 ( .A(n35610), .B(n12801), .X(n12798) );
  nor_x1_sg U49174 ( .A(n34404), .B(n40953), .X(n12801) );
  nand_x1_sg U49175 ( .A(n12806), .B(n32397), .X(n12805) );
  nor_x1_sg U49176 ( .A(n35609), .B(n12807), .X(n12804) );
  nor_x1_sg U49177 ( .A(n31997), .B(n40952), .X(n12807) );
  nand_x1_sg U49178 ( .A(n12812), .B(n32390), .X(n12811) );
  nor_x1_sg U49179 ( .A(n35601), .B(n12813), .X(n12810) );
  nor_x1_sg U49180 ( .A(n30857), .B(n40951), .X(n12813) );
  nand_x1_sg U49181 ( .A(n12818), .B(n32387), .X(n12817) );
  nor_x1_sg U49182 ( .A(n35608), .B(n12819), .X(n12816) );
  nor_x1_sg U49183 ( .A(n31752), .B(n42704), .X(n12819) );
  nand_x1_sg U49184 ( .A(n12824), .B(n34563), .X(n12823) );
  nor_x1_sg U49185 ( .A(n35607), .B(n12825), .X(n12822) );
  nor_x1_sg U49186 ( .A(n30113), .B(n42705), .X(n12825) );
  nand_x1_sg U49187 ( .A(n12830), .B(n32395), .X(n12829) );
  nor_x1_sg U49188 ( .A(n35603), .B(n12831), .X(n12828) );
  nor_x1_sg U49189 ( .A(n12717), .B(n40950), .X(n12831) );
  nand_x1_sg U49190 ( .A(n12846), .B(n30143), .X(n12845) );
  nor_x1_sg U49191 ( .A(n35503), .B(n12847), .X(n12844) );
  nor_x1_sg U49192 ( .A(n31998), .B(n41084), .X(n12847) );
  nand_x1_sg U49193 ( .A(n12852), .B(n32390), .X(n12851) );
  nor_x1_sg U49194 ( .A(n35593), .B(n12853), .X(n12850) );
  nor_x1_sg U49195 ( .A(n34405), .B(n41083), .X(n12853) );
  nand_x1_sg U49196 ( .A(n12864), .B(n30142), .X(n12863) );
  nor_x1_sg U49197 ( .A(n35592), .B(n12865), .X(n12862) );
  nor_x1_sg U49198 ( .A(n30113), .B(n42588), .X(n12865) );
  nand_x1_sg U49199 ( .A(n12876), .B(n32396), .X(n12875) );
  nor_x1_sg U49200 ( .A(n35591), .B(n12877), .X(n12874) );
  nor_x1_sg U49201 ( .A(n31752), .B(n41081), .X(n12877) );
  nand_x1_sg U49202 ( .A(n12882), .B(n32388), .X(n12881) );
  nor_x1_sg U49203 ( .A(n35590), .B(n12883), .X(n12880) );
  nor_x1_sg U49204 ( .A(n30857), .B(n41080), .X(n12883) );
  nand_x1_sg U49205 ( .A(n12888), .B(n32398), .X(n12887) );
  nor_x1_sg U49206 ( .A(n35506), .B(n12889), .X(n12886) );
  nor_x1_sg U49207 ( .A(n34403), .B(n41079), .X(n12889) );
  nand_x1_sg U49208 ( .A(n12894), .B(n32398), .X(n12893) );
  nor_x1_sg U49209 ( .A(n35589), .B(n12895), .X(n12892) );
  nor_x1_sg U49210 ( .A(n31996), .B(n42590), .X(n12895) );
  nand_x1_sg U49211 ( .A(n12900), .B(n32391), .X(n12899) );
  nor_x1_sg U49212 ( .A(n35588), .B(n12901), .X(n12898) );
  nor_x1_sg U49213 ( .A(n34404), .B(n42591), .X(n12901) );
  nand_x1_sg U49214 ( .A(n12906), .B(n32395), .X(n12905) );
  nor_x1_sg U49215 ( .A(n35513), .B(n12907), .X(n12904) );
  nor_x1_sg U49216 ( .A(n31996), .B(n41078), .X(n12907) );
  nand_x1_sg U49217 ( .A(n12912), .B(n34561), .X(n12911) );
  nor_x1_sg U49218 ( .A(n35587), .B(n12913), .X(n12910) );
  nor_x1_sg U49219 ( .A(n34406), .B(n41077), .X(n12913) );
  nand_x1_sg U49220 ( .A(n12918), .B(n32395), .X(n12917) );
  nor_x1_sg U49221 ( .A(n35586), .B(n12919), .X(n12916) );
  nor_x1_sg U49222 ( .A(n30113), .B(n42592), .X(n12919) );
  nand_x1_sg U49223 ( .A(n12924), .B(n34562), .X(n12923) );
  nor_x1_sg U49224 ( .A(n35505), .B(n12925), .X(n12922) );
  nor_x1_sg U49225 ( .A(n34405), .B(n42593), .X(n12925) );
  nand_x1_sg U49226 ( .A(n12930), .B(n34560), .X(n12929) );
  nor_x1_sg U49227 ( .A(n35585), .B(n12931), .X(n12928) );
  nor_x1_sg U49228 ( .A(n31752), .B(n41076), .X(n12931) );
  nand_x1_sg U49229 ( .A(n12936), .B(n32391), .X(n12935) );
  nor_x1_sg U49230 ( .A(n35584), .B(n12937), .X(n12934) );
  nor_x1_sg U49231 ( .A(n31997), .B(n41075), .X(n12937) );
  nand_x1_sg U49232 ( .A(n12942), .B(n34561), .X(n12941) );
  nor_x1_sg U49233 ( .A(n35512), .B(n12943), .X(n12940) );
  nor_x1_sg U49234 ( .A(n30857), .B(n41074), .X(n12943) );
  nand_x1_sg U49235 ( .A(n12960), .B(n32393), .X(n12959) );
  nor_x1_sg U49236 ( .A(n35583), .B(n12961), .X(n12958) );
  nor_x1_sg U49237 ( .A(n34403), .B(n41073), .X(n12961) );
  nor_x1_sg U49238 ( .A(n13365), .B(n13366), .X(n13363) );
  nor_x1_sg U49239 ( .A(n35128), .B(n31371), .X(n13366) );
  nor_x1_sg U49240 ( .A(n31769), .B(n40973), .X(n13365) );
  nor_x1_sg U49241 ( .A(n13385), .B(n13386), .X(n13383) );
  nor_x1_sg U49242 ( .A(n42682), .B(n31797), .X(n13386) );
  nor_x1_sg U49243 ( .A(n31329), .B(n42674), .X(n13385) );
  nor_x1_sg U49244 ( .A(n13403), .B(n13404), .X(n13401) );
  nor_x1_sg U49245 ( .A(n35124), .B(n34276), .X(n13404) );
  nor_x1_sg U49246 ( .A(n29713), .B(n40969), .X(n13403) );
  nor_x1_sg U49247 ( .A(n13421), .B(n13422), .X(n13419) );
  nor_x1_sg U49248 ( .A(n42685), .B(n34277), .X(n13422) );
  nor_x1_sg U49249 ( .A(n30348), .B(n42677), .X(n13421) );
  nor_x1_sg U49250 ( .A(n13439), .B(n13440), .X(n13437) );
  nor_x1_sg U49251 ( .A(n42686), .B(n34275), .X(n13440) );
  nor_x1_sg U49252 ( .A(n31770), .B(n42678), .X(n13439) );
  nor_x1_sg U49253 ( .A(n13457), .B(n13458), .X(n13455) );
  nor_x1_sg U49254 ( .A(n35119), .B(n29727), .X(n13458) );
  nor_x1_sg U49255 ( .A(n31329), .B(n40964), .X(n13457) );
  nor_x1_sg U49256 ( .A(n13475), .B(n13476), .X(n13473) );
  nor_x1_sg U49257 ( .A(n42689), .B(n31372), .X(n13476) );
  nor_x1_sg U49258 ( .A(n34344), .B(n42681), .X(n13475) );
  nor_x1_sg U49259 ( .A(n13500), .B(n13501), .X(n13498) );
  nor_x1_sg U49260 ( .A(n35152), .B(n31372), .X(n13501) );
  nor_x1_sg U49261 ( .A(n31329), .B(n41095), .X(n13500) );
  nor_x1_sg U49262 ( .A(n13534), .B(n13535), .X(n13532) );
  nor_x1_sg U49263 ( .A(n35148), .B(n31371), .X(n13535) );
  nor_x1_sg U49264 ( .A(n31769), .B(n41091), .X(n13534) );
  nor_x1_sg U49265 ( .A(n13552), .B(n13553), .X(n13550) );
  nor_x1_sg U49266 ( .A(n35147), .B(n34275), .X(n13553) );
  nor_x1_sg U49267 ( .A(n34344), .B(n41090), .X(n13552) );
  nor_x1_sg U49268 ( .A(n13570), .B(n13571), .X(n13568) );
  nor_x1_sg U49269 ( .A(n42577), .B(n34274), .X(n13571) );
  nor_x1_sg U49270 ( .A(n30104), .B(n42569), .X(n13570) );
  nor_x1_sg U49271 ( .A(n13588), .B(n13589), .X(n13586) );
  nor_x1_sg U49272 ( .A(n35143), .B(n31797), .X(n13589) );
  nor_x1_sg U49273 ( .A(n34346), .B(n41086), .X(n13588) );
  nor_x1_sg U49274 ( .A(n13604), .B(n13605), .X(n13602) );
  nor_x1_sg U49275 ( .A(n35142), .B(n31798), .X(n13605) );
  nor_x1_sg U49276 ( .A(n31329), .B(n41085), .X(n13604) );
  nor_x1_sg U49277 ( .A(n13373), .B(n13374), .X(n13371) );
  nor_x1_sg U49278 ( .A(n35127), .B(n34274), .X(n13374) );
  nor_x1_sg U49279 ( .A(n13368), .B(n40972), .X(n13373) );
  nor_x1_sg U49280 ( .A(n13379), .B(n13380), .X(n13377) );
  nor_x1_sg U49281 ( .A(n35126), .B(n31798), .X(n13380) );
  nor_x1_sg U49282 ( .A(n34345), .B(n40971), .X(n13379) );
  nor_x1_sg U49283 ( .A(n13391), .B(n13392), .X(n13389) );
  nor_x1_sg U49284 ( .A(n42683), .B(n29727), .X(n13392) );
  nor_x1_sg U49285 ( .A(n34345), .B(n42675), .X(n13391) );
  nor_x1_sg U49286 ( .A(n13397), .B(n13398), .X(n13395) );
  nor_x1_sg U49287 ( .A(n35125), .B(n30090), .X(n13398) );
  nor_x1_sg U49288 ( .A(n31330), .B(n40970), .X(n13397) );
  nor_x1_sg U49289 ( .A(n13409), .B(n13410), .X(n13407) );
  nor_x1_sg U49290 ( .A(n35123), .B(n31372), .X(n13410) );
  nor_x1_sg U49291 ( .A(n34346), .B(n40968), .X(n13409) );
  nor_x1_sg U49292 ( .A(n13415), .B(n13416), .X(n13413) );
  nor_x1_sg U49293 ( .A(n42684), .B(n34277), .X(n13416) );
  nor_x1_sg U49294 ( .A(n30104), .B(n42676), .X(n13415) );
  nor_x1_sg U49295 ( .A(n13427), .B(n13428), .X(n13425) );
  nor_x1_sg U49296 ( .A(n35122), .B(n30320), .X(n13428) );
  nor_x1_sg U49297 ( .A(n34347), .B(n40967), .X(n13427) );
  nor_x1_sg U49298 ( .A(n13433), .B(n13434), .X(n13431) );
  nor_x1_sg U49299 ( .A(n35121), .B(n31372), .X(n13434) );
  nor_x1_sg U49300 ( .A(n34347), .B(n40966), .X(n13433) );
  nor_x1_sg U49301 ( .A(n13445), .B(n13446), .X(n13443) );
  nor_x1_sg U49302 ( .A(n42687), .B(n31371), .X(n13446) );
  nor_x1_sg U49303 ( .A(n30104), .B(n42679), .X(n13445) );
  nor_x1_sg U49304 ( .A(n13451), .B(n13452), .X(n13449) );
  nor_x1_sg U49305 ( .A(n35120), .B(n31797), .X(n13452) );
  nor_x1_sg U49306 ( .A(n31770), .B(n40965), .X(n13451) );
  nor_x1_sg U49307 ( .A(n13463), .B(n13464), .X(n13461) );
  nor_x1_sg U49308 ( .A(n35118), .B(n34275), .X(n13464) );
  nor_x1_sg U49309 ( .A(n34347), .B(n40963), .X(n13463) );
  nor_x1_sg U49310 ( .A(n13469), .B(n13470), .X(n13467) );
  nor_x1_sg U49311 ( .A(n42688), .B(n13367), .X(n13470) );
  nor_x1_sg U49312 ( .A(n30348), .B(n42680), .X(n13469) );
  nor_x1_sg U49313 ( .A(n13481), .B(n13482), .X(n13479) );
  nor_x1_sg U49314 ( .A(n35117), .B(n30320), .X(n13482) );
  nor_x1_sg U49315 ( .A(n34347), .B(n40962), .X(n13481) );
  nor_x1_sg U49316 ( .A(n13494), .B(n13495), .X(n13492) );
  nor_x1_sg U49317 ( .A(n35153), .B(n34277), .X(n13495) );
  nor_x1_sg U49318 ( .A(n31769), .B(n41096), .X(n13494) );
  nor_x1_sg U49319 ( .A(n13511), .B(n13512), .X(n13509) );
  nor_x1_sg U49320 ( .A(n42572), .B(n34277), .X(n13512) );
  nor_x1_sg U49321 ( .A(n29713), .B(n42564), .X(n13511) );
  nor_x1_sg U49322 ( .A(n13522), .B(n13523), .X(n13520) );
  nor_x1_sg U49323 ( .A(n35150), .B(n31798), .X(n13523) );
  nor_x1_sg U49324 ( .A(n34346), .B(n41093), .X(n13522) );
  nor_x1_sg U49325 ( .A(n13528), .B(n13529), .X(n13526) );
  nor_x1_sg U49326 ( .A(n35149), .B(n34276), .X(n13529) );
  nor_x1_sg U49327 ( .A(n30348), .B(n41092), .X(n13528) );
  nor_x1_sg U49328 ( .A(n13540), .B(n13541), .X(n13538) );
  nor_x1_sg U49329 ( .A(n42574), .B(n34274), .X(n13541) );
  nor_x1_sg U49330 ( .A(n31330), .B(n42566), .X(n13540) );
  nor_x1_sg U49331 ( .A(n13546), .B(n13547), .X(n13544) );
  nor_x1_sg U49332 ( .A(n42575), .B(n34275), .X(n13547) );
  nor_x1_sg U49333 ( .A(n34345), .B(n42567), .X(n13546) );
  nor_x1_sg U49334 ( .A(n13558), .B(n13559), .X(n13556) );
  nor_x1_sg U49335 ( .A(n35146), .B(n31798), .X(n13559) );
  nor_x1_sg U49336 ( .A(n31330), .B(n41089), .X(n13558) );
  nor_x1_sg U49337 ( .A(n13564), .B(n13565), .X(n13562) );
  nor_x1_sg U49338 ( .A(n42576), .B(n31797), .X(n13565) );
  nor_x1_sg U49339 ( .A(n31330), .B(n42568), .X(n13564) );
  nor_x1_sg U49340 ( .A(n13576), .B(n13577), .X(n13574) );
  nor_x1_sg U49341 ( .A(n35145), .B(n34276), .X(n13577) );
  nor_x1_sg U49342 ( .A(n34345), .B(n41088), .X(n13576) );
  nor_x1_sg U49343 ( .A(n13582), .B(n13583), .X(n13580) );
  nor_x1_sg U49344 ( .A(n35144), .B(n30090), .X(n13583) );
  nor_x1_sg U49345 ( .A(n31769), .B(n41087), .X(n13582) );
  nor_x1_sg U49346 ( .A(n14752), .B(n41282), .X(n14725) );
  inv_x1_sg U49347 ( .A(n14753), .X(n41282) );
  nor_x1_sg U49348 ( .A(n34418), .B(n41102), .X(n14752) );
  nor_x1_sg U49349 ( .A(n14129), .B(n41270), .X(n14102) );
  inv_x1_sg U49350 ( .A(n14130), .X(n41270) );
  nor_x1_sg U49351 ( .A(n30851), .B(n40979), .X(n14129) );
  nor_x1_sg U49352 ( .A(n14160), .B(n41271), .X(n14133) );
  inv_x1_sg U49353 ( .A(n14161), .X(n41271) );
  nor_x1_sg U49354 ( .A(n30115), .B(n40978), .X(n14160) );
  nor_x1_sg U49355 ( .A(n13818), .B(n41264), .X(n13785) );
  inv_x1_sg U49356 ( .A(n13819), .X(n41264) );
  nor_x1_sg U49357 ( .A(n30115), .B(n40985), .X(n13818) );
  nor_x1_sg U49358 ( .A(n13850), .B(n41265), .X(n13823) );
  inv_x1_sg U49359 ( .A(n13851), .X(n41265) );
  nor_x1_sg U49360 ( .A(n30115), .B(n40984), .X(n13850) );
  nor_x1_sg U49361 ( .A(n13881), .B(n41266), .X(n13854) );
  inv_x1_sg U49362 ( .A(n13882), .X(n41266) );
  nor_x1_sg U49363 ( .A(n34417), .B(n40983), .X(n13881) );
  nor_x1_sg U49364 ( .A(n13912), .B(n13913), .X(n13885) );
  nor_x1_sg U49365 ( .A(n31984), .B(n42658), .X(n13912) );
  nor_x1_sg U49366 ( .A(n32515), .B(n42666), .X(n13913) );
  nor_x1_sg U49367 ( .A(n13943), .B(n13944), .X(n13916) );
  nor_x1_sg U49368 ( .A(n35634), .B(n42659), .X(n13943) );
  nor_x1_sg U49369 ( .A(n32514), .B(n42667), .X(n13944) );
  nor_x1_sg U49370 ( .A(n13974), .B(n41267), .X(n13947) );
  inv_x1_sg U49371 ( .A(n13975), .X(n41267) );
  nor_x1_sg U49372 ( .A(n30850), .B(n40982), .X(n13974) );
  nor_x1_sg U49373 ( .A(n14005), .B(n41268), .X(n13978) );
  inv_x1_sg U49374 ( .A(n14006), .X(n41268) );
  nor_x1_sg U49375 ( .A(n34417), .B(n40981), .X(n14005) );
  nor_x1_sg U49376 ( .A(n14036), .B(n41269), .X(n14009) );
  inv_x1_sg U49377 ( .A(n14037), .X(n41269) );
  nor_x1_sg U49378 ( .A(n34420), .B(n40980), .X(n14036) );
  nor_x1_sg U49379 ( .A(n14067), .B(n14068), .X(n14040) );
  nor_x1_sg U49380 ( .A(n30851), .B(n42660), .X(n14067) );
  nor_x1_sg U49381 ( .A(n32512), .B(n42668), .X(n14068) );
  nor_x1_sg U49382 ( .A(n14098), .B(n14099), .X(n14071) );
  nor_x1_sg U49383 ( .A(n31981), .B(n42661), .X(n14098) );
  nor_x1_sg U49384 ( .A(n32512), .B(n42669), .X(n14099) );
  nor_x1_sg U49385 ( .A(n14315), .B(n41274), .X(n14288) );
  inv_x1_sg U49386 ( .A(n14316), .X(n41274) );
  nor_x1_sg U49387 ( .A(n34418), .B(n40975), .X(n14315) );
  nor_x1_sg U49388 ( .A(n14346), .B(n14347), .X(n14319) );
  nor_x1_sg U49389 ( .A(n34417), .B(n42664), .X(n14346) );
  nor_x1_sg U49390 ( .A(n32514), .B(n42672), .X(n14347) );
  nor_x1_sg U49391 ( .A(n14377), .B(n14378), .X(n14350) );
  nor_x1_sg U49392 ( .A(n30115), .B(n42665), .X(n14377) );
  nor_x1_sg U49393 ( .A(n32515), .B(n42673), .X(n14378) );
  nor_x1_sg U49394 ( .A(n14408), .B(n41275), .X(n14381) );
  inv_x1_sg U49395 ( .A(n14409), .X(n41275) );
  nor_x1_sg U49396 ( .A(n34419), .B(n40974), .X(n14408) );
  nor_x1_sg U49397 ( .A(n14440), .B(n41276), .X(n14413) );
  inv_x1_sg U49398 ( .A(n14441), .X(n41276) );
  nor_x1_sg U49399 ( .A(n31981), .B(n41108), .X(n14440) );
  nor_x1_sg U49400 ( .A(n14471), .B(n41277), .X(n14444) );
  inv_x1_sg U49401 ( .A(n14472), .X(n41277) );
  nor_x1_sg U49402 ( .A(n31983), .B(n41107), .X(n14471) );
  nor_x1_sg U49403 ( .A(n14504), .B(n41278), .X(n14475) );
  inv_x1_sg U49404 ( .A(n14505), .X(n41278) );
  nor_x1_sg U49405 ( .A(n30851), .B(n41106), .X(n14504) );
  nor_x1_sg U49406 ( .A(n14535), .B(n14536), .X(n14508) );
  nor_x1_sg U49407 ( .A(n31982), .B(n42548), .X(n14535) );
  nor_x1_sg U49408 ( .A(n32513), .B(n42556), .X(n14536) );
  nor_x1_sg U49409 ( .A(n14597), .B(n41279), .X(n14570) );
  inv_x1_sg U49410 ( .A(n14598), .X(n41279) );
  nor_x1_sg U49411 ( .A(n35634), .B(n41105), .X(n14597) );
  nor_x1_sg U49412 ( .A(n14628), .B(n41280), .X(n14601) );
  inv_x1_sg U49413 ( .A(n14629), .X(n41280) );
  nor_x1_sg U49414 ( .A(n31982), .B(n41104), .X(n14628) );
  nor_x1_sg U49415 ( .A(n14659), .B(n41281), .X(n14632) );
  inv_x1_sg U49416 ( .A(n14660), .X(n41281) );
  nor_x1_sg U49417 ( .A(n31982), .B(n41103), .X(n14659) );
  nor_x1_sg U49418 ( .A(n14690), .B(n14691), .X(n14663) );
  nor_x1_sg U49419 ( .A(n31984), .B(n42550), .X(n14690) );
  nor_x1_sg U49420 ( .A(n32513), .B(n42558), .X(n14691) );
  nor_x1_sg U49421 ( .A(n14721), .B(n14722), .X(n14694) );
  nor_x1_sg U49422 ( .A(n34418), .B(n42551), .X(n14721) );
  nor_x1_sg U49423 ( .A(n32512), .B(n42559), .X(n14722) );
  nor_x1_sg U49424 ( .A(n14783), .B(n41283), .X(n14756) );
  inv_x1_sg U49425 ( .A(n14784), .X(n41283) );
  nor_x1_sg U49426 ( .A(n34419), .B(n41101), .X(n14783) );
  nor_x1_sg U49427 ( .A(n14814), .B(n14815), .X(n14787) );
  nor_x1_sg U49428 ( .A(n34420), .B(n42552), .X(n14814) );
  nor_x1_sg U49429 ( .A(n32512), .B(n42560), .X(n14815) );
  nor_x1_sg U49430 ( .A(n14845), .B(n14846), .X(n14818) );
  nor_x1_sg U49431 ( .A(n34419), .B(n42553), .X(n14845) );
  nor_x1_sg U49432 ( .A(n32514), .B(n42561), .X(n14846) );
  nor_x1_sg U49433 ( .A(n14876), .B(n41284), .X(n14849) );
  inv_x1_sg U49434 ( .A(n14877), .X(n41284) );
  nor_x1_sg U49435 ( .A(n31982), .B(n41100), .X(n14876) );
  nor_x1_sg U49436 ( .A(n14907), .B(n41285), .X(n14880) );
  inv_x1_sg U49437 ( .A(n14908), .X(n41285) );
  nor_x1_sg U49438 ( .A(n34419), .B(n41099), .X(n14907) );
  nor_x1_sg U49439 ( .A(n14938), .B(n41286), .X(n14911) );
  inv_x1_sg U49440 ( .A(n14939), .X(n41286) );
  nor_x1_sg U49441 ( .A(n34418), .B(n41098), .X(n14938) );
  nor_x1_sg U49442 ( .A(n14969), .B(n14970), .X(n14942) );
  nor_x1_sg U49443 ( .A(n31983), .B(n42554), .X(n14969) );
  nor_x1_sg U49444 ( .A(n32513), .B(n42562), .X(n14970) );
  nor_x1_sg U49445 ( .A(n15000), .B(n15001), .X(n14973) );
  nor_x1_sg U49446 ( .A(n31984), .B(n42555), .X(n15000) );
  nor_x1_sg U49447 ( .A(n32514), .B(n42563), .X(n15001) );
  nor_x1_sg U49448 ( .A(n15031), .B(n41287), .X(n15004) );
  inv_x1_sg U49449 ( .A(n15032), .X(n41287) );
  nor_x1_sg U49450 ( .A(n30850), .B(n41097), .X(n15031) );
  nor_x1_sg U49451 ( .A(n14191), .B(n14192), .X(n14164) );
  nor_x1_sg U49452 ( .A(n30850), .B(n42662), .X(n14191) );
  nor_x1_sg U49453 ( .A(n32515), .B(n42670), .X(n14192) );
  nor_x1_sg U49454 ( .A(n14222), .B(n14223), .X(n14195) );
  nor_x1_sg U49455 ( .A(n31983), .B(n42663), .X(n14222) );
  nor_x1_sg U49456 ( .A(n32515), .B(n42671), .X(n14223) );
  nor_x1_sg U49457 ( .A(n14566), .B(n14567), .X(n14539) );
  nor_x1_sg U49458 ( .A(n34417), .B(n42549), .X(n14566) );
  nor_x1_sg U49459 ( .A(n32513), .B(n42557), .X(n14567) );
  nor_x1_sg U49460 ( .A(n14253), .B(n41272), .X(n14226) );
  inv_x1_sg U49461 ( .A(n14254), .X(n41272) );
  nor_x1_sg U49462 ( .A(n34420), .B(n40977), .X(n14253) );
  nor_x1_sg U49463 ( .A(n14284), .B(n41273), .X(n14257) );
  inv_x1_sg U49464 ( .A(n14285), .X(n41273) );
  nor_x1_sg U49465 ( .A(n31981), .B(n40976), .X(n14284) );
  nand_x1_sg U49466 ( .A(n35460), .B(n32001), .X(n15167) );
  nand_x1_sg U49467 ( .A(n34262), .B(n42750), .X(n13911) );
  nand_x1_sg U49468 ( .A(n30311), .B(n42751), .X(n13942) );
  nand_x1_sg U49469 ( .A(n34260), .B(n42752), .X(n14066) );
  nand_x1_sg U49470 ( .A(n31380), .B(n42753), .X(n14097) );
  nand_x1_sg U49471 ( .A(n30313), .B(n42754), .X(n14190) );
  nand_x1_sg U49472 ( .A(n34260), .B(n42755), .X(n14221) );
  nand_x1_sg U49473 ( .A(n31381), .B(n42756), .X(n14345) );
  nand_x1_sg U49474 ( .A(n30313), .B(n42757), .X(n14376) );
  nand_x1_sg U49475 ( .A(n30087), .B(n42637), .X(n14689) );
  nand_x1_sg U49476 ( .A(n31381), .B(n42638), .X(n14720) );
  nand_x1_sg U49477 ( .A(n30311), .B(n42639), .X(n14813) );
  nand_x1_sg U49478 ( .A(n34261), .B(n42640), .X(n14844) );
  nand_x1_sg U49479 ( .A(n34261), .B(n42642), .X(n14937) );
  nand_x1_sg U49480 ( .A(n15068), .B(n15070), .X(n15069) );
  nand_x1_sg U49481 ( .A(n15204), .B(n15206), .X(n15205) );
  nor_x1_sg U49482 ( .A(n12614), .B(n12615), .X(n12612) );
  nor_x1_sg U49483 ( .A(n12616), .B(n31882), .X(n12615) );
  nand_x1_sg U49484 ( .A(n12705), .B(n12613), .X(n12704) );
  nor_x1_sg U49485 ( .A(n12706), .B(n12707), .X(n12705) );
  nor_x1_sg U49486 ( .A(n12708), .B(n32004), .X(n12707) );
  inv_x1_sg U49487 ( .A(n11567), .X(n41167) );
  inv_x1_sg U49488 ( .A(n11581), .X(n41181) );
  inv_x1_sg U49489 ( .A(n11537), .X(n41143) );
  inv_x1_sg U49490 ( .A(n11538), .X(n41144) );
  inv_x1_sg U49491 ( .A(n11541), .X(n41147) );
  inv_x1_sg U49492 ( .A(n11544), .X(n41150) );
  inv_x1_sg U49493 ( .A(n11547), .X(n41153) );
  inv_x1_sg U49494 ( .A(n11550), .X(n41156) );
  inv_x1_sg U49495 ( .A(n11551), .X(n41157) );
  inv_x1_sg U49496 ( .A(n11552), .X(n41158) );
  inv_x1_sg U49497 ( .A(n11555), .X(n41161) );
  inv_x1_sg U49498 ( .A(n11556), .X(n41162) );
  inv_x1_sg U49499 ( .A(n11563), .X(n41163) );
  inv_x1_sg U49500 ( .A(n11564), .X(n41164) );
  inv_x1_sg U49501 ( .A(n11570), .X(n41170) );
  inv_x1_sg U49502 ( .A(n11573), .X(n41173) );
  inv_x1_sg U49503 ( .A(n11576), .X(n41176) );
  inv_x1_sg U49504 ( .A(n11577), .X(n41177) );
  inv_x1_sg U49505 ( .A(n11578), .X(n41178) );
  inv_x1_sg U49506 ( .A(n11582), .X(n41182) );
  inv_x1_sg U49507 ( .A(n11565), .X(n41165) );
  inv_x1_sg U49508 ( .A(n11580), .X(n41180) );
  inv_x1_sg U49509 ( .A(n11539), .X(n41145) );
  inv_x1_sg U49510 ( .A(n11540), .X(n41146) );
  inv_x1_sg U49511 ( .A(n11542), .X(n41148) );
  inv_x1_sg U49512 ( .A(n11543), .X(n41149) );
  inv_x1_sg U49513 ( .A(n11545), .X(n41151) );
  inv_x1_sg U49514 ( .A(n11546), .X(n41152) );
  inv_x1_sg U49515 ( .A(n11548), .X(n41154) );
  inv_x1_sg U49516 ( .A(n11549), .X(n41155) );
  inv_x1_sg U49517 ( .A(n11553), .X(n41159) );
  inv_x1_sg U49518 ( .A(n11554), .X(n41160) );
  inv_x1_sg U49519 ( .A(n11566), .X(n41166) );
  inv_x1_sg U49520 ( .A(n11568), .X(n41168) );
  inv_x1_sg U49521 ( .A(n11569), .X(n41169) );
  inv_x1_sg U49522 ( .A(n11571), .X(n41171) );
  inv_x1_sg U49523 ( .A(n11572), .X(n41172) );
  inv_x1_sg U49524 ( .A(n11574), .X(n41174) );
  inv_x1_sg U49525 ( .A(n11575), .X(n41175) );
  inv_x1_sg U49526 ( .A(n11579), .X(n41179) );
  inv_x1_sg U49527 ( .A(n11618), .X(n41208) );
  inv_x1_sg U49528 ( .A(n11632), .X(n41222) );
  inv_x1_sg U49529 ( .A(n11587), .X(n41184) );
  inv_x1_sg U49530 ( .A(n11588), .X(n41185) );
  inv_x1_sg U49531 ( .A(n11591), .X(n41188) );
  inv_x1_sg U49532 ( .A(n11594), .X(n41191) );
  inv_x1_sg U49533 ( .A(n11597), .X(n41194) );
  inv_x1_sg U49534 ( .A(n11600), .X(n41197) );
  inv_x1_sg U49535 ( .A(n11601), .X(n41198) );
  inv_x1_sg U49536 ( .A(n11602), .X(n41199) );
  inv_x1_sg U49537 ( .A(n11605), .X(n41202) );
  inv_x1_sg U49538 ( .A(n11606), .X(n41203) );
  inv_x1_sg U49539 ( .A(n11614), .X(n41204) );
  inv_x1_sg U49540 ( .A(n11615), .X(n41205) );
  inv_x1_sg U49541 ( .A(n11616), .X(n41206) );
  inv_x1_sg U49542 ( .A(n11621), .X(n41211) );
  inv_x1_sg U49543 ( .A(n11624), .X(n41214) );
  inv_x1_sg U49544 ( .A(n11627), .X(n41217) );
  inv_x1_sg U49545 ( .A(n11628), .X(n41218) );
  inv_x1_sg U49546 ( .A(n11629), .X(n41219) );
  inv_x1_sg U49547 ( .A(n11631), .X(n41221) );
  inv_x1_sg U49548 ( .A(n11633), .X(n41223) );
  inv_x1_sg U49549 ( .A(n11589), .X(n41186) );
  inv_x1_sg U49550 ( .A(n11590), .X(n41187) );
  inv_x1_sg U49551 ( .A(n11592), .X(n41189) );
  inv_x1_sg U49552 ( .A(n11593), .X(n41190) );
  inv_x1_sg U49553 ( .A(n11595), .X(n41192) );
  inv_x1_sg U49554 ( .A(n11596), .X(n41193) );
  inv_x1_sg U49555 ( .A(n11598), .X(n41195) );
  inv_x1_sg U49556 ( .A(n11599), .X(n41196) );
  inv_x1_sg U49557 ( .A(n11603), .X(n41200) );
  inv_x1_sg U49558 ( .A(n11604), .X(n41201) );
  inv_x1_sg U49559 ( .A(n11617), .X(n41207) );
  inv_x1_sg U49560 ( .A(n11619), .X(n41209) );
  inv_x1_sg U49561 ( .A(n11620), .X(n41210) );
  inv_x1_sg U49562 ( .A(n11622), .X(n41212) );
  inv_x1_sg U49563 ( .A(n11623), .X(n41213) );
  inv_x1_sg U49564 ( .A(n11625), .X(n41215) );
  inv_x1_sg U49565 ( .A(n11626), .X(n41216) );
  inv_x1_sg U49566 ( .A(n11630), .X(n41220) );
  inv_x1_sg U49567 ( .A(n11642), .X(n41224) );
  inv_x1_sg U49568 ( .A(n11643), .X(n41225) );
  inv_x1_sg U49569 ( .A(n11644), .X(n41226) );
  inv_x1_sg U49570 ( .A(n11645), .X(n41227) );
  inv_x1_sg U49571 ( .A(n11646), .X(n41228) );
  inv_x1_sg U49572 ( .A(n11647), .X(n41229) );
  inv_x1_sg U49573 ( .A(n11648), .X(n41230) );
  inv_x1_sg U49574 ( .A(n11649), .X(n41231) );
  inv_x1_sg U49575 ( .A(n11650), .X(n41232) );
  inv_x1_sg U49576 ( .A(n11651), .X(n41233) );
  inv_x1_sg U49577 ( .A(n11652), .X(n41234) );
  inv_x1_sg U49578 ( .A(n11653), .X(n41235) );
  inv_x1_sg U49579 ( .A(n11654), .X(n41236) );
  inv_x1_sg U49580 ( .A(n11655), .X(n41237) );
  inv_x1_sg U49581 ( .A(n11656), .X(n41238) );
  inv_x1_sg U49582 ( .A(n11657), .X(n41239) );
  inv_x1_sg U49583 ( .A(n11658), .X(n41240) );
  inv_x1_sg U49584 ( .A(n11659), .X(n41241) );
  inv_x1_sg U49585 ( .A(n11660), .X(n41242) );
  inv_x1_sg U49586 ( .A(n11661), .X(n41243) );
  inv_x1_sg U49587 ( .A(n11668), .X(n41244) );
  inv_x1_sg U49588 ( .A(n11669), .X(n41245) );
  inv_x1_sg U49589 ( .A(n11670), .X(n41246) );
  inv_x1_sg U49590 ( .A(n11671), .X(n41247) );
  inv_x1_sg U49591 ( .A(n11672), .X(n41248) );
  inv_x1_sg U49592 ( .A(n11673), .X(n41249) );
  inv_x1_sg U49593 ( .A(n11674), .X(n41250) );
  inv_x1_sg U49594 ( .A(n11675), .X(n41251) );
  inv_x1_sg U49595 ( .A(n11676), .X(n41252) );
  inv_x1_sg U49596 ( .A(n11677), .X(n41253) );
  inv_x1_sg U49597 ( .A(n11678), .X(n41254) );
  inv_x1_sg U49598 ( .A(n11679), .X(n41255) );
  inv_x1_sg U49599 ( .A(n11680), .X(n41256) );
  inv_x1_sg U49600 ( .A(n11681), .X(n41257) );
  inv_x1_sg U49601 ( .A(n11682), .X(n41258) );
  inv_x1_sg U49602 ( .A(n11683), .X(n41259) );
  inv_x1_sg U49603 ( .A(n11684), .X(n41260) );
  inv_x1_sg U49604 ( .A(n11685), .X(n41261) );
  inv_x1_sg U49605 ( .A(n11686), .X(n41262) );
  inv_x1_sg U49606 ( .A(n11687), .X(n41263) );
  inv_x1_sg U49607 ( .A(n11690), .X(n41419) );
  inv_x1_sg U49608 ( .A(n11691), .X(n41420) );
  inv_x1_sg U49609 ( .A(n11692), .X(n41421) );
  inv_x1_sg U49610 ( .A(n11693), .X(n41422) );
  inv_x1_sg U49611 ( .A(n11694), .X(n41423) );
  inv_x1_sg U49612 ( .A(n11695), .X(n41424) );
  inv_x1_sg U49613 ( .A(n11696), .X(n41425) );
  inv_x1_sg U49614 ( .A(n11697), .X(n41426) );
  inv_x1_sg U49615 ( .A(n11698), .X(n41427) );
  inv_x1_sg U49616 ( .A(n11699), .X(n41428) );
  inv_x1_sg U49617 ( .A(n11700), .X(n41429) );
  inv_x1_sg U49618 ( .A(n11701), .X(n41430) );
  inv_x1_sg U49619 ( .A(n11702), .X(n41431) );
  inv_x1_sg U49620 ( .A(n11703), .X(n41432) );
  inv_x1_sg U49621 ( .A(n11704), .X(n41433) );
  inv_x1_sg U49622 ( .A(n11705), .X(n41434) );
  inv_x1_sg U49623 ( .A(n11706), .X(n41435) );
  inv_x1_sg U49624 ( .A(n11707), .X(n41436) );
  inv_x1_sg U49625 ( .A(n11708), .X(n41437) );
  inv_x1_sg U49626 ( .A(n11709), .X(n41438) );
  inv_x1_sg U49627 ( .A(n11717), .X(n41439) );
  inv_x1_sg U49628 ( .A(n11718), .X(n41440) );
  inv_x1_sg U49629 ( .A(n11719), .X(n41441) );
  inv_x1_sg U49630 ( .A(n11720), .X(n41442) );
  inv_x1_sg U49631 ( .A(n11721), .X(n41443) );
  inv_x1_sg U49632 ( .A(n11722), .X(n41444) );
  inv_x1_sg U49633 ( .A(n11723), .X(n41445) );
  inv_x1_sg U49634 ( .A(n11724), .X(n41446) );
  inv_x1_sg U49635 ( .A(n11725), .X(n41447) );
  inv_x1_sg U49636 ( .A(n11726), .X(n41448) );
  inv_x1_sg U49637 ( .A(n11727), .X(n41449) );
  inv_x1_sg U49638 ( .A(n11728), .X(n41450) );
  inv_x1_sg U49639 ( .A(n11729), .X(n41451) );
  inv_x1_sg U49640 ( .A(n11730), .X(n41452) );
  inv_x1_sg U49641 ( .A(n11731), .X(n41453) );
  inv_x1_sg U49642 ( .A(n11732), .X(n41454) );
  inv_x1_sg U49643 ( .A(n11733), .X(n41455) );
  inv_x1_sg U49644 ( .A(n11734), .X(n41456) );
  inv_x1_sg U49645 ( .A(n11735), .X(n41457) );
  inv_x1_sg U49646 ( .A(n11736), .X(n41458) );
  inv_x1_sg U49647 ( .A(n11743), .X(n41459) );
  inv_x1_sg U49648 ( .A(n11744), .X(n41460) );
  inv_x1_sg U49649 ( .A(n11745), .X(n41461) );
  inv_x1_sg U49650 ( .A(n11746), .X(n41462) );
  inv_x1_sg U49651 ( .A(n11747), .X(n41463) );
  inv_x1_sg U49652 ( .A(n11748), .X(n41464) );
  inv_x1_sg U49653 ( .A(n11749), .X(n41465) );
  inv_x1_sg U49654 ( .A(n11750), .X(n41466) );
  inv_x1_sg U49655 ( .A(n11751), .X(n41467) );
  inv_x1_sg U49656 ( .A(n11752), .X(n41468) );
  inv_x1_sg U49657 ( .A(n11753), .X(n41469) );
  inv_x1_sg U49658 ( .A(n11754), .X(n41470) );
  inv_x1_sg U49659 ( .A(n11755), .X(n41471) );
  inv_x1_sg U49660 ( .A(n11756), .X(n41472) );
  inv_x1_sg U49661 ( .A(n11757), .X(n41473) );
  inv_x1_sg U49662 ( .A(n11758), .X(n41474) );
  inv_x1_sg U49663 ( .A(n11759), .X(n41475) );
  inv_x1_sg U49664 ( .A(n11760), .X(n41476) );
  inv_x1_sg U49665 ( .A(n11761), .X(n41477) );
  inv_x1_sg U49666 ( .A(n11762), .X(n41478) );
  inv_x1_sg U49667 ( .A(n11771), .X(n41479) );
  inv_x1_sg U49668 ( .A(n11772), .X(n41480) );
  inv_x1_sg U49669 ( .A(n11773), .X(n41481) );
  inv_x1_sg U49670 ( .A(n11774), .X(n41482) );
  inv_x1_sg U49671 ( .A(n11775), .X(n41483) );
  inv_x1_sg U49672 ( .A(n11776), .X(n41484) );
  inv_x1_sg U49673 ( .A(n11777), .X(n41485) );
  inv_x1_sg U49674 ( .A(n11778), .X(n41486) );
  inv_x1_sg U49675 ( .A(n11779), .X(n41487) );
  inv_x1_sg U49676 ( .A(n11780), .X(n41488) );
  inv_x1_sg U49677 ( .A(n11781), .X(n41489) );
  inv_x1_sg U49678 ( .A(n11782), .X(n41490) );
  inv_x1_sg U49679 ( .A(n11783), .X(n41491) );
  inv_x1_sg U49680 ( .A(n11784), .X(n41492) );
  inv_x1_sg U49681 ( .A(n11785), .X(n41493) );
  inv_x1_sg U49682 ( .A(n11786), .X(n41494) );
  inv_x1_sg U49683 ( .A(n11787), .X(n41495) );
  inv_x1_sg U49684 ( .A(n11788), .X(n41496) );
  inv_x1_sg U49685 ( .A(n11789), .X(n41497) );
  inv_x1_sg U49686 ( .A(n11790), .X(n41498) );
  nand_x1_sg U49687 ( .A(n30287), .B(n42724), .X(n14059) );
  nor_x1_sg U49688 ( .A(n14060), .B(n14061), .X(n14058) );
  nand_x1_sg U49689 ( .A(n30285), .B(n42725), .X(n14090) );
  nor_x1_sg U49690 ( .A(n14091), .B(n14092), .X(n14089) );
  nand_x1_sg U49691 ( .A(n31414), .B(n42726), .X(n14183) );
  nor_x1_sg U49692 ( .A(n14184), .B(n14185), .X(n14182) );
  nand_x1_sg U49693 ( .A(n34204), .B(n42727), .X(n14214) );
  nor_x1_sg U49694 ( .A(n14215), .B(n14216), .X(n14213) );
  nor_x1_sg U49695 ( .A(n33036), .B(n13703), .X(\shifter_0/n6713 ) );
  nor_x1_sg U49696 ( .A(n29998), .B(n13707), .X(\shifter_0/n6709 ) );
  nor_x1_sg U49697 ( .A(n33033), .B(n13711), .X(\shifter_0/n6705 ) );
  nor_x1_sg U49698 ( .A(n33035), .B(n13714), .X(\shifter_0/n6701 ) );
  nor_x1_sg U49699 ( .A(n33034), .B(n13718), .X(\shifter_0/n6697 ) );
  nor_x1_sg U49700 ( .A(n33036), .B(n13721), .X(\shifter_0/n6693 ) );
  nor_x1_sg U49701 ( .A(n33034), .B(n13725), .X(\shifter_0/n6689 ) );
  nor_x1_sg U49702 ( .A(n33033), .B(n13729), .X(\shifter_0/n6685 ) );
  nor_x1_sg U49703 ( .A(n33034), .B(n13733), .X(\shifter_0/n6681 ) );
  nor_x1_sg U49704 ( .A(n33035), .B(n13737), .X(\shifter_0/n6677 ) );
  nor_x1_sg U49705 ( .A(n33034), .B(n13741), .X(\shifter_0/n6673 ) );
  nor_x1_sg U49706 ( .A(n29998), .B(n13745), .X(\shifter_0/n6669 ) );
  nor_x1_sg U49707 ( .A(n33035), .B(n13749), .X(\shifter_0/n6665 ) );
  nor_x1_sg U49708 ( .A(n33033), .B(n13753), .X(\shifter_0/n6661 ) );
  nor_x1_sg U49709 ( .A(n35241), .B(n13757), .X(\shifter_0/n6657 ) );
  nor_x1_sg U49710 ( .A(n33033), .B(n13761), .X(\shifter_0/n6653 ) );
  nor_x1_sg U49711 ( .A(n35241), .B(n13765), .X(\shifter_0/n6649 ) );
  nor_x1_sg U49712 ( .A(n33036), .B(n13769), .X(\shifter_0/n6645 ) );
  nor_x1_sg U49713 ( .A(n33036), .B(n13772), .X(\shifter_0/n6641 ) );
  nor_x1_sg U49714 ( .A(n33035), .B(n13775), .X(\shifter_0/n6637 ) );
  nor_x1_sg U49715 ( .A(n33014), .B(n13616), .X(\shifter_0/n6793 ) );
  nor_x1_sg U49716 ( .A(n30002), .B(n13621), .X(\shifter_0/n6789 ) );
  nor_x1_sg U49717 ( .A(n33015), .B(n13625), .X(\shifter_0/n6785 ) );
  nor_x1_sg U49718 ( .A(n33013), .B(n13629), .X(\shifter_0/n6781 ) );
  nor_x1_sg U49719 ( .A(n33016), .B(n13633), .X(\shifter_0/n6777 ) );
  nor_x1_sg U49720 ( .A(n33014), .B(n13637), .X(\shifter_0/n6773 ) );
  nor_x1_sg U49721 ( .A(n33014), .B(n13641), .X(\shifter_0/n6769 ) );
  nor_x1_sg U49722 ( .A(n33015), .B(n13645), .X(\shifter_0/n6765 ) );
  nor_x1_sg U49723 ( .A(n33015), .B(n13649), .X(\shifter_0/n6761 ) );
  nor_x1_sg U49724 ( .A(n30002), .B(n13653), .X(\shifter_0/n6757 ) );
  nor_x1_sg U49725 ( .A(n33016), .B(n13657), .X(\shifter_0/n6753 ) );
  nor_x1_sg U49726 ( .A(n33016), .B(n13661), .X(\shifter_0/n6749 ) );
  nor_x1_sg U49727 ( .A(n33016), .B(n13665), .X(\shifter_0/n6745 ) );
  nor_x1_sg U49728 ( .A(n33013), .B(n13669), .X(\shifter_0/n6741 ) );
  nor_x1_sg U49729 ( .A(n35245), .B(n13673), .X(\shifter_0/n6737 ) );
  nor_x1_sg U49730 ( .A(n33013), .B(n13677), .X(\shifter_0/n6733 ) );
  nor_x1_sg U49731 ( .A(n35245), .B(n13681), .X(\shifter_0/n6729 ) );
  nor_x1_sg U49732 ( .A(n33015), .B(n13685), .X(\shifter_0/n6725 ) );
  nor_x1_sg U49733 ( .A(n33014), .B(n13689), .X(\shifter_0/n6721 ) );
  nor_x1_sg U49734 ( .A(n33013), .B(n13693), .X(\shifter_0/n6717 ) );
  nor_x1_sg U49735 ( .A(n30000), .B(n13228), .X(\shifter_0/n7113 ) );
  nor_x1_sg U49736 ( .A(n33023), .B(n13231), .X(\shifter_0/n7109 ) );
  nor_x1_sg U49737 ( .A(n35243), .B(n13234), .X(\shifter_0/n7105 ) );
  nor_x1_sg U49738 ( .A(n33025), .B(n13237), .X(\shifter_0/n7101 ) );
  nor_x1_sg U49739 ( .A(n33026), .B(n13240), .X(\shifter_0/n7097 ) );
  nor_x1_sg U49740 ( .A(n33024), .B(n13243), .X(\shifter_0/n7093 ) );
  nor_x1_sg U49741 ( .A(n33026), .B(n13246), .X(\shifter_0/n7089 ) );
  nor_x1_sg U49742 ( .A(n33026), .B(n13249), .X(\shifter_0/n7085 ) );
  nor_x1_sg U49743 ( .A(n33026), .B(n13252), .X(\shifter_0/n7081 ) );
  nor_x1_sg U49744 ( .A(n33025), .B(n13255), .X(\shifter_0/n7077 ) );
  nor_x1_sg U49745 ( .A(n33023), .B(n13258), .X(\shifter_0/n7073 ) );
  nor_x1_sg U49746 ( .A(n30000), .B(n13261), .X(\shifter_0/n7069 ) );
  nor_x1_sg U49747 ( .A(n33024), .B(n13264), .X(\shifter_0/n7065 ) );
  nor_x1_sg U49748 ( .A(n33023), .B(n13267), .X(\shifter_0/n7061 ) );
  nor_x1_sg U49749 ( .A(n33023), .B(n13270), .X(\shifter_0/n7057 ) );
  nor_x1_sg U49750 ( .A(n33024), .B(n13273), .X(\shifter_0/n7053 ) );
  nor_x1_sg U49751 ( .A(n35243), .B(n13276), .X(\shifter_0/n7049 ) );
  nor_x1_sg U49752 ( .A(n33024), .B(n13279), .X(\shifter_0/n7045 ) );
  nor_x1_sg U49753 ( .A(n33025), .B(n13282), .X(\shifter_0/n7041 ) );
  nor_x1_sg U49754 ( .A(n33025), .B(n13285), .X(\shifter_0/n7037 ) );
  nor_x1_sg U49755 ( .A(n32999), .B(n13294), .X(\shifter_0/n7033 ) );
  nor_x1_sg U49756 ( .A(n33000), .B(n13297), .X(\shifter_0/n7029 ) );
  nor_x1_sg U49757 ( .A(n32999), .B(n13300), .X(\shifter_0/n7025 ) );
  nor_x1_sg U49758 ( .A(n33000), .B(n13304), .X(\shifter_0/n7021 ) );
  nor_x1_sg U49759 ( .A(n32998), .B(n13307), .X(\shifter_0/n7017 ) );
  nor_x1_sg U49760 ( .A(n33000), .B(n13311), .X(\shifter_0/n7013 ) );
  nor_x1_sg U49761 ( .A(n35406), .B(n13314), .X(\shifter_0/n7009 ) );
  nor_x1_sg U49762 ( .A(n29992), .B(n13317), .X(\shifter_0/n7005 ) );
  nor_x1_sg U49763 ( .A(n32999), .B(n13320), .X(\shifter_0/n7001 ) );
  nor_x1_sg U49764 ( .A(n32998), .B(n13323), .X(\shifter_0/n6997 ) );
  nor_x1_sg U49765 ( .A(n33000), .B(n13326), .X(\shifter_0/n6993 ) );
  nor_x1_sg U49766 ( .A(n32998), .B(n13329), .X(\shifter_0/n6989 ) );
  nor_x1_sg U49767 ( .A(n29992), .B(n13332), .X(\shifter_0/n6985 ) );
  nor_x1_sg U49768 ( .A(n35406), .B(n13335), .X(\shifter_0/n6981 ) );
  nor_x1_sg U49769 ( .A(n33001), .B(n13338), .X(\shifter_0/n6977 ) );
  nor_x1_sg U49770 ( .A(n33001), .B(n13341), .X(\shifter_0/n6973 ) );
  nor_x1_sg U49771 ( .A(n32999), .B(n13344), .X(\shifter_0/n6969 ) );
  nor_x1_sg U49772 ( .A(n32998), .B(n13347), .X(\shifter_0/n6965 ) );
  nor_x1_sg U49773 ( .A(n33001), .B(n13351), .X(\shifter_0/n6961 ) );
  nor_x1_sg U49774 ( .A(n33001), .B(n13355), .X(\shifter_0/n6957 ) );
  nand_x1_sg U49775 ( .A(n13301), .B(n14477), .X(n14476) );
  nand_x1_sg U49776 ( .A(n31404), .B(n14478), .X(n14477) );
  nor_x1_sg U49777 ( .A(n14479), .B(n14480), .X(n14478) );
  nand_x1_sg U49778 ( .A(n13308), .B(n14541), .X(n14540) );
  nand_x1_sg U49779 ( .A(n34221), .B(n14542), .X(n14541) );
  nor_x1_sg U49780 ( .A(n14543), .B(n14544), .X(n14542) );
  nand_x1_sg U49781 ( .A(n13348), .B(n14944), .X(n14943) );
  nand_x1_sg U49782 ( .A(n34222), .B(n14945), .X(n14944) );
  nor_x1_sg U49783 ( .A(n14946), .B(n14947), .X(n14945) );
  nand_x1_sg U49784 ( .A(n13352), .B(n14975), .X(n14974) );
  nand_x1_sg U49785 ( .A(n34221), .B(n14976), .X(n14975) );
  nor_x1_sg U49786 ( .A(n14977), .B(n14978), .X(n14976) );
  nor_x1_sg U49787 ( .A(n33039), .B(n11800), .X(\shifter_0/n8073 ) );
  nor_x1_sg U49788 ( .A(n33753), .B(n11803), .X(\shifter_0/n8069 ) );
  nor_x1_sg U49789 ( .A(n33038), .B(n11805), .X(\shifter_0/n8065 ) );
  nor_x1_sg U49790 ( .A(n33040), .B(n11807), .X(\shifter_0/n8061 ) );
  nor_x1_sg U49791 ( .A(n33040), .B(n11809), .X(\shifter_0/n8057 ) );
  nor_x1_sg U49792 ( .A(n33038), .B(n11811), .X(\shifter_0/n8053 ) );
  nor_x1_sg U49793 ( .A(n33040), .B(n11813), .X(\shifter_0/n8049 ) );
  nor_x1_sg U49794 ( .A(n35409), .B(n11815), .X(\shifter_0/n8045 ) );
  nor_x1_sg U49795 ( .A(n33039), .B(n11817), .X(\shifter_0/n8041 ) );
  nor_x1_sg U49796 ( .A(n33039), .B(n11819), .X(\shifter_0/n8037 ) );
  nor_x1_sg U49797 ( .A(n30008), .B(n11821), .X(\shifter_0/n8033 ) );
  nor_x1_sg U49798 ( .A(n33040), .B(n11823), .X(\shifter_0/n8029 ) );
  nor_x1_sg U49799 ( .A(n30009), .B(n11825), .X(\shifter_0/n8025 ) );
  nor_x1_sg U49800 ( .A(n30009), .B(n11827), .X(\shifter_0/n8021 ) );
  nor_x1_sg U49801 ( .A(n33039), .B(n11829), .X(\shifter_0/n8017 ) );
  nor_x1_sg U49802 ( .A(n35409), .B(n11831), .X(\shifter_0/n8013 ) );
  nor_x1_sg U49803 ( .A(n35409), .B(n11833), .X(\shifter_0/n8009 ) );
  nor_x1_sg U49804 ( .A(n33038), .B(n11835), .X(\shifter_0/n8005 ) );
  nor_x1_sg U49805 ( .A(n33038), .B(n11837), .X(\shifter_0/n8001 ) );
  nor_x1_sg U49806 ( .A(n30008), .B(n11839), .X(\shifter_0/n7997 ) );
  nor_x1_sg U49807 ( .A(n33011), .B(n11848), .X(\shifter_0/n7993 ) );
  nor_x1_sg U49808 ( .A(n33009), .B(n11851), .X(\shifter_0/n7989 ) );
  nor_x1_sg U49809 ( .A(n35246), .B(n11853), .X(\shifter_0/n7985 ) );
  nor_x1_sg U49810 ( .A(n33008), .B(n11855), .X(\shifter_0/n7981 ) );
  nor_x1_sg U49811 ( .A(n33009), .B(n11857), .X(\shifter_0/n7977 ) );
  nor_x1_sg U49812 ( .A(n30006), .B(n11859), .X(\shifter_0/n7973 ) );
  nor_x1_sg U49813 ( .A(n30006), .B(n11861), .X(\shifter_0/n7969 ) );
  nor_x1_sg U49814 ( .A(n33010), .B(n11863), .X(\shifter_0/n7965 ) );
  nor_x1_sg U49815 ( .A(n33011), .B(n11865), .X(\shifter_0/n7961 ) );
  nor_x1_sg U49816 ( .A(n33008), .B(n11867), .X(\shifter_0/n7957 ) );
  nor_x1_sg U49817 ( .A(n33010), .B(n11869), .X(\shifter_0/n7953 ) );
  nor_x1_sg U49818 ( .A(n33010), .B(n11871), .X(\shifter_0/n7949 ) );
  nor_x1_sg U49819 ( .A(n35246), .B(n11873), .X(\shifter_0/n7945 ) );
  nor_x1_sg U49820 ( .A(n33011), .B(n11875), .X(\shifter_0/n7941 ) );
  nor_x1_sg U49821 ( .A(n33009), .B(n11877), .X(\shifter_0/n7937 ) );
  nor_x1_sg U49822 ( .A(n33008), .B(n11879), .X(\shifter_0/n7933 ) );
  nor_x1_sg U49823 ( .A(n33011), .B(n11881), .X(\shifter_0/n7929 ) );
  nor_x1_sg U49824 ( .A(n33008), .B(n11883), .X(\shifter_0/n7925 ) );
  nor_x1_sg U49825 ( .A(n33009), .B(n11885), .X(\shifter_0/n7921 ) );
  nor_x1_sg U49826 ( .A(n33010), .B(n11887), .X(\shifter_0/n7917 ) );
  nor_x1_sg U49827 ( .A(n35614), .B(n12974), .X(\shifter_0/n7273 ) );
  nor_x1_sg U49828 ( .A(n12975), .B(n33288), .X(n12974) );
  nor_x1_sg U49829 ( .A(n33802), .B(n12972), .X(n12975) );
  nor_x1_sg U49830 ( .A(n35561), .B(n12981), .X(\shifter_0/n7269 ) );
  nor_x1_sg U49831 ( .A(n12982), .B(n33288), .X(n12981) );
  nor_x1_sg U49832 ( .A(n30985), .B(n12980), .X(n12982) );
  nor_x1_sg U49833 ( .A(n35613), .B(n12987), .X(\shifter_0/n7265 ) );
  nor_x1_sg U49834 ( .A(n12988), .B(n33288), .X(n12987) );
  nor_x1_sg U49835 ( .A(n30986), .B(n12986), .X(n12988) );
  nor_x1_sg U49836 ( .A(n35509), .B(n12993), .X(\shifter_0/n7261 ) );
  nor_x1_sg U49837 ( .A(n12994), .B(n29913), .X(n12993) );
  nor_x1_sg U49838 ( .A(n30986), .B(n12992), .X(n12994) );
  nor_x1_sg U49839 ( .A(n35604), .B(n12999), .X(\shifter_0/n7257 ) );
  nor_x1_sg U49840 ( .A(n13000), .B(n33287), .X(n12999) );
  nor_x1_sg U49841 ( .A(n33758), .B(n12998), .X(n13000) );
  nor_x1_sg U49842 ( .A(n35619), .B(n13005), .X(\shifter_0/n7253 ) );
  nor_x1_sg U49843 ( .A(n13006), .B(n33285), .X(n13005) );
  nor_x1_sg U49844 ( .A(n33802), .B(n13004), .X(n13006) );
  nor_x1_sg U49845 ( .A(n35514), .B(n13011), .X(\shifter_0/n7249 ) );
  nor_x1_sg U49846 ( .A(n13012), .B(n33285), .X(n13011) );
  nor_x1_sg U49847 ( .A(n35410), .B(n13010), .X(n13012) );
  nor_x1_sg U49848 ( .A(n35618), .B(n13017), .X(\shifter_0/n7245 ) );
  nor_x1_sg U49849 ( .A(n13018), .B(n29913), .X(n13017) );
  nor_x1_sg U49850 ( .A(n33802), .B(n13016), .X(n13018) );
  nor_x1_sg U49851 ( .A(n35612), .B(n13023), .X(\shifter_0/n7241 ) );
  nor_x1_sg U49852 ( .A(n13024), .B(n29913), .X(n13023) );
  nor_x1_sg U49853 ( .A(n33800), .B(n13022), .X(n13024) );
  nor_x1_sg U49854 ( .A(n35617), .B(n13029), .X(\shifter_0/n7237 ) );
  nor_x1_sg U49855 ( .A(n13030), .B(n33286), .X(n13029) );
  nor_x1_sg U49856 ( .A(n33800), .B(n13028), .X(n13030) );
  nor_x1_sg U49857 ( .A(n35602), .B(n13035), .X(\shifter_0/n7233 ) );
  nor_x1_sg U49858 ( .A(n13036), .B(n33288), .X(n13035) );
  nor_x1_sg U49859 ( .A(n33801), .B(n13034), .X(n13036) );
  nor_x1_sg U49860 ( .A(n35616), .B(n13041), .X(\shifter_0/n7229 ) );
  nor_x1_sg U49861 ( .A(n13042), .B(n33287), .X(n13041) );
  nor_x1_sg U49862 ( .A(n35410), .B(n13040), .X(n13042) );
  nor_x1_sg U49863 ( .A(n35611), .B(n13047), .X(\shifter_0/n7225 ) );
  nor_x1_sg U49864 ( .A(n13048), .B(n33285), .X(n13047) );
  nor_x1_sg U49865 ( .A(n33800), .B(n13046), .X(n13048) );
  nor_x1_sg U49866 ( .A(n35615), .B(n13053), .X(\shifter_0/n7221 ) );
  nor_x1_sg U49867 ( .A(n13054), .B(n33286), .X(n13053) );
  nor_x1_sg U49868 ( .A(n33801), .B(n13052), .X(n13054) );
  nor_x1_sg U49869 ( .A(n35610), .B(n13059), .X(\shifter_0/n7217 ) );
  nor_x1_sg U49870 ( .A(n13060), .B(n33286), .X(n13059) );
  nor_x1_sg U49871 ( .A(n30986), .B(n13058), .X(n13060) );
  nor_x1_sg U49872 ( .A(n35609), .B(n13065), .X(\shifter_0/n7213 ) );
  nor_x1_sg U49873 ( .A(n13066), .B(n33287), .X(n13065) );
  nor_x1_sg U49874 ( .A(n33800), .B(n13064), .X(n13066) );
  nor_x1_sg U49875 ( .A(n35601), .B(n13071), .X(\shifter_0/n7209 ) );
  nor_x1_sg U49876 ( .A(n13072), .B(n29913), .X(n13071) );
  nor_x1_sg U49877 ( .A(n33801), .B(n13070), .X(n13072) );
  nor_x1_sg U49878 ( .A(n35608), .B(n13077), .X(\shifter_0/n7205 ) );
  nor_x1_sg U49879 ( .A(n13078), .B(n33287), .X(n13077) );
  nor_x1_sg U49880 ( .A(n33802), .B(n13076), .X(n13078) );
  nor_x1_sg U49881 ( .A(n35607), .B(n13083), .X(\shifter_0/n7201 ) );
  nor_x1_sg U49882 ( .A(n13084), .B(n33285), .X(n13083) );
  nor_x1_sg U49883 ( .A(n33801), .B(n13082), .X(n13084) );
  nor_x1_sg U49884 ( .A(n35603), .B(n13089), .X(\shifter_0/n7197 ) );
  nor_x1_sg U49885 ( .A(n13090), .B(n33286), .X(n13089) );
  nor_x1_sg U49886 ( .A(n30985), .B(n13088), .X(n13090) );
  nor_x1_sg U49887 ( .A(n35503), .B(n13105), .X(\shifter_0/n7193 ) );
  nor_x1_sg U49888 ( .A(n13106), .B(n33870), .X(n13105) );
  nor_x1_sg U49889 ( .A(n32919), .B(n13103), .X(n13106) );
  nor_x1_sg U49890 ( .A(n35593), .B(n13112), .X(\shifter_0/n7189 ) );
  nor_x1_sg U49891 ( .A(n13113), .B(n33871), .X(n13112) );
  nor_x1_sg U49892 ( .A(n29774), .B(n13111), .X(n13113) );
  nor_x1_sg U49893 ( .A(n35592), .B(n13123), .X(\shifter_0/n7181 ) );
  nor_x1_sg U49894 ( .A(n13124), .B(n30944), .X(n13123) );
  nor_x1_sg U49895 ( .A(n32919), .B(n13122), .X(n13124) );
  nor_x1_sg U49896 ( .A(n35591), .B(n13134), .X(\shifter_0/n7173 ) );
  nor_x1_sg U49897 ( .A(n13135), .B(n33871), .X(n13134) );
  nor_x1_sg U49898 ( .A(n32917), .B(n13133), .X(n13135) );
  nor_x1_sg U49899 ( .A(n35590), .B(n13140), .X(\shifter_0/n7169 ) );
  nor_x1_sg U49900 ( .A(n13141), .B(n33873), .X(n13140) );
  nor_x1_sg U49901 ( .A(n32918), .B(n13139), .X(n13141) );
  nor_x1_sg U49902 ( .A(n35506), .B(n13146), .X(\shifter_0/n7165 ) );
  nor_x1_sg U49903 ( .A(n13147), .B(n33872), .X(n13146) );
  nor_x1_sg U49904 ( .A(n32918), .B(n13145), .X(n13147) );
  nor_x1_sg U49905 ( .A(n35589), .B(n13152), .X(\shifter_0/n7161 ) );
  nor_x1_sg U49906 ( .A(n13153), .B(n33872), .X(n13152) );
  nor_x1_sg U49907 ( .A(n32918), .B(n13151), .X(n13153) );
  nor_x1_sg U49908 ( .A(n35588), .B(n13158), .X(\shifter_0/n7157 ) );
  nor_x1_sg U49909 ( .A(n13159), .B(n33871), .X(n13158) );
  nor_x1_sg U49910 ( .A(n32918), .B(n13157), .X(n13159) );
  nor_x1_sg U49911 ( .A(n35513), .B(n13164), .X(\shifter_0/n7153 ) );
  nor_x1_sg U49912 ( .A(n13165), .B(n30944), .X(n13164) );
  nor_x1_sg U49913 ( .A(n29774), .B(n13163), .X(n13165) );
  nor_x1_sg U49914 ( .A(n35587), .B(n13170), .X(\shifter_0/n7149 ) );
  nor_x1_sg U49915 ( .A(n13171), .B(n33870), .X(n13170) );
  nor_x1_sg U49916 ( .A(n32916), .B(n13169), .X(n13171) );
  nor_x1_sg U49917 ( .A(n35586), .B(n13176), .X(\shifter_0/n7145 ) );
  nor_x1_sg U49918 ( .A(n13177), .B(n30943), .X(n13176) );
  nor_x1_sg U49919 ( .A(n32919), .B(n13175), .X(n13177) );
  nor_x1_sg U49920 ( .A(n35505), .B(n13182), .X(\shifter_0/n7141 ) );
  nor_x1_sg U49921 ( .A(n13183), .B(n30943), .X(n13182) );
  nor_x1_sg U49922 ( .A(n32917), .B(n13181), .X(n13183) );
  nor_x1_sg U49923 ( .A(n35585), .B(n13188), .X(\shifter_0/n7137 ) );
  nor_x1_sg U49924 ( .A(n13189), .B(n33872), .X(n13188) );
  nor_x1_sg U49925 ( .A(n32916), .B(n13187), .X(n13189) );
  nor_x1_sg U49926 ( .A(n35584), .B(n13194), .X(\shifter_0/n7133 ) );
  nor_x1_sg U49927 ( .A(n13195), .B(n33870), .X(n13194) );
  nor_x1_sg U49928 ( .A(n32916), .B(n13193), .X(n13195) );
  nor_x1_sg U49929 ( .A(n35512), .B(n13200), .X(\shifter_0/n7129 ) );
  nor_x1_sg U49930 ( .A(n13201), .B(n33873), .X(n13200) );
  nor_x1_sg U49931 ( .A(n29774), .B(n13199), .X(n13201) );
  nor_x1_sg U49932 ( .A(n35583), .B(n13216), .X(\shifter_0/n7117 ) );
  nor_x1_sg U49933 ( .A(n13217), .B(n33873), .X(n13216) );
  nor_x1_sg U49934 ( .A(n32919), .B(n13215), .X(n13217) );
  nor_x1_sg U49935 ( .A(n30018), .B(n31204), .X(\filter_0/n6284 ) );
  nand_x1_sg U49936 ( .A(n30308), .B(n35116), .X(n13814) );
  nand_x1_sg U49937 ( .A(n34256), .B(n35115), .X(n13848) );
  nand_x1_sg U49938 ( .A(n34255), .B(n42766), .X(n13879) );
  nand_x1_sg U49939 ( .A(n34255), .B(n42767), .X(n13910) );
  nand_x1_sg U49940 ( .A(n30310), .B(n35114), .X(n13941) );
  nand_x1_sg U49941 ( .A(n34256), .B(n42768), .X(n13972) );
  nand_x1_sg U49942 ( .A(n31383), .B(n42769), .X(n14003) );
  nand_x1_sg U49943 ( .A(n34257), .B(n35113), .X(n14034) );
  nand_x1_sg U49944 ( .A(n30086), .B(n42774), .X(n14313) );
  nand_x1_sg U49945 ( .A(n30310), .B(n42775), .X(n14344) );
  nand_x1_sg U49946 ( .A(n34256), .B(n35108), .X(n14375) );
  nand_x1_sg U49947 ( .A(n31802), .B(n35107), .X(n14406) );
  nand_x1_sg U49948 ( .A(n34257), .B(n35138), .X(n14438) );
  nand_x1_sg U49949 ( .A(n31384), .B(n35137), .X(n14469) );
  nand_x1_sg U49950 ( .A(n30308), .B(n42650), .X(n14533) );
  nand_x1_sg U49951 ( .A(n34256), .B(n42651), .X(n14595) );
  nand_x1_sg U49952 ( .A(n34254), .B(n42652), .X(n14626) );
  nand_x1_sg U49953 ( .A(n34257), .B(n35135), .X(n14657) );
  nand_x1_sg U49954 ( .A(n30308), .B(n42653), .X(n14688) );
  nand_x1_sg U49955 ( .A(n31384), .B(n42654), .X(n14719) );
  nand_x1_sg U49956 ( .A(n34254), .B(n35134), .X(n14750) );
  nand_x1_sg U49957 ( .A(n30308), .B(n42655), .X(n14781) );
  nand_x1_sg U49958 ( .A(n31383), .B(n42656), .X(n14812) );
  nand_x1_sg U49959 ( .A(n34254), .B(n35133), .X(n14843) );
  nand_x1_sg U49960 ( .A(n31802), .B(n35132), .X(n14874) );
  nand_x1_sg U49961 ( .A(n30086), .B(n35131), .X(n14905) );
  nand_x1_sg U49962 ( .A(n30086), .B(n42657), .X(n14936) );
  nand_x1_sg U49963 ( .A(n30310), .B(n35129), .X(n15029) );
  nand_x1_sg U49964 ( .A(n31384), .B(n42770), .X(n14065) );
  nand_x1_sg U49965 ( .A(n31383), .B(n42771), .X(n14096) );
  nand_x1_sg U49966 ( .A(n31802), .B(n35112), .X(n14127) );
  nand_x1_sg U49967 ( .A(n34257), .B(n42772), .X(n14158) );
  nand_x1_sg U49968 ( .A(n31802), .B(n42773), .X(n14189) );
  nand_x1_sg U49969 ( .A(n34254), .B(n35111), .X(n14220) );
  nand_x1_sg U49970 ( .A(n31383), .B(n35110), .X(n14251) );
  nand_x1_sg U49971 ( .A(n34255), .B(n35109), .X(n14282) );
  nor_x1_sg U49972 ( .A(n31850), .B(n11690), .X(\shifter_0/n8393 ) );
  nor_x1_sg U49973 ( .A(n30058), .B(n11691), .X(\shifter_0/n8389 ) );
  nor_x1_sg U49974 ( .A(n34125), .B(n11692), .X(\shifter_0/n8385 ) );
  nor_x1_sg U49975 ( .A(n31461), .B(n11693), .X(\shifter_0/n8381 ) );
  nor_x1_sg U49976 ( .A(n34126), .B(n11694), .X(\shifter_0/n8377 ) );
  nor_x1_sg U49977 ( .A(n31461), .B(n11695), .X(\shifter_0/n8373 ) );
  nor_x1_sg U49978 ( .A(n30057), .B(n11696), .X(\shifter_0/n8369 ) );
  nor_x1_sg U49979 ( .A(n30058), .B(n11697), .X(\shifter_0/n8365 ) );
  nor_x1_sg U49980 ( .A(n31851), .B(n11698), .X(\shifter_0/n8361 ) );
  nor_x1_sg U49981 ( .A(n34127), .B(n11699), .X(\shifter_0/n8357 ) );
  nor_x1_sg U49982 ( .A(n30058), .B(n11700), .X(\shifter_0/n8353 ) );
  nor_x1_sg U49983 ( .A(n34124), .B(n11701), .X(\shifter_0/n8349 ) );
  nor_x1_sg U49984 ( .A(n34125), .B(n11702), .X(\shifter_0/n8345 ) );
  nor_x1_sg U49985 ( .A(n31851), .B(n11703), .X(\shifter_0/n8341 ) );
  nor_x1_sg U49986 ( .A(n34126), .B(n11704), .X(\shifter_0/n8337 ) );
  nor_x1_sg U49987 ( .A(n34124), .B(n11705), .X(\shifter_0/n8333 ) );
  nor_x1_sg U49988 ( .A(n34125), .B(n11706), .X(\shifter_0/n8329 ) );
  nor_x1_sg U49989 ( .A(n31462), .B(n11707), .X(\shifter_0/n8325 ) );
  nor_x1_sg U49990 ( .A(n30057), .B(n11708), .X(\shifter_0/n8321 ) );
  nor_x1_sg U49991 ( .A(n31851), .B(n11709), .X(\shifter_0/n8317 ) );
  nor_x1_sg U49992 ( .A(n34118), .B(n11717), .X(\shifter_0/n8313 ) );
  nor_x1_sg U49993 ( .A(n34116), .B(n11718), .X(\shifter_0/n8309 ) );
  nor_x1_sg U49994 ( .A(n30052), .B(n11719), .X(\shifter_0/n8305 ) );
  nor_x1_sg U49995 ( .A(n30051), .B(n11720), .X(\shifter_0/n8301 ) );
  nor_x1_sg U49996 ( .A(n30051), .B(n11721), .X(\shifter_0/n8297 ) );
  nor_x1_sg U49997 ( .A(n31467), .B(n11722), .X(\shifter_0/n8293 ) );
  nor_x1_sg U49998 ( .A(n34116), .B(n11723), .X(\shifter_0/n8289 ) );
  nor_x1_sg U49999 ( .A(n31468), .B(n11724), .X(\shifter_0/n8285 ) );
  nor_x1_sg U50000 ( .A(n34119), .B(n11725), .X(\shifter_0/n8281 ) );
  nor_x1_sg U50001 ( .A(n31854), .B(n11726), .X(\shifter_0/n8277 ) );
  nor_x1_sg U50002 ( .A(n31467), .B(n11727), .X(\shifter_0/n8273 ) );
  nor_x1_sg U50003 ( .A(n31855), .B(n11728), .X(\shifter_0/n8269 ) );
  nor_x1_sg U50004 ( .A(n34117), .B(n11729), .X(\shifter_0/n8265 ) );
  nor_x1_sg U50005 ( .A(n34117), .B(n11730), .X(\shifter_0/n8261 ) );
  nor_x1_sg U50006 ( .A(n34119), .B(n11731), .X(\shifter_0/n8257 ) );
  nor_x1_sg U50007 ( .A(n31854), .B(n11732), .X(\shifter_0/n8253 ) );
  nor_x1_sg U50008 ( .A(n31855), .B(n11733), .X(\shifter_0/n8249 ) );
  nor_x1_sg U50009 ( .A(n34119), .B(n11734), .X(\shifter_0/n8245 ) );
  nor_x1_sg U50010 ( .A(n34118), .B(n11735), .X(\shifter_0/n8241 ) );
  nor_x1_sg U50011 ( .A(n30051), .B(n11736), .X(\shifter_0/n8237 ) );
  nor_x1_sg U50012 ( .A(n30049), .B(n11743), .X(\shifter_0/n8233 ) );
  nor_x1_sg U50013 ( .A(n34115), .B(n11744), .X(\shifter_0/n8229 ) );
  nor_x1_sg U50014 ( .A(n31470), .B(n11745), .X(\shifter_0/n8225 ) );
  nor_x1_sg U50015 ( .A(n34114), .B(n11746), .X(\shifter_0/n8221 ) );
  nor_x1_sg U50016 ( .A(n31857), .B(n11747), .X(\shifter_0/n8217 ) );
  nor_x1_sg U50017 ( .A(n30049), .B(n11748), .X(\shifter_0/n8213 ) );
  nor_x1_sg U50018 ( .A(n30049), .B(n11749), .X(\shifter_0/n8209 ) );
  nor_x1_sg U50019 ( .A(n34115), .B(n11750), .X(\shifter_0/n8205 ) );
  nor_x1_sg U50020 ( .A(n30048), .B(n11751), .X(\shifter_0/n8201 ) );
  nor_x1_sg U50021 ( .A(n34112), .B(n11752), .X(\shifter_0/n8197 ) );
  nor_x1_sg U50022 ( .A(n34114), .B(n11753), .X(\shifter_0/n8193 ) );
  nor_x1_sg U50023 ( .A(n34113), .B(n11754), .X(\shifter_0/n8189 ) );
  nor_x1_sg U50024 ( .A(n31470), .B(n11755), .X(\shifter_0/n8185 ) );
  nor_x1_sg U50025 ( .A(n34112), .B(n11756), .X(\shifter_0/n8181 ) );
  nor_x1_sg U50026 ( .A(n31857), .B(n11757), .X(\shifter_0/n8177 ) );
  nor_x1_sg U50027 ( .A(n31856), .B(n11758), .X(\shifter_0/n8173 ) );
  nor_x1_sg U50028 ( .A(n31471), .B(n11759), .X(\shifter_0/n8169 ) );
  nor_x1_sg U50029 ( .A(n31856), .B(n11760), .X(\shifter_0/n8165 ) );
  nor_x1_sg U50030 ( .A(n34112), .B(n11761), .X(\shifter_0/n8161 ) );
  nor_x1_sg U50031 ( .A(n31857), .B(n11762), .X(\shifter_0/n8157 ) );
  nor_x1_sg U50032 ( .A(n30055), .B(n11771), .X(\shifter_0/n8153 ) );
  nor_x1_sg U50033 ( .A(n30055), .B(n11772), .X(\shifter_0/n8149 ) );
  nor_x1_sg U50034 ( .A(n34120), .B(n11773), .X(\shifter_0/n8145 ) );
  nor_x1_sg U50035 ( .A(n31852), .B(n11774), .X(\shifter_0/n8141 ) );
  nor_x1_sg U50036 ( .A(n34122), .B(n11775), .X(\shifter_0/n8137 ) );
  nor_x1_sg U50037 ( .A(n31853), .B(n11776), .X(\shifter_0/n8133 ) );
  nor_x1_sg U50038 ( .A(n31853), .B(n11777), .X(\shifter_0/n8129 ) );
  nor_x1_sg U50039 ( .A(n30055), .B(n11778), .X(\shifter_0/n8125 ) );
  nor_x1_sg U50040 ( .A(n30055), .B(n11779), .X(\shifter_0/n8121 ) );
  nor_x1_sg U50041 ( .A(n31852), .B(n11780), .X(\shifter_0/n8117 ) );
  nor_x1_sg U50042 ( .A(n31853), .B(n11781), .X(\shifter_0/n8113 ) );
  nor_x1_sg U50043 ( .A(n31465), .B(n11782), .X(\shifter_0/n8109 ) );
  nor_x1_sg U50044 ( .A(n34120), .B(n11783), .X(\shifter_0/n8105 ) );
  nor_x1_sg U50045 ( .A(n30054), .B(n11784), .X(\shifter_0/n8101 ) );
  nor_x1_sg U50046 ( .A(n30054), .B(n11785), .X(\shifter_0/n8097 ) );
  nor_x1_sg U50047 ( .A(n34121), .B(n11786), .X(\shifter_0/n8093 ) );
  nor_x1_sg U50048 ( .A(n31465), .B(n11787), .X(\shifter_0/n8089 ) );
  nor_x1_sg U50049 ( .A(n34122), .B(n11788), .X(\shifter_0/n8085 ) );
  nor_x1_sg U50050 ( .A(n34121), .B(n11789), .X(\shifter_0/n8081 ) );
  nor_x1_sg U50051 ( .A(n34123), .B(n11790), .X(\shifter_0/n8077 ) );
  nand_x1_sg U50052 ( .A(n31378), .B(n42742), .X(n13901) );
  nand_x1_sg U50053 ( .A(n30089), .B(n42758), .X(n13902) );
  nand_x1_sg U50054 ( .A(n30314), .B(n42743), .X(n13932) );
  nand_x1_sg U50055 ( .A(n34270), .B(n42759), .X(n13933) );
  nand_x1_sg U50056 ( .A(n34266), .B(n42744), .X(n14056) );
  nand_x1_sg U50057 ( .A(n34270), .B(n42760), .X(n14057) );
  nand_x1_sg U50058 ( .A(n31377), .B(n42745), .X(n14087) );
  nand_x1_sg U50059 ( .A(n30317), .B(n42761), .X(n14088) );
  nand_x1_sg U50060 ( .A(n34264), .B(n42746), .X(n14180) );
  nand_x1_sg U50061 ( .A(n34269), .B(n42762), .X(n14181) );
  nand_x1_sg U50062 ( .A(n34267), .B(n42747), .X(n14211) );
  nand_x1_sg U50063 ( .A(n34271), .B(n42763), .X(n14212) );
  nand_x1_sg U50064 ( .A(n31800), .B(n42748), .X(n14335) );
  nand_x1_sg U50065 ( .A(n34272), .B(n42764), .X(n14336) );
  nand_x1_sg U50066 ( .A(n34265), .B(n42749), .X(n14366) );
  nand_x1_sg U50067 ( .A(n31799), .B(n42765), .X(n14367) );
  nand_x1_sg U50068 ( .A(n34267), .B(n42630), .X(n14679) );
  nand_x1_sg U50069 ( .A(n34271), .B(n42644), .X(n14680) );
  nand_x1_sg U50070 ( .A(n30316), .B(n42631), .X(n14710) );
  nand_x1_sg U50071 ( .A(n34271), .B(n42645), .X(n14711) );
  nand_x1_sg U50072 ( .A(n30314), .B(n42632), .X(n14803) );
  nand_x1_sg U50073 ( .A(n34270), .B(n42646), .X(n14804) );
  nand_x1_sg U50074 ( .A(n30316), .B(n42633), .X(n14834) );
  nand_x1_sg U50075 ( .A(n34272), .B(n42647), .X(n14835) );
  nand_x1_sg U50076 ( .A(n34267), .B(n42635), .X(n14927) );
  nand_x1_sg U50077 ( .A(n30319), .B(n42649), .X(n14928) );
  nor_x1_sg U50078 ( .A(n42766), .B(n31755), .X(\shifter_0/n6466 ) );
  nor_x1_sg U50079 ( .A(n42767), .B(n34379), .X(\shifter_0/n6462 ) );
  nor_x1_sg U50080 ( .A(n42768), .B(n30111), .X(\shifter_0/n6454 ) );
  nor_x1_sg U50081 ( .A(n42769), .B(n34382), .X(\shifter_0/n6450 ) );
  nor_x1_sg U50082 ( .A(n42770), .B(n34380), .X(\shifter_0/n6442 ) );
  nor_x1_sg U50083 ( .A(n42771), .B(n31308), .X(\shifter_0/n6438 ) );
  nor_x1_sg U50084 ( .A(n42772), .B(n34379), .X(\shifter_0/n6430 ) );
  nor_x1_sg U50085 ( .A(n42773), .B(n34381), .X(\shifter_0/n6426 ) );
  nor_x1_sg U50086 ( .A(n42774), .B(n30362), .X(\shifter_0/n6410 ) );
  nor_x1_sg U50087 ( .A(n42775), .B(n34379), .X(\shifter_0/n6406 ) );
  nor_x1_sg U50088 ( .A(n31764), .B(n11587), .X(\shifter_0/n8713 ) );
  nor_x1_sg U50089 ( .A(n31320), .B(n11588), .X(\shifter_0/n8709 ) );
  nor_x1_sg U50090 ( .A(n31320), .B(n11589), .X(\shifter_0/n8705 ) );
  nor_x1_sg U50091 ( .A(n30354), .B(n11590), .X(\shifter_0/n8701 ) );
  nor_x1_sg U50092 ( .A(n31321), .B(n11591), .X(\shifter_0/n8697 ) );
  nor_x1_sg U50093 ( .A(n34362), .B(n11592), .X(\shifter_0/n8693 ) );
  nor_x1_sg U50094 ( .A(n34360), .B(n11593), .X(\shifter_0/n8689 ) );
  nor_x1_sg U50095 ( .A(n31763), .B(n11594), .X(\shifter_0/n8685 ) );
  nor_x1_sg U50096 ( .A(n34361), .B(n11595), .X(\shifter_0/n8681 ) );
  nor_x1_sg U50097 ( .A(n31763), .B(n11596), .X(\shifter_0/n8677 ) );
  nor_x1_sg U50098 ( .A(n31321), .B(n11597), .X(\shifter_0/n8673 ) );
  nor_x1_sg U50099 ( .A(n30354), .B(n11598), .X(\shifter_0/n8669 ) );
  nor_x1_sg U50100 ( .A(n30354), .B(n11599), .X(\shifter_0/n8665 ) );
  nor_x1_sg U50101 ( .A(n34360), .B(n11600), .X(\shifter_0/n8661 ) );
  nor_x1_sg U50102 ( .A(n31321), .B(n11601), .X(\shifter_0/n8657 ) );
  nor_x1_sg U50103 ( .A(n34360), .B(n11602), .X(\shifter_0/n8653 ) );
  nor_x1_sg U50104 ( .A(n11586), .B(n11603), .X(\shifter_0/n8649 ) );
  nor_x1_sg U50105 ( .A(n34362), .B(n11604), .X(\shifter_0/n8645 ) );
  nor_x1_sg U50106 ( .A(n34359), .B(n11605), .X(\shifter_0/n8641 ) );
  nor_x1_sg U50107 ( .A(n31763), .B(n11606), .X(\shifter_0/n8637 ) );
  nor_x1_sg U50108 ( .A(n11536), .B(n11537), .X(\shifter_0/n8873 ) );
  nor_x1_sg U50109 ( .A(n31762), .B(n11538), .X(\shifter_0/n8869 ) );
  nor_x1_sg U50110 ( .A(n34364), .B(n11539), .X(\shifter_0/n8865 ) );
  nor_x1_sg U50111 ( .A(n29709), .B(n11540), .X(\shifter_0/n8861 ) );
  nor_x1_sg U50112 ( .A(n34364), .B(n11541), .X(\shifter_0/n8857 ) );
  nor_x1_sg U50113 ( .A(n30108), .B(n11542), .X(\shifter_0/n8853 ) );
  nor_x1_sg U50114 ( .A(n31318), .B(n11543), .X(\shifter_0/n8849 ) );
  nor_x1_sg U50115 ( .A(n30108), .B(n11544), .X(\shifter_0/n8845 ) );
  nor_x1_sg U50116 ( .A(n31762), .B(n11545), .X(\shifter_0/n8841 ) );
  nor_x1_sg U50117 ( .A(n34366), .B(n11546), .X(\shifter_0/n8837 ) );
  nor_x1_sg U50118 ( .A(n31318), .B(n11547), .X(\shifter_0/n8833 ) );
  nor_x1_sg U50119 ( .A(n31318), .B(n11548), .X(\shifter_0/n8829 ) );
  nor_x1_sg U50120 ( .A(n31317), .B(n11549), .X(\shifter_0/n8825 ) );
  nor_x1_sg U50121 ( .A(n34367), .B(n11550), .X(\shifter_0/n8821 ) );
  nor_x1_sg U50122 ( .A(n34364), .B(n11551), .X(\shifter_0/n8817 ) );
  nor_x1_sg U50123 ( .A(n31317), .B(n11552), .X(\shifter_0/n8813 ) );
  nor_x1_sg U50124 ( .A(n29709), .B(n11553), .X(\shifter_0/n8809 ) );
  nor_x1_sg U50125 ( .A(n34367), .B(n11554), .X(\shifter_0/n8805 ) );
  nor_x1_sg U50126 ( .A(n30356), .B(n11555), .X(\shifter_0/n8801 ) );
  nor_x1_sg U50127 ( .A(n31761), .B(n11556), .X(\shifter_0/n8797 ) );
  nor_x1_sg U50128 ( .A(n34355), .B(n11563), .X(\shifter_0/n8793 ) );
  nor_x1_sg U50129 ( .A(n34356), .B(n11564), .X(\shifter_0/n8789 ) );
  nor_x1_sg U50130 ( .A(n34354), .B(n11565), .X(\shifter_0/n8785 ) );
  nor_x1_sg U50131 ( .A(n31323), .B(n11566), .X(\shifter_0/n8781 ) );
  nor_x1_sg U50132 ( .A(n31765), .B(n11567), .X(\shifter_0/n8777 ) );
  nor_x1_sg U50133 ( .A(n34357), .B(n11568), .X(\shifter_0/n8773 ) );
  nor_x1_sg U50134 ( .A(n30352), .B(n11569), .X(\shifter_0/n8769 ) );
  nor_x1_sg U50135 ( .A(n31324), .B(n11570), .X(\shifter_0/n8765 ) );
  nor_x1_sg U50136 ( .A(n31323), .B(n11571), .X(\shifter_0/n8761 ) );
  nor_x1_sg U50137 ( .A(n11562), .B(n11572), .X(\shifter_0/n8757 ) );
  nor_x1_sg U50138 ( .A(n34357), .B(n11573), .X(\shifter_0/n8753 ) );
  nor_x1_sg U50139 ( .A(n31765), .B(n11574), .X(\shifter_0/n8749 ) );
  nor_x1_sg U50140 ( .A(n31323), .B(n11575), .X(\shifter_0/n8745 ) );
  nor_x1_sg U50141 ( .A(n30106), .B(n11576), .X(\shifter_0/n8741 ) );
  nor_x1_sg U50142 ( .A(n31766), .B(n11577), .X(\shifter_0/n8737 ) );
  nor_x1_sg U50143 ( .A(n31324), .B(n11578), .X(\shifter_0/n8733 ) );
  nor_x1_sg U50144 ( .A(n31766), .B(n11579), .X(\shifter_0/n8729 ) );
  nor_x1_sg U50145 ( .A(n31766), .B(n11580), .X(\shifter_0/n8725 ) );
  nor_x1_sg U50146 ( .A(n34354), .B(n11581), .X(\shifter_0/n8721 ) );
  nor_x1_sg U50147 ( .A(n31765), .B(n11582), .X(\shifter_0/n8717 ) );
  nor_x1_sg U50148 ( .A(n35116), .B(n30111), .X(\shifter_0/n6474 ) );
  nor_x1_sg U50149 ( .A(n35115), .B(n31756), .X(\shifter_0/n6470 ) );
  nor_x1_sg U50150 ( .A(n35114), .B(n31309), .X(\shifter_0/n6458 ) );
  nor_x1_sg U50151 ( .A(n35113), .B(n31755), .X(\shifter_0/n6446 ) );
  nor_x1_sg U50152 ( .A(n35112), .B(n31309), .X(\shifter_0/n6434 ) );
  nor_x1_sg U50153 ( .A(n35111), .B(n31308), .X(\shifter_0/n6422 ) );
  nor_x1_sg U50154 ( .A(n35110), .B(n29706), .X(\shifter_0/n6418 ) );
  nor_x1_sg U50155 ( .A(n35109), .B(n30111), .X(\shifter_0/n6414 ) );
  nor_x1_sg U50156 ( .A(n35108), .B(n31755), .X(\shifter_0/n6402 ) );
  nor_x1_sg U50157 ( .A(n35107), .B(n34380), .X(\shifter_0/n6398 ) );
  nor_x1_sg U50158 ( .A(n34216), .B(n41564), .X(\shifter_0/n7594 ) );
  inv_x1_sg U50159 ( .A(n12528), .X(n41564) );
  nor_x1_sg U50160 ( .A(n34214), .B(n12528), .X(\shifter_0/n7593 ) );
  nor_x1_sg U50161 ( .A(n31816), .B(n41565), .X(\shifter_0/n7590 ) );
  inv_x1_sg U50162 ( .A(n12534), .X(n41565) );
  nor_x1_sg U50163 ( .A(n34216), .B(n12534), .X(\shifter_0/n7589 ) );
  nor_x1_sg U50164 ( .A(n29733), .B(n41566), .X(\shifter_0/n7586 ) );
  inv_x1_sg U50165 ( .A(n12538), .X(n41566) );
  nor_x1_sg U50166 ( .A(n31407), .B(n12538), .X(\shifter_0/n7585 ) );
  nor_x1_sg U50167 ( .A(n31407), .B(n41567), .X(\shifter_0/n7582 ) );
  inv_x1_sg U50168 ( .A(n12542), .X(n41567) );
  nor_x1_sg U50169 ( .A(n34217), .B(n12542), .X(\shifter_0/n7581 ) );
  nor_x1_sg U50170 ( .A(n31408), .B(n41574), .X(\shifter_0/n7554 ) );
  inv_x1_sg U50171 ( .A(n12570), .X(n41574) );
  nor_x1_sg U50172 ( .A(n34215), .B(n12570), .X(\shifter_0/n7553 ) );
  nor_x1_sg U50173 ( .A(n29733), .B(n41575), .X(\shifter_0/n7550 ) );
  inv_x1_sg U50174 ( .A(n12574), .X(n41575) );
  nor_x1_sg U50175 ( .A(n34216), .B(n12574), .X(\shifter_0/n7549 ) );
  nor_x1_sg U50176 ( .A(n30078), .B(n41578), .X(\shifter_0/n7538 ) );
  inv_x1_sg U50177 ( .A(n12586), .X(n41578) );
  nor_x1_sg U50178 ( .A(n34214), .B(n12586), .X(\shifter_0/n7537 ) );
  nor_x1_sg U50179 ( .A(n31407), .B(n41579), .X(\shifter_0/n7534 ) );
  inv_x1_sg U50180 ( .A(n12590), .X(n41579) );
  nor_x1_sg U50181 ( .A(n31815), .B(n12590), .X(\shifter_0/n7533 ) );
  nor_x1_sg U50182 ( .A(n31816), .B(n41580), .X(\shifter_0/n7530 ) );
  inv_x1_sg U50183 ( .A(n12594), .X(n41580) );
  nor_x1_sg U50184 ( .A(n30290), .B(n12594), .X(\shifter_0/n7529 ) );
  nor_x1_sg U50185 ( .A(n30078), .B(n41581), .X(\shifter_0/n7526 ) );
  inv_x1_sg U50186 ( .A(n12598), .X(n41581) );
  nor_x1_sg U50187 ( .A(n31815), .B(n12598), .X(\shifter_0/n7525 ) );
  nor_x1_sg U50188 ( .A(n35645), .B(n41582), .X(\shifter_0/n7522 ) );
  inv_x1_sg U50189 ( .A(n12602), .X(n41582) );
  nor_x1_sg U50190 ( .A(n34217), .B(n12602), .X(\shifter_0/n7521 ) );
  nor_x1_sg U50191 ( .A(n31408), .B(n41583), .X(\shifter_0/n7518 ) );
  inv_x1_sg U50192 ( .A(n12606), .X(n41583) );
  nor_x1_sg U50193 ( .A(n31407), .B(n12606), .X(\shifter_0/n7517 ) );
  nor_x1_sg U50194 ( .A(n31410), .B(n41584), .X(\shifter_0/n7514 ) );
  inv_x1_sg U50195 ( .A(n12619), .X(n41584) );
  nor_x1_sg U50196 ( .A(n34212), .B(n12619), .X(\shifter_0/n7513 ) );
  nor_x1_sg U50197 ( .A(n34210), .B(n41585), .X(\shifter_0/n7510 ) );
  inv_x1_sg U50198 ( .A(n12623), .X(n41585) );
  nor_x1_sg U50199 ( .A(n30077), .B(n12623), .X(\shifter_0/n7509 ) );
  nor_x1_sg U50200 ( .A(n31411), .B(n41586), .X(\shifter_0/n7506 ) );
  inv_x1_sg U50201 ( .A(n12627), .X(n41586) );
  nor_x1_sg U50202 ( .A(n30077), .B(n12627), .X(\shifter_0/n7505 ) );
  nor_x1_sg U50203 ( .A(n31817), .B(n41587), .X(\shifter_0/n7502 ) );
  inv_x1_sg U50204 ( .A(n12632), .X(n41587) );
  nor_x1_sg U50205 ( .A(n34212), .B(n12632), .X(\shifter_0/n7501 ) );
  nor_x1_sg U50206 ( .A(n30288), .B(n41594), .X(\shifter_0/n7474 ) );
  inv_x1_sg U50207 ( .A(n12661), .X(n41594) );
  nor_x1_sg U50208 ( .A(n29734), .B(n12661), .X(\shifter_0/n7473 ) );
  nor_x1_sg U50209 ( .A(n30077), .B(n41595), .X(\shifter_0/n7470 ) );
  inv_x1_sg U50210 ( .A(n12665), .X(n41595) );
  nor_x1_sg U50211 ( .A(n31411), .B(n12665), .X(\shifter_0/n7469 ) );
  nor_x1_sg U50212 ( .A(n34209), .B(n41598), .X(\shifter_0/n7458 ) );
  inv_x1_sg U50213 ( .A(n12677), .X(n41598) );
  nor_x1_sg U50214 ( .A(n34211), .B(n12677), .X(\shifter_0/n7457 ) );
  nor_x1_sg U50215 ( .A(n35644), .B(n41599), .X(\shifter_0/n7454 ) );
  inv_x1_sg U50216 ( .A(n12681), .X(n41599) );
  nor_x1_sg U50217 ( .A(n31818), .B(n12681), .X(\shifter_0/n7453 ) );
  nor_x1_sg U50218 ( .A(n29734), .B(n41600), .X(\shifter_0/n7450 ) );
  inv_x1_sg U50219 ( .A(n12685), .X(n41600) );
  nor_x1_sg U50220 ( .A(n34210), .B(n12685), .X(\shifter_0/n7449 ) );
  nor_x1_sg U50221 ( .A(n34210), .B(n41601), .X(\shifter_0/n7446 ) );
  inv_x1_sg U50222 ( .A(n12689), .X(n41601) );
  nor_x1_sg U50223 ( .A(n31817), .B(n12689), .X(\shifter_0/n7445 ) );
  nor_x1_sg U50224 ( .A(n31410), .B(n41602), .X(\shifter_0/n7442 ) );
  inv_x1_sg U50225 ( .A(n12694), .X(n41602) );
  nor_x1_sg U50226 ( .A(n34209), .B(n12694), .X(\shifter_0/n7441 ) );
  nor_x1_sg U50227 ( .A(n31818), .B(n41603), .X(\shifter_0/n7438 ) );
  inv_x1_sg U50228 ( .A(n12699), .X(n41603) );
  nor_x1_sg U50229 ( .A(n30288), .B(n12699), .X(\shifter_0/n7437 ) );
  nor_x1_sg U50230 ( .A(n30017), .B(n15057), .X(\filter_0/n6312 ) );
  nor_x1_sg U50231 ( .A(n33965), .B(n15062), .X(\filter_0/n6308 ) );
  nor_x1_sg U50232 ( .A(n33964), .B(n15076), .X(\filter_0/n6301 ) );
  nor_x1_sg U50233 ( .A(n33965), .B(n15158), .X(\filter_0/n6292 ) );
  nor_x1_sg U50234 ( .A(n31650), .B(n15162), .X(\filter_0/n6288 ) );
  nor_x1_sg U50235 ( .A(n30017), .B(n15193), .X(\filter_0/n4996 ) );
  nor_x1_sg U50236 ( .A(n33965), .B(n15198), .X(\filter_0/n4992 ) );
  nor_x1_sg U50237 ( .A(n31651), .B(n15212), .X(\filter_0/n4985 ) );
  nor_x1_sg U50238 ( .A(n34376), .B(n11614), .X(\shifter_0/n8633 ) );
  nor_x1_sg U50239 ( .A(n34374), .B(n11615), .X(\shifter_0/n8629 ) );
  nor_x1_sg U50240 ( .A(n31758), .B(n11616), .X(\shifter_0/n8625 ) );
  nor_x1_sg U50241 ( .A(n34375), .B(n11617), .X(\shifter_0/n8621 ) );
  nor_x1_sg U50242 ( .A(n31312), .B(n11618), .X(\shifter_0/n8617 ) );
  nor_x1_sg U50243 ( .A(n31311), .B(n11619), .X(\shifter_0/n8613 ) );
  nor_x1_sg U50244 ( .A(n31757), .B(n11620), .X(\shifter_0/n8609 ) );
  nor_x1_sg U50245 ( .A(n31312), .B(n11621), .X(\shifter_0/n8605 ) );
  nor_x1_sg U50246 ( .A(n29707), .B(n11625), .X(\shifter_0/n8589 ) );
  nor_x1_sg U50247 ( .A(n34375), .B(n11626), .X(\shifter_0/n8585 ) );
  nor_x1_sg U50248 ( .A(n30110), .B(n11627), .X(\shifter_0/n8581 ) );
  nor_x1_sg U50249 ( .A(n29707), .B(n11628), .X(\shifter_0/n8577 ) );
  nor_x1_sg U50250 ( .A(n31311), .B(n11629), .X(\shifter_0/n8573 ) );
  nor_x1_sg U50251 ( .A(n31758), .B(n11630), .X(\shifter_0/n8569 ) );
  nor_x1_sg U50252 ( .A(n34377), .B(n11631), .X(\shifter_0/n8565 ) );
  nor_x1_sg U50253 ( .A(n34377), .B(n11632), .X(\shifter_0/n8561 ) );
  nor_x1_sg U50254 ( .A(n30110), .B(n11633), .X(\shifter_0/n8557 ) );
  nor_x1_sg U50255 ( .A(n34279), .B(n11668), .X(\shifter_0/n8473 ) );
  nor_x1_sg U50256 ( .A(n31795), .B(n11669), .X(\shifter_0/n8469 ) );
  nor_x1_sg U50257 ( .A(n29726), .B(n11670), .X(\shifter_0/n8465 ) );
  nor_x1_sg U50258 ( .A(n34280), .B(n11671), .X(\shifter_0/n8461 ) );
  nor_x1_sg U50259 ( .A(n34281), .B(n11672), .X(\shifter_0/n8457 ) );
  nor_x1_sg U50260 ( .A(n34279), .B(n11673), .X(\shifter_0/n8453 ) );
  nor_x1_sg U50261 ( .A(n31369), .B(n11674), .X(\shifter_0/n8449 ) );
  nor_x1_sg U50262 ( .A(n34282), .B(n11675), .X(\shifter_0/n8445 ) );
  nor_x1_sg U50263 ( .A(n30091), .B(n11679), .X(\shifter_0/n8429 ) );
  nor_x1_sg U50264 ( .A(n31369), .B(n11680), .X(\shifter_0/n8425 ) );
  nor_x1_sg U50265 ( .A(n31369), .B(n11681), .X(\shifter_0/n8421 ) );
  nor_x1_sg U50266 ( .A(n34279), .B(n11682), .X(\shifter_0/n8417 ) );
  nor_x1_sg U50267 ( .A(n34280), .B(n11683), .X(\shifter_0/n8413 ) );
  nor_x1_sg U50268 ( .A(n31368), .B(n11684), .X(\shifter_0/n8409 ) );
  nor_x1_sg U50269 ( .A(n34282), .B(n11685), .X(\shifter_0/n8405 ) );
  nor_x1_sg U50270 ( .A(n30322), .B(n11686), .X(\shifter_0/n8401 ) );
  nor_x1_sg U50271 ( .A(n31369), .B(n11687), .X(\shifter_0/n8397 ) );
  nor_x1_sg U50272 ( .A(n34286), .B(n35138), .X(\shifter_0/n6394 ) );
  nor_x1_sg U50273 ( .A(n30324), .B(n35137), .X(\shifter_0/n8950 ) );
  nor_x1_sg U50274 ( .A(n31366), .B(n35136), .X(\shifter_0/n8946 ) );
  nor_x1_sg U50275 ( .A(n34284), .B(n42650), .X(\shifter_0/n8942 ) );
  nor_x1_sg U50276 ( .A(n34286), .B(n42651), .X(\shifter_0/n8934 ) );
  nor_x1_sg U50277 ( .A(n30092), .B(n42652), .X(\shifter_0/n8930 ) );
  nor_x1_sg U50278 ( .A(n30324), .B(n35135), .X(\shifter_0/n8926 ) );
  nor_x1_sg U50279 ( .A(n31794), .B(n42653), .X(\shifter_0/n8922 ) );
  nor_x1_sg U50280 ( .A(n34284), .B(n42654), .X(\shifter_0/n8918 ) );
  nor_x1_sg U50281 ( .A(n31793), .B(n42655), .X(\shifter_0/n8910 ) );
  nor_x1_sg U50282 ( .A(n34285), .B(n42656), .X(\shifter_0/n8906 ) );
  nor_x1_sg U50283 ( .A(n30092), .B(n35133), .X(\shifter_0/n8902 ) );
  nor_x1_sg U50284 ( .A(n30092), .B(n35132), .X(\shifter_0/n8898 ) );
  nor_x1_sg U50285 ( .A(n34287), .B(n35131), .X(\shifter_0/n8894 ) );
  nor_x1_sg U50286 ( .A(n31366), .B(n42657), .X(\shifter_0/n8890 ) );
  nor_x1_sg U50287 ( .A(n31365), .B(n35130), .X(\shifter_0/n8886 ) );
  nor_x1_sg U50288 ( .A(n34287), .B(n35129), .X(\shifter_0/n8878 ) );
  nor_x1_sg U50289 ( .A(n31759), .B(n11642), .X(\shifter_0/n8553 ) );
  nor_x1_sg U50290 ( .A(n31760), .B(n11643), .X(\shifter_0/n8549 ) );
  nor_x1_sg U50291 ( .A(n31314), .B(n11644), .X(\shifter_0/n8545 ) );
  nor_x1_sg U50292 ( .A(n29708), .B(n11645), .X(\shifter_0/n8541 ) );
  nor_x1_sg U50293 ( .A(n30109), .B(n11646), .X(\shifter_0/n8537 ) );
  nor_x1_sg U50294 ( .A(n30358), .B(n11647), .X(\shifter_0/n8533 ) );
  nor_x1_sg U50295 ( .A(n34369), .B(n11648), .X(\shifter_0/n8529 ) );
  nor_x1_sg U50296 ( .A(n31760), .B(n11649), .X(\shifter_0/n8525 ) );
  nor_x1_sg U50297 ( .A(n34371), .B(n11653), .X(\shifter_0/n8509 ) );
  nor_x1_sg U50298 ( .A(n34371), .B(n11654), .X(\shifter_0/n8505 ) );
  nor_x1_sg U50299 ( .A(n34369), .B(n11655), .X(\shifter_0/n8501 ) );
  nor_x1_sg U50300 ( .A(n34372), .B(n11656), .X(\shifter_0/n8497 ) );
  nor_x1_sg U50301 ( .A(n34372), .B(n11657), .X(\shifter_0/n8493 ) );
  nor_x1_sg U50302 ( .A(n31315), .B(n11658), .X(\shifter_0/n8489 ) );
  nor_x1_sg U50303 ( .A(n34372), .B(n11659), .X(\shifter_0/n8485 ) );
  nor_x1_sg U50304 ( .A(n34370), .B(n11660), .X(\shifter_0/n8481 ) );
  nor_x1_sg U50305 ( .A(n34369), .B(n11661), .X(\shifter_0/n8477 ) );
  nor_x1_sg U50306 ( .A(n34215), .B(n41572), .X(\shifter_0/n7562 ) );
  inv_x1_sg U50307 ( .A(n12562), .X(n41572) );
  nor_x1_sg U50308 ( .A(n30290), .B(n12562), .X(\shifter_0/n7561 ) );
  nor_x1_sg U50309 ( .A(n31816), .B(n41573), .X(\shifter_0/n7558 ) );
  inv_x1_sg U50310 ( .A(n12566), .X(n41573) );
  nor_x1_sg U50311 ( .A(n34214), .B(n12566), .X(\shifter_0/n7557 ) );
  nor_x1_sg U50312 ( .A(n31408), .B(n41576), .X(\shifter_0/n7546 ) );
  inv_x1_sg U50313 ( .A(n12578), .X(n41576) );
  nor_x1_sg U50314 ( .A(n34217), .B(n12578), .X(\shifter_0/n7545 ) );
  nor_x1_sg U50315 ( .A(n34214), .B(n41577), .X(\shifter_0/n7542 ) );
  inv_x1_sg U50316 ( .A(n12582), .X(n41577) );
  nor_x1_sg U50317 ( .A(n34217), .B(n12582), .X(\shifter_0/n7541 ) );
  nor_x1_sg U50318 ( .A(n31818), .B(n41592), .X(\shifter_0/n7482 ) );
  inv_x1_sg U50319 ( .A(n12653), .X(n41592) );
  nor_x1_sg U50320 ( .A(n31410), .B(n12653), .X(\shifter_0/n7481 ) );
  nor_x1_sg U50321 ( .A(n31817), .B(n41593), .X(\shifter_0/n7478 ) );
  inv_x1_sg U50322 ( .A(n12657), .X(n41593) );
  nor_x1_sg U50323 ( .A(n34212), .B(n12657), .X(\shifter_0/n7477 ) );
  nor_x1_sg U50324 ( .A(n34209), .B(n41596), .X(\shifter_0/n7466 ) );
  inv_x1_sg U50325 ( .A(n12669), .X(n41596) );
  nor_x1_sg U50326 ( .A(n31411), .B(n12669), .X(\shifter_0/n7465 ) );
  nor_x1_sg U50327 ( .A(n31410), .B(n41597), .X(\shifter_0/n7462 ) );
  inv_x1_sg U50328 ( .A(n12673), .X(n41597) );
  nor_x1_sg U50329 ( .A(n31817), .B(n12673), .X(\shifter_0/n7461 ) );
  nor_x1_sg U50330 ( .A(n34376), .B(n11623), .X(\shifter_0/n8597 ) );
  nor_x1_sg U50331 ( .A(n34374), .B(n11624), .X(\shifter_0/n8593 ) );
  nor_x1_sg U50332 ( .A(n34279), .B(n11677), .X(\shifter_0/n8437 ) );
  nor_x1_sg U50333 ( .A(n31368), .B(n11678), .X(\shifter_0/n8433 ) );
  nor_x1_sg U50334 ( .A(n34372), .B(n11651), .X(\shifter_0/n8517 ) );
  nor_x1_sg U50335 ( .A(n30109), .B(n11652), .X(\shifter_0/n8513 ) );
  nor_x1_sg U50336 ( .A(n31815), .B(n41568), .X(\shifter_0/n7578 ) );
  inv_x1_sg U50337 ( .A(n12546), .X(n41568) );
  nor_x1_sg U50338 ( .A(n31815), .B(n12546), .X(\shifter_0/n7577 ) );
  nor_x1_sg U50339 ( .A(n30290), .B(n41569), .X(\shifter_0/n7574 ) );
  inv_x1_sg U50340 ( .A(n12550), .X(n41569) );
  nor_x1_sg U50341 ( .A(n34215), .B(n12550), .X(\shifter_0/n7573 ) );
  nor_x1_sg U50342 ( .A(n31816), .B(n41570), .X(\shifter_0/n7570 ) );
  inv_x1_sg U50343 ( .A(n12554), .X(n41570) );
  nor_x1_sg U50344 ( .A(n30078), .B(n12554), .X(\shifter_0/n7569 ) );
  nor_x1_sg U50345 ( .A(n31408), .B(n41571), .X(\shifter_0/n7566 ) );
  inv_x1_sg U50346 ( .A(n12558), .X(n41571) );
  nor_x1_sg U50347 ( .A(n34215), .B(n12558), .X(\shifter_0/n7565 ) );
  nor_x1_sg U50348 ( .A(n34212), .B(n41588), .X(\shifter_0/n7498 ) );
  inv_x1_sg U50349 ( .A(n12636), .X(n41588) );
  nor_x1_sg U50350 ( .A(n34211), .B(n12636), .X(\shifter_0/n7497 ) );
  nor_x1_sg U50351 ( .A(n31818), .B(n41589), .X(\shifter_0/n7494 ) );
  inv_x1_sg U50352 ( .A(n12641), .X(n41589) );
  nor_x1_sg U50353 ( .A(n34211), .B(n12641), .X(\shifter_0/n7493 ) );
  nor_x1_sg U50354 ( .A(n30288), .B(n41590), .X(\shifter_0/n7490 ) );
  inv_x1_sg U50355 ( .A(n12645), .X(n41590) );
  nor_x1_sg U50356 ( .A(n34210), .B(n12645), .X(\shifter_0/n7489 ) );
  nor_x1_sg U50357 ( .A(n34209), .B(n41591), .X(\shifter_0/n7486 ) );
  inv_x1_sg U50358 ( .A(n12649), .X(n41591) );
  nor_x1_sg U50359 ( .A(n31411), .B(n12649), .X(\shifter_0/n7485 ) );
  nor_x1_sg U50360 ( .A(n34375), .B(n11622), .X(\shifter_0/n8601 ) );
  nor_x1_sg U50361 ( .A(n34280), .B(n11676), .X(\shifter_0/n8441 ) );
  nor_x1_sg U50362 ( .A(n31365), .B(n35134), .X(\shifter_0/n8914 ) );
  nor_x1_sg U50363 ( .A(n31314), .B(n11650), .X(\shifter_0/n8521 ) );
  nor_x1_sg U50364 ( .A(n15207), .B(n33966), .X(\filter_0/n4988 ) );
  nor_x1_sg U50365 ( .A(n15208), .B(n15209), .X(n15207) );
  nor_x1_sg U50366 ( .A(n31878), .B(n30543), .X(n15209) );
  nor_x1_sg U50367 ( .A(n35096), .B(n15206), .X(n15208) );
  nor_x1_sg U50368 ( .A(n15066), .B(n30018), .X(\filter_0/n6305 ) );
  nor_x1_sg U50369 ( .A(n42403), .B(n15067), .X(n15066) );
  nor_x1_sg U50370 ( .A(n35269), .B(n15068), .X(n15067) );
  nor_x1_sg U50371 ( .A(n15085), .B(n42383), .X(n15084) );
  nor_x1_sg U50372 ( .A(n15221), .B(n42384), .X(n15220) );
  nor_x1_sg U50373 ( .A(n42406), .B(n31650), .X(\filter_0/n6313 ) );
  inv_x1_sg U50374 ( .A(n15057), .X(n42406) );
  nor_x1_sg U50375 ( .A(n42405), .B(n30017), .X(\filter_0/n6309 ) );
  inv_x1_sg U50376 ( .A(n15062), .X(n42405) );
  nor_x1_sg U50377 ( .A(n42401), .B(n31651), .X(\filter_0/n6300 ) );
  inv_x1_sg U50378 ( .A(n15076), .X(n42401) );
  nor_x1_sg U50379 ( .A(n42376), .B(n33966), .X(\filter_0/n6293 ) );
  inv_x1_sg U50380 ( .A(n15158), .X(n42376) );
  nor_x1_sg U50381 ( .A(n42366), .B(n31650), .X(\filter_0/n6289 ) );
  inv_x1_sg U50382 ( .A(n15162), .X(n42366) );
  nor_x1_sg U50383 ( .A(n42396), .B(n30018), .X(\filter_0/n4997 ) );
  inv_x1_sg U50384 ( .A(n15193), .X(n42396) );
  nor_x1_sg U50385 ( .A(n42398), .B(n31651), .X(\filter_0/n4993 ) );
  inv_x1_sg U50386 ( .A(n15198), .X(n42398) );
  nor_x1_sg U50387 ( .A(n42400), .B(n31650), .X(\filter_0/n4984 ) );
  inv_x1_sg U50388 ( .A(n15212), .X(n42400) );
  nand_x1_sg U50389 ( .A(n30569), .B(n32913), .X(n13100) );
  nand_x1_sg U50390 ( .A(n30946), .B(n13103), .X(n13101) );
  nand_x1_sg U50391 ( .A(n30565), .B(n32912), .X(n13109) );
  nand_x1_sg U50392 ( .A(n33867), .B(n13111), .X(n13110) );
  nand_x1_sg U50393 ( .A(n33866), .B(n13117), .X(n13116) );
  nand_x1_sg U50394 ( .A(n33870), .B(n12448), .X(n13115) );
  nand_x1_sg U50395 ( .A(n30583), .B(n32914), .X(n13120) );
  nand_x1_sg U50396 ( .A(n33865), .B(n13122), .X(n13121) );
  nand_x1_sg U50397 ( .A(n30947), .B(n35453), .X(n13127) );
  nand_x1_sg U50398 ( .A(n33873), .B(n12457), .X(n13126) );
  nand_x1_sg U50399 ( .A(n30582), .B(n32914), .X(n13131) );
  nand_x1_sg U50400 ( .A(n33867), .B(n13133), .X(n13132) );
  nand_x1_sg U50401 ( .A(n30581), .B(n32911), .X(n13137) );
  nand_x1_sg U50402 ( .A(n30947), .B(n13139), .X(n13138) );
  nand_x1_sg U50403 ( .A(n30567), .B(n32912), .X(n13143) );
  nand_x1_sg U50404 ( .A(n30946), .B(n13145), .X(n13144) );
  nand_x1_sg U50405 ( .A(n30580), .B(n32911), .X(n13149) );
  nand_x1_sg U50406 ( .A(n33867), .B(n13151), .X(n13150) );
  nand_x1_sg U50407 ( .A(n30579), .B(n32913), .X(n13155) );
  nand_x1_sg U50408 ( .A(n33868), .B(n13157), .X(n13156) );
  nand_x1_sg U50409 ( .A(n30573), .B(n32913), .X(n13161) );
  nand_x1_sg U50410 ( .A(n33868), .B(n13163), .X(n13162) );
  nand_x1_sg U50411 ( .A(n30578), .B(n32914), .X(n13167) );
  nand_x1_sg U50412 ( .A(n33865), .B(n13169), .X(n13168) );
  nand_x1_sg U50413 ( .A(n30577), .B(n29773), .X(n13173) );
  nand_x1_sg U50414 ( .A(n33865), .B(n13175), .X(n13174) );
  nand_x1_sg U50415 ( .A(n30574), .B(n32913), .X(n13179) );
  nand_x1_sg U50416 ( .A(n30947), .B(n13181), .X(n13180) );
  nand_x1_sg U50417 ( .A(n30576), .B(n32911), .X(n13185) );
  nand_x1_sg U50418 ( .A(n30946), .B(n13187), .X(n13186) );
  nand_x1_sg U50419 ( .A(n30575), .B(n32912), .X(n13191) );
  nand_x1_sg U50420 ( .A(n33867), .B(n13193), .X(n13192) );
  nand_x1_sg U50421 ( .A(n30570), .B(n32914), .X(n13197) );
  nand_x1_sg U50422 ( .A(n30947), .B(n13199), .X(n13198) );
  nand_x1_sg U50423 ( .A(n30946), .B(n13205), .X(n13204) );
  nand_x1_sg U50424 ( .A(n33872), .B(n12510), .X(n13203) );
  nand_x1_sg U50425 ( .A(n33866), .B(n13210), .X(n13209) );
  nand_x1_sg U50426 ( .A(n30944), .B(n12515), .X(n13208) );
  nand_x1_sg U50427 ( .A(n30568), .B(n32912), .X(n13213) );
  nand_x1_sg U50428 ( .A(n33868), .B(n13215), .X(n13214) );
  nand_x1_sg U50429 ( .A(n41139), .B(n33877), .X(n12449) );
  nand_x1_sg U50430 ( .A(n33861), .B(n35141), .X(n12450) );
  nand_x1_sg U50431 ( .A(n41141), .B(n30940), .X(n12511) );
  nand_x1_sg U50432 ( .A(n30950), .B(n35140), .X(n12512) );
  nand_x1_sg U50433 ( .A(n41142), .B(n33876), .X(n12516) );
  nand_x1_sg U50434 ( .A(n33861), .B(n35139), .X(n12517) );
  nand_x1_sg U50435 ( .A(n30551), .B(n30988), .X(n12969) );
  nand_x1_sg U50436 ( .A(n33276), .B(n12972), .X(n12970) );
  nand_x1_sg U50437 ( .A(n30566), .B(n33762), .X(n12978) );
  nand_x1_sg U50438 ( .A(n33275), .B(n12980), .X(n12979) );
  nand_x1_sg U50439 ( .A(n30571), .B(n33761), .X(n12990) );
  nand_x1_sg U50440 ( .A(n33275), .B(n12992), .X(n12991) );
  nand_x1_sg U50441 ( .A(n30559), .B(n33759), .X(n12996) );
  nand_x1_sg U50442 ( .A(n33275), .B(n12998), .X(n12997) );
  nand_x1_sg U50443 ( .A(n30572), .B(n33760), .X(n13008) );
  nand_x1_sg U50444 ( .A(n33276), .B(n13010), .X(n13009) );
  nand_x1_sg U50445 ( .A(n30547), .B(n33760), .X(n13014) );
  nand_x1_sg U50446 ( .A(n33277), .B(n13016), .X(n13015) );
  nand_x1_sg U50447 ( .A(n30548), .B(n33760), .X(n13026) );
  nand_x1_sg U50448 ( .A(n33276), .B(n13028), .X(n13027) );
  nand_x1_sg U50449 ( .A(n30561), .B(n33799), .X(n13032) );
  nand_x1_sg U50450 ( .A(n33278), .B(n13034), .X(n13033) );
  nand_x1_sg U50451 ( .A(n30554), .B(n33762), .X(n13044) );
  nand_x1_sg U50452 ( .A(n29909), .B(n13046), .X(n13045) );
  nand_x1_sg U50453 ( .A(n30550), .B(n33759), .X(n13050) );
  nand_x1_sg U50454 ( .A(n33276), .B(n13052), .X(n13051) );
  nand_x1_sg U50455 ( .A(n30556), .B(n33761), .X(n13062) );
  nand_x1_sg U50456 ( .A(n29909), .B(n13064), .X(n13063) );
  nand_x1_sg U50457 ( .A(n30562), .B(n33762), .X(n13068) );
  nand_x1_sg U50458 ( .A(n33278), .B(n13070), .X(n13069) );
  nand_x1_sg U50459 ( .A(n30558), .B(n33759), .X(n13080) );
  nand_x1_sg U50460 ( .A(n33278), .B(n13082), .X(n13081) );
  nand_x1_sg U50461 ( .A(n30560), .B(n30988), .X(n13086) );
  nand_x1_sg U50462 ( .A(n33277), .B(n13088), .X(n13087) );
  nand_x1_sg U50463 ( .A(n30552), .B(n33759), .X(n12984) );
  nand_x1_sg U50464 ( .A(n33278), .B(n12986), .X(n12985) );
  nand_x1_sg U50465 ( .A(n30546), .B(n33762), .X(n13002) );
  nand_x1_sg U50466 ( .A(n29909), .B(n13004), .X(n13003) );
  nand_x1_sg U50467 ( .A(n30553), .B(n33761), .X(n13020) );
  nand_x1_sg U50468 ( .A(n33277), .B(n13022), .X(n13021) );
  nand_x1_sg U50469 ( .A(n30549), .B(n33761), .X(n13038) );
  nand_x1_sg U50470 ( .A(n33275), .B(n13040), .X(n13039) );
  nand_x1_sg U50471 ( .A(n30555), .B(n30988), .X(n13056) );
  nand_x1_sg U50472 ( .A(n29909), .B(n13058), .X(n13057) );
  nand_x1_sg U50473 ( .A(n30557), .B(n30988), .X(n13074) );
  nand_x1_sg U50474 ( .A(n33277), .B(n13076), .X(n13075) );
  nand_x1_sg U50475 ( .A(n33757), .B(n11803), .X(n11802) );
  nand_x1_sg U50476 ( .A(n33757), .B(n11807), .X(n11806) );
  nand_x1_sg U50477 ( .A(n33757), .B(n11811), .X(n11810) );
  nand_x1_sg U50478 ( .A(n33755), .B(n11815), .X(n11814) );
  nand_x1_sg U50479 ( .A(n33754), .B(n11819), .X(n11818) );
  nand_x1_sg U50480 ( .A(n33756), .B(n11823), .X(n11822) );
  nand_x1_sg U50481 ( .A(n30989), .B(n11827), .X(n11826) );
  nand_x1_sg U50482 ( .A(n30990), .B(n11851), .X(n11850) );
  nand_x1_sg U50483 ( .A(n33751), .B(n11855), .X(n11854) );
  nand_x1_sg U50484 ( .A(n33751), .B(n11859), .X(n11858) );
  nand_x1_sg U50485 ( .A(n35652), .B(n11863), .X(n11862) );
  nand_x1_sg U50486 ( .A(n30007), .B(n11867), .X(n11866) );
  nand_x1_sg U50487 ( .A(n33752), .B(n11871), .X(n11870) );
  nand_x1_sg U50488 ( .A(n33751), .B(n11875), .X(n11874) );
  nand_x1_sg U50489 ( .A(n33754), .B(n11805), .X(n11804) );
  nand_x1_sg U50490 ( .A(n33755), .B(n11809), .X(n11808) );
  nand_x1_sg U50491 ( .A(n30010), .B(n11813), .X(n11812) );
  nand_x1_sg U50492 ( .A(n33756), .B(n11817), .X(n11816) );
  nand_x1_sg U50493 ( .A(n30010), .B(n11821), .X(n11820) );
  nand_x1_sg U50494 ( .A(n30989), .B(n11825), .X(n11824) );
  nand_x1_sg U50495 ( .A(n30989), .B(n11829), .X(n11828) );
  nand_x1_sg U50496 ( .A(n30989), .B(n11831), .X(n11830) );
  nand_x1_sg U50497 ( .A(n33754), .B(n11833), .X(n11832) );
  nand_x1_sg U50498 ( .A(n33757), .B(n11835), .X(n11834) );
  nand_x1_sg U50499 ( .A(n33754), .B(n11837), .X(n11836) );
  nand_x1_sg U50500 ( .A(n33756), .B(n11839), .X(n11838) );
  nand_x1_sg U50501 ( .A(n33752), .B(n11853), .X(n11852) );
  nand_x1_sg U50502 ( .A(n30990), .B(n11857), .X(n11856) );
  nand_x1_sg U50503 ( .A(n33752), .B(n11861), .X(n11860) );
  nand_x1_sg U50504 ( .A(n33751), .B(n11865), .X(n11864) );
  nand_x1_sg U50505 ( .A(n30990), .B(n11869), .X(n11868) );
  nand_x1_sg U50506 ( .A(n30007), .B(n11873), .X(n11872) );
  nand_x1_sg U50507 ( .A(n33750), .B(n11877), .X(n11876) );
  nand_x1_sg U50508 ( .A(n33752), .B(n11879), .X(n11878) );
  nand_x1_sg U50509 ( .A(n33750), .B(n11881), .X(n11880) );
  nand_x1_sg U50510 ( .A(n30990), .B(n11883), .X(n11882) );
  nand_x1_sg U50511 ( .A(n30007), .B(n11885), .X(n11884) );
  nand_x1_sg U50512 ( .A(n30007), .B(n11887), .X(n11886) );
  nand_x1_sg U50513 ( .A(n33734), .B(n13231), .X(n13230) );
  nand_x1_sg U50514 ( .A(n33733), .B(n13243), .X(n13242) );
  nand_x1_sg U50515 ( .A(n30994), .B(n13249), .X(n13248) );
  nand_x1_sg U50516 ( .A(n35639), .B(n13255), .X(n13254) );
  nand_x1_sg U50517 ( .A(n33637), .B(n13297), .X(n13296) );
  nand_x1_sg U50518 ( .A(n35621), .B(n13311), .X(n13310) );
  nand_x1_sg U50519 ( .A(n33636), .B(n13317), .X(n13316) );
  nand_x1_sg U50520 ( .A(n31000), .B(n13323), .X(n13322) );
  nand_x1_sg U50521 ( .A(n33735), .B(n13228), .X(n13226) );
  nand_x1_sg U50522 ( .A(n33734), .B(n13234), .X(n13233) );
  nand_x1_sg U50523 ( .A(n30001), .B(n13240), .X(n13239) );
  nand_x1_sg U50524 ( .A(n33735), .B(n13246), .X(n13245) );
  nand_x1_sg U50525 ( .A(n30001), .B(n13252), .X(n13251) );
  nand_x1_sg U50526 ( .A(n30994), .B(n13258), .X(n13257) );
  nand_x1_sg U50527 ( .A(n30994), .B(n13264), .X(n13263) );
  nand_x1_sg U50528 ( .A(n35639), .B(n13270), .X(n13269) );
  nand_x1_sg U50529 ( .A(n33733), .B(n13273), .X(n13272) );
  nand_x1_sg U50530 ( .A(n33734), .B(n13276), .X(n13275) );
  nand_x1_sg U50531 ( .A(n33734), .B(n13279), .X(n13278) );
  nand_x1_sg U50532 ( .A(n30001), .B(n13282), .X(n13281) );
  nand_x1_sg U50533 ( .A(n29993), .B(n13294), .X(n13292) );
  nand_x1_sg U50534 ( .A(n29993), .B(n13300), .X(n13299) );
  nand_x1_sg U50535 ( .A(n29993), .B(n13307), .X(n13306) );
  nand_x1_sg U50536 ( .A(n33636), .B(n13314), .X(n13313) );
  nand_x1_sg U50537 ( .A(n31000), .B(n13320), .X(n13319) );
  nand_x1_sg U50538 ( .A(n31000), .B(n13326), .X(n13325) );
  nand_x1_sg U50539 ( .A(n31000), .B(n13332), .X(n13331) );
  nand_x1_sg U50540 ( .A(n33636), .B(n13338), .X(n13337) );
  nand_x1_sg U50541 ( .A(n33637), .B(n13341), .X(n13340) );
  nand_x1_sg U50542 ( .A(n33635), .B(n13344), .X(n13343) );
  nand_x1_sg U50543 ( .A(n33635), .B(n13347), .X(n13346) );
  nand_x1_sg U50544 ( .A(n33637), .B(n13351), .X(n13350) );
  nand_x1_sg U50545 ( .A(n33739), .B(n13621), .X(n13620) );
  nand_x1_sg U50546 ( .A(n30003), .B(n13637), .X(n13636) );
  nand_x1_sg U50547 ( .A(n30993), .B(n13645), .X(n13644) );
  nand_x1_sg U50548 ( .A(n33737), .B(n13653), .X(n13652) );
  nand_x1_sg U50549 ( .A(n33738), .B(n13616), .X(n13614) );
  nand_x1_sg U50550 ( .A(n33739), .B(n13625), .X(n13624) );
  nand_x1_sg U50551 ( .A(n33738), .B(n13633), .X(n13632) );
  nand_x1_sg U50552 ( .A(n30003), .B(n13641), .X(n13640) );
  nand_x1_sg U50553 ( .A(n30003), .B(n13649), .X(n13648) );
  nand_x1_sg U50554 ( .A(n30993), .B(n13657), .X(n13656) );
  nand_x1_sg U50555 ( .A(n30993), .B(n13665), .X(n13664) );
  nand_x1_sg U50556 ( .A(n33739), .B(n13673), .X(n13672) );
  nand_x1_sg U50557 ( .A(n35637), .B(n13677), .X(n13676) );
  nand_x1_sg U50558 ( .A(n33738), .B(n13681), .X(n13680) );
  nand_x1_sg U50559 ( .A(n30003), .B(n13685), .X(n13684) );
  nand_x1_sg U50560 ( .A(n35637), .B(n13689), .X(n13688) );
  nand_x1_sg U50561 ( .A(n33725), .B(n13707), .X(n13706) );
  nand_x1_sg U50562 ( .A(n33725), .B(n13721), .X(n13720) );
  nand_x1_sg U50563 ( .A(n29999), .B(n13729), .X(n13728) );
  nand_x1_sg U50564 ( .A(n29999), .B(n13737), .X(n13736) );
  nand_x1_sg U50565 ( .A(n29999), .B(n13703), .X(n13701) );
  nand_x1_sg U50566 ( .A(n33724), .B(n13711), .X(n13710) );
  nand_x1_sg U50567 ( .A(n30996), .B(n13718), .X(n13717) );
  nand_x1_sg U50568 ( .A(n33726), .B(n13725), .X(n13724) );
  nand_x1_sg U50569 ( .A(n35636), .B(n13733), .X(n13732) );
  nand_x1_sg U50570 ( .A(n33725), .B(n13741), .X(n13740) );
  nand_x1_sg U50571 ( .A(n35636), .B(n13749), .X(n13748) );
  nand_x1_sg U50572 ( .A(n29999), .B(n13757), .X(n13756) );
  nand_x1_sg U50573 ( .A(n30996), .B(n13761), .X(n13760) );
  nand_x1_sg U50574 ( .A(n33724), .B(n13765), .X(n13764) );
  nand_x1_sg U50575 ( .A(n30996), .B(n13769), .X(n13768) );
  nand_x1_sg U50576 ( .A(n33725), .B(n13772), .X(n13771) );
  nand_x1_sg U50577 ( .A(n11800), .B(n33756), .X(n11799) );
  nand_x1_sg U50578 ( .A(n11848), .B(n35652), .X(n11847) );
  nand_x1_sg U50579 ( .A(\shifter_0/n9407 ), .B(n31226), .X(n21953) );
  nand_x1_sg U50580 ( .A(oi_4[15]), .B(n32629), .X(n21954) );
  nand_x1_sg U50581 ( .A(\shifter_0/n9406 ), .B(n30226), .X(n21955) );
  nand_x1_sg U50582 ( .A(oi_4[14]), .B(n34794), .X(n21956) );
  nand_x1_sg U50583 ( .A(\shifter_0/n9405 ), .B(n31554), .X(n21957) );
  nand_x1_sg U50584 ( .A(oi_4[13]), .B(n32550), .X(n21958) );
  nand_x1_sg U50585 ( .A(\shifter_0/n9035 ), .B(n33206), .X(n18891) );
  nand_x1_sg U50586 ( .A(oi_13[3]), .B(n34953), .X(n18892) );
  nand_x1_sg U50587 ( .A(\shifter_0/n9034 ), .B(n33171), .X(n18893) );
  nand_x1_sg U50588 ( .A(oi_13[2]), .B(n34496), .X(n18894) );
  nand_x1_sg U50589 ( .A(\shifter_0/n9033 ), .B(n31537), .X(n18895) );
  nand_x1_sg U50590 ( .A(oi_13[1]), .B(n30795), .X(n18896) );
  nand_x1_sg U50591 ( .A(\shifter_0/n8963 ), .B(n33159), .X(n18955) );
  nand_x1_sg U50592 ( .A(oi_15[11]), .B(n34792), .X(n18956) );
  nand_x1_sg U50593 ( .A(\shifter_0/n8962 ), .B(n33180), .X(n18957) );
  nand_x1_sg U50594 ( .A(oi_15[10]), .B(n32587), .X(n18958) );
  nand_x1_sg U50595 ( .A(\shifter_0/n8961 ), .B(n35004), .X(n18959) );
  nand_x1_sg U50596 ( .A(oi_15[9]), .B(n34794), .X(n18960) );
  nand_x1_sg U50597 ( .A(\shifter_0/n9335 ), .B(n33216), .X(n19211) );
  nand_x1_sg U50598 ( .A(ow_5[3]), .B(n34499), .X(n19212) );
  nand_x1_sg U50599 ( .A(\shifter_0/n9334 ), .B(n33180), .X(n19213) );
  nand_x1_sg U50600 ( .A(ow_5[2]), .B(n32582), .X(n19214) );
  nand_x1_sg U50601 ( .A(\shifter_0/n9333 ), .B(n31551), .X(n19215) );
  nand_x1_sg U50602 ( .A(ow_5[1]), .B(n32563), .X(n19216) );
  nand_x1_sg U50603 ( .A(\shifter_0/n9058 ), .B(n33164), .X(n19485) );
  nand_x1_sg U50604 ( .A(ow_12[6]), .B(n32581), .X(n19486) );
  nand_x1_sg U50605 ( .A(\shifter_0/n9057 ), .B(n33156), .X(n19487) );
  nand_x1_sg U50606 ( .A(ow_12[5]), .B(n32624), .X(n19488) );
  nand_x1_sg U50607 ( .A(\shifter_0/n9056 ), .B(n33172), .X(n19489) );
  nand_x1_sg U50608 ( .A(ow_12[4]), .B(n32586), .X(n19490) );
  nand_x1_sg U50609 ( .A(\shifter_0/n9583 ), .B(n29849), .X(n21761) );
  nand_x1_sg U50610 ( .A(ow_15[11]), .B(n34952), .X(n21762) );
  nand_x1_sg U50611 ( .A(\shifter_0/n9582 ), .B(n29845), .X(n21763) );
  nand_x1_sg U50612 ( .A(ow_15[10]), .B(n32627), .X(n21764) );
  nand_x1_sg U50613 ( .A(\shifter_0/n9581 ), .B(n31221), .X(n21765) );
  nand_x1_sg U50614 ( .A(ow_15[9]), .B(n34778), .X(n21766) );
  nand_x1_sg U50615 ( .A(\shifter_0/n9519 ), .B(n33138), .X(n21849) );
  nand_x1_sg U50616 ( .A(oi_1[7]), .B(n34766), .X(n21850) );
  nand_x1_sg U50617 ( .A(\shifter_0/n9518 ), .B(n33203), .X(n21851) );
  nand_x1_sg U50618 ( .A(oi_1[6]), .B(n32625), .X(n21852) );
  nand_x1_sg U50619 ( .A(\shifter_0/n9517 ), .B(n33189), .X(n21853) );
  nand_x1_sg U50620 ( .A(oi_1[5]), .B(n32567), .X(n21854) );
  nand_x1_sg U50621 ( .A(\shifter_0/n9159 ), .B(n30970), .X(n18761) );
  nand_x1_sg U50622 ( .A(oi_10[7]), .B(n30799), .X(n18762) );
  nand_x1_sg U50623 ( .A(\shifter_0/n9158 ), .B(n34985), .X(n18765) );
  nand_x1_sg U50624 ( .A(oi_10[6]), .B(n34764), .X(n18766) );
  nand_x1_sg U50625 ( .A(\shifter_0/n9157 ), .B(n29853), .X(n18767) );
  nand_x1_sg U50626 ( .A(oi_10[5]), .B(n34948), .X(n18768) );
  nand_x1_sg U50627 ( .A(\shifter_0/n9191 ), .B(n33150), .X(n19339) );
  nand_x1_sg U50628 ( .A(ow_9[19]), .B(n32095), .X(n19340) );
  nand_x1_sg U50629 ( .A(\shifter_0/n9190 ), .B(n33170), .X(n19341) );
  nand_x1_sg U50630 ( .A(ow_9[18]), .B(n32628), .X(n19342) );
  nand_x1_sg U50631 ( .A(\shifter_0/n9189 ), .B(n34974), .X(n19343) );
  nand_x1_sg U50632 ( .A(ow_9[17]), .B(n31932), .X(n19344) );
  nand_x1_sg U50633 ( .A(\shifter_0/n9580 ), .B(n34994), .X(n21767) );
  nand_x1_sg U50634 ( .A(ow_15[8]), .B(n32549), .X(n21768) );
  nand_x1_sg U50635 ( .A(\shifter_0/n9579 ), .B(n33184), .X(n21769) );
  nand_x1_sg U50636 ( .A(ow_15[7]), .B(n34761), .X(n21770) );
  nand_x1_sg U50637 ( .A(\shifter_0/n9578 ), .B(n33143), .X(n21771) );
  nand_x1_sg U50638 ( .A(ow_15[6]), .B(n34955), .X(n21772) );
  nand_x1_sg U50639 ( .A(\shifter_0/n9577 ), .B(n29863), .X(n21773) );
  nand_x1_sg U50640 ( .A(ow_15[5]), .B(n32584), .X(n21774) );
  nand_x1_sg U50641 ( .A(\shifter_0/n9576 ), .B(n31227), .X(n21775) );
  nand_x1_sg U50642 ( .A(ow_15[4]), .B(n32569), .X(n21776) );
  nand_x1_sg U50643 ( .A(\shifter_0/n9575 ), .B(n33135), .X(n21777) );
  nand_x1_sg U50644 ( .A(ow_15[3]), .B(n34764), .X(n21778) );
  nand_x1_sg U50645 ( .A(\shifter_0/n9574 ), .B(n34982), .X(n21779) );
  nand_x1_sg U50646 ( .A(ow_15[2]), .B(n32623), .X(n21780) );
  nand_x1_sg U50647 ( .A(\shifter_0/n9573 ), .B(n33201), .X(n21781) );
  nand_x1_sg U50648 ( .A(ow_15[1]), .B(n32598), .X(n21782) );
  nand_x1_sg U50649 ( .A(\shifter_0/n9572 ), .B(n31536), .X(n21783) );
  nand_x1_sg U50650 ( .A(ow_15[0]), .B(n32588), .X(n21784) );
  nand_x1_sg U50651 ( .A(\shifter_0/n9571 ), .B(n33173), .X(n21785) );
  nand_x1_sg U50652 ( .A(oi_0[19]), .B(n32556), .X(n21786) );
  nand_x1_sg U50653 ( .A(\shifter_0/n9570 ), .B(n34980), .X(n21787) );
  nand_x1_sg U50654 ( .A(oi_0[18]), .B(n32558), .X(n21788) );
  nand_x1_sg U50655 ( .A(\shifter_0/n9569 ), .B(n33177), .X(n21789) );
  nand_x1_sg U50656 ( .A(oi_0[17]), .B(n32551), .X(n21790) );
  nand_x1_sg U50657 ( .A(\shifter_0/n9568 ), .B(n29842), .X(n21791) );
  nand_x1_sg U50658 ( .A(oi_0[16]), .B(n32568), .X(n21792) );
  nand_x1_sg U50659 ( .A(\shifter_0/n9567 ), .B(n33212), .X(n21793) );
  nand_x1_sg U50660 ( .A(oi_0[15]), .B(n30799), .X(n21794) );
  nand_x1_sg U50661 ( .A(\shifter_0/n9566 ), .B(n31546), .X(n21795) );
  nand_x1_sg U50662 ( .A(oi_0[14]), .B(n34764), .X(n21796) );
  nand_x1_sg U50663 ( .A(\shifter_0/n9565 ), .B(n33175), .X(n21797) );
  nand_x1_sg U50664 ( .A(oi_0[13]), .B(n30657), .X(n21798) );
  nand_x1_sg U50665 ( .A(\shifter_0/n9564 ), .B(n35006), .X(n21799) );
  nand_x1_sg U50666 ( .A(oi_0[12]), .B(n32561), .X(n21800) );
  nand_x1_sg U50667 ( .A(\shifter_0/n9563 ), .B(n31542), .X(n21801) );
  nand_x1_sg U50668 ( .A(oi_0[11]), .B(n30796), .X(n21802) );
  nand_x1_sg U50669 ( .A(\shifter_0/n9562 ), .B(n33155), .X(n21803) );
  nand_x1_sg U50670 ( .A(oi_0[10]), .B(n30661), .X(n21804) );
  nand_x1_sg U50671 ( .A(\shifter_0/n9561 ), .B(n33161), .X(n21805) );
  nand_x1_sg U50672 ( .A(oi_0[9]), .B(n32577), .X(n21806) );
  nand_x1_sg U50673 ( .A(\shifter_0/n9560 ), .B(n33199), .X(n21807) );
  nand_x1_sg U50674 ( .A(oi_0[8]), .B(n34777), .X(n21808) );
  nand_x1_sg U50675 ( .A(\shifter_0/n9559 ), .B(n34977), .X(n21809) );
  nand_x1_sg U50676 ( .A(oi_0[7]), .B(n32551), .X(n21810) );
  nand_x1_sg U50677 ( .A(\shifter_0/n9558 ), .B(n33155), .X(n21811) );
  nand_x1_sg U50678 ( .A(oi_0[6]), .B(n32611), .X(n21812) );
  nand_x1_sg U50679 ( .A(\shifter_0/n9557 ), .B(n33187), .X(n21813) );
  nand_x1_sg U50680 ( .A(oi_0[5]), .B(n32548), .X(n21814) );
  nand_x1_sg U50681 ( .A(\shifter_0/n9556 ), .B(n30238), .X(n21815) );
  nand_x1_sg U50682 ( .A(oi_0[4]), .B(n32618), .X(n21816) );
  nand_x1_sg U50683 ( .A(\shifter_0/n9555 ), .B(n29851), .X(n21817) );
  nand_x1_sg U50684 ( .A(oi_0[3]), .B(n34794), .X(n21818) );
  nand_x1_sg U50685 ( .A(\shifter_0/n9554 ), .B(n31535), .X(n21819) );
  nand_x1_sg U50686 ( .A(oi_0[2]), .B(n34496), .X(n21820) );
  nand_x1_sg U50687 ( .A(\shifter_0/n9553 ), .B(n33145), .X(n21821) );
  nand_x1_sg U50688 ( .A(oi_0[1]), .B(n32603), .X(n21822) );
  nand_x1_sg U50689 ( .A(\shifter_0/n9552 ), .B(n34987), .X(n21823) );
  nand_x1_sg U50690 ( .A(oi_0[0]), .B(n30648), .X(n21824) );
  nand_x1_sg U50691 ( .A(\shifter_0/n9516 ), .B(n29867), .X(n21855) );
  nand_x1_sg U50692 ( .A(oi_1[4]), .B(n34493), .X(n21856) );
  nand_x1_sg U50693 ( .A(\shifter_0/n9515 ), .B(n31219), .X(n21857) );
  nand_x1_sg U50694 ( .A(oi_1[3]), .B(n32100), .X(n21858) );
  nand_x1_sg U50695 ( .A(\shifter_0/n9514 ), .B(n31222), .X(n21859) );
  nand_x1_sg U50696 ( .A(oi_1[2]), .B(n32589), .X(n21860) );
  nand_x1_sg U50697 ( .A(\shifter_0/n9513 ), .B(n31552), .X(n21861) );
  nand_x1_sg U50698 ( .A(oi_1[1]), .B(n30657), .X(n21862) );
  nand_x1_sg U50699 ( .A(\shifter_0/n9512 ), .B(n30970), .X(n21863) );
  nand_x1_sg U50700 ( .A(oi_1[0]), .B(n30653), .X(n21864) );
  nand_x1_sg U50701 ( .A(\shifter_0/n9491 ), .B(n31561), .X(n21865) );
  nand_x1_sg U50702 ( .A(oi_2[19]), .B(n32621), .X(n21866) );
  nand_x1_sg U50703 ( .A(\shifter_0/n9490 ), .B(n31541), .X(n21867) );
  nand_x1_sg U50704 ( .A(oi_2[18]), .B(n32598), .X(n21868) );
  nand_x1_sg U50705 ( .A(\shifter_0/n9489 ), .B(n33170), .X(n21869) );
  nand_x1_sg U50706 ( .A(oi_2[17]), .B(n34769), .X(n21870) );
  nand_x1_sg U50707 ( .A(\shifter_0/n9488 ), .B(n33157), .X(n21871) );
  nand_x1_sg U50708 ( .A(oi_2[16]), .B(n30673), .X(n21872) );
  nand_x1_sg U50709 ( .A(\shifter_0/n9487 ), .B(n33162), .X(n21873) );
  nand_x1_sg U50710 ( .A(oi_2[15]), .B(n32621), .X(n21874) );
  nand_x1_sg U50711 ( .A(\shifter_0/n9486 ), .B(n31542), .X(n21875) );
  nand_x1_sg U50712 ( .A(oi_2[14]), .B(n32569), .X(n21876) );
  nand_x1_sg U50713 ( .A(\shifter_0/n9485 ), .B(n33220), .X(n21877) );
  nand_x1_sg U50714 ( .A(oi_2[13]), .B(n34494), .X(n21878) );
  nand_x1_sg U50715 ( .A(\shifter_0/n9484 ), .B(n33176), .X(n21879) );
  nand_x1_sg U50716 ( .A(oi_2[12]), .B(n32621), .X(n21880) );
  nand_x1_sg U50717 ( .A(\shifter_0/n9483 ), .B(n33213), .X(n21881) );
  nand_x1_sg U50718 ( .A(oi_2[11]), .B(n32577), .X(n21882) );
  nand_x1_sg U50719 ( .A(\shifter_0/n9482 ), .B(n33180), .X(n21883) );
  nand_x1_sg U50720 ( .A(oi_2[10]), .B(n32611), .X(n21884) );
  nand_x1_sg U50721 ( .A(\shifter_0/n9481 ), .B(n30233), .X(n21885) );
  nand_x1_sg U50722 ( .A(oi_2[9]), .B(n32577), .X(n21886) );
  nand_x1_sg U50723 ( .A(\shifter_0/n9480 ), .B(n33197), .X(n21887) );
  nand_x1_sg U50724 ( .A(oi_2[8]), .B(n32604), .X(n21888) );
  nand_x1_sg U50725 ( .A(\shifter_0/n9439 ), .B(n33207), .X(n21929) );
  nand_x1_sg U50726 ( .A(oi_3[7]), .B(n32625), .X(n21930) );
  nand_x1_sg U50727 ( .A(\shifter_0/n9438 ), .B(n33188), .X(n21931) );
  nand_x1_sg U50728 ( .A(oi_3[6]), .B(n30796), .X(n21932) );
  nand_x1_sg U50729 ( .A(\shifter_0/n9437 ), .B(n34988), .X(n21933) );
  nand_x1_sg U50730 ( .A(oi_3[5]), .B(n32624), .X(n21934) );
  nand_x1_sg U50731 ( .A(\shifter_0/n9436 ), .B(n30234), .X(n21935) );
  nand_x1_sg U50732 ( .A(oi_3[4]), .B(n32549), .X(n21936) );
  nand_x1_sg U50733 ( .A(\shifter_0/n9435 ), .B(n33827), .X(n21937) );
  nand_x1_sg U50734 ( .A(oi_3[3]), .B(n32558), .X(n21938) );
  nand_x1_sg U50735 ( .A(\shifter_0/n9434 ), .B(n31540), .X(n21939) );
  nand_x1_sg U50736 ( .A(oi_3[2]), .B(n32586), .X(n21940) );
  nand_x1_sg U50737 ( .A(\shifter_0/n9433 ), .B(n29864), .X(n21941) );
  nand_x1_sg U50738 ( .A(oi_3[1]), .B(n32593), .X(n21942) );
  nand_x1_sg U50739 ( .A(\shifter_0/n9432 ), .B(n34986), .X(n21943) );
  nand_x1_sg U50740 ( .A(oi_3[0]), .B(n32600), .X(n21944) );
  nand_x1_sg U50741 ( .A(\shifter_0/n9411 ), .B(n33164), .X(n21945) );
  nand_x1_sg U50742 ( .A(oi_4[19]), .B(n30795), .X(n21946) );
  nand_x1_sg U50743 ( .A(\shifter_0/n9410 ), .B(n33211), .X(n21947) );
  nand_x1_sg U50744 ( .A(oi_4[18]), .B(n34759), .X(n21948) );
  nand_x1_sg U50745 ( .A(\shifter_0/n9409 ), .B(n29860), .X(n21949) );
  nand_x1_sg U50746 ( .A(oi_4[17]), .B(n34774), .X(n21950) );
  nand_x1_sg U50747 ( .A(\shifter_0/n9408 ), .B(n29844), .X(n21951) );
  nand_x1_sg U50748 ( .A(oi_4[16]), .B(n32604), .X(n21952) );
  nand_x1_sg U50749 ( .A(\shifter_0/n9355 ), .B(n34975), .X(n22017) );
  nand_x1_sg U50750 ( .A(oi_5[3]), .B(n32552), .X(n22018) );
  nand_x1_sg U50751 ( .A(\shifter_0/n9354 ), .B(n33218), .X(n22019) );
  nand_x1_sg U50752 ( .A(oi_5[2]), .B(n34794), .X(n22020) );
  nand_x1_sg U50753 ( .A(\shifter_0/n9353 ), .B(n33180), .X(n22021) );
  nand_x1_sg U50754 ( .A(oi_5[1]), .B(n32098), .X(n22022) );
  nand_x1_sg U50755 ( .A(\shifter_0/n9352 ), .B(n31547), .X(n22023) );
  nand_x1_sg U50756 ( .A(oi_5[0]), .B(n30674), .X(n22024) );
  nand_x1_sg U50757 ( .A(\shifter_0/n9331 ), .B(n31536), .X(n22025) );
  nand_x1_sg U50758 ( .A(oi_6[19]), .B(n32553), .X(n22026) );
  nand_x1_sg U50759 ( .A(\shifter_0/n9330 ), .B(n31222), .X(n22027) );
  nand_x1_sg U50760 ( .A(oi_6[18]), .B(n32562), .X(n22028) );
  nand_x1_sg U50761 ( .A(\shifter_0/n9329 ), .B(n33214), .X(n22029) );
  nand_x1_sg U50762 ( .A(oi_6[17]), .B(n34771), .X(n22030) );
  nand_x1_sg U50763 ( .A(\shifter_0/n9328 ), .B(n35005), .X(n22031) );
  nand_x1_sg U50764 ( .A(oi_6[16]), .B(n32100), .X(n22032) );
  nand_x1_sg U50765 ( .A(\shifter_0/n9327 ), .B(n29853), .X(n22033) );
  nand_x1_sg U50766 ( .A(oi_6[15]), .B(n34783), .X(n22034) );
  nand_x1_sg U50767 ( .A(\shifter_0/n9326 ), .B(n30222), .X(n22035) );
  nand_x1_sg U50768 ( .A(oi_6[14]), .B(n32617), .X(n22036) );
  nand_x1_sg U50769 ( .A(\shifter_0/n9325 ), .B(n33145), .X(n22037) );
  nand_x1_sg U50770 ( .A(oi_6[13]), .B(n34495), .X(n22038) );
  nand_x1_sg U50771 ( .A(\shifter_0/n9324 ), .B(n35009), .X(n22039) );
  nand_x1_sg U50772 ( .A(oi_6[12]), .B(n32632), .X(n22040) );
  nand_x1_sg U50773 ( .A(\shifter_0/n9323 ), .B(n31561), .X(n22041) );
  nand_x1_sg U50774 ( .A(oi_6[11]), .B(n34763), .X(n22042) );
  nand_x1_sg U50775 ( .A(\shifter_0/n9322 ), .B(n33185), .X(n22043) );
  nand_x1_sg U50776 ( .A(oi_6[10]), .B(n32561), .X(n22044) );
  nand_x1_sg U50777 ( .A(\shifter_0/n9321 ), .B(n30224), .X(n22045) );
  nand_x1_sg U50778 ( .A(oi_6[9]), .B(n32605), .X(n22046) );
  nand_x1_sg U50779 ( .A(\shifter_0/n9320 ), .B(n35008), .X(n22047) );
  nand_x1_sg U50780 ( .A(oi_6[8]), .B(n34758), .X(n22048) );
  nand_x1_sg U50781 ( .A(\shifter_0/n9279 ), .B(n35008), .X(n22089) );
  nand_x1_sg U50782 ( .A(oi_7[7]), .B(n32620), .X(n22090) );
  nand_x1_sg U50783 ( .A(\shifter_0/n9278 ), .B(n33141), .X(n22091) );
  nand_x1_sg U50784 ( .A(oi_7[6]), .B(n32587), .X(n22092) );
  nand_x1_sg U50785 ( .A(\shifter_0/n9277 ), .B(n33140), .X(n22093) );
  nand_x1_sg U50786 ( .A(oi_7[5]), .B(n32582), .X(n22094) );
  nand_x1_sg U50787 ( .A(\shifter_0/n9276 ), .B(n33190), .X(n22095) );
  nand_x1_sg U50788 ( .A(oi_7[4]), .B(n30796), .X(n22096) );
  nand_x1_sg U50789 ( .A(\shifter_0/n9275 ), .B(n30227), .X(n22097) );
  nand_x1_sg U50790 ( .A(oi_7[3]), .B(n32588), .X(n22098) );
  nand_x1_sg U50791 ( .A(\shifter_0/n9274 ), .B(n34984), .X(n22099) );
  nand_x1_sg U50792 ( .A(oi_7[2]), .B(n34947), .X(n22100) );
  nand_x1_sg U50793 ( .A(\shifter_0/n9273 ), .B(n33153), .X(n22101) );
  nand_x1_sg U50794 ( .A(oi_7[1]), .B(n34787), .X(n22102) );
  nand_x1_sg U50795 ( .A(\shifter_0/n9272 ), .B(n34996), .X(n22103) );
  nand_x1_sg U50796 ( .A(oi_7[0]), .B(n32605), .X(n22104) );
  nand_x1_sg U50797 ( .A(\shifter_0/n9251 ), .B(n34998), .X(n22105) );
  nand_x1_sg U50798 ( .A(oi_8[19]), .B(n32582), .X(n22106) );
  nand_x1_sg U50799 ( .A(\shifter_0/n9250 ), .B(n29864), .X(n22107) );
  nand_x1_sg U50800 ( .A(oi_8[18]), .B(n32598), .X(n22108) );
  nand_x1_sg U50801 ( .A(\shifter_0/n9249 ), .B(n33133), .X(n22109) );
  nand_x1_sg U50802 ( .A(oi_8[17]), .B(n32565), .X(n22110) );
  nand_x1_sg U50803 ( .A(\shifter_0/n9248 ), .B(n33168), .X(n22111) );
  nand_x1_sg U50804 ( .A(oi_8[16]), .B(n31930), .X(n22112) );
  nand_x1_sg U50805 ( .A(\shifter_0/n9247 ), .B(n33161), .X(n22113) );
  nand_x1_sg U50806 ( .A(oi_8[15]), .B(n30660), .X(n22114) );
  nand_x1_sg U50807 ( .A(\shifter_0/n9246 ), .B(n33191), .X(n22115) );
  nand_x1_sg U50808 ( .A(oi_8[14]), .B(n34788), .X(n22116) );
  nand_x1_sg U50809 ( .A(\shifter_0/n9245 ), .B(n30220), .X(n22117) );
  nand_x1_sg U50810 ( .A(oi_8[13]), .B(n32589), .X(n22118) );
  nand_x1_sg U50811 ( .A(\shifter_0/n9244 ), .B(n33218), .X(n22119) );
  nand_x1_sg U50812 ( .A(oi_8[12]), .B(n30798), .X(n22120) );
  nand_x1_sg U50813 ( .A(\shifter_0/n9243 ), .B(n33826), .X(n22121) );
  nand_x1_sg U50814 ( .A(oi_8[11]), .B(n32096), .X(n22122) );
  nand_x1_sg U50815 ( .A(\shifter_0/n9242 ), .B(n31536), .X(n22123) );
  nand_x1_sg U50816 ( .A(oi_8[10]), .B(n30676), .X(n22124) );
  nand_x1_sg U50817 ( .A(\shifter_0/n9241 ), .B(n34974), .X(n22125) );
  nand_x1_sg U50818 ( .A(oi_8[9]), .B(n34789), .X(n22126) );
  nand_x1_sg U50819 ( .A(\shifter_0/n9240 ), .B(n33220), .X(n22127) );
  nand_x1_sg U50820 ( .A(oi_8[8]), .B(n32632), .X(n22128) );
  nand_x1_sg U50821 ( .A(\shifter_0/n9239 ), .B(n30223), .X(n22129) );
  nand_x1_sg U50822 ( .A(oi_8[7]), .B(n32618), .X(n22130) );
  nand_x1_sg U50823 ( .A(\shifter_0/n9238 ), .B(n33207), .X(n22131) );
  nand_x1_sg U50824 ( .A(oi_8[6]), .B(n34494), .X(n22132) );
  nand_x1_sg U50825 ( .A(\shifter_0/n9237 ), .B(n34999), .X(n22133) );
  nand_x1_sg U50826 ( .A(oi_8[5]), .B(n32560), .X(n22134) );
  nand_x1_sg U50827 ( .A(\shifter_0/n9236 ), .B(n33168), .X(n22135) );
  nand_x1_sg U50828 ( .A(oi_8[4]), .B(n30649), .X(n22136) );
  nand_x1_sg U50829 ( .A(\shifter_0/n9235 ), .B(n33132), .X(n22137) );
  nand_x1_sg U50830 ( .A(oi_8[3]), .B(n31930), .X(n22138) );
  nand_x1_sg U50831 ( .A(\shifter_0/n9234 ), .B(n30226), .X(n22139) );
  nand_x1_sg U50832 ( .A(oi_8[2]), .B(n30661), .X(n22140) );
  nand_x1_sg U50833 ( .A(\shifter_0/n9233 ), .B(n33155), .X(n22141) );
  nand_x1_sg U50834 ( .A(oi_8[1]), .B(n34772), .X(n22142) );
  nand_x1_sg U50835 ( .A(\shifter_0/n9232 ), .B(n33154), .X(n22143) );
  nand_x1_sg U50836 ( .A(oi_8[0]), .B(n32608), .X(n22144) );
  nand_x1_sg U50837 ( .A(\shifter_0/n9211 ), .B(n34979), .X(n22145) );
  nand_x1_sg U50838 ( .A(oi_9[19]), .B(n32550), .X(n22146) );
  nand_x1_sg U50839 ( .A(\shifter_0/n9210 ), .B(n30230), .X(n22147) );
  nand_x1_sg U50840 ( .A(oi_9[18]), .B(n32552), .X(n22148) );
  nand_x1_sg U50841 ( .A(\shifter_0/n9209 ), .B(n30970), .X(n22149) );
  nand_x1_sg U50842 ( .A(oi_9[17]), .B(n32627), .X(n22150) );
  nand_x1_sg U50843 ( .A(\shifter_0/n9208 ), .B(n34998), .X(n22151) );
  nand_x1_sg U50844 ( .A(oi_9[16]), .B(n34784), .X(n22152) );
  nand_x1_sg U50845 ( .A(\shifter_0/n9207 ), .B(n35004), .X(n22153) );
  nand_x1_sg U50846 ( .A(oi_9[15]), .B(n30676), .X(n22154) );
  nand_x1_sg U50847 ( .A(\shifter_0/n9206 ), .B(n33184), .X(n22155) );
  nand_x1_sg U50848 ( .A(oi_9[14]), .B(n34786), .X(n22156) );
  nand_x1_sg U50849 ( .A(\shifter_0/n9205 ), .B(n33188), .X(n22157) );
  nand_x1_sg U50850 ( .A(oi_9[13]), .B(n34945), .X(n22158) );
  nand_x1_sg U50851 ( .A(\shifter_0/n9204 ), .B(n29839), .X(n22159) );
  nand_x1_sg U50852 ( .A(oi_9[12]), .B(n34758), .X(n22160) );
  nand_x1_sg U50853 ( .A(\shifter_0/n9203 ), .B(n34976), .X(n22161) );
  nand_x1_sg U50854 ( .A(oi_9[11]), .B(n30652), .X(n22162) );
  nand_x1_sg U50855 ( .A(\shifter_0/n9202 ), .B(n35004), .X(n22163) );
  nand_x1_sg U50856 ( .A(oi_9[10]), .B(n32628), .X(n22164) );
  nand_x1_sg U50857 ( .A(\shifter_0/n9201 ), .B(n35000), .X(n22165) );
  nand_x1_sg U50858 ( .A(oi_9[9]), .B(n34946), .X(n22166) );
  nand_x1_sg U50859 ( .A(\shifter_0/n9200 ), .B(n33185), .X(n22167) );
  nand_x1_sg U50860 ( .A(oi_9[8]), .B(n34778), .X(n22168) );
  nand_x1_sg U50861 ( .A(\shifter_0/n9199 ), .B(n29842), .X(n22169) );
  nand_x1_sg U50862 ( .A(oi_9[7]), .B(n34788), .X(n22170) );
  nand_x1_sg U50863 ( .A(\shifter_0/n9198 ), .B(n33171), .X(n22171) );
  nand_x1_sg U50864 ( .A(oi_9[6]), .B(n32567), .X(n22172) );
  nand_x1_sg U50865 ( .A(\shifter_0/n9197 ), .B(n29849), .X(n22173) );
  nand_x1_sg U50866 ( .A(oi_9[5]), .B(n30659), .X(n22174) );
  nand_x1_sg U50867 ( .A(\shifter_0/n9196 ), .B(n33147), .X(n22175) );
  nand_x1_sg U50868 ( .A(oi_9[4]), .B(n30610), .X(n22176) );
  nand_x1_sg U50869 ( .A(\shifter_0/n9195 ), .B(n35003), .X(n22177) );
  nand_x1_sg U50870 ( .A(oi_9[3]), .B(n32557), .X(n22178) );
  nand_x1_sg U50871 ( .A(\shifter_0/n9194 ), .B(n35000), .X(n22179) );
  nand_x1_sg U50872 ( .A(oi_9[2]), .B(n32094), .X(n22180) );
  nand_x1_sg U50873 ( .A(\shifter_0/n9193 ), .B(n31538), .X(n22181) );
  nand_x1_sg U50874 ( .A(oi_9[1]), .B(n34793), .X(n22182) );
  nand_x1_sg U50875 ( .A(\shifter_0/n9192 ), .B(n33165), .X(n22183) );
  nand_x1_sg U50876 ( .A(oi_9[0]), .B(n34947), .X(n22184) );
  nand_x1_sg U50877 ( .A(\shifter_0/n9171 ), .B(n31553), .X(n22185) );
  nand_x1_sg U50878 ( .A(oi_10[19]), .B(n32596), .X(n22186) );
  nand_x1_sg U50879 ( .A(\shifter_0/n9170 ), .B(n29860), .X(n22187) );
  nand_x1_sg U50880 ( .A(oi_10[18]), .B(n32598), .X(n22188) );
  nand_x1_sg U50881 ( .A(\shifter_0/n9169 ), .B(n31551), .X(n22189) );
  nand_x1_sg U50882 ( .A(oi_10[17]), .B(n34763), .X(n22190) );
  nand_x1_sg U50883 ( .A(\shifter_0/n9168 ), .B(n33140), .X(n22191) );
  nand_x1_sg U50884 ( .A(oi_10[16]), .B(n31929), .X(n22192) );
  nand_x1_sg U50885 ( .A(\shifter_0/n9167 ), .B(n33137), .X(n22193) );
  nand_x1_sg U50886 ( .A(oi_10[15]), .B(n34766), .X(n22194) );
  nand_x1_sg U50887 ( .A(\shifter_0/n9166 ), .B(n29863), .X(n22195) );
  nand_x1_sg U50888 ( .A(oi_10[14]), .B(n32568), .X(n22196) );
  nand_x1_sg U50889 ( .A(\shifter_0/n9165 ), .B(n33209), .X(n22197) );
  nand_x1_sg U50890 ( .A(oi_10[13]), .B(n32546), .X(n22198) );
  nand_x1_sg U50891 ( .A(\shifter_0/n9164 ), .B(n29850), .X(n22199) );
  nand_x1_sg U50892 ( .A(oi_10[12]), .B(n32563), .X(n22200) );
  nand_x1_sg U50893 ( .A(\shifter_0/n9163 ), .B(n33189), .X(n22201) );
  nand_x1_sg U50894 ( .A(oi_10[11]), .B(n32612), .X(n22202) );
  nand_x1_sg U50895 ( .A(\shifter_0/n9162 ), .B(n33135), .X(n22203) );
  nand_x1_sg U50896 ( .A(oi_10[10]), .B(n32570), .X(n22204) );
  nand_x1_sg U50897 ( .A(\shifter_0/n9161 ), .B(n33190), .X(n22205) );
  nand_x1_sg U50898 ( .A(oi_10[9]), .B(n34954), .X(n22206) );
  nand_x1_sg U50899 ( .A(\shifter_0/n9160 ), .B(n31223), .X(n22207) );
  nand_x1_sg U50900 ( .A(oi_10[8]), .B(n32633), .X(n22208) );
  nand_x1_sg U50901 ( .A(\shifter_0/n9156 ), .B(n33175), .X(n18769) );
  nand_x1_sg U50902 ( .A(oi_10[4]), .B(n32616), .X(n18770) );
  nand_x1_sg U50903 ( .A(\shifter_0/n9155 ), .B(n33218), .X(n18771) );
  nand_x1_sg U50904 ( .A(oi_10[3]), .B(n32579), .X(n18772) );
  nand_x1_sg U50905 ( .A(\shifter_0/n9154 ), .B(n33156), .X(n18773) );
  nand_x1_sg U50906 ( .A(oi_10[2]), .B(n32580), .X(n18774) );
  nand_x1_sg U50907 ( .A(\shifter_0/n9153 ), .B(n31555), .X(n18775) );
  nand_x1_sg U50908 ( .A(oi_10[1]), .B(n34762), .X(n18776) );
  nand_x1_sg U50909 ( .A(\shifter_0/n9152 ), .B(n34995), .X(n18777) );
  nand_x1_sg U50910 ( .A(oi_10[0]), .B(n32096), .X(n18778) );
  nand_x1_sg U50911 ( .A(\shifter_0/n9131 ), .B(n33144), .X(n18779) );
  nand_x1_sg U50912 ( .A(oi_11[19]), .B(n32099), .X(n18780) );
  nand_x1_sg U50913 ( .A(\shifter_0/n9130 ), .B(n33220), .X(n18781) );
  nand_x1_sg U50914 ( .A(oi_11[18]), .B(n32555), .X(n18782) );
  nand_x1_sg U50915 ( .A(\shifter_0/n9129 ), .B(n33825), .X(n18783) );
  nand_x1_sg U50916 ( .A(oi_11[17]), .B(n30669), .X(n18784) );
  nand_x1_sg U50917 ( .A(\shifter_0/n9128 ), .B(n31535), .X(n18785) );
  nand_x1_sg U50918 ( .A(oi_11[16]), .B(n32616), .X(n18786) );
  nand_x1_sg U50919 ( .A(\shifter_0/n9127 ), .B(n31548), .X(n18787) );
  nand_x1_sg U50920 ( .A(oi_11[15]), .B(n32610), .X(n18788) );
  nand_x1_sg U50921 ( .A(\shifter_0/n9126 ), .B(n33149), .X(n18789) );
  nand_x1_sg U50922 ( .A(oi_11[14]), .B(n30661), .X(n18790) );
  nand_x1_sg U50923 ( .A(\shifter_0/n9125 ), .B(n33171), .X(n18791) );
  nand_x1_sg U50924 ( .A(oi_11[13]), .B(n32586), .X(n18792) );
  nand_x1_sg U50925 ( .A(\shifter_0/n9124 ), .B(n33196), .X(n18793) );
  nand_x1_sg U50926 ( .A(oi_11[12]), .B(n32548), .X(n18794) );
  nand_x1_sg U50927 ( .A(\shifter_0/n9123 ), .B(n33212), .X(n18795) );
  nand_x1_sg U50928 ( .A(oi_11[11]), .B(n32557), .X(n18796) );
  nand_x1_sg U50929 ( .A(\shifter_0/n9122 ), .B(n33163), .X(n18797) );
  nand_x1_sg U50930 ( .A(oi_11[10]), .B(n31932), .X(n18798) );
  nand_x1_sg U50931 ( .A(\shifter_0/n9121 ), .B(n33189), .X(n18799) );
  nand_x1_sg U50932 ( .A(oi_11[9]), .B(n30795), .X(n18800) );
  nand_x1_sg U50933 ( .A(\shifter_0/n9120 ), .B(n34981), .X(n18801) );
  nand_x1_sg U50934 ( .A(oi_11[8]), .B(n34498), .X(n18802) );
  nand_x1_sg U50935 ( .A(\shifter_0/n9079 ), .B(n33153), .X(n18843) );
  nand_x1_sg U50936 ( .A(oi_12[7]), .B(n30678), .X(n18844) );
  nand_x1_sg U50937 ( .A(\shifter_0/n9078 ), .B(n31225), .X(n18845) );
  nand_x1_sg U50938 ( .A(oi_12[6]), .B(n32563), .X(n18846) );
  nand_x1_sg U50939 ( .A(\shifter_0/n9077 ), .B(n33160), .X(n18847) );
  nand_x1_sg U50940 ( .A(oi_12[5]), .B(n32600), .X(n18848) );
  nand_x1_sg U50941 ( .A(\shifter_0/n9076 ), .B(n31226), .X(n18849) );
  nand_x1_sg U50942 ( .A(oi_12[4]), .B(n32573), .X(n18850) );
  nand_x1_sg U50943 ( .A(\shifter_0/n9075 ), .B(n35000), .X(n18851) );
  nand_x1_sg U50944 ( .A(oi_12[3]), .B(n30665), .X(n18852) );
  nand_x1_sg U50945 ( .A(\shifter_0/n9074 ), .B(n31538), .X(n18853) );
  nand_x1_sg U50946 ( .A(oi_12[2]), .B(n32604), .X(n18854) );
  nand_x1_sg U50947 ( .A(\shifter_0/n9073 ), .B(n33145), .X(n18855) );
  nand_x1_sg U50948 ( .A(oi_12[1]), .B(n32560), .X(n18856) );
  nand_x1_sg U50949 ( .A(\shifter_0/n9072 ), .B(n33209), .X(n18857) );
  nand_x1_sg U50950 ( .A(oi_12[0]), .B(n32603), .X(n18858) );
  nand_x1_sg U50951 ( .A(\shifter_0/n9051 ), .B(n35005), .X(n18859) );
  nand_x1_sg U50952 ( .A(oi_13[19]), .B(n34773), .X(n18860) );
  nand_x1_sg U50953 ( .A(\shifter_0/n9050 ), .B(n31222), .X(n18861) );
  nand_x1_sg U50954 ( .A(oi_13[18]), .B(n30667), .X(n18862) );
  nand_x1_sg U50955 ( .A(\shifter_0/n9049 ), .B(n33215), .X(n18863) );
  nand_x1_sg U50956 ( .A(oi_13[17]), .B(n34788), .X(n18864) );
  nand_x1_sg U50957 ( .A(\shifter_0/n9048 ), .B(n29864), .X(n18865) );
  nand_x1_sg U50958 ( .A(oi_13[16]), .B(n32561), .X(n18866) );
  nand_x1_sg U50959 ( .A(\shifter_0/n9047 ), .B(n33196), .X(n18867) );
  nand_x1_sg U50960 ( .A(oi_13[15]), .B(n34757), .X(n18868) );
  nand_x1_sg U50961 ( .A(\shifter_0/n9046 ), .B(n29845), .X(n18869) );
  nand_x1_sg U50962 ( .A(oi_13[14]), .B(n32588), .X(n18870) );
  nand_x1_sg U50963 ( .A(\shifter_0/n9045 ), .B(n33191), .X(n18871) );
  nand_x1_sg U50964 ( .A(oi_13[13]), .B(n34793), .X(n18872) );
  nand_x1_sg U50965 ( .A(\shifter_0/n9044 ), .B(n31223), .X(n18873) );
  nand_x1_sg U50966 ( .A(oi_13[12]), .B(n32620), .X(n18874) );
  nand_x1_sg U50967 ( .A(\shifter_0/n9043 ), .B(n33192), .X(n18875) );
  nand_x1_sg U50968 ( .A(oi_13[11]), .B(n34500), .X(n18876) );
  nand_x1_sg U50969 ( .A(\shifter_0/n9042 ), .B(n30231), .X(n18877) );
  nand_x1_sg U50970 ( .A(oi_13[10]), .B(n32585), .X(n18878) );
  nand_x1_sg U50971 ( .A(\shifter_0/n9041 ), .B(n34998), .X(n18879) );
  nand_x1_sg U50972 ( .A(oi_13[9]), .B(n32612), .X(n18880) );
  nand_x1_sg U50973 ( .A(\shifter_0/n9040 ), .B(n33219), .X(n18881) );
  nand_x1_sg U50974 ( .A(oi_13[8]), .B(n32552), .X(n18882) );
  nand_x1_sg U50975 ( .A(\shifter_0/n9039 ), .B(n34989), .X(n18883) );
  nand_x1_sg U50976 ( .A(oi_13[7]), .B(n32553), .X(n18884) );
  nand_x1_sg U50977 ( .A(\shifter_0/n9038 ), .B(n30231), .X(n18885) );
  nand_x1_sg U50978 ( .A(oi_13[6]), .B(n32615), .X(n18886) );
  nand_x1_sg U50979 ( .A(\shifter_0/n9037 ), .B(n35006), .X(n18887) );
  nand_x1_sg U50980 ( .A(oi_13[5]), .B(n34498), .X(n18888) );
  nand_x1_sg U50981 ( .A(\shifter_0/n9036 ), .B(n31537), .X(n18889) );
  nand_x1_sg U50982 ( .A(oi_13[4]), .B(n32576), .X(n18890) );
  nand_x1_sg U50983 ( .A(\shifter_0/n8966 ), .B(n33187), .X(n18949) );
  nand_x1_sg U50984 ( .A(oi_15[14]), .B(n30677), .X(n18950) );
  nand_x1_sg U50985 ( .A(\shifter_0/n8965 ), .B(n29856), .X(n18951) );
  nand_x1_sg U50986 ( .A(oi_15[13]), .B(n34772), .X(n18952) );
  nand_x1_sg U50987 ( .A(\shifter_0/n8964 ), .B(n33167), .X(n18953) );
  nand_x1_sg U50988 ( .A(oi_15[12]), .B(n32098), .X(n18954) );
  nand_x1_sg U50989 ( .A(\shifter_0/n9499 ), .B(n33137), .X(n19043) );
  nand_x1_sg U50990 ( .A(ow_1[7]), .B(n34953), .X(n19044) );
  nand_x1_sg U50991 ( .A(\shifter_0/n9498 ), .B(n33197), .X(n19045) );
  nand_x1_sg U50992 ( .A(ow_1[6]), .B(n34782), .X(n19046) );
  nand_x1_sg U50993 ( .A(\shifter_0/n9497 ), .B(n31548), .X(n19047) );
  nand_x1_sg U50994 ( .A(ow_1[5]), .B(n34951), .X(n19048) );
  nand_x1_sg U50995 ( .A(\shifter_0/n9496 ), .B(n31555), .X(n19049) );
  nand_x1_sg U50996 ( .A(ow_1[4]), .B(n34766), .X(n19050) );
  nand_x1_sg U50997 ( .A(\shifter_0/n9495 ), .B(n33213), .X(n19051) );
  nand_x1_sg U50998 ( .A(ow_1[3]), .B(n30648), .X(n19052) );
  nand_x1_sg U50999 ( .A(\shifter_0/n9494 ), .B(n29856), .X(n19053) );
  nand_x1_sg U51000 ( .A(ow_1[2]), .B(n32605), .X(n19054) );
  nand_x1_sg U51001 ( .A(\shifter_0/n9493 ), .B(n34997), .X(n19055) );
  nand_x1_sg U51002 ( .A(ow_1[1]), .B(n32587), .X(n19056) );
  nand_x1_sg U51003 ( .A(\shifter_0/n9492 ), .B(n34998), .X(n19057) );
  nand_x1_sg U51004 ( .A(ow_1[0]), .B(n32628), .X(n19058) );
  nand_x1_sg U51005 ( .A(\shifter_0/n9471 ), .B(n33150), .X(n19059) );
  nand_x1_sg U51006 ( .A(ow_2[19]), .B(n34767), .X(n19060) );
  nand_x1_sg U51007 ( .A(\shifter_0/n9470 ), .B(n33825), .X(n19061) );
  nand_x1_sg U51008 ( .A(ow_2[18]), .B(n34501), .X(n19062) );
  nand_x1_sg U51009 ( .A(\shifter_0/n9469 ), .B(n30224), .X(n19063) );
  nand_x1_sg U51010 ( .A(ow_2[17]), .B(n32541), .X(n19064) );
  nand_x1_sg U51011 ( .A(\shifter_0/n9468 ), .B(n33152), .X(n19065) );
  nand_x1_sg U51012 ( .A(ow_2[16]), .B(n32574), .X(n19066) );
  nand_x1_sg U51013 ( .A(\shifter_0/n9467 ), .B(n31223), .X(n19067) );
  nand_x1_sg U51014 ( .A(ow_2[15]), .B(n30124), .X(n19068) );
  nand_x1_sg U51015 ( .A(\shifter_0/n9466 ), .B(n34994), .X(n19069) );
  nand_x1_sg U51016 ( .A(ow_2[14]), .B(n32610), .X(n19070) );
  nand_x1_sg U51017 ( .A(\shifter_0/n9465 ), .B(n33206), .X(n19071) );
  nand_x1_sg U51018 ( .A(ow_2[13]), .B(n32608), .X(n19072) );
  nand_x1_sg U51019 ( .A(\shifter_0/n9464 ), .B(n31551), .X(n19073) );
  nand_x1_sg U51020 ( .A(ow_2[12]), .B(n32627), .X(n19074) );
  nand_x1_sg U51021 ( .A(\shifter_0/n9463 ), .B(n34997), .X(n19075) );
  nand_x1_sg U51022 ( .A(ow_2[11]), .B(n30647), .X(n19076) );
  nand_x1_sg U51023 ( .A(\shifter_0/n9462 ), .B(n33826), .X(n19077) );
  nand_x1_sg U51024 ( .A(ow_2[10]), .B(n30214), .X(n19078) );
  nand_x1_sg U51025 ( .A(\shifter_0/n9461 ), .B(n33147), .X(n19079) );
  nand_x1_sg U51026 ( .A(ow_2[9]), .B(n32616), .X(n19080) );
  nand_x1_sg U51027 ( .A(\shifter_0/n9460 ), .B(n29853), .X(n19081) );
  nand_x1_sg U51028 ( .A(ow_2[8]), .B(n32601), .X(n19082) );
  nand_x1_sg U51029 ( .A(\shifter_0/n9419 ), .B(n33172), .X(n19123) );
  nand_x1_sg U51030 ( .A(ow_3[7]), .B(n34949), .X(n19124) );
  nand_x1_sg U51031 ( .A(\shifter_0/n9418 ), .B(n30971), .X(n19125) );
  nand_x1_sg U51032 ( .A(ow_3[6]), .B(n34946), .X(n19126) );
  nand_x1_sg U51033 ( .A(\shifter_0/n9417 ), .B(n30238), .X(n19127) );
  nand_x1_sg U51034 ( .A(ow_3[5]), .B(n30651), .X(n19128) );
  nand_x1_sg U51035 ( .A(\shifter_0/n9416 ), .B(n33824), .X(n19129) );
  nand_x1_sg U51036 ( .A(ow_3[4]), .B(n30678), .X(n19130) );
  nand_x1_sg U51037 ( .A(\shifter_0/n9415 ), .B(n33202), .X(n19131) );
  nand_x1_sg U51038 ( .A(ow_3[3]), .B(n32094), .X(n19132) );
  nand_x1_sg U51039 ( .A(\shifter_0/n9414 ), .B(n34982), .X(n19133) );
  nand_x1_sg U51040 ( .A(ow_3[2]), .B(n34495), .X(n19134) );
  nand_x1_sg U51041 ( .A(\shifter_0/n9413 ), .B(n31561), .X(n19135) );
  nand_x1_sg U51042 ( .A(ow_3[1]), .B(n30647), .X(n19136) );
  nand_x1_sg U51043 ( .A(\shifter_0/n9412 ), .B(n34977), .X(n19137) );
  nand_x1_sg U51044 ( .A(ow_3[0]), .B(n30798), .X(n19138) );
  nand_x1_sg U51045 ( .A(\shifter_0/n9391 ), .B(n33179), .X(n19139) );
  nand_x1_sg U51046 ( .A(ow_4[19]), .B(n30678), .X(n19140) );
  nand_x1_sg U51047 ( .A(\shifter_0/n9390 ), .B(n33148), .X(n19141) );
  nand_x1_sg U51048 ( .A(ow_4[18]), .B(n34781), .X(n19142) );
  nand_x1_sg U51049 ( .A(\shifter_0/n9389 ), .B(n29847), .X(n19143) );
  nand_x1_sg U51050 ( .A(ow_4[17]), .B(n34781), .X(n19144) );
  nand_x1_sg U51051 ( .A(\shifter_0/n9388 ), .B(n33202), .X(n19145) );
  nand_x1_sg U51052 ( .A(ow_4[16]), .B(n32576), .X(n19146) );
  nand_x1_sg U51053 ( .A(\shifter_0/n9387 ), .B(n29844), .X(n19147) );
  nand_x1_sg U51054 ( .A(ow_4[15]), .B(n30652), .X(n19148) );
  nand_x1_sg U51055 ( .A(\shifter_0/n9386 ), .B(n31546), .X(n19149) );
  nand_x1_sg U51056 ( .A(ow_4[14]), .B(n32609), .X(n19150) );
  nand_x1_sg U51057 ( .A(\shifter_0/n9385 ), .B(n33194), .X(n19151) );
  nand_x1_sg U51058 ( .A(ow_4[13]), .B(n32622), .X(n19152) );
  nand_x1_sg U51059 ( .A(\shifter_0/n9384 ), .B(n31223), .X(n19153) );
  nand_x1_sg U51060 ( .A(ow_4[12]), .B(n32613), .X(n19154) );
  nand_x1_sg U51061 ( .A(\shifter_0/n9383 ), .B(n33196), .X(n19155) );
  nand_x1_sg U51062 ( .A(ow_4[11]), .B(n31929), .X(n19156) );
  nand_x1_sg U51063 ( .A(\shifter_0/n9382 ), .B(n33204), .X(n19157) );
  nand_x1_sg U51064 ( .A(ow_4[10]), .B(n34774), .X(n19158) );
  nand_x1_sg U51065 ( .A(\shifter_0/n9381 ), .B(n29846), .X(n19159) );
  nand_x1_sg U51066 ( .A(ow_4[9]), .B(n32549), .X(n19160) );
  nand_x1_sg U51067 ( .A(\shifter_0/n9380 ), .B(n33165), .X(n19161) );
  nand_x1_sg U51068 ( .A(ow_4[8]), .B(n34768), .X(n19162) );
  nand_x1_sg U51069 ( .A(\shifter_0/n9339 ), .B(n33172), .X(n19203) );
  nand_x1_sg U51070 ( .A(ow_5[7]), .B(n32540), .X(n19204) );
  nand_x1_sg U51071 ( .A(\shifter_0/n9338 ), .B(n33138), .X(n19205) );
  nand_x1_sg U51072 ( .A(ow_5[6]), .B(n32560), .X(n19206) );
  nand_x1_sg U51073 ( .A(\shifter_0/n9337 ), .B(n33153), .X(n19207) );
  nand_x1_sg U51074 ( .A(ow_5[5]), .B(n32540), .X(n19208) );
  nand_x1_sg U51075 ( .A(\shifter_0/n9336 ), .B(n33170), .X(n19209) );
  nand_x1_sg U51076 ( .A(ow_5[4]), .B(n32624), .X(n19210) );
  nand_x1_sg U51077 ( .A(\shifter_0/n9263 ), .B(n33153), .X(n19275) );
  nand_x1_sg U51078 ( .A(ow_7[11]), .B(n30674), .X(n19276) );
  nand_x1_sg U51079 ( .A(\shifter_0/n9262 ), .B(n31220), .X(n19277) );
  nand_x1_sg U51080 ( .A(ow_7[10]), .B(n32610), .X(n19278) );
  nand_x1_sg U51081 ( .A(\shifter_0/n9261 ), .B(n29850), .X(n19279) );
  nand_x1_sg U51082 ( .A(ow_7[9]), .B(n32098), .X(n19280) );
  nand_x1_sg U51083 ( .A(\shifter_0/n9260 ), .B(n33147), .X(n19281) );
  nand_x1_sg U51084 ( .A(ow_7[8]), .B(n34773), .X(n19282) );
  nand_x1_sg U51085 ( .A(\shifter_0/n9259 ), .B(n33206), .X(n19283) );
  nand_x1_sg U51086 ( .A(ow_7[7]), .B(n32608), .X(n19284) );
  nand_x1_sg U51087 ( .A(\shifter_0/n9258 ), .B(n34989), .X(n19285) );
  nand_x1_sg U51088 ( .A(ow_7[6]), .B(n32599), .X(n19286) );
  nand_x1_sg U51089 ( .A(\shifter_0/n9257 ), .B(n34984), .X(n19287) );
  nand_x1_sg U51090 ( .A(ow_7[5]), .B(n34771), .X(n19288) );
  nand_x1_sg U51091 ( .A(\shifter_0/n9256 ), .B(n29847), .X(n19289) );
  nand_x1_sg U51092 ( .A(ow_7[4]), .B(n34761), .X(n19290) );
  nand_x1_sg U51093 ( .A(\shifter_0/n9255 ), .B(n34984), .X(n19291) );
  nand_x1_sg U51094 ( .A(ow_7[3]), .B(n32555), .X(n19292) );
  nand_x1_sg U51095 ( .A(\shifter_0/n9254 ), .B(n34995), .X(n19293) );
  nand_x1_sg U51096 ( .A(ow_7[2]), .B(n31931), .X(n19294) );
  nand_x1_sg U51097 ( .A(\shifter_0/n9253 ), .B(n29864), .X(n19295) );
  nand_x1_sg U51098 ( .A(ow_7[1]), .B(n32603), .X(n19296) );
  nand_x1_sg U51099 ( .A(\shifter_0/n9252 ), .B(n33141), .X(n19297) );
  nand_x1_sg U51100 ( .A(ow_7[0]), .B(n30676), .X(n19298) );
  nand_x1_sg U51101 ( .A(\shifter_0/n9231 ), .B(n29839), .X(n19299) );
  nand_x1_sg U51102 ( .A(ow_8[19]), .B(n32592), .X(n19300) );
  nand_x1_sg U51103 ( .A(\shifter_0/n9230 ), .B(n34975), .X(n19301) );
  nand_x1_sg U51104 ( .A(ow_8[18]), .B(n30796), .X(n19302) );
  nand_x1_sg U51105 ( .A(\shifter_0/n9229 ), .B(n34980), .X(n19303) );
  nand_x1_sg U51106 ( .A(ow_8[17]), .B(n32615), .X(n19304) );
  nand_x1_sg U51107 ( .A(\shifter_0/n9228 ), .B(n29857), .X(n19305) );
  nand_x1_sg U51108 ( .A(ow_8[16]), .B(n32580), .X(n19306) );
  nand_x1_sg U51109 ( .A(\shifter_0/n9227 ), .B(n33175), .X(n19307) );
  nand_x1_sg U51110 ( .A(ow_8[15]), .B(n32099), .X(n19308) );
  nand_x1_sg U51111 ( .A(\shifter_0/n9226 ), .B(n29844), .X(n19309) );
  nand_x1_sg U51112 ( .A(ow_8[14]), .B(n32610), .X(n19310) );
  nand_x1_sg U51113 ( .A(\shifter_0/n9225 ), .B(n33159), .X(n19311) );
  nand_x1_sg U51114 ( .A(ow_8[13]), .B(n32568), .X(n19312) );
  nand_x1_sg U51115 ( .A(\shifter_0/n9224 ), .B(n33143), .X(n19313) );
  nand_x1_sg U51116 ( .A(ow_8[12]), .B(n32095), .X(n19314) );
  nand_x1_sg U51117 ( .A(\shifter_0/n9223 ), .B(n35007), .X(n19315) );
  nand_x1_sg U51118 ( .A(ow_8[11]), .B(n32630), .X(n19316) );
  nand_x1_sg U51119 ( .A(\shifter_0/n9222 ), .B(n33188), .X(n19317) );
  nand_x1_sg U51120 ( .A(ow_8[10]), .B(n32574), .X(n19318) );
  nand_x1_sg U51121 ( .A(\shifter_0/n9221 ), .B(n33177), .X(n19319) );
  nand_x1_sg U51122 ( .A(ow_8[9]), .B(n30677), .X(n19320) );
  nand_x1_sg U51123 ( .A(\shifter_0/n9220 ), .B(n30233), .X(n19321) );
  nand_x1_sg U51124 ( .A(ow_8[8]), .B(n32544), .X(n19322) );
  nand_x1_sg U51125 ( .A(\shifter_0/n9219 ), .B(n33208), .X(n19323) );
  nand_x1_sg U51126 ( .A(ow_8[7]), .B(n34767), .X(n19324) );
  nand_x1_sg U51127 ( .A(\shifter_0/n9218 ), .B(n29857), .X(n19325) );
  nand_x1_sg U51128 ( .A(ow_8[6]), .B(n32634), .X(n19326) );
  nand_x1_sg U51129 ( .A(\shifter_0/n9217 ), .B(n33154), .X(n19327) );
  nand_x1_sg U51130 ( .A(ow_8[5]), .B(n34946), .X(n19328) );
  nand_x1_sg U51131 ( .A(\shifter_0/n9216 ), .B(n33142), .X(n19329) );
  nand_x1_sg U51132 ( .A(ow_8[4]), .B(n32567), .X(n19330) );
  nand_x1_sg U51133 ( .A(\shifter_0/n9215 ), .B(n33201), .X(n19331) );
  nand_x1_sg U51134 ( .A(ow_8[3]), .B(n32099), .X(n19332) );
  nand_x1_sg U51135 ( .A(\shifter_0/n9214 ), .B(n34976), .X(n19333) );
  nand_x1_sg U51136 ( .A(ow_8[2]), .B(n32596), .X(n19334) );
  nand_x1_sg U51137 ( .A(\shifter_0/n9213 ), .B(n33132), .X(n19335) );
  nand_x1_sg U51138 ( .A(ow_8[1]), .B(n32569), .X(n19336) );
  nand_x1_sg U51139 ( .A(\shifter_0/n9212 ), .B(n33133), .X(n19337) );
  nand_x1_sg U51140 ( .A(ow_8[0]), .B(n32634), .X(n19338) );
  nand_x1_sg U51141 ( .A(\shifter_0/n9188 ), .B(n33191), .X(n19345) );
  nand_x1_sg U51142 ( .A(ow_9[16]), .B(n30651), .X(n19346) );
  nand_x1_sg U51143 ( .A(\shifter_0/n9187 ), .B(n34979), .X(n19347) );
  nand_x1_sg U51144 ( .A(ow_9[15]), .B(n32606), .X(n19348) );
  nand_x1_sg U51145 ( .A(\shifter_0/n9186 ), .B(n30971), .X(n19349) );
  nand_x1_sg U51146 ( .A(ow_9[14]), .B(n34776), .X(n19350) );
  nand_x1_sg U51147 ( .A(\shifter_0/n9185 ), .B(n31534), .X(n19351) );
  nand_x1_sg U51148 ( .A(ow_9[13]), .B(n30660), .X(n19352) );
  nand_x1_sg U51149 ( .A(\shifter_0/n9184 ), .B(n33195), .X(n19353) );
  nand_x1_sg U51150 ( .A(ow_9[12]), .B(n34783), .X(n19354) );
  nand_x1_sg U51151 ( .A(\shifter_0/n9183 ), .B(n34988), .X(n19355) );
  nand_x1_sg U51152 ( .A(ow_9[11]), .B(n32577), .X(n19356) );
  nand_x1_sg U51153 ( .A(\shifter_0/n9182 ), .B(n33203), .X(n19357) );
  nand_x1_sg U51154 ( .A(ow_9[10]), .B(n34498), .X(n19358) );
  nand_x1_sg U51155 ( .A(\shifter_0/n9181 ), .B(n33209), .X(n19359) );
  nand_x1_sg U51156 ( .A(ow_9[9]), .B(n32629), .X(n19360) );
  nand_x1_sg U51157 ( .A(\shifter_0/n9180 ), .B(n33162), .X(n19361) );
  nand_x1_sg U51158 ( .A(ow_9[8]), .B(n32599), .X(n19362) );
  nand_x1_sg U51159 ( .A(\shifter_0/n9139 ), .B(n34983), .X(n19403) );
  nand_x1_sg U51160 ( .A(ow_10[7]), .B(n30214), .X(n19404) );
  nand_x1_sg U51161 ( .A(\shifter_0/n9138 ), .B(n33160), .X(n19405) );
  nand_x1_sg U51162 ( .A(ow_10[6]), .B(n32579), .X(n19406) );
  nand_x1_sg U51163 ( .A(\shifter_0/n9137 ), .B(n34986), .X(n19407) );
  nand_x1_sg U51164 ( .A(ow_10[5]), .B(n32621), .X(n19408) );
  nand_x1_sg U51165 ( .A(\shifter_0/n9136 ), .B(n34997), .X(n19409) );
  nand_x1_sg U51166 ( .A(ow_10[4]), .B(n32593), .X(n19410) );
  nand_x1_sg U51167 ( .A(\shifter_0/n9135 ), .B(n33160), .X(n19411) );
  nand_x1_sg U51168 ( .A(ow_10[3]), .B(n30608), .X(n19412) );
  nand_x1_sg U51169 ( .A(\shifter_0/n9134 ), .B(n33216), .X(n19413) );
  nand_x1_sg U51170 ( .A(ow_10[2]), .B(n34793), .X(n19414) );
  nand_x1_sg U51171 ( .A(\shifter_0/n9133 ), .B(n33195), .X(n19415) );
  nand_x1_sg U51172 ( .A(ow_10[1]), .B(n30674), .X(n19416) );
  nand_x1_sg U51173 ( .A(\shifter_0/n9132 ), .B(n34977), .X(n19417) );
  nand_x1_sg U51174 ( .A(ow_10[0]), .B(n34784), .X(n19418) );
  nand_x1_sg U51175 ( .A(\shifter_0/n9111 ), .B(n33135), .X(n19419) );
  nand_x1_sg U51176 ( .A(ow_11[19]), .B(n32572), .X(n19420) );
  nand_x1_sg U51177 ( .A(\shifter_0/n9110 ), .B(n29843), .X(n19421) );
  nand_x1_sg U51178 ( .A(ow_11[18]), .B(n34763), .X(n19422) );
  nand_x1_sg U51179 ( .A(\shifter_0/n9109 ), .B(n33142), .X(n19423) );
  nand_x1_sg U51180 ( .A(ow_11[17]), .B(n32095), .X(n19424) );
  nand_x1_sg U51181 ( .A(\shifter_0/n9108 ), .B(n30236), .X(n19425) );
  nand_x1_sg U51182 ( .A(ow_11[16]), .B(n32613), .X(n19426) );
  nand_x1_sg U51183 ( .A(\shifter_0/n9107 ), .B(n33148), .X(n19427) );
  nand_x1_sg U51184 ( .A(ow_11[15]), .B(n30608), .X(n19428) );
  nand_x1_sg U51185 ( .A(\shifter_0/n9106 ), .B(n34996), .X(n19429) );
  nand_x1_sg U51186 ( .A(ow_11[14]), .B(n32592), .X(n19430) );
  nand_x1_sg U51187 ( .A(\shifter_0/n9105 ), .B(n33163), .X(n19431) );
  nand_x1_sg U51188 ( .A(ow_11[13]), .B(n34953), .X(n19432) );
  nand_x1_sg U51189 ( .A(\shifter_0/n9104 ), .B(n33208), .X(n19433) );
  nand_x1_sg U51190 ( .A(ow_11[12]), .B(n32575), .X(n19434) );
  nand_x1_sg U51191 ( .A(\shifter_0/n9103 ), .B(n31554), .X(n19435) );
  nand_x1_sg U51192 ( .A(ow_11[11]), .B(n32615), .X(n19436) );
  nand_x1_sg U51193 ( .A(\shifter_0/n9102 ), .B(n31535), .X(n19437) );
  nand_x1_sg U51194 ( .A(ow_11[10]), .B(n34779), .X(n19438) );
  nand_x1_sg U51195 ( .A(\shifter_0/n9101 ), .B(n29857), .X(n19439) );
  nand_x1_sg U51196 ( .A(ow_11[9]), .B(n32617), .X(n19440) );
  nand_x1_sg U51197 ( .A(\shifter_0/n9100 ), .B(n29850), .X(n19441) );
  nand_x1_sg U51198 ( .A(ow_11[8]), .B(n32581), .X(n19442) );
  nand_x1_sg U51199 ( .A(\shifter_0/n9059 ), .B(n33194), .X(n19483) );
  nand_x1_sg U51200 ( .A(ow_12[7]), .B(n31931), .X(n19484) );
  nand_x1_sg U51201 ( .A(\shifter_0/n9591 ), .B(n30223), .X(n21745) );
  nand_x1_sg U51202 ( .A(ow_15[19]), .B(n32597), .X(n21746) );
  nand_x1_sg U51203 ( .A(\shifter_0/n9590 ), .B(n31543), .X(n21747) );
  nand_x1_sg U51204 ( .A(ow_15[18]), .B(n34792), .X(n21748) );
  nand_x1_sg U51205 ( .A(\shifter_0/n9589 ), .B(n30227), .X(n21749) );
  nand_x1_sg U51206 ( .A(ow_15[17]), .B(n32597), .X(n21750) );
  nand_x1_sg U51207 ( .A(\shifter_0/n9588 ), .B(n33207), .X(n21751) );
  nand_x1_sg U51208 ( .A(ow_15[16]), .B(n34778), .X(n21752) );
  nand_x1_sg U51209 ( .A(\shifter_0/n9587 ), .B(n33213), .X(n21753) );
  nand_x1_sg U51210 ( .A(ow_15[15]), .B(n32545), .X(n21754) );
  nand_x1_sg U51211 ( .A(\shifter_0/n9586 ), .B(n31543), .X(n21755) );
  nand_x1_sg U51212 ( .A(ow_15[14]), .B(n32585), .X(n21756) );
  nand_x1_sg U51213 ( .A(\shifter_0/n9585 ), .B(n33218), .X(n21757) );
  nand_x1_sg U51214 ( .A(ow_15[13]), .B(n34761), .X(n21758) );
  nand_x1_sg U51215 ( .A(\shifter_0/n9584 ), .B(n34985), .X(n21759) );
  nand_x1_sg U51216 ( .A(ow_15[12]), .B(n32620), .X(n21760) );
  nand_x1_sg U51217 ( .A(\shifter_0/n9531 ), .B(n35007), .X(n21825) );
  nand_x1_sg U51218 ( .A(oi_1[19]), .B(n34782), .X(n21826) );
  nand_x1_sg U51219 ( .A(\shifter_0/n9530 ), .B(n29863), .X(n21827) );
  nand_x1_sg U51220 ( .A(oi_1[18]), .B(n32594), .X(n21828) );
  nand_x1_sg U51221 ( .A(\shifter_0/n9529 ), .B(n31560), .X(n21829) );
  nand_x1_sg U51222 ( .A(oi_1[17]), .B(n32600), .X(n21830) );
  nand_x1_sg U51223 ( .A(\shifter_0/n9528 ), .B(n30227), .X(n21831) );
  nand_x1_sg U51224 ( .A(oi_1[16]), .B(n30676), .X(n21832) );
  nand_x1_sg U51225 ( .A(\shifter_0/n9527 ), .B(n31547), .X(n21833) );
  nand_x1_sg U51226 ( .A(oi_1[15]), .B(n32630), .X(n21834) );
  nand_x1_sg U51227 ( .A(\shifter_0/n9526 ), .B(n31549), .X(n21835) );
  nand_x1_sg U51228 ( .A(oi_1[14]), .B(n32570), .X(n21836) );
  nand_x1_sg U51229 ( .A(\shifter_0/n9525 ), .B(n35009), .X(n21837) );
  nand_x1_sg U51230 ( .A(oi_1[13]), .B(n32594), .X(n21838) );
  nand_x1_sg U51231 ( .A(\shifter_0/n9524 ), .B(n29856), .X(n21839) );
  nand_x1_sg U51232 ( .A(oi_1[12]), .B(n30655), .X(n21840) );
  nand_x1_sg U51233 ( .A(\shifter_0/n9523 ), .B(n33195), .X(n21841) );
  nand_x1_sg U51234 ( .A(oi_1[11]), .B(n32099), .X(n21842) );
  nand_x1_sg U51235 ( .A(\shifter_0/n9522 ), .B(n33135), .X(n21843) );
  nand_x1_sg U51236 ( .A(oi_1[10]), .B(n34499), .X(n21844) );
  nand_x1_sg U51237 ( .A(\shifter_0/n9521 ), .B(n33187), .X(n21845) );
  nand_x1_sg U51238 ( .A(oi_1[9]), .B(n32552), .X(n21846) );
  nand_x1_sg U51239 ( .A(\shifter_0/n9520 ), .B(n33216), .X(n21847) );
  nand_x1_sg U51240 ( .A(oi_1[8]), .B(n34776), .X(n21848) );
  nand_x1_sg U51241 ( .A(\shifter_0/n9404 ), .B(n33156), .X(n21959) );
  nand_x1_sg U51242 ( .A(oi_4[12]), .B(n34778), .X(n21960) );
  nand_x1_sg U51243 ( .A(\shifter_0/n9403 ), .B(n30220), .X(n21961) );
  nand_x1_sg U51244 ( .A(oi_4[11]), .B(n34783), .X(n21962) );
  nand_x1_sg U51245 ( .A(\shifter_0/n9402 ), .B(n31560), .X(n21963) );
  nand_x1_sg U51246 ( .A(oi_4[10]), .B(n32575), .X(n21964) );
  nand_x1_sg U51247 ( .A(\shifter_0/n9401 ), .B(n33166), .X(n21965) );
  nand_x1_sg U51248 ( .A(oi_4[9]), .B(n32094), .X(n21966) );
  nand_x1_sg U51249 ( .A(\shifter_0/n9400 ), .B(n31546), .X(n21967) );
  nand_x1_sg U51250 ( .A(oi_4[8]), .B(n32599), .X(n21968) );
  nand_x1_sg U51251 ( .A(\shifter_0/n9359 ), .B(n33144), .X(n22009) );
  nand_x1_sg U51252 ( .A(oi_5[7]), .B(n32600), .X(n22010) );
  nand_x1_sg U51253 ( .A(\shifter_0/n9358 ), .B(n30219), .X(n22011) );
  nand_x1_sg U51254 ( .A(oi_5[6]), .B(n32591), .X(n22012) );
  nand_x1_sg U51255 ( .A(\shifter_0/n9357 ), .B(n33149), .X(n22013) );
  nand_x1_sg U51256 ( .A(oi_5[5]), .B(n32579), .X(n22014) );
  nand_x1_sg U51257 ( .A(\shifter_0/n9356 ), .B(n35002), .X(n22015) );
  nand_x1_sg U51258 ( .A(oi_5[4]), .B(n32576), .X(n22016) );
  nand_x1_sg U51259 ( .A(\shifter_0/n9032 ), .B(n31536), .X(n18897) );
  nand_x1_sg U51260 ( .A(oi_13[0]), .B(n30663), .X(n18898) );
  nand_x1_sg U51261 ( .A(\shifter_0/n9011 ), .B(n33183), .X(n18899) );
  nand_x1_sg U51262 ( .A(oi_14[19]), .B(n32630), .X(n18900) );
  nand_x1_sg U51263 ( .A(\shifter_0/n9010 ), .B(n33215), .X(n18901) );
  nand_x1_sg U51264 ( .A(oi_14[18]), .B(n32584), .X(n18902) );
  nand_x1_sg U51265 ( .A(\shifter_0/n9009 ), .B(n31543), .X(n18903) );
  nand_x1_sg U51266 ( .A(oi_14[17]), .B(n32543), .X(n18904) );
  nand_x1_sg U51267 ( .A(\shifter_0/n9008 ), .B(n31224), .X(n18905) );
  nand_x1_sg U51268 ( .A(oi_14[16]), .B(n30651), .X(n18906) );
  nand_x1_sg U51269 ( .A(\shifter_0/n9007 ), .B(n33152), .X(n18907) );
  nand_x1_sg U51270 ( .A(oi_14[15]), .B(n32620), .X(n18908) );
  nand_x1_sg U51271 ( .A(\shifter_0/n9006 ), .B(n29839), .X(n18909) );
  nand_x1_sg U51272 ( .A(oi_14[14]), .B(n32611), .X(n18910) );
  nand_x1_sg U51273 ( .A(\shifter_0/n9005 ), .B(n31554), .X(n18911) );
  nand_x1_sg U51274 ( .A(oi_14[13]), .B(n34495), .X(n18912) );
  nand_x1_sg U51275 ( .A(\shifter_0/n9004 ), .B(n33132), .X(n18913) );
  nand_x1_sg U51276 ( .A(oi_14[12]), .B(n32597), .X(n18914) );
  nand_x1_sg U51277 ( .A(\shifter_0/n9003 ), .B(n30230), .X(n18915) );
  nand_x1_sg U51278 ( .A(oi_14[11]), .B(n34768), .X(n18916) );
  nand_x1_sg U51279 ( .A(\shifter_0/n9002 ), .B(n30234), .X(n18917) );
  nand_x1_sg U51280 ( .A(oi_14[10]), .B(n32608), .X(n18918) );
  nand_x1_sg U51281 ( .A(\shifter_0/n9001 ), .B(n31550), .X(n18919) );
  nand_x1_sg U51282 ( .A(oi_14[9]), .B(n32572), .X(n18920) );
  nand_x1_sg U51283 ( .A(\shifter_0/n9000 ), .B(n33161), .X(n18921) );
  nand_x1_sg U51284 ( .A(oi_14[8]), .B(n34948), .X(n18922) );
  nand_x1_sg U51285 ( .A(\shifter_0/n8999 ), .B(n33216), .X(n18923) );
  nand_x1_sg U51286 ( .A(oi_14[7]), .B(n32546), .X(n18924) );
  nand_x1_sg U51287 ( .A(\shifter_0/n8998 ), .B(n33165), .X(n18925) );
  nand_x1_sg U51288 ( .A(oi_14[6]), .B(n32617), .X(n18926) );
  nand_x1_sg U51289 ( .A(\shifter_0/n8997 ), .B(n31550), .X(n18927) );
  nand_x1_sg U51290 ( .A(oi_14[5]), .B(n32564), .X(n18928) );
  nand_x1_sg U51291 ( .A(\shifter_0/n8996 ), .B(n33221), .X(n18929) );
  nand_x1_sg U51292 ( .A(oi_14[4]), .B(n32096), .X(n18930) );
  nand_x1_sg U51293 ( .A(\shifter_0/n8995 ), .B(n34981), .X(n18931) );
  nand_x1_sg U51294 ( .A(oi_14[3]), .B(n32546), .X(n18932) );
  nand_x1_sg U51295 ( .A(\shifter_0/n8994 ), .B(n33177), .X(n18933) );
  nand_x1_sg U51296 ( .A(oi_14[2]), .B(n32555), .X(n18934) );
  nand_x1_sg U51297 ( .A(\shifter_0/n8993 ), .B(n29845), .X(n18935) );
  nand_x1_sg U51298 ( .A(oi_14[1]), .B(n34764), .X(n18936) );
  nand_x1_sg U51299 ( .A(\shifter_0/n8992 ), .B(n33187), .X(n18937) );
  nand_x1_sg U51300 ( .A(oi_14[0]), .B(n32545), .X(n18938) );
  nand_x1_sg U51301 ( .A(\shifter_0/n8971 ), .B(n33175), .X(n18939) );
  nand_x1_sg U51302 ( .A(oi_15[19]), .B(n30647), .X(n18940) );
  nand_x1_sg U51303 ( .A(\shifter_0/n8970 ), .B(n33133), .X(n18941) );
  nand_x1_sg U51304 ( .A(oi_15[18]), .B(n34954), .X(n18942) );
  nand_x1_sg U51305 ( .A(\shifter_0/n8969 ), .B(n33136), .X(n18943) );
  nand_x1_sg U51306 ( .A(oi_15[17]), .B(n32634), .X(n18944) );
  nand_x1_sg U51307 ( .A(\shifter_0/n8968 ), .B(n33215), .X(n18945) );
  nand_x1_sg U51308 ( .A(oi_15[16]), .B(n32617), .X(n18946) );
  nand_x1_sg U51309 ( .A(\shifter_0/n8967 ), .B(n34978), .X(n18947) );
  nand_x1_sg U51310 ( .A(oi_15[15]), .B(n34786), .X(n18948) );
  nand_x1_sg U51311 ( .A(\shifter_0/n8960 ), .B(n33183), .X(n18961) );
  nand_x1_sg U51312 ( .A(oi_15[8]), .B(n32624), .X(n18962) );
  nand_x1_sg U51313 ( .A(\shifter_0/n8959 ), .B(n31539), .X(n18963) );
  nand_x1_sg U51314 ( .A(oi_15[7]), .B(n30668), .X(n18964) );
  nand_x1_sg U51315 ( .A(\shifter_0/n8958 ), .B(n33199), .X(n18965) );
  nand_x1_sg U51316 ( .A(oi_15[6]), .B(n30656), .X(n18966) );
  nand_x1_sg U51317 ( .A(\shifter_0/n8957 ), .B(n31555), .X(n18967) );
  nand_x1_sg U51318 ( .A(oi_15[5]), .B(n34756), .X(n18968) );
  nand_x1_sg U51319 ( .A(\shifter_0/n8956 ), .B(n29863), .X(n18969) );
  nand_x1_sg U51320 ( .A(oi_15[4]), .B(n30652), .X(n18970) );
  nand_x1_sg U51321 ( .A(\shifter_0/n8955 ), .B(n33170), .X(n18971) );
  nand_x1_sg U51322 ( .A(oi_15[3]), .B(n32625), .X(n18972) );
  nand_x1_sg U51323 ( .A(\shifter_0/n8954 ), .B(n34983), .X(n18973) );
  nand_x1_sg U51324 ( .A(oi_15[2]), .B(n32603), .X(n18974) );
  nand_x1_sg U51325 ( .A(\shifter_0/n8953 ), .B(n33149), .X(n18975) );
  nand_x1_sg U51326 ( .A(oi_15[1]), .B(n34769), .X(n18976) );
  nand_x1_sg U51327 ( .A(\shifter_0/n8952 ), .B(n33827), .X(n18977) );
  nand_x1_sg U51328 ( .A(oi_15[0]), .B(n32541), .X(n18978) );
  nand_x1_sg U51329 ( .A(\shifter_0/n9551 ), .B(n33201), .X(n18979) );
  nand_x1_sg U51330 ( .A(ow_0[19]), .B(n34789), .X(n18980) );
  nand_x1_sg U51331 ( .A(\shifter_0/n9550 ), .B(n33826), .X(n18981) );
  nand_x1_sg U51332 ( .A(ow_0[18]), .B(n32594), .X(n18982) );
  nand_x1_sg U51333 ( .A(\shifter_0/n9549 ), .B(n30224), .X(n18983) );
  nand_x1_sg U51334 ( .A(ow_0[17]), .B(n32615), .X(n18984) );
  nand_x1_sg U51335 ( .A(\shifter_0/n9548 ), .B(n31539), .X(n18985) );
  nand_x1_sg U51336 ( .A(ow_0[16]), .B(n30667), .X(n18986) );
  nand_x1_sg U51337 ( .A(\shifter_0/n9547 ), .B(n33211), .X(n18987) );
  nand_x1_sg U51338 ( .A(ow_0[15]), .B(n32635), .X(n18988) );
  nand_x1_sg U51339 ( .A(\shifter_0/n9546 ), .B(n33211), .X(n18989) );
  nand_x1_sg U51340 ( .A(ow_0[14]), .B(n32585), .X(n18990) );
  nand_x1_sg U51341 ( .A(\shifter_0/n9545 ), .B(n31539), .X(n18991) );
  nand_x1_sg U51342 ( .A(ow_0[13]), .B(n32560), .X(n18992) );
  nand_x1_sg U51343 ( .A(\shifter_0/n9544 ), .B(n35002), .X(n18993) );
  nand_x1_sg U51344 ( .A(ow_0[12]), .B(n32612), .X(n18994) );
  nand_x1_sg U51345 ( .A(\shifter_0/n9543 ), .B(n34995), .X(n18995) );
  nand_x1_sg U51346 ( .A(ow_0[11]), .B(n34779), .X(n18996) );
  nand_x1_sg U51347 ( .A(\shifter_0/n9542 ), .B(n33140), .X(n18997) );
  nand_x1_sg U51348 ( .A(ow_0[10]), .B(n32593), .X(n18998) );
  nand_x1_sg U51349 ( .A(\shifter_0/n9541 ), .B(n33166), .X(n18999) );
  nand_x1_sg U51350 ( .A(ow_0[9]), .B(n34757), .X(n19000) );
  nand_x1_sg U51351 ( .A(\shifter_0/n9540 ), .B(n33167), .X(n19001) );
  nand_x1_sg U51352 ( .A(ow_0[8]), .B(n32540), .X(n19002) );
  nand_x1_sg U51353 ( .A(\shifter_0/n9332 ), .B(n33208), .X(n19217) );
  nand_x1_sg U51354 ( .A(ow_5[0]), .B(n34951), .X(n19218) );
  nand_x1_sg U51355 ( .A(\shifter_0/n9311 ), .B(n31221), .X(n19219) );
  nand_x1_sg U51356 ( .A(ow_6[19]), .B(n30649), .X(n19220) );
  nand_x1_sg U51357 ( .A(\shifter_0/n9310 ), .B(n33141), .X(n19221) );
  nand_x1_sg U51358 ( .A(ow_6[18]), .B(n31929), .X(n19222) );
  nand_x1_sg U51359 ( .A(\shifter_0/n9309 ), .B(n34988), .X(n19223) );
  nand_x1_sg U51360 ( .A(ow_6[17]), .B(n34789), .X(n19224) );
  nand_x1_sg U51361 ( .A(\shifter_0/n9308 ), .B(n34984), .X(n19225) );
  nand_x1_sg U51362 ( .A(ow_6[16]), .B(n32623), .X(n19226) );
  nand_x1_sg U51363 ( .A(\shifter_0/n9307 ), .B(n33141), .X(n19227) );
  nand_x1_sg U51364 ( .A(ow_6[15]), .B(n32540), .X(n19228) );
  nand_x1_sg U51365 ( .A(\shifter_0/n9306 ), .B(n31547), .X(n19229) );
  nand_x1_sg U51366 ( .A(ow_6[14]), .B(n30798), .X(n19230) );
  nand_x1_sg U51367 ( .A(\shifter_0/n9305 ), .B(n31535), .X(n19231) );
  nand_x1_sg U51368 ( .A(ow_6[13]), .B(n32623), .X(n19232) );
  nand_x1_sg U51369 ( .A(\shifter_0/n9304 ), .B(n33214), .X(n19233) );
  nand_x1_sg U51370 ( .A(ow_6[12]), .B(n32570), .X(n19234) );
  nand_x1_sg U51371 ( .A(\shifter_0/n9303 ), .B(n33148), .X(n19235) );
  nand_x1_sg U51372 ( .A(ow_6[11]), .B(n30677), .X(n19236) );
  nand_x1_sg U51373 ( .A(\shifter_0/n9302 ), .B(n34975), .X(n19237) );
  nand_x1_sg U51374 ( .A(ow_6[10]), .B(n34777), .X(n19238) );
  nand_x1_sg U51375 ( .A(\shifter_0/n9301 ), .B(n33826), .X(n19239) );
  nand_x1_sg U51376 ( .A(ow_6[9]), .B(n32630), .X(n19240) );
  nand_x1_sg U51377 ( .A(\shifter_0/n9300 ), .B(n33199), .X(n19241) );
  nand_x1_sg U51378 ( .A(ow_6[8]), .B(n32606), .X(n19242) );
  nand_x1_sg U51379 ( .A(\shifter_0/n9299 ), .B(n30219), .X(n19243) );
  nand_x1_sg U51380 ( .A(ow_6[7]), .B(n32606), .X(n19244) );
  nand_x1_sg U51381 ( .A(\shifter_0/n9298 ), .B(n33147), .X(n19245) );
  nand_x1_sg U51382 ( .A(ow_6[6]), .B(n34498), .X(n19246) );
  nand_x1_sg U51383 ( .A(\shifter_0/n9297 ), .B(n33137), .X(n19247) );
  nand_x1_sg U51384 ( .A(ow_6[5]), .B(n32568), .X(n19248) );
  nand_x1_sg U51385 ( .A(\shifter_0/n9296 ), .B(n31220), .X(n19249) );
  nand_x1_sg U51386 ( .A(ow_6[4]), .B(n34758), .X(n19250) );
  nand_x1_sg U51387 ( .A(\shifter_0/n9295 ), .B(n33200), .X(n19251) );
  nand_x1_sg U51388 ( .A(ow_6[3]), .B(n34768), .X(n19252) );
  nand_x1_sg U51389 ( .A(\shifter_0/n9294 ), .B(n33220), .X(n19253) );
  nand_x1_sg U51390 ( .A(ow_6[2]), .B(n32579), .X(n19254) );
  nand_x1_sg U51391 ( .A(\shifter_0/n9293 ), .B(n31546), .X(n19255) );
  nand_x1_sg U51392 ( .A(ow_6[1]), .B(n34949), .X(n19256) );
  nand_x1_sg U51393 ( .A(\shifter_0/n9292 ), .B(n34996), .X(n19257) );
  nand_x1_sg U51394 ( .A(ow_6[0]), .B(n34499), .X(n19258) );
  nand_x1_sg U51395 ( .A(\shifter_0/n9271 ), .B(n33173), .X(n19259) );
  nand_x1_sg U51396 ( .A(ow_7[19]), .B(n34952), .X(n19260) );
  nand_x1_sg U51397 ( .A(\shifter_0/n9270 ), .B(n33221), .X(n19261) );
  nand_x1_sg U51398 ( .A(ow_7[18]), .B(n32632), .X(n19262) );
  nand_x1_sg U51399 ( .A(\shifter_0/n9269 ), .B(n29842), .X(n19263) );
  nand_x1_sg U51400 ( .A(ow_7[17]), .B(n30664), .X(n19264) );
  nand_x1_sg U51401 ( .A(\shifter_0/n9268 ), .B(n33197), .X(n19265) );
  nand_x1_sg U51402 ( .A(ow_7[16]), .B(n32100), .X(n19266) );
  nand_x1_sg U51403 ( .A(\shifter_0/n9267 ), .B(n35005), .X(n19267) );
  nand_x1_sg U51404 ( .A(ow_7[15]), .B(n34500), .X(n19268) );
  nand_x1_sg U51405 ( .A(\shifter_0/n9266 ), .B(n31561), .X(n19269) );
  nand_x1_sg U51406 ( .A(ow_7[14]), .B(n34954), .X(n19270) );
  nand_x1_sg U51407 ( .A(\shifter_0/n9265 ), .B(n29846), .X(n19271) );
  nand_x1_sg U51408 ( .A(ow_7[13]), .B(n34952), .X(n19272) );
  nand_x1_sg U51409 ( .A(\shifter_0/n9264 ), .B(n33194), .X(n19273) );
  nand_x1_sg U51410 ( .A(ow_7[12]), .B(n32550), .X(n19274) );
  nand_x1_sg U51411 ( .A(\shifter_0/n9055 ), .B(n31225), .X(n19491) );
  nand_x1_sg U51412 ( .A(ow_12[3]), .B(n30610), .X(n19492) );
  nand_x1_sg U51413 ( .A(\shifter_0/n9054 ), .B(n34997), .X(n19493) );
  nand_x1_sg U51414 ( .A(ow_12[2]), .B(n31931), .X(n19494) );
  nand_x1_sg U51415 ( .A(\shifter_0/n9053 ), .B(n31560), .X(n19495) );
  nand_x1_sg U51416 ( .A(ow_12[1]), .B(n30647), .X(n19496) );
  nand_x1_sg U51417 ( .A(\shifter_0/n9052 ), .B(n33211), .X(n19497) );
  nand_x1_sg U51418 ( .A(ow_12[0]), .B(n32591), .X(n19498) );
  nand_x1_sg U51419 ( .A(\shifter_0/n9031 ), .B(n34986), .X(n19499) );
  nand_x1_sg U51420 ( .A(ow_13[19]), .B(n34501), .X(n19500) );
  nand_x1_sg U51421 ( .A(\shifter_0/n9030 ), .B(n33204), .X(n19501) );
  nand_x1_sg U51422 ( .A(ow_13[18]), .B(n30659), .X(n19502) );
  nand_x1_sg U51423 ( .A(\shifter_0/n9029 ), .B(n29867), .X(n19503) );
  nand_x1_sg U51424 ( .A(ow_13[17]), .B(n32596), .X(n19504) );
  nand_x1_sg U51425 ( .A(\shifter_0/n9028 ), .B(n35008), .X(n19505) );
  nand_x1_sg U51426 ( .A(ow_13[16]), .B(n34777), .X(n19506) );
  nand_x1_sg U51427 ( .A(\shifter_0/n9027 ), .B(n35001), .X(n19507) );
  nand_x1_sg U51428 ( .A(ow_13[15]), .B(n34791), .X(n19508) );
  nand_x1_sg U51429 ( .A(\shifter_0/n9026 ), .B(n33138), .X(n19509) );
  nand_x1_sg U51430 ( .A(ow_13[14]), .B(n34500), .X(n19510) );
  nand_x1_sg U51431 ( .A(\shifter_0/n9025 ), .B(n31551), .X(n19511) );
  nand_x1_sg U51432 ( .A(ow_13[13]), .B(n32550), .X(n19512) );
  nand_x1_sg U51433 ( .A(\shifter_0/n9024 ), .B(n34987), .X(n19513) );
  nand_x1_sg U51434 ( .A(ow_13[12]), .B(n34793), .X(n19514) );
  nand_x1_sg U51435 ( .A(\shifter_0/n9023 ), .B(n33827), .X(n19515) );
  nand_x1_sg U51436 ( .A(ow_13[11]), .B(n32613), .X(n19516) );
  nand_x1_sg U51437 ( .A(\shifter_0/n9022 ), .B(n31543), .X(n19517) );
  nand_x1_sg U51438 ( .A(ow_13[10]), .B(n30667), .X(n19518) );
  nand_x1_sg U51439 ( .A(\shifter_0/n9021 ), .B(n33164), .X(n19519) );
  nand_x1_sg U51440 ( .A(ow_13[9]), .B(n34759), .X(n19520) );
  nand_x1_sg U51441 ( .A(\shifter_0/n9020 ), .B(n34978), .X(n19521) );
  nand_x1_sg U51442 ( .A(ow_13[8]), .B(n32596), .X(n19522) );
  nand_x1_sg U51443 ( .A(\shifter_0/n8979 ), .B(n31224), .X(n19563) );
  nand_x1_sg U51444 ( .A(ow_14[7]), .B(n34762), .X(n19564) );
  nand_x1_sg U51445 ( .A(\shifter_0/n8978 ), .B(n33221), .X(n19565) );
  nand_x1_sg U51446 ( .A(ow_14[6]), .B(n34955), .X(n19566) );
  nand_x1_sg U51447 ( .A(\shifter_0/n8977 ), .B(n31547), .X(n19567) );
  nand_x1_sg U51448 ( .A(ow_14[5]), .B(n34787), .X(n19568) );
  nand_x1_sg U51449 ( .A(\shifter_0/n8976 ), .B(n34977), .X(n19569) );
  nand_x1_sg U51450 ( .A(ow_14[4]), .B(n32095), .X(n19570) );
  nand_x1_sg U51451 ( .A(\shifter_0/n8975 ), .B(n33219), .X(n19571) );
  nand_x1_sg U51452 ( .A(ow_14[3]), .B(n34779), .X(n19572) );
  nand_x1_sg U51453 ( .A(\shifter_0/n8974 ), .B(n33185), .X(n19573) );
  nand_x1_sg U51454 ( .A(ow_14[2]), .B(n32100), .X(n19574) );
  nand_x1_sg U51455 ( .A(\shifter_0/n8973 ), .B(n33202), .X(n19575) );
  nand_x1_sg U51456 ( .A(ow_14[1]), .B(n30673), .X(n19576) );
  nand_x1_sg U51457 ( .A(\shifter_0/n8972 ), .B(n33179), .X(n19577) );
  nand_x1_sg U51458 ( .A(ow_14[0]), .B(n32587), .X(n19578) );
  nand_x1_sg U51459 ( .A(\shifter_0/n9015 ), .B(n34980), .X(n19531) );
  nand_x1_sg U51460 ( .A(ow_13[3]), .B(n34501), .X(n19532) );
  nand_x1_sg U51461 ( .A(\shifter_0/n9014 ), .B(n33200), .X(n19533) );
  nand_x1_sg U51462 ( .A(ow_13[2]), .B(n32570), .X(n19534) );
  nand_x1_sg U51463 ( .A(\shifter_0/n9013 ), .B(n33142), .X(n19535) );
  nand_x1_sg U51464 ( .A(ow_13[1]), .B(n32562), .X(n19536) );
  nand_x1_sg U51465 ( .A(\shifter_0/n9283 ), .B(n33209), .X(n22081) );
  nand_x1_sg U51466 ( .A(oi_7[11]), .B(n34493), .X(n22082) );
  nand_x1_sg U51467 ( .A(\shifter_0/n9282 ), .B(n33824), .X(n22083) );
  nand_x1_sg U51468 ( .A(oi_7[10]), .B(n32563), .X(n22084) );
  nand_x1_sg U51469 ( .A(\shifter_0/n9281 ), .B(n29851), .X(n22085) );
  nand_x1_sg U51470 ( .A(oi_7[9]), .B(n32612), .X(n22086) );
  nand_x1_sg U51471 ( .A(\shifter_0/n9511 ), .B(n34989), .X(n19019) );
  nand_x1_sg U51472 ( .A(ow_1[19]), .B(n34946), .X(n19020) );
  nand_x1_sg U51473 ( .A(\shifter_0/n9510 ), .B(n33191), .X(n19021) );
  nand_x1_sg U51474 ( .A(ow_1[18]), .B(n32543), .X(n19022) );
  nand_x1_sg U51475 ( .A(\shifter_0/n9509 ), .B(n33200), .X(n19023) );
  nand_x1_sg U51476 ( .A(ow_1[17]), .B(n30653), .X(n19024) );
  nand_x1_sg U51477 ( .A(\shifter_0/n9456 ), .B(n31541), .X(n19089) );
  nand_x1_sg U51478 ( .A(ow_2[4]), .B(n32599), .X(n19090) );
  nand_x1_sg U51479 ( .A(\shifter_0/n9455 ), .B(n33189), .X(n19091) );
  nand_x1_sg U51480 ( .A(ow_2[3]), .B(n32594), .X(n19092) );
  nand_x1_sg U51481 ( .A(\shifter_0/n9454 ), .B(n31552), .X(n19093) );
  nand_x1_sg U51482 ( .A(ow_2[2]), .B(n32564), .X(n19094) );
  nand_x1_sg U51483 ( .A(\shifter_0/n9479 ), .B(n31219), .X(n21889) );
  nand_x1_sg U51484 ( .A(oi_2[7]), .B(n32541), .X(n21890) );
  nand_x1_sg U51485 ( .A(\shifter_0/n9478 ), .B(n33143), .X(n21891) );
  nand_x1_sg U51486 ( .A(oi_2[6]), .B(n34783), .X(n21892) );
  nand_x1_sg U51487 ( .A(\shifter_0/n9477 ), .B(n33150), .X(n21893) );
  nand_x1_sg U51488 ( .A(oi_2[5]), .B(n32634), .X(n21894) );
  nand_x1_sg U51489 ( .A(\shifter_0/n9476 ), .B(n31540), .X(n21895) );
  nand_x1_sg U51490 ( .A(oi_2[4]), .B(n32541), .X(n21896) );
  nand_x1_sg U51491 ( .A(\shifter_0/n9475 ), .B(n33156), .X(n21897) );
  nand_x1_sg U51492 ( .A(oi_2[3]), .B(n34496), .X(n21898) );
  nand_x1_sg U51493 ( .A(\shifter_0/n9474 ), .B(n33184), .X(n21899) );
  nand_x1_sg U51494 ( .A(oi_2[2]), .B(n34784), .X(n21900) );
  nand_x1_sg U51495 ( .A(\shifter_0/n9473 ), .B(n31221), .X(n21901) );
  nand_x1_sg U51496 ( .A(oi_2[1]), .B(n32586), .X(n21902) );
  nand_x1_sg U51497 ( .A(\shifter_0/n9472 ), .B(n33154), .X(n21903) );
  nand_x1_sg U51498 ( .A(oi_2[0]), .B(n31932), .X(n21904) );
  nand_x1_sg U51499 ( .A(\shifter_0/n9451 ), .B(n33825), .X(n21905) );
  nand_x1_sg U51500 ( .A(oi_3[19]), .B(n34773), .X(n21906) );
  nand_x1_sg U51501 ( .A(\shifter_0/n9450 ), .B(n31226), .X(n21907) );
  nand_x1_sg U51502 ( .A(oi_3[18]), .B(n31929), .X(n21908) );
  nand_x1_sg U51503 ( .A(\shifter_0/n9449 ), .B(n33183), .X(n21909) );
  nand_x1_sg U51504 ( .A(oi_3[17]), .B(n34791), .X(n21910) );
  nand_x1_sg U51505 ( .A(\shifter_0/n9448 ), .B(n33152), .X(n21911) );
  nand_x1_sg U51506 ( .A(oi_3[16]), .B(n30668), .X(n21912) );
  nand_x1_sg U51507 ( .A(\shifter_0/n9447 ), .B(n31538), .X(n21913) );
  nand_x1_sg U51508 ( .A(oi_3[15]), .B(n34786), .X(n21914) );
  nand_x1_sg U51509 ( .A(\shifter_0/n9446 ), .B(n31534), .X(n21915) );
  nand_x1_sg U51510 ( .A(oi_3[14]), .B(n32556), .X(n21916) );
  nand_x1_sg U51511 ( .A(\shifter_0/n9445 ), .B(n35006), .X(n21917) );
  nand_x1_sg U51512 ( .A(oi_3[13]), .B(n32574), .X(n21918) );
  nand_x1_sg U51513 ( .A(\shifter_0/n9444 ), .B(n29857), .X(n21919) );
  nand_x1_sg U51514 ( .A(oi_3[12]), .B(n30669), .X(n21920) );
  nand_x1_sg U51515 ( .A(\shifter_0/n9443 ), .B(n33177), .X(n21921) );
  nand_x1_sg U51516 ( .A(oi_3[11]), .B(n32635), .X(n21922) );
  nand_x1_sg U51517 ( .A(\shifter_0/n9442 ), .B(n35001), .X(n21923) );
  nand_x1_sg U51518 ( .A(oi_3[10]), .B(n30673), .X(n21924) );
  nand_x1_sg U51519 ( .A(\shifter_0/n9441 ), .B(n31541), .X(n21925) );
  nand_x1_sg U51520 ( .A(oi_3[9]), .B(n32556), .X(n21926) );
  nand_x1_sg U51521 ( .A(\shifter_0/n9440 ), .B(n33188), .X(n21927) );
  nand_x1_sg U51522 ( .A(oi_3[8]), .B(n30655), .X(n21928) );
  nand_x1_sg U51523 ( .A(\shifter_0/n9319 ), .B(n33157), .X(n22049) );
  nand_x1_sg U51524 ( .A(oi_6[7]), .B(n30665), .X(n22050) );
  nand_x1_sg U51525 ( .A(\shifter_0/n9318 ), .B(n31224), .X(n22051) );
  nand_x1_sg U51526 ( .A(oi_6[6]), .B(n34791), .X(n22052) );
  nand_x1_sg U51527 ( .A(\shifter_0/n9317 ), .B(n30970), .X(n22053) );
  nand_x1_sg U51528 ( .A(oi_6[5]), .B(n30673), .X(n22054) );
  nand_x1_sg U51529 ( .A(\shifter_0/n9316 ), .B(n33168), .X(n22055) );
  nand_x1_sg U51530 ( .A(oi_6[4]), .B(n34769), .X(n22056) );
  nand_x1_sg U51531 ( .A(\shifter_0/n9315 ), .B(n33163), .X(n22057) );
  nand_x1_sg U51532 ( .A(oi_6[3]), .B(n30608), .X(n22058) );
  nand_x1_sg U51533 ( .A(\shifter_0/n9314 ), .B(n33185), .X(n22059) );
  nand_x1_sg U51534 ( .A(oi_6[2]), .B(n32551), .X(n22060) );
  nand_x1_sg U51535 ( .A(\shifter_0/n9313 ), .B(n33214), .X(n22061) );
  nand_x1_sg U51536 ( .A(oi_6[1]), .B(n32601), .X(n22062) );
  nand_x1_sg U51537 ( .A(\shifter_0/n9312 ), .B(n33197), .X(n22063) );
  nand_x1_sg U51538 ( .A(oi_6[0]), .B(n32584), .X(n22064) );
  nand_x1_sg U51539 ( .A(\shifter_0/n9291 ), .B(n30222), .X(n22065) );
  nand_x1_sg U51540 ( .A(oi_7[19]), .B(n32565), .X(n22066) );
  nand_x1_sg U51541 ( .A(\shifter_0/n9290 ), .B(n33190), .X(n22067) );
  nand_x1_sg U51542 ( .A(oi_7[18]), .B(n34493), .X(n22068) );
  nand_x1_sg U51543 ( .A(\shifter_0/n9289 ), .B(n33182), .X(n22069) );
  nand_x1_sg U51544 ( .A(oi_7[17]), .B(n32548), .X(n22070) );
  nand_x1_sg U51545 ( .A(\shifter_0/n9288 ), .B(n33212), .X(n22071) );
  nand_x1_sg U51546 ( .A(oi_7[16]), .B(n30667), .X(n22072) );
  nand_x1_sg U51547 ( .A(\shifter_0/n9287 ), .B(n29846), .X(n22073) );
  nand_x1_sg U51548 ( .A(oi_7[15]), .B(n32553), .X(n22074) );
  nand_x1_sg U51549 ( .A(\shifter_0/n9286 ), .B(n33219), .X(n22075) );
  nand_x1_sg U51550 ( .A(oi_7[14]), .B(n32588), .X(n22076) );
  nand_x1_sg U51551 ( .A(\shifter_0/n9285 ), .B(n34985), .X(n22077) );
  nand_x1_sg U51552 ( .A(oi_7[13]), .B(n32562), .X(n22078) );
  nand_x1_sg U51553 ( .A(\shifter_0/n9284 ), .B(n31225), .X(n22079) );
  nand_x1_sg U51554 ( .A(oi_7[12]), .B(n30664), .X(n22080) );
  nand_x1_sg U51555 ( .A(\shifter_0/n9280 ), .B(n31227), .X(n22087) );
  nand_x1_sg U51556 ( .A(oi_7[8]), .B(n32562), .X(n22088) );
  nand_x1_sg U51557 ( .A(\shifter_0/n9119 ), .B(n33182), .X(n18803) );
  nand_x1_sg U51558 ( .A(oi_11[7]), .B(n32629), .X(n18804) );
  nand_x1_sg U51559 ( .A(\shifter_0/n9118 ), .B(n31560), .X(n18805) );
  nand_x1_sg U51560 ( .A(oi_11[6]), .B(n30653), .X(n18806) );
  nand_x1_sg U51561 ( .A(\shifter_0/n9117 ), .B(n30971), .X(n18807) );
  nand_x1_sg U51562 ( .A(oi_11[5]), .B(n32558), .X(n18808) );
  nand_x1_sg U51563 ( .A(\shifter_0/n9116 ), .B(n34996), .X(n18809) );
  nand_x1_sg U51564 ( .A(oi_11[4]), .B(n34948), .X(n18810) );
  nand_x1_sg U51565 ( .A(\shifter_0/n9115 ), .B(n29845), .X(n18811) );
  nand_x1_sg U51566 ( .A(oi_11[3]), .B(n32581), .X(n18812) );
  nand_x1_sg U51567 ( .A(\shifter_0/n9114 ), .B(n31553), .X(n18813) );
  nand_x1_sg U51568 ( .A(oi_11[2]), .B(n32591), .X(n18814) );
  nand_x1_sg U51569 ( .A(\shifter_0/n9113 ), .B(n33162), .X(n18815) );
  nand_x1_sg U51570 ( .A(oi_11[1]), .B(n34945), .X(n18816) );
  nand_x1_sg U51571 ( .A(\shifter_0/n9112 ), .B(n34981), .X(n18817) );
  nand_x1_sg U51572 ( .A(oi_11[0]), .B(n32564), .X(n18818) );
  nand_x1_sg U51573 ( .A(\shifter_0/n9091 ), .B(n33172), .X(n18819) );
  nand_x1_sg U51574 ( .A(oi_12[19]), .B(n31930), .X(n18820) );
  nand_x1_sg U51575 ( .A(\shifter_0/n9090 ), .B(n33182), .X(n18821) );
  nand_x1_sg U51576 ( .A(oi_12[18]), .B(n30656), .X(n18822) );
  nand_x1_sg U51577 ( .A(\shifter_0/n9089 ), .B(n33145), .X(n18823) );
  nand_x1_sg U51578 ( .A(oi_12[17]), .B(n30674), .X(n18824) );
  nand_x1_sg U51579 ( .A(\shifter_0/n9088 ), .B(n33179), .X(n18825) );
  nand_x1_sg U51580 ( .A(oi_12[16]), .B(n32584), .X(n18826) );
  nand_x1_sg U51581 ( .A(\shifter_0/n9087 ), .B(n31539), .X(n18827) );
  nand_x1_sg U51582 ( .A(oi_12[15]), .B(n34952), .X(n18828) );
  nand_x1_sg U51583 ( .A(\shifter_0/n9086 ), .B(n29842), .X(n18829) );
  nand_x1_sg U51584 ( .A(oi_12[14]), .B(n30648), .X(n18830) );
  nand_x1_sg U51585 ( .A(\shifter_0/n9085 ), .B(n33195), .X(n18831) );
  nand_x1_sg U51586 ( .A(oi_12[13]), .B(n30655), .X(n18832) );
  nand_x1_sg U51587 ( .A(\shifter_0/n9084 ), .B(n31552), .X(n18833) );
  nand_x1_sg U51588 ( .A(oi_12[12]), .B(n30610), .X(n18834) );
  nand_x1_sg U51589 ( .A(\shifter_0/n9083 ), .B(n34989), .X(n18835) );
  nand_x1_sg U51590 ( .A(oi_12[11]), .B(n32628), .X(n18836) );
  nand_x1_sg U51591 ( .A(\shifter_0/n9082 ), .B(n33163), .X(n18837) );
  nand_x1_sg U51592 ( .A(oi_12[10]), .B(n32543), .X(n18838) );
  nand_x1_sg U51593 ( .A(\shifter_0/n9081 ), .B(n33182), .X(n18839) );
  nand_x1_sg U51594 ( .A(oi_12[9]), .B(n32576), .X(n18840) );
  nand_x1_sg U51595 ( .A(\shifter_0/n9080 ), .B(n31220), .X(n18841) );
  nand_x1_sg U51596 ( .A(oi_12[8]), .B(n32544), .X(n18842) );
  nand_x1_sg U51597 ( .A(\shifter_0/n9508 ), .B(n33142), .X(n19025) );
  nand_x1_sg U51598 ( .A(ow_1[16]), .B(n32565), .X(n19026) );
  nand_x1_sg U51599 ( .A(\shifter_0/n9507 ), .B(n33164), .X(n19027) );
  nand_x1_sg U51600 ( .A(ow_1[15]), .B(n34792), .X(n19028) );
  nand_x1_sg U51601 ( .A(\shifter_0/n9506 ), .B(n33184), .X(n19029) );
  nand_x1_sg U51602 ( .A(ow_1[14]), .B(n30664), .X(n19030) );
  nand_x1_sg U51603 ( .A(\shifter_0/n9505 ), .B(n35009), .X(n19031) );
  nand_x1_sg U51604 ( .A(ow_1[13]), .B(n30125), .X(n19032) );
  nand_x1_sg U51605 ( .A(\shifter_0/n9504 ), .B(n30231), .X(n19033) );
  nand_x1_sg U51606 ( .A(ow_1[12]), .B(n34955), .X(n19034) );
  nand_x1_sg U51607 ( .A(\shifter_0/n9503 ), .B(n35001), .X(n19035) );
  nand_x1_sg U51608 ( .A(ow_1[11]), .B(n32545), .X(n19036) );
  nand_x1_sg U51609 ( .A(\shifter_0/n9502 ), .B(n33176), .X(n19037) );
  nand_x1_sg U51610 ( .A(ow_1[10]), .B(n34788), .X(n19038) );
  nand_x1_sg U51611 ( .A(\shifter_0/n9501 ), .B(n33154), .X(n19039) );
  nand_x1_sg U51612 ( .A(ow_1[9]), .B(n34949), .X(n19040) );
  nand_x1_sg U51613 ( .A(\shifter_0/n9500 ), .B(n33173), .X(n19041) );
  nand_x1_sg U51614 ( .A(ow_1[8]), .B(n32592), .X(n19042) );
  nand_x1_sg U51615 ( .A(\shifter_0/n9453 ), .B(n33206), .X(n19095) );
  nand_x1_sg U51616 ( .A(ow_2[1]), .B(n34787), .X(n19096) );
  nand_x1_sg U51617 ( .A(\shifter_0/n9452 ), .B(n33162), .X(n19097) );
  nand_x1_sg U51618 ( .A(ow_2[0]), .B(n31931), .X(n19098) );
  nand_x1_sg U51619 ( .A(\shifter_0/n9431 ), .B(n31221), .X(n19099) );
  nand_x1_sg U51620 ( .A(ow_3[19]), .B(n32581), .X(n19100) );
  nand_x1_sg U51621 ( .A(\shifter_0/n9430 ), .B(n31226), .X(n19101) );
  nand_x1_sg U51622 ( .A(ow_3[18]), .B(n32591), .X(n19102) );
  nand_x1_sg U51623 ( .A(\shifter_0/n9429 ), .B(n29867), .X(n19103) );
  nand_x1_sg U51624 ( .A(ow_3[17]), .B(n30663), .X(n19104) );
  nand_x1_sg U51625 ( .A(\shifter_0/n9428 ), .B(n33221), .X(n19105) );
  nand_x1_sg U51626 ( .A(ow_3[16]), .B(n32564), .X(n19106) );
  nand_x1_sg U51627 ( .A(\shifter_0/n9427 ), .B(n33201), .X(n19107) );
  nand_x1_sg U51628 ( .A(ow_3[15]), .B(n32544), .X(n19108) );
  nand_x1_sg U51629 ( .A(\shifter_0/n9426 ), .B(n29843), .X(n19109) );
  nand_x1_sg U51630 ( .A(ow_3[14]), .B(n30659), .X(n19110) );
  nand_x1_sg U51631 ( .A(\shifter_0/n9425 ), .B(n31549), .X(n19111) );
  nand_x1_sg U51632 ( .A(ow_3[13]), .B(n34756), .X(n19112) );
  nand_x1_sg U51633 ( .A(\shifter_0/n9424 ), .B(n31553), .X(n19113) );
  nand_x1_sg U51634 ( .A(ow_3[12]), .B(n32549), .X(n19114) );
  nand_x1_sg U51635 ( .A(\shifter_0/n9423 ), .B(n33166), .X(n19115) );
  nand_x1_sg U51636 ( .A(ow_3[11]), .B(n32569), .X(n19116) );
  nand_x1_sg U51637 ( .A(\shifter_0/n9422 ), .B(n31219), .X(n19117) );
  nand_x1_sg U51638 ( .A(ow_3[10]), .B(n32609), .X(n19118) );
  nand_x1_sg U51639 ( .A(\shifter_0/n9421 ), .B(n33138), .X(n19119) );
  nand_x1_sg U51640 ( .A(ow_3[9]), .B(n30657), .X(n19120) );
  nand_x1_sg U51641 ( .A(\shifter_0/n9420 ), .B(n33149), .X(n19121) );
  nand_x1_sg U51642 ( .A(ow_3[8]), .B(n30663), .X(n19122) );
  nand_x1_sg U51643 ( .A(\shifter_0/n9379 ), .B(n33159), .X(n19163) );
  nand_x1_sg U51644 ( .A(ow_4[7]), .B(n30665), .X(n19164) );
  nand_x1_sg U51645 ( .A(\shifter_0/n9378 ), .B(n35001), .X(n19165) );
  nand_x1_sg U51646 ( .A(ow_4[6]), .B(n32575), .X(n19166) );
  nand_x1_sg U51647 ( .A(\shifter_0/n9377 ), .B(n31537), .X(n19167) );
  nand_x1_sg U51648 ( .A(ow_4[5]), .B(n34500), .X(n19168) );
  nand_x1_sg U51649 ( .A(\shifter_0/n9376 ), .B(n33157), .X(n19169) );
  nand_x1_sg U51650 ( .A(ow_4[4]), .B(n32543), .X(n19170) );
  nand_x1_sg U51651 ( .A(\shifter_0/n9375 ), .B(n33178), .X(n19171) );
  nand_x1_sg U51652 ( .A(ow_4[3]), .B(n30799), .X(n19172) );
  nand_x1_sg U51653 ( .A(\shifter_0/n9374 ), .B(n33137), .X(n19173) );
  nand_x1_sg U51654 ( .A(ow_4[2]), .B(n34494), .X(n19174) );
  nand_x1_sg U51655 ( .A(\shifter_0/n9373 ), .B(n35008), .X(n19175) );
  nand_x1_sg U51656 ( .A(ow_4[1]), .B(n30660), .X(n19176) );
  nand_x1_sg U51657 ( .A(\shifter_0/n9372 ), .B(n33200), .X(n19177) );
  nand_x1_sg U51658 ( .A(ow_4[0]), .B(n31932), .X(n19178) );
  nand_x1_sg U51659 ( .A(\shifter_0/n9351 ), .B(n33143), .X(n19179) );
  nand_x1_sg U51660 ( .A(ow_5[19]), .B(n32597), .X(n19180) );
  nand_x1_sg U51661 ( .A(\shifter_0/n9350 ), .B(n31549), .X(n19181) );
  nand_x1_sg U51662 ( .A(ow_5[18]), .B(n34947), .X(n19182) );
  nand_x1_sg U51663 ( .A(\shifter_0/n9349 ), .B(n33178), .X(n19183) );
  nand_x1_sg U51664 ( .A(ow_5[17]), .B(n32575), .X(n19184) );
  nand_x1_sg U51665 ( .A(\shifter_0/n9348 ), .B(n33150), .X(n19185) );
  nand_x1_sg U51666 ( .A(ow_5[16]), .B(n34776), .X(n19186) );
  nand_x1_sg U51667 ( .A(\shifter_0/n9347 ), .B(n29851), .X(n19187) );
  nand_x1_sg U51668 ( .A(ow_5[15]), .B(n32561), .X(n19188) );
  nand_x1_sg U51669 ( .A(\shifter_0/n9346 ), .B(n31537), .X(n19189) );
  nand_x1_sg U51670 ( .A(ow_5[14]), .B(n30655), .X(n19190) );
  nand_x1_sg U51671 ( .A(\shifter_0/n9345 ), .B(n31534), .X(n19191) );
  nand_x1_sg U51672 ( .A(ow_5[13]), .B(n34951), .X(n19192) );
  nand_x1_sg U51673 ( .A(\shifter_0/n9344 ), .B(n34988), .X(n19193) );
  nand_x1_sg U51674 ( .A(ow_5[12]), .B(n30669), .X(n19194) );
  nand_x1_sg U51675 ( .A(\shifter_0/n9343 ), .B(n31222), .X(n19195) );
  nand_x1_sg U51676 ( .A(ow_5[11]), .B(n32629), .X(n19196) );
  nand_x1_sg U51677 ( .A(\shifter_0/n9342 ), .B(n34999), .X(n19197) );
  nand_x1_sg U51678 ( .A(ow_5[10]), .B(n32546), .X(n19198) );
  nand_x1_sg U51679 ( .A(\shifter_0/n9341 ), .B(n31224), .X(n19199) );
  nand_x1_sg U51680 ( .A(ow_5[9]), .B(n32622), .X(n19200) );
  nand_x1_sg U51681 ( .A(\shifter_0/n9340 ), .B(n33214), .X(n19201) );
  nand_x1_sg U51682 ( .A(ow_5[8]), .B(n34493), .X(n19202) );
  nand_x1_sg U51683 ( .A(\shifter_0/n9179 ), .B(n34982), .X(n19363) );
  nand_x1_sg U51684 ( .A(ow_9[7]), .B(n32558), .X(n19364) );
  nand_x1_sg U51685 ( .A(\shifter_0/n9178 ), .B(n31550), .X(n19365) );
  nand_x1_sg U51686 ( .A(ow_9[6]), .B(n32605), .X(n19366) );
  nand_x1_sg U51687 ( .A(\shifter_0/n9177 ), .B(n34987), .X(n19367) );
  nand_x1_sg U51688 ( .A(ow_9[5]), .B(n30656), .X(n19368) );
  nand_x1_sg U51689 ( .A(\shifter_0/n9176 ), .B(n33171), .X(n19369) );
  nand_x1_sg U51690 ( .A(ow_9[4]), .B(n34763), .X(n19370) );
  nand_x1_sg U51691 ( .A(\shifter_0/n9175 ), .B(n33148), .X(n19371) );
  nand_x1_sg U51692 ( .A(ow_9[3]), .B(n30795), .X(n19372) );
  nand_x1_sg U51693 ( .A(\shifter_0/n9174 ), .B(n29860), .X(n19373) );
  nand_x1_sg U51694 ( .A(ow_9[2]), .B(n32572), .X(n19374) );
  nand_x1_sg U51695 ( .A(\shifter_0/n9173 ), .B(n29844), .X(n19375) );
  nand_x1_sg U51696 ( .A(ow_9[1]), .B(n32609), .X(n19376) );
  nand_x1_sg U51697 ( .A(\shifter_0/n9172 ), .B(n33132), .X(n19377) );
  nand_x1_sg U51698 ( .A(ow_9[0]), .B(n34501), .X(n19378) );
  nand_x1_sg U51699 ( .A(\shifter_0/n9151 ), .B(n31548), .X(n19379) );
  nand_x1_sg U51700 ( .A(ow_10[19]), .B(n32551), .X(n19380) );
  nand_x1_sg U51701 ( .A(\shifter_0/n9150 ), .B(n34980), .X(n19381) );
  nand_x1_sg U51702 ( .A(ow_10[18]), .B(n32557), .X(n19382) );
  nand_x1_sg U51703 ( .A(\shifter_0/n9149 ), .B(n33165), .X(n19383) );
  nand_x1_sg U51704 ( .A(ow_10[17]), .B(n31930), .X(n19384) );
  nand_x1_sg U51705 ( .A(\shifter_0/n9148 ), .B(n33199), .X(n19385) );
  nand_x1_sg U51706 ( .A(ow_10[16]), .B(n32616), .X(n19386) );
  nand_x1_sg U51707 ( .A(\shifter_0/n9147 ), .B(n34987), .X(n19387) );
  nand_x1_sg U51708 ( .A(ow_10[15]), .B(n30125), .X(n19388) );
  nand_x1_sg U51709 ( .A(\shifter_0/n9146 ), .B(n33178), .X(n19389) );
  nand_x1_sg U51710 ( .A(ow_10[14]), .B(n34772), .X(n19390) );
  nand_x1_sg U51711 ( .A(\shifter_0/n9145 ), .B(n33155), .X(n19391) );
  nand_x1_sg U51712 ( .A(ow_10[13]), .B(n32096), .X(n19392) );
  nand_x1_sg U51713 ( .A(\shifter_0/n9144 ), .B(n33136), .X(n19393) );
  nand_x1_sg U51714 ( .A(ow_10[12]), .B(n32627), .X(n19394) );
  nand_x1_sg U51715 ( .A(\shifter_0/n9143 ), .B(n31540), .X(n19395) );
  nand_x1_sg U51716 ( .A(ow_10[11]), .B(n32544), .X(n19396) );
  nand_x1_sg U51717 ( .A(\shifter_0/n9142 ), .B(n33219), .X(n19397) );
  nand_x1_sg U51718 ( .A(ow_10[10]), .B(n30124), .X(n19398) );
  nand_x1_sg U51719 ( .A(\shifter_0/n9141 ), .B(n33133), .X(n19399) );
  nand_x1_sg U51720 ( .A(ow_10[9]), .B(n30651), .X(n19400) );
  nand_x1_sg U51721 ( .A(\shifter_0/n9140 ), .B(n33212), .X(n19401) );
  nand_x1_sg U51722 ( .A(ow_10[8]), .B(n32557), .X(n19402) );
  nand_x1_sg U51723 ( .A(\shifter_0/n9099 ), .B(n33827), .X(n19443) );
  nand_x1_sg U51724 ( .A(ow_11[7]), .B(n34496), .X(n19444) );
  nand_x1_sg U51725 ( .A(\shifter_0/n9098 ), .B(n34976), .X(n19445) );
  nand_x1_sg U51726 ( .A(ow_11[6]), .B(n32585), .X(n19446) );
  nand_x1_sg U51727 ( .A(\shifter_0/n9097 ), .B(n35003), .X(n19447) );
  nand_x1_sg U51728 ( .A(ow_11[5]), .B(n32623), .X(n19448) );
  nand_x1_sg U51729 ( .A(\shifter_0/n9096 ), .B(n33192), .X(n19449) );
  nand_x1_sg U51730 ( .A(ow_11[4]), .B(n34781), .X(n19450) );
  nand_x1_sg U51731 ( .A(\shifter_0/n9095 ), .B(n31553), .X(n19451) );
  nand_x1_sg U51732 ( .A(ow_11[3]), .B(n32573), .X(n19452) );
  nand_x1_sg U51733 ( .A(\shifter_0/n9094 ), .B(n35004), .X(n19453) );
  nand_x1_sg U51734 ( .A(ow_11[2]), .B(n32582), .X(n19454) );
  nand_x1_sg U51735 ( .A(\shifter_0/n9093 ), .B(n33161), .X(n19455) );
  nand_x1_sg U51736 ( .A(ow_11[1]), .B(n32580), .X(n19456) );
  nand_x1_sg U51737 ( .A(\shifter_0/n9092 ), .B(n33166), .X(n19457) );
  nand_x1_sg U51738 ( .A(ow_11[0]), .B(n32618), .X(n19458) );
  nand_x1_sg U51739 ( .A(\shifter_0/n9071 ), .B(n29839), .X(n19459) );
  nand_x1_sg U51740 ( .A(ow_12[19]), .B(n34784), .X(n19460) );
  nand_x1_sg U51741 ( .A(\shifter_0/n9070 ), .B(n31540), .X(n19461) );
  nand_x1_sg U51742 ( .A(ow_12[18]), .B(n32601), .X(n19462) );
  nand_x1_sg U51743 ( .A(\shifter_0/n9069 ), .B(n33178), .X(n19463) );
  nand_x1_sg U51744 ( .A(ow_12[17]), .B(n30668), .X(n19464) );
  nand_x1_sg U51745 ( .A(\shifter_0/n9068 ), .B(n31541), .X(n19465) );
  nand_x1_sg U51746 ( .A(ow_12[16]), .B(n32565), .X(n19466) );
  nand_x1_sg U51747 ( .A(\shifter_0/n9067 ), .B(n33204), .X(n19467) );
  nand_x1_sg U51748 ( .A(ow_12[15]), .B(n32574), .X(n19468) );
  nand_x1_sg U51749 ( .A(\shifter_0/n9066 ), .B(n33159), .X(n19469) );
  nand_x1_sg U51750 ( .A(ow_12[14]), .B(n34768), .X(n19470) );
  nand_x1_sg U51751 ( .A(\shifter_0/n9065 ), .B(n35007), .X(n19471) );
  nand_x1_sg U51752 ( .A(ow_12[13]), .B(n32633), .X(n19472) );
  nand_x1_sg U51753 ( .A(\shifter_0/n9064 ), .B(n29856), .X(n19473) );
  nand_x1_sg U51754 ( .A(ow_12[12]), .B(n32573), .X(n19474) );
  nand_x1_sg U51755 ( .A(\shifter_0/n9063 ), .B(n30223), .X(n19475) );
  nand_x1_sg U51756 ( .A(ow_12[11]), .B(n32622), .X(n19476) );
  nand_x1_sg U51757 ( .A(\shifter_0/n9062 ), .B(n31552), .X(n19477) );
  nand_x1_sg U51758 ( .A(ow_12[10]), .B(n30214), .X(n19478) );
  nand_x1_sg U51759 ( .A(\shifter_0/n9061 ), .B(n31227), .X(n19479) );
  nand_x1_sg U51760 ( .A(ow_12[9]), .B(n32555), .X(n19480) );
  nand_x1_sg U51761 ( .A(\shifter_0/n9060 ), .B(n33203), .X(n19481) );
  nand_x1_sg U51762 ( .A(ow_12[8]), .B(n32633), .X(n19482) );
  nand_x1_sg U51763 ( .A(\shifter_0/n9018 ), .B(n33160), .X(n19525) );
  nand_x1_sg U51764 ( .A(ow_13[6]), .B(n34767), .X(n19526) );
  nand_x1_sg U51765 ( .A(\shifter_0/n9017 ), .B(n33136), .X(n19527) );
  nand_x1_sg U51766 ( .A(ow_13[5]), .B(n34495), .X(n19528) );
  nand_x1_sg U51767 ( .A(\shifter_0/n9016 ), .B(n31542), .X(n19529) );
  nand_x1_sg U51768 ( .A(ow_13[4]), .B(n30663), .X(n19530) );
  nand_x1_sg U51769 ( .A(\shifter_0/n9399 ), .B(n29867), .X(n21969) );
  nand_x1_sg U51770 ( .A(oi_4[7]), .B(n34773), .X(n21970) );
  nand_x1_sg U51771 ( .A(\shifter_0/n9398 ), .B(n33208), .X(n21971) );
  nand_x1_sg U51772 ( .A(oi_4[6]), .B(n32545), .X(n21972) );
  nand_x1_sg U51773 ( .A(\shifter_0/n9397 ), .B(n33203), .X(n21973) );
  nand_x1_sg U51774 ( .A(oi_4[5]), .B(n32632), .X(n21974) );
  nand_x1_sg U51775 ( .A(\shifter_0/n9396 ), .B(n33179), .X(n21975) );
  nand_x1_sg U51776 ( .A(oi_4[4]), .B(n32633), .X(n21976) );
  nand_x1_sg U51777 ( .A(\shifter_0/n9395 ), .B(n33192), .X(n21977) );
  nand_x1_sg U51778 ( .A(oi_4[3]), .B(n34759), .X(n21978) );
  nand_x1_sg U51779 ( .A(\shifter_0/n9394 ), .B(n29851), .X(n21979) );
  nand_x1_sg U51780 ( .A(oi_4[2]), .B(n32553), .X(n21980) );
  nand_x1_sg U51781 ( .A(\shifter_0/n9393 ), .B(n33183), .X(n21981) );
  nand_x1_sg U51782 ( .A(oi_4[1]), .B(n34771), .X(n21982) );
  nand_x1_sg U51783 ( .A(\shifter_0/n9392 ), .B(n33176), .X(n21983) );
  nand_x1_sg U51784 ( .A(oi_4[0]), .B(n32589), .X(n21984) );
  nand_x1_sg U51785 ( .A(\shifter_0/n9371 ), .B(n33207), .X(n21985) );
  nand_x1_sg U51786 ( .A(oi_5[19]), .B(n32622), .X(n21986) );
  nand_x1_sg U51787 ( .A(\shifter_0/n9370 ), .B(n33194), .X(n21987) );
  nand_x1_sg U51788 ( .A(oi_5[18]), .B(n32611), .X(n21988) );
  nand_x1_sg U51789 ( .A(\shifter_0/n9369 ), .B(n33204), .X(n21989) );
  nand_x1_sg U51790 ( .A(oi_5[17]), .B(n34782), .X(n21990) );
  nand_x1_sg U51791 ( .A(\shifter_0/n9368 ), .B(n31548), .X(n21991) );
  nand_x1_sg U51792 ( .A(oi_5[16]), .B(n34758), .X(n21992) );
  nand_x1_sg U51793 ( .A(\shifter_0/n9367 ), .B(n29846), .X(n21993) );
  nand_x1_sg U51794 ( .A(oi_5[15]), .B(n34759), .X(n21994) );
  nand_x1_sg U51795 ( .A(\shifter_0/n9366 ), .B(n33167), .X(n21995) );
  nand_x1_sg U51796 ( .A(oi_5[14]), .B(n32572), .X(n21996) );
  nand_x1_sg U51797 ( .A(\shifter_0/n9365 ), .B(n34981), .X(n21997) );
  nand_x1_sg U51798 ( .A(oi_5[13]), .B(n32556), .X(n21998) );
  nand_x1_sg U51799 ( .A(\shifter_0/n9364 ), .B(n33192), .X(n21999) );
  nand_x1_sg U51800 ( .A(oi_5[12]), .B(n32604), .X(n22000) );
  nand_x1_sg U51801 ( .A(\shifter_0/n9363 ), .B(n35005), .X(n22001) );
  nand_x1_sg U51802 ( .A(oi_5[11]), .B(n30659), .X(n22002) );
  nand_x1_sg U51803 ( .A(\shifter_0/n9362 ), .B(n31542), .X(n22003) );
  nand_x1_sg U51804 ( .A(oi_5[10]), .B(n32573), .X(n22004) );
  nand_x1_sg U51805 ( .A(\shifter_0/n9361 ), .B(n33824), .X(n22005) );
  nand_x1_sg U51806 ( .A(oi_5[9]), .B(n32635), .X(n22006) );
  nand_x1_sg U51807 ( .A(\shifter_0/n9360 ), .B(n33152), .X(n22007) );
  nand_x1_sg U51808 ( .A(oi_5[8]), .B(n32548), .X(n22008) );
  nand_x1_sg U51809 ( .A(\shifter_0/n9539 ), .B(n33144), .X(n19003) );
  nand_x1_sg U51810 ( .A(ow_0[7]), .B(n32606), .X(n19004) );
  nand_x1_sg U51811 ( .A(\shifter_0/n9538 ), .B(n31555), .X(n19005) );
  nand_x1_sg U51812 ( .A(ow_0[6]), .B(n34757), .X(n19006) );
  nand_x1_sg U51813 ( .A(\shifter_0/n9537 ), .B(n31538), .X(n19007) );
  nand_x1_sg U51814 ( .A(ow_0[5]), .B(n32567), .X(n19008) );
  nand_x1_sg U51815 ( .A(\shifter_0/n9536 ), .B(n31549), .X(n19009) );
  nand_x1_sg U51816 ( .A(ow_0[4]), .B(n32618), .X(n19010) );
  nand_x1_sg U51817 ( .A(\shifter_0/n9535 ), .B(n33213), .X(n19011) );
  nand_x1_sg U51818 ( .A(ow_0[3]), .B(n34762), .X(n19012) );
  nand_x1_sg U51819 ( .A(\shifter_0/n9534 ), .B(n33196), .X(n19013) );
  nand_x1_sg U51820 ( .A(ow_0[2]), .B(n32635), .X(n19014) );
  nand_x1_sg U51821 ( .A(\shifter_0/n9533 ), .B(n29847), .X(n19015) );
  nand_x1_sg U51822 ( .A(ow_0[1]), .B(n32601), .X(n19016) );
  nand_x1_sg U51823 ( .A(\shifter_0/n9532 ), .B(n33140), .X(n19017) );
  nand_x1_sg U51824 ( .A(ow_0[0]), .B(n34789), .X(n19018) );
  nand_x1_sg U51825 ( .A(\shifter_0/n9459 ), .B(n33173), .X(n19083) );
  nand_x1_sg U51826 ( .A(ow_2[7]), .B(n32094), .X(n19084) );
  nand_x1_sg U51827 ( .A(\shifter_0/n9458 ), .B(n33168), .X(n19085) );
  nand_x1_sg U51828 ( .A(ow_2[6]), .B(n32609), .X(n19086) );
  nand_x1_sg U51829 ( .A(\shifter_0/n9457 ), .B(n29853), .X(n19087) );
  nand_x1_sg U51830 ( .A(ow_2[5]), .B(n34756), .X(n19088) );
  nand_x1_sg U51831 ( .A(\shifter_0/n9019 ), .B(n33202), .X(n19523) );
  nand_x1_sg U51832 ( .A(ow_13[7]), .B(n34774), .X(n19524) );
  nand_x1_sg U51833 ( .A(\shifter_0/n9012 ), .B(n34979), .X(n19537) );
  nand_x1_sg U51834 ( .A(ow_13[0]), .B(n32098), .X(n19538) );
  nand_x1_sg U51835 ( .A(\shifter_0/n8991 ), .B(n33190), .X(n19539) );
  nand_x1_sg U51836 ( .A(ow_14[19]), .B(n34779), .X(n19540) );
  nand_x1_sg U51837 ( .A(\shifter_0/n8990 ), .B(n31554), .X(n19541) );
  nand_x1_sg U51838 ( .A(ow_14[18]), .B(n34769), .X(n19542) );
  nand_x1_sg U51839 ( .A(\shifter_0/n8989 ), .B(n29850), .X(n19543) );
  nand_x1_sg U51840 ( .A(ow_14[17]), .B(n32593), .X(n19544) );
  nand_x1_sg U51841 ( .A(\shifter_0/n8988 ), .B(n33176), .X(n19545) );
  nand_x1_sg U51842 ( .A(ow_14[16]), .B(n30799), .X(n19546) );
  nand_x1_sg U51843 ( .A(\shifter_0/n8987 ), .B(n33215), .X(n19547) );
  nand_x1_sg U51844 ( .A(ow_14[15]), .B(n30649), .X(n19548) );
  nand_x1_sg U51845 ( .A(\shifter_0/n8986 ), .B(n35009), .X(n19549) );
  nand_x1_sg U51846 ( .A(ow_14[14]), .B(n32580), .X(n19550) );
  nand_x1_sg U51847 ( .A(\shifter_0/n8985 ), .B(n29847), .X(n19551) );
  nand_x1_sg U51848 ( .A(ow_14[13]), .B(n34945), .X(n19552) );
  nand_x1_sg U51849 ( .A(\shifter_0/n8984 ), .B(n30236), .X(n19553) );
  nand_x1_sg U51850 ( .A(ow_14[12]), .B(n34774), .X(n19554) );
  nand_x1_sg U51851 ( .A(\shifter_0/n8983 ), .B(n31225), .X(n19555) );
  nand_x1_sg U51852 ( .A(ow_14[11]), .B(n32592), .X(n19556) );
  nand_x1_sg U51853 ( .A(\shifter_0/n8982 ), .B(n33136), .X(n19557) );
  nand_x1_sg U51854 ( .A(ow_14[10]), .B(n32589), .X(n19558) );
  nand_x1_sg U51855 ( .A(\shifter_0/n8981 ), .B(n33157), .X(n19559) );
  nand_x1_sg U51856 ( .A(ow_14[9]), .B(n30798), .X(n19560) );
  nand_x1_sg U51857 ( .A(\shifter_0/n8980 ), .B(n29860), .X(n19561) );
  nand_x1_sg U51858 ( .A(ow_14[8]), .B(n32625), .X(n19562) );
  nor_x1_sg U51859 ( .A(n35457), .B(n26196), .X(n26195) );
  nand_x1_sg U51860 ( .A(n42414), .B(output_taken), .X(n26196) );
  inv_x1_sg U51861 ( .A(state[0]), .X(n42414) );
  nand_x1_sg U51862 ( .A(reg_iii_2[4]), .B(n32775), .X(n26004) );
  nand_x1_sg U51863 ( .A(reg_ii_2[4]), .B(n32837), .X(n26005) );
  nand_x1_sg U51864 ( .A(reg_iii_2[5]), .B(n31926), .X(n26006) );
  nand_x1_sg U51865 ( .A(reg_ii_2[5]), .B(n30859), .X(n26007) );
  nand_x1_sg U51866 ( .A(reg_iii_2[7]), .B(n32239), .X(n26010) );
  nand_x1_sg U51867 ( .A(reg_ii_2[7]), .B(n35233), .X(n26011) );
  nand_x1_sg U51868 ( .A(reg_iii_2[8]), .B(n32018), .X(n26012) );
  nand_x1_sg U51869 ( .A(reg_ii_2[8]), .B(n30874), .X(n26013) );
  nand_x1_sg U51870 ( .A(reg_iii_2[10]), .B(n31727), .X(n26016) );
  nand_x1_sg U51871 ( .A(reg_ii_2[10]), .B(n34724), .X(n26017) );
  nand_x1_sg U51872 ( .A(reg_iii_2[11]), .B(n30014), .X(n26018) );
  nand_x1_sg U51873 ( .A(reg_ii_2[11]), .B(n35344), .X(n26019) );
  nand_x1_sg U51874 ( .A(reg_iii_2[13]), .B(n31639), .X(n26022) );
  nand_x1_sg U51875 ( .A(reg_ii_2[13]), .B(n31096), .X(n26023) );
  nand_x1_sg U51876 ( .A(reg_iii_2[14]), .B(n31634), .X(n26024) );
  nand_x1_sg U51877 ( .A(reg_ii_2[14]), .B(n31097), .X(n26025) );
  nand_x1_sg U51878 ( .A(reg_iii_2[16]), .B(n32010), .X(n26028) );
  nand_x1_sg U51879 ( .A(reg_ii_2[16]), .B(n35217), .X(n26029) );
  nand_x1_sg U51880 ( .A(reg_iii_2[17]), .B(n32450), .X(n26030) );
  nand_x1_sg U51881 ( .A(reg_ii_2[17]), .B(n32840), .X(n26031) );
  nand_x1_sg U51882 ( .A(reg_iii_2[19]), .B(n32248), .X(n26034) );
  nand_x1_sg U51883 ( .A(reg_ii_2[19]), .B(n32753), .X(n26035) );
  nand_x1_sg U51884 ( .A(reg_iii_4[0]), .B(n32216), .X(n26154) );
  nand_x1_sg U51885 ( .A(reg_ii_4[0]), .B(n31672), .X(n26155) );
  nand_x1_sg U51886 ( .A(reg_iii_4[1]), .B(n32011), .X(n26156) );
  nand_x1_sg U51887 ( .A(reg_ii_4[1]), .B(n35200), .X(n26157) );
  nand_x1_sg U51888 ( .A(reg_iii_4[3]), .B(n32333), .X(n26160) );
  nand_x1_sg U51889 ( .A(reg_ii_4[3]), .B(n35237), .X(n26161) );
  nand_x1_sg U51890 ( .A(reg_iii_4[4]), .B(n32010), .X(n26162) );
  nand_x1_sg U51891 ( .A(reg_ii_4[4]), .B(n32744), .X(n26163) );
  nand_x1_sg U51892 ( .A(reg_iii_4[6]), .B(n32496), .X(n26166) );
  nand_x1_sg U51893 ( .A(reg_ii_4[6]), .B(n30866), .X(n26167) );
  nand_x1_sg U51894 ( .A(reg_iii_4[7]), .B(n34580), .X(n26168) );
  nand_x1_sg U51895 ( .A(reg_ii_4[7]), .B(n32753), .X(n26169) );
  nand_x1_sg U51896 ( .A(reg_iii_4[9]), .B(n32246), .X(n26172) );
  nand_x1_sg U51897 ( .A(reg_ii_4[9]), .B(n35191), .X(n26173) );
  nand_x1_sg U51898 ( .A(reg_iii_4[10]), .B(n32456), .X(n26174) );
  nand_x1_sg U51899 ( .A(reg_ii_4[10]), .B(n32442), .X(n26175) );
  nand_x1_sg U51900 ( .A(reg_iii_4[12]), .B(n34566), .X(n26178) );
  nand_x1_sg U51901 ( .A(reg_ii_4[12]), .B(n30866), .X(n26179) );
  nand_x1_sg U51902 ( .A(reg_iii_4[13]), .B(n34653), .X(n26180) );
  nand_x1_sg U51903 ( .A(reg_ii_4[13]), .B(n35221), .X(n26181) );
  nand_x1_sg U51904 ( .A(reg_iii_4[15]), .B(n32453), .X(n26184) );
  nand_x1_sg U51905 ( .A(reg_ii_4[15]), .B(n35161), .X(n26185) );
  nand_x1_sg U51906 ( .A(reg_iii_4[16]), .B(n31716), .X(n26186) );
  nand_x1_sg U51907 ( .A(reg_ii_4[16]), .B(n35330), .X(n26187) );
  nand_x1_sg U51908 ( .A(reg_iii_4[18]), .B(n32156), .X(n26190) );
  nand_x1_sg U51909 ( .A(reg_ii_4[18]), .B(n32742), .X(n26191) );
  nand_x1_sg U51910 ( .A(reg_iii_4[19]), .B(n32777), .X(n26192) );
  nand_x1_sg U51911 ( .A(reg_ii_4[19]), .B(n35200), .X(n26193) );
  nand_x1_sg U51912 ( .A(reg_iii_5[0]), .B(n32856), .X(n25440) );
  nand_x1_sg U51913 ( .A(reg_ii_5[0]), .B(n35215), .X(n25441) );
  nand_x1_sg U51914 ( .A(reg_iii_5[1]), .B(n31636), .X(n25442) );
  nand_x1_sg U51915 ( .A(reg_ii_5[1]), .B(n30718), .X(n25443) );
  nand_x1_sg U51916 ( .A(reg_iii_5[3]), .B(n31643), .X(n25446) );
  nand_x1_sg U51917 ( .A(reg_ii_5[3]), .B(n30868), .X(n25447) );
  nand_x1_sg U51918 ( .A(reg_iii_5[4]), .B(n31924), .X(n25448) );
  nand_x1_sg U51919 ( .A(reg_ii_5[4]), .B(n33996), .X(n25449) );
  nand_x1_sg U51920 ( .A(reg_iii_5[6]), .B(n32455), .X(n25452) );
  nand_x1_sg U51921 ( .A(reg_ii_5[6]), .B(n35163), .X(n25453) );
  nand_x1_sg U51922 ( .A(reg_iii_5[7]), .B(n32251), .X(n25454) );
  nand_x1_sg U51923 ( .A(reg_ii_5[7]), .B(n30877), .X(n25455) );
  nand_x1_sg U51924 ( .A(reg_iii_5[9]), .B(n33977), .X(n25458) );
  nand_x1_sg U51925 ( .A(reg_ii_5[9]), .B(n32724), .X(n25459) );
  nand_x1_sg U51926 ( .A(reg_iii_5[10]), .B(n32019), .X(n25460) );
  nand_x1_sg U51927 ( .A(reg_ii_5[10]), .B(n31060), .X(n25461) );
  nand_x1_sg U51928 ( .A(reg_iii_5[12]), .B(n32856), .X(n25464) );
  nand_x1_sg U51929 ( .A(reg_ii_5[12]), .B(n33997), .X(n25465) );
  nand_x1_sg U51930 ( .A(reg_iii_5[13]), .B(n31897), .X(n25466) );
  nand_x1_sg U51931 ( .A(reg_ii_5[13]), .B(n35186), .X(n25467) );
  nand_x1_sg U51932 ( .A(reg_iii_5[15]), .B(n34553), .X(n25470) );
  nand_x1_sg U51933 ( .A(reg_ii_5[15]), .B(n35091), .X(n25471) );
  nand_x1_sg U51934 ( .A(reg_iii_5[16]), .B(n32163), .X(n25472) );
  nand_x1_sg U51935 ( .A(reg_ii_5[16]), .B(n35084), .X(n25473) );
  nand_x1_sg U51936 ( .A(reg_iii_5[18]), .B(n32354), .X(n25476) );
  nand_x1_sg U51937 ( .A(reg_ii_5[18]), .B(n31092), .X(n25477) );
  nand_x1_sg U51938 ( .A(reg_iii_5[19]), .B(n32857), .X(n25478) );
  nand_x1_sg U51939 ( .A(reg_ii_5[19]), .B(n35370), .X(n25479) );
  nand_x1_sg U51940 ( .A(reg_iii_6[17]), .B(n31645), .X(n25554) );
  nand_x1_sg U51941 ( .A(reg_ii_6[17]), .B(n30863), .X(n25555) );
  nand_x1_sg U51942 ( .A(reg_iii_6[18]), .B(n31515), .X(n25556) );
  nand_x1_sg U51943 ( .A(reg_ii_6[18]), .B(n31092), .X(n25557) );
  nand_x1_sg U51944 ( .A(reg_iii_7[1]), .B(n30155), .X(n25602) );
  nand_x1_sg U51945 ( .A(reg_ii_7[1]), .B(n30747), .X(n25603) );
  nand_x1_sg U51946 ( .A(reg_iii_7[2]), .B(n30916), .X(n25604) );
  nand_x1_sg U51947 ( .A(reg_ii_7[2]), .B(n31031), .X(n25605) );
  nand_x1_sg U51948 ( .A(reg_iii_7[4]), .B(n31634), .X(n25608) );
  nand_x1_sg U51949 ( .A(reg_ii_7[4]), .B(n35345), .X(n25609) );
  nand_x1_sg U51950 ( .A(reg_iii_7[5]), .B(n31724), .X(n25610) );
  nand_x1_sg U51951 ( .A(reg_ii_7[5]), .B(n35377), .X(n25611) );
  nand_x1_sg U51952 ( .A(reg_iii_7[7]), .B(n32046), .X(n25614) );
  nand_x1_sg U51953 ( .A(reg_ii_7[7]), .B(n30595), .X(n25615) );
  nand_x1_sg U51954 ( .A(reg_iii_7[8]), .B(n31728), .X(n25616) );
  nand_x1_sg U51955 ( .A(reg_ii_7[8]), .B(n35403), .X(n25617) );
  nand_x1_sg U51956 ( .A(reg_iii_8[1]), .B(n31721), .X(n25682) );
  nand_x1_sg U51957 ( .A(reg_ii_8[1]), .B(n32842), .X(n25683) );
  nand_x1_sg U51958 ( .A(reg_iii_8[3]), .B(n34851), .X(n25686) );
  nand_x1_sg U51959 ( .A(reg_ii_8[3]), .B(n33996), .X(n25687) );
  nand_x1_sg U51960 ( .A(reg_iii_8[4]), .B(n32327), .X(n25688) );
  nand_x1_sg U51961 ( .A(reg_ii_8[4]), .B(n32835), .X(n25689) );
  nand_x1_sg U51962 ( .A(reg_iii_8[6]), .B(n32303), .X(n25692) );
  nand_x1_sg U51963 ( .A(reg_ii_8[6]), .B(n35396), .X(n25693) );
  nand_x1_sg U51964 ( .A(reg_iii_8[7]), .B(n31642), .X(n25694) );
  nand_x1_sg U51965 ( .A(reg_ii_8[7]), .B(n34001), .X(n25695) );
  nand_x1_sg U51966 ( .A(reg_iii_8[9]), .B(n32246), .X(n25698) );
  nand_x1_sg U51967 ( .A(reg_ii_8[9]), .B(n30889), .X(n25699) );
  nand_x1_sg U51968 ( .A(reg_iii_8[10]), .B(n32451), .X(n25700) );
  nand_x1_sg U51969 ( .A(reg_ii_8[10]), .B(n30882), .X(n25701) );
  nand_x1_sg U51970 ( .A(reg_iii_8[12]), .B(n34653), .X(n25704) );
  nand_x1_sg U51971 ( .A(reg_ii_8[12]), .B(n35327), .X(n25705) );
  nand_x1_sg U51972 ( .A(reg_iii_8[13]), .B(n35080), .X(n25706) );
  nand_x1_sg U51973 ( .A(reg_ii_8[13]), .B(n31025), .X(n25707) );
  nand_x1_sg U51974 ( .A(reg_iii_8[15]), .B(n35078), .X(n25710) );
  nand_x1_sg U51975 ( .A(reg_ii_8[15]), .B(n31029), .X(n25711) );
  nand_x1_sg U51976 ( .A(reg_iii_8[16]), .B(n32340), .X(n25712) );
  nand_x1_sg U51977 ( .A(reg_ii_8[16]), .B(n35090), .X(n25713) );
  nand_x1_sg U51978 ( .A(reg_iii_8[18]), .B(n30014), .X(n25716) );
  nand_x1_sg U51979 ( .A(reg_ii_8[18]), .B(n30587), .X(n25717) );
  nand_x1_sg U51980 ( .A(reg_iii_8[19]), .B(n32036), .X(n25718) );
  nand_x1_sg U51981 ( .A(reg_ii_8[19]), .B(n35404), .X(n25719) );
  nand_x1_sg U51982 ( .A(reg_iii_11[0]), .B(n32378), .X(n25124) );
  nand_x1_sg U51983 ( .A(reg_ii_11[0]), .B(n30874), .X(n25125) );
  nand_x1_sg U51984 ( .A(reg_iii_11[2]), .B(n32030), .X(n25128) );
  nand_x1_sg U51985 ( .A(reg_ii_11[2]), .B(n31058), .X(n25129) );
  nand_x1_sg U51986 ( .A(reg_iii_11[3]), .B(n34940), .X(n25130) );
  nand_x1_sg U51987 ( .A(reg_ii_11[3]), .B(n30877), .X(n25131) );
  nand_x1_sg U51988 ( .A(reg_iii_11[5]), .B(n33952), .X(n25134) );
  nand_x1_sg U51989 ( .A(reg_ii_11[5]), .B(n32716), .X(n25135) );
  nand_x1_sg U51990 ( .A(reg_iii_11[6]), .B(n31894), .X(n25136) );
  nand_x1_sg U51991 ( .A(reg_ii_11[6]), .B(n31097), .X(n25137) );
  nand_x1_sg U51992 ( .A(reg_iii_11[8]), .B(n32403), .X(n25140) );
  nand_x1_sg U51993 ( .A(reg_ii_11[8]), .B(n32726), .X(n25141) );
  nand_x1_sg U51994 ( .A(reg_iii_11[9]), .B(n33971), .X(n25142) );
  nand_x1_sg U51995 ( .A(reg_ii_11[9]), .B(n34667), .X(n25143) );
  nand_x1_sg U51996 ( .A(reg_iii_11[11]), .B(n31723), .X(n25146) );
  nand_x1_sg U51997 ( .A(reg_ii_11[11]), .B(n32440), .X(n25147) );
  nand_x1_sg U51998 ( .A(reg_iii_11[12]), .B(n31640), .X(n25148) );
  nand_x1_sg U51999 ( .A(reg_ii_11[12]), .B(n35173), .X(n25149) );
  nand_x1_sg U52000 ( .A(reg_iii_11[14]), .B(n32372), .X(n25152) );
  nand_x1_sg U52001 ( .A(reg_ii_11[14]), .B(n30903), .X(n25153) );
  nand_x1_sg U52002 ( .A(reg_iii_11[15]), .B(n31503), .X(n25154) );
  nand_x1_sg U52003 ( .A(reg_ii_11[15]), .B(n35336), .X(n25155) );
  nand_x1_sg U52004 ( .A(reg_iii_11[17]), .B(n33950), .X(n25158) );
  nand_x1_sg U52005 ( .A(reg_ii_11[17]), .B(n32757), .X(n25159) );
  nand_x1_sg U52006 ( .A(reg_iii_11[18]), .B(n32150), .X(n25160) );
  nand_x1_sg U52007 ( .A(reg_ii_11[18]), .B(n34719), .X(n25161) );
  nand_x1_sg U52008 ( .A(reg_www_2[0]), .B(n31890), .X(n24888) );
  nand_x1_sg U52009 ( .A(reg_ww_2[0]), .B(n30722), .X(n24889) );
  nand_x1_sg U52010 ( .A(reg_www_2[1]), .B(n32344), .X(n24890) );
  nand_x1_sg U52011 ( .A(reg_ww_2[1]), .B(n32714), .X(n24891) );
  nand_x1_sg U52012 ( .A(reg_www_2[3]), .B(n34650), .X(n24894) );
  nand_x1_sg U52013 ( .A(reg_ww_2[3]), .B(n35327), .X(n24895) );
  nand_x1_sg U52014 ( .A(reg_www_2[4]), .B(n31630), .X(n24896) );
  nand_x1_sg U52015 ( .A(reg_ww_2[4]), .B(n32729), .X(n24897) );
  nand_x1_sg U52016 ( .A(reg_www_2[6]), .B(n32141), .X(n24900) );
  nand_x1_sg U52017 ( .A(reg_ww_2[6]), .B(n35240), .X(n24901) );
  nand_x1_sg U52018 ( .A(reg_www_2[7]), .B(n31924), .X(n24902) );
  nand_x1_sg U52019 ( .A(reg_ww_2[7]), .B(n30724), .X(n24903) );
  nand_x1_sg U52020 ( .A(reg_www_2[9]), .B(n32406), .X(n24906) );
  nand_x1_sg U52021 ( .A(reg_ww_2[9]), .B(n35404), .X(n24907) );
  nand_x1_sg U52022 ( .A(reg_www_2[10]), .B(n32495), .X(n24908) );
  nand_x1_sg U52023 ( .A(reg_ww_2[10]), .B(n30868), .X(n24909) );
  nand_x1_sg U52024 ( .A(reg_www_2[12]), .B(n32316), .X(n24912) );
  nand_x1_sg U52025 ( .A(reg_ww_2[12]), .B(n30897), .X(n24913) );
  nand_x1_sg U52026 ( .A(reg_www_3[9]), .B(n30914), .X(n24978) );
  nand_x1_sg U52027 ( .A(reg_ww_3[9]), .B(n35207), .X(n24979) );
  nand_x1_sg U52028 ( .A(reg_www_3[10]), .B(n32315), .X(n24980) );
  nand_x1_sg U52029 ( .A(reg_ww_3[10]), .B(n31096), .X(n24981) );
  nand_x1_sg U52030 ( .A(reg_www_3[12]), .B(n32357), .X(n24984) );
  nand_x1_sg U52031 ( .A(reg_ww_3[12]), .B(n35189), .X(n24985) );
  nand_x1_sg U52032 ( .A(reg_www_3[13]), .B(n32163), .X(n24986) );
  nand_x1_sg U52033 ( .A(reg_ww_3[13]), .B(n35224), .X(n24987) );
  nand_x1_sg U52034 ( .A(reg_www_3[15]), .B(n31892), .X(n24990) );
  nand_x1_sg U52035 ( .A(reg_ww_3[15]), .B(n32742), .X(n24991) );
  nand_x1_sg U52036 ( .A(reg_www_3[16]), .B(n31724), .X(n24992) );
  nand_x1_sg U52037 ( .A(reg_ww_3[16]), .B(n29767), .X(n24993) );
  nand_x1_sg U52038 ( .A(reg_www_3[18]), .B(n31497), .X(n24996) );
  nand_x1_sg U52039 ( .A(reg_ww_3[18]), .B(n31033), .X(n24997) );
  nand_x1_sg U52040 ( .A(reg_www_3[19]), .B(n31505), .X(n24998) );
  nand_x1_sg U52041 ( .A(reg_ww_3[19]), .B(n35225), .X(n24999) );
  nand_x1_sg U52042 ( .A(reg_www_4[12]), .B(n32019), .X(n24276) );
  nand_x1_sg U52043 ( .A(reg_ww_4[12]), .B(n35359), .X(n24277) );
  nand_x1_sg U52044 ( .A(reg_www_4[13]), .B(n33972), .X(n24278) );
  nand_x1_sg U52045 ( .A(reg_ww_4[13]), .B(n32711), .X(n24279) );
  nand_x1_sg U52046 ( .A(reg_www_4[15]), .B(n32374), .X(n24282) );
  nand_x1_sg U52047 ( .A(reg_ww_4[15]), .B(n30879), .X(n24283) );
  nand_x1_sg U52048 ( .A(reg_www_4[16]), .B(n32856), .X(n24284) );
  nand_x1_sg U52049 ( .A(reg_ww_4[16]), .B(n32738), .X(n24285) );
  nand_x1_sg U52050 ( .A(reg_www_4[18]), .B(n32364), .X(n24288) );
  nand_x1_sg U52051 ( .A(reg_ww_4[18]), .B(n30872), .X(n24289) );
  nand_x1_sg U52052 ( .A(reg_www_4[19]), .B(n32046), .X(n24290) );
  nand_x1_sg U52053 ( .A(reg_ww_4[19]), .B(n35371), .X(n24291) );
  nand_x1_sg U52054 ( .A(reg_www_5[0]), .B(n35080), .X(n24332) );
  nand_x1_sg U52055 ( .A(reg_ww_5[0]), .B(n35342), .X(n24333) );
  nand_x1_sg U52056 ( .A(reg_www_5[2]), .B(n32040), .X(n24336) );
  nand_x1_sg U52057 ( .A(reg_ww_5[2]), .B(n35377), .X(n24337) );
  nand_x1_sg U52058 ( .A(reg_www_6[1]), .B(n32332), .X(n24414) );
  nand_x1_sg U52059 ( .A(reg_ww_6[1]), .B(n35205), .X(n24415) );
  nand_x1_sg U52060 ( .A(reg_www_6[2]), .B(n32215), .X(n24416) );
  nand_x1_sg U52061 ( .A(reg_ww_6[2]), .B(n32762), .X(n24417) );
  nand_x1_sg U52062 ( .A(reg_www_6[4]), .B(n32323), .X(n24420) );
  nand_x1_sg U52063 ( .A(reg_ww_6[4]), .B(n35341), .X(n24421) );
  nand_x1_sg U52064 ( .A(reg_www_6[5]), .B(n34940), .X(n24422) );
  nand_x1_sg U52065 ( .A(reg_ww_6[5]), .B(n30591), .X(n24423) );
  nand_x1_sg U52066 ( .A(reg_www_6[7]), .B(n32361), .X(n24426) );
  nand_x1_sg U52067 ( .A(reg_ww_6[7]), .B(n32749), .X(n24427) );
  nand_x1_sg U52068 ( .A(reg_www_6[8]), .B(n30170), .X(n24428) );
  nand_x1_sg U52069 ( .A(reg_ww_6[8]), .B(n30870), .X(n24429) );
  nand_x1_sg U52070 ( .A(reg_www_6[10]), .B(n32141), .X(n24432) );
  nand_x1_sg U52071 ( .A(reg_ww_6[10]), .B(n35348), .X(n24433) );
  nand_x1_sg U52072 ( .A(reg_www_6[11]), .B(n34650), .X(n24434) );
  nand_x1_sg U52073 ( .A(reg_ww_6[11]), .B(n30861), .X(n24435) );
  nand_x1_sg U52074 ( .A(reg_www_6[13]), .B(n32300), .X(n24438) );
  nand_x1_sg U52075 ( .A(reg_ww_6[13]), .B(n32440), .X(n24439) );
  nand_x1_sg U52076 ( .A(reg_www_6[14]), .B(n32149), .X(n24440) );
  nand_x1_sg U52077 ( .A(reg_ww_6[14]), .B(n30171), .X(n24441) );
  nand_x1_sg U52078 ( .A(reg_www_6[16]), .B(n32227), .X(n24444) );
  nand_x1_sg U52079 ( .A(reg_ww_6[16]), .B(n34004), .X(n24445) );
  nand_x1_sg U52080 ( .A(reg_www_6[17]), .B(n32249), .X(n24446) );
  nand_x1_sg U52081 ( .A(reg_ww_6[17]), .B(n31035), .X(n24447) );
  nand_x1_sg U52082 ( .A(reg_www_6[19]), .B(n34849), .X(n24450) );
  nand_x1_sg U52083 ( .A(reg_ww_6[19]), .B(n32756), .X(n24451) );
  nand_x1_sg U52084 ( .A(reg_www_7[19]), .B(n31743), .X(n24530) );
  nand_x1_sg U52085 ( .A(reg_ww_7[19]), .B(n30878), .X(n24531) );
  nand_x1_sg U52086 ( .A(reg_www_8[1]), .B(n31924), .X(n24564) );
  nand_x1_sg U52087 ( .A(reg_ww_8[1]), .B(n35327), .X(n24565) );
  nand_x1_sg U52088 ( .A(reg_www_8[2]), .B(n31505), .X(n24566) );
  nand_x1_sg U52089 ( .A(reg_ww_8[2]), .B(n35362), .X(n24567) );
  nand_x1_sg U52090 ( .A(reg_www_8[4]), .B(n32498), .X(n24570) );
  nand_x1_sg U52091 ( .A(reg_ww_8[4]), .B(n34712), .X(n24571) );
  nand_x1_sg U52092 ( .A(reg_www_8[5]), .B(n32342), .X(n24572) );
  nand_x1_sg U52093 ( .A(reg_ww_8[5]), .B(n30717), .X(n24573) );
  nand_x1_sg U52094 ( .A(reg_www_8[7]), .B(n32364), .X(n24576) );
  nand_x1_sg U52095 ( .A(reg_ww_8[7]), .B(n30872), .X(n24577) );
  nand_x1_sg U52096 ( .A(reg_www_8[8]), .B(n32323), .X(n24578) );
  nand_x1_sg U52097 ( .A(reg_ww_8[8]), .B(n30726), .X(n24579) );
  nand_x1_sg U52098 ( .A(reg_www_8[10]), .B(n32032), .X(n24582) );
  nand_x1_sg U52099 ( .A(reg_ww_8[10]), .B(n32757), .X(n24583) );
  nand_x1_sg U52100 ( .A(reg_www_8[11]), .B(n32774), .X(n24584) );
  nand_x1_sg U52101 ( .A(reg_ww_8[11]), .B(n30717), .X(n24585) );
  nand_x1_sg U52102 ( .A(reg_www_8[13]), .B(n34847), .X(n24588) );
  nand_x1_sg U52103 ( .A(reg_ww_8[13]), .B(n31096), .X(n24589) );
  nand_x1_sg U52104 ( .A(reg_www_8[14]), .B(n31648), .X(n24590) );
  nand_x1_sg U52105 ( .A(reg_ww_8[14]), .B(n30726), .X(n24591) );
  nand_x1_sg U52106 ( .A(reg_www_9[0]), .B(n32252), .X(n23856) );
  nand_x1_sg U52107 ( .A(reg_ww_9[0]), .B(n30748), .X(n23857) );
  nand_x1_sg U52108 ( .A(reg_www_9[1]), .B(n32854), .X(n23858) );
  nand_x1_sg U52109 ( .A(reg_ww_9[1]), .B(n35341), .X(n23859) );
  nand_x1_sg U52110 ( .A(reg_www_9[3]), .B(n32333), .X(n23862) );
  nand_x1_sg U52111 ( .A(reg_ww_9[3]), .B(n30891), .X(n23863) );
  nand_x1_sg U52112 ( .A(reg_www_9[4]), .B(n32236), .X(n23864) );
  nand_x1_sg U52113 ( .A(reg_ww_9[4]), .B(n34708), .X(n23865) );
  nand_x1_sg U52114 ( .A(reg_www_9[6]), .B(n32044), .X(n23868) );
  nand_x1_sg U52115 ( .A(reg_ww_9[6]), .B(n32731), .X(n23869) );
  nand_x1_sg U52116 ( .A(reg_www_9[7]), .B(n32244), .X(n23870) );
  nand_x1_sg U52117 ( .A(reg_ww_9[7]), .B(n32748), .X(n23871) );
  nand_x1_sg U52118 ( .A(reg_www_9[9]), .B(n32400), .X(n23874) );
  nand_x1_sg U52119 ( .A(reg_ww_9[9]), .B(n31207), .X(n23875) );
  nand_x1_sg U52120 ( .A(reg_www_9[10]), .B(n32771), .X(n23876) );
  nand_x1_sg U52121 ( .A(reg_ww_9[10]), .B(n32442), .X(n23877) );
  nand_x1_sg U52122 ( .A(reg_www_9[12]), .B(n32775), .X(n23880) );
  nand_x1_sg U52123 ( .A(reg_ww_9[12]), .B(n35197), .X(n23881) );
  nand_x1_sg U52124 ( .A(reg_www_9[13]), .B(n31906), .X(n23882) );
  nand_x1_sg U52125 ( .A(reg_ww_9[13]), .B(n30865), .X(n23883) );
  nand_x1_sg U52126 ( .A(reg_www_9[15]), .B(n32385), .X(n23886) );
  nand_x1_sg U52127 ( .A(reg_ww_9[15]), .B(n34095), .X(n23887) );
  nand_x1_sg U52128 ( .A(reg_www_9[16]), .B(n32325), .X(n23888) );
  nand_x1_sg U52129 ( .A(reg_ww_9[16]), .B(n30897), .X(n23889) );
  nand_x1_sg U52130 ( .A(reg_www_10[9]), .B(n31901), .X(n23954) );
  nand_x1_sg U52131 ( .A(reg_ww_10[9]), .B(n30174), .X(n23955) );
  nand_x1_sg U52132 ( .A(reg_www_10[11]), .B(n32340), .X(n23958) );
  nand_x1_sg U52133 ( .A(reg_ww_10[11]), .B(n32840), .X(n23959) );
  nand_x1_sg U52134 ( .A(reg_www_10[12]), .B(n32146), .X(n23960) );
  nand_x1_sg U52135 ( .A(reg_ww_10[12]), .B(n35160), .X(n23961) );
  nand_x1_sg U52136 ( .A(reg_www_10[14]), .B(n34895), .X(n23964) );
  nand_x1_sg U52137 ( .A(reg_ww_10[14]), .B(n32733), .X(n23965) );
  nand_x1_sg U52138 ( .A(reg_www_10[15]), .B(n32215), .X(n23966) );
  nand_x1_sg U52139 ( .A(reg_ww_10[15]), .B(n30887), .X(n23967) );
  nand_x1_sg U52140 ( .A(reg_www_10[17]), .B(n31733), .X(n23970) );
  nand_x1_sg U52141 ( .A(reg_ww_10[17]), .B(n30879), .X(n23971) );
  nand_x1_sg U52142 ( .A(reg_www_10[18]), .B(n31646), .X(n23972) );
  nand_x1_sg U52143 ( .A(reg_ww_10[18]), .B(n30709), .X(n23973) );
  nand_x1_sg U52144 ( .A(reg_www_14[7]), .B(n32246), .X(n23700) );
  nand_x1_sg U52145 ( .A(reg_ww_14[7]), .B(n32709), .X(n23701) );
  nand_x1_sg U52146 ( .A(reg_www_14[8]), .B(n34572), .X(n23702) );
  nand_x1_sg U52147 ( .A(reg_ww_14[8]), .B(n35359), .X(n23703) );
  nand_x1_sg U52148 ( .A(reg_www_14[10]), .B(n31905), .X(n23706) );
  nand_x1_sg U52149 ( .A(reg_ww_14[10]), .B(n34668), .X(n23707) );
  nand_x1_sg U52150 ( .A(reg_www_14[11]), .B(n31739), .X(n23708) );
  nand_x1_sg U52151 ( .A(reg_ww_14[11]), .B(n35380), .X(n23709) );
  nand_x1_sg U52152 ( .A(reg_www_14[13]), .B(n32164), .X(n23712) );
  nand_x1_sg U52153 ( .A(reg_ww_14[13]), .B(n31092), .X(n23713) );
  nand_x1_sg U52154 ( .A(reg_www_14[14]), .B(n32165), .X(n23714) );
  nand_x1_sg U52155 ( .A(reg_ww_14[14]), .B(n35398), .X(n23715) );
  nand_x1_sg U52156 ( .A(reg_www_14[16]), .B(n31908), .X(n23718) );
  nand_x1_sg U52157 ( .A(reg_ww_14[16]), .B(n35094), .X(n23719) );
  nand_x1_sg U52158 ( .A(reg_www_14[17]), .B(n32374), .X(n23720) );
  nand_x1_sg U52159 ( .A(reg_ww_14[17]), .B(n35329), .X(n23721) );
  nand_x1_sg U52160 ( .A(reg_www_14[19]), .B(n34697), .X(n23724) );
  nand_x1_sg U52161 ( .A(reg_ww_14[19]), .B(n35345), .X(n23725) );
  nand_x1_sg U52162 ( .A(reg_iii_2[3]), .B(n33967), .X(n26002) );
  nand_x1_sg U52163 ( .A(reg_ii_2[3]), .B(n35085), .X(n26003) );
  nand_x1_sg U52164 ( .A(reg_iii_2[6]), .B(n31908), .X(n26008) );
  nand_x1_sg U52165 ( .A(reg_ii_2[6]), .B(n32733), .X(n26009) );
  nand_x1_sg U52166 ( .A(reg_iii_2[9]), .B(n31712), .X(n26014) );
  nand_x1_sg U52167 ( .A(reg_ii_2[9]), .B(n32835), .X(n26015) );
  nand_x1_sg U52168 ( .A(reg_iii_2[12]), .B(n33943), .X(n26020) );
  nand_x1_sg U52169 ( .A(reg_ii_2[12]), .B(n32740), .X(n26021) );
  nand_x1_sg U52170 ( .A(reg_iii_2[15]), .B(n32036), .X(n26026) );
  nand_x1_sg U52171 ( .A(reg_ii_2[15]), .B(n32832), .X(n26027) );
  nand_x1_sg U52172 ( .A(reg_iii_2[18]), .B(n31633), .X(n26032) );
  nand_x1_sg U52173 ( .A(reg_ii_2[18]), .B(n30897), .X(n26033) );
  nand_x1_sg U52174 ( .A(reg_iii_4[2]), .B(n32373), .X(n26158) );
  nand_x1_sg U52175 ( .A(reg_ii_4[2]), .B(n32767), .X(n26159) );
  nand_x1_sg U52176 ( .A(reg_iii_4[5]), .B(n32247), .X(n26164) );
  nand_x1_sg U52177 ( .A(reg_ii_4[5]), .B(n32744), .X(n26165) );
  nand_x1_sg U52178 ( .A(reg_iii_4[8]), .B(n31727), .X(n26170) );
  nand_x1_sg U52179 ( .A(reg_ii_4[8]), .B(n30895), .X(n26171) );
  nand_x1_sg U52180 ( .A(reg_iii_4[11]), .B(n32034), .X(n26176) );
  nand_x1_sg U52181 ( .A(reg_ii_4[11]), .B(n30713), .X(n26177) );
  nand_x1_sg U52182 ( .A(reg_iii_4[14]), .B(n32310), .X(n26182) );
  nand_x1_sg U52183 ( .A(reg_ii_4[14]), .B(n32721), .X(n26183) );
  nand_x1_sg U52184 ( .A(reg_iii_4[17]), .B(n32340), .X(n26188) );
  nand_x1_sg U52185 ( .A(reg_ii_4[17]), .B(n30902), .X(n26189) );
  nand_x1_sg U52186 ( .A(reg_iii_5[2]), .B(n32356), .X(n25444) );
  nand_x1_sg U52187 ( .A(reg_ii_5[2]), .B(n32711), .X(n25445) );
  nand_x1_sg U52188 ( .A(reg_iii_5[5]), .B(n32455), .X(n25450) );
  nand_x1_sg U52189 ( .A(reg_ii_5[5]), .B(n32750), .X(n25451) );
  nand_x1_sg U52190 ( .A(reg_iii_5[8]), .B(n32429), .X(n25456) );
  nand_x1_sg U52191 ( .A(reg_ii_5[8]), .B(n35228), .X(n25457) );
  nand_x1_sg U52192 ( .A(reg_iii_5[11]), .B(n31901), .X(n25462) );
  nand_x1_sg U52193 ( .A(reg_ii_5[11]), .B(n30884), .X(n25463) );
  nand_x1_sg U52194 ( .A(reg_iii_5[14]), .B(n31497), .X(n25468) );
  nand_x1_sg U52195 ( .A(reg_ii_5[14]), .B(n35094), .X(n25469) );
  nand_x1_sg U52196 ( .A(reg_iii_5[17]), .B(n31906), .X(n25474) );
  nand_x1_sg U52197 ( .A(reg_ii_5[17]), .B(n32737), .X(n25475) );
  nand_x1_sg U52198 ( .A(reg_iii_6[19]), .B(n31711), .X(n25558) );
  nand_x1_sg U52199 ( .A(reg_ii_6[19]), .B(n31490), .X(n25559) );
  nand_x1_sg U52200 ( .A(reg_iii_7[0]), .B(n32042), .X(n25600) );
  nand_x1_sg U52201 ( .A(reg_ii_7[0]), .B(n30864), .X(n25601) );
  nand_x1_sg U52202 ( .A(reg_iii_7[3]), .B(n32344), .X(n25606) );
  nand_x1_sg U52203 ( .A(reg_ii_7[3]), .B(n34005), .X(n25607) );
  nand_x1_sg U52204 ( .A(reg_iii_7[6]), .B(n32151), .X(n25612) );
  nand_x1_sg U52205 ( .A(reg_ii_7[6]), .B(n32745), .X(n25613) );
  nand_x1_sg U52206 ( .A(reg_iii_8[2]), .B(n32031), .X(n25684) );
  nand_x1_sg U52207 ( .A(reg_ii_8[2]), .B(n31027), .X(n25685) );
  nand_x1_sg U52208 ( .A(reg_iii_8[5]), .B(n32775), .X(n25690) );
  nand_x1_sg U52209 ( .A(reg_ii_8[5]), .B(n32752), .X(n25691) );
  nand_x1_sg U52210 ( .A(reg_iii_8[8]), .B(n32379), .X(n25696) );
  nand_x1_sg U52211 ( .A(reg_ii_8[8]), .B(n34713), .X(n25697) );
  nand_x1_sg U52212 ( .A(reg_iii_8[11]), .B(n32428), .X(n25702) );
  nand_x1_sg U52213 ( .A(reg_ii_8[11]), .B(n32760), .X(n25703) );
  nand_x1_sg U52214 ( .A(reg_iii_8[14]), .B(n31909), .X(n25708) );
  nand_x1_sg U52215 ( .A(reg_ii_8[14]), .B(n35083), .X(n25709) );
  nand_x1_sg U52216 ( .A(reg_iii_8[17]), .B(n31513), .X(n25714) );
  nand_x1_sg U52217 ( .A(reg_ii_8[17]), .B(n31025), .X(n25715) );
  nand_x1_sg U52218 ( .A(reg_iii_11[1]), .B(n31725), .X(n25126) );
  nand_x1_sg U52219 ( .A(reg_ii_11[1]), .B(n35339), .X(n25127) );
  nand_x1_sg U52220 ( .A(reg_iii_11[4]), .B(n34698), .X(n25132) );
  nand_x1_sg U52221 ( .A(reg_ii_11[4]), .B(n30863), .X(n25133) );
  nand_x1_sg U52222 ( .A(reg_iii_11[7]), .B(n32283), .X(n25138) );
  nand_x1_sg U52223 ( .A(reg_ii_11[7]), .B(n30867), .X(n25139) );
  nand_x1_sg U52224 ( .A(reg_iii_11[10]), .B(n32281), .X(n25144) );
  nand_x1_sg U52225 ( .A(reg_ii_11[10]), .B(n34042), .X(n25145) );
  nand_x1_sg U52226 ( .A(reg_iii_11[13]), .B(n32038), .X(n25150) );
  nand_x1_sg U52227 ( .A(reg_ii_11[13]), .B(n30709), .X(n25151) );
  nand_x1_sg U52228 ( .A(reg_iii_11[16]), .B(n30611), .X(n25156) );
  nand_x1_sg U52229 ( .A(reg_ii_11[16]), .B(n32760), .X(n25157) );
  nand_x1_sg U52230 ( .A(reg_iii_11[19]), .B(n33942), .X(n25162) );
  nand_x1_sg U52231 ( .A(reg_ii_11[19]), .B(n35326), .X(n25163) );
  nand_x1_sg U52232 ( .A(reg_www_2[2]), .B(n31737), .X(n24892) );
  nand_x1_sg U52233 ( .A(reg_ww_2[2]), .B(n35356), .X(n24893) );
  nand_x1_sg U52234 ( .A(reg_www_2[5]), .B(n33951), .X(n24898) );
  nand_x1_sg U52235 ( .A(reg_ww_2[5]), .B(n32732), .X(n24899) );
  nand_x1_sg U52236 ( .A(reg_www_2[8]), .B(n33953), .X(n24904) );
  nand_x1_sg U52237 ( .A(reg_ww_2[8]), .B(n32728), .X(n24905) );
  nand_x1_sg U52238 ( .A(reg_www_2[11]), .B(n32857), .X(n24910) );
  nand_x1_sg U52239 ( .A(reg_ww_2[11]), .B(n30892), .X(n24911) );
  nand_x1_sg U52240 ( .A(reg_www_3[11]), .B(n34570), .X(n24982) );
  nand_x1_sg U52241 ( .A(reg_ww_3[11]), .B(n32728), .X(n24983) );
  nand_x1_sg U52242 ( .A(reg_www_3[14]), .B(n33968), .X(n24988) );
  nand_x1_sg U52243 ( .A(reg_ww_3[14]), .B(n35187), .X(n24989) );
  nand_x1_sg U52244 ( .A(reg_www_3[17]), .B(n32242), .X(n24994) );
  nand_x1_sg U52245 ( .A(reg_ww_3[17]), .B(n35329), .X(n24995) );
  nand_x1_sg U52246 ( .A(reg_www_4[11]), .B(n31898), .X(n24274) );
  nand_x1_sg U52247 ( .A(reg_ww_4[11]), .B(n30863), .X(n24275) );
  nand_x1_sg U52248 ( .A(reg_www_4[14]), .B(n34582), .X(n24280) );
  nand_x1_sg U52249 ( .A(reg_ww_4[14]), .B(n30891), .X(n24281) );
  nand_x1_sg U52250 ( .A(reg_www_4[17]), .B(n32035), .X(n24286) );
  nand_x1_sg U52251 ( .A(reg_ww_4[17]), .B(n35339), .X(n24287) );
  nand_x1_sg U52252 ( .A(reg_www_5[1]), .B(n32042), .X(n24334) );
  nand_x1_sg U52253 ( .A(reg_ww_5[1]), .B(n32837), .X(n24335) );
  nand_x1_sg U52254 ( .A(reg_www_6[0]), .B(n32772), .X(n24412) );
  nand_x1_sg U52255 ( .A(reg_ww_6[0]), .B(n30172), .X(n24413) );
  nand_x1_sg U52256 ( .A(reg_www_6[3]), .B(n32333), .X(n24418) );
  nand_x1_sg U52257 ( .A(reg_ww_6[3]), .B(n31027), .X(n24419) );
  nand_x1_sg U52258 ( .A(reg_www_6[6]), .B(n31900), .X(n24424) );
  nand_x1_sg U52259 ( .A(reg_ww_6[6]), .B(n35182), .X(n24425) );
  nand_x1_sg U52260 ( .A(reg_www_6[9]), .B(n32376), .X(n24430) );
  nand_x1_sg U52261 ( .A(reg_ww_6[9]), .B(n35171), .X(n24431) );
  nand_x1_sg U52262 ( .A(reg_www_6[12]), .B(n32327), .X(n24436) );
  nand_x1_sg U52263 ( .A(reg_ww_6[12]), .B(n35335), .X(n24437) );
  nand_x1_sg U52264 ( .A(reg_www_6[15]), .B(n34850), .X(n24442) );
  nand_x1_sg U52265 ( .A(reg_ww_6[15]), .B(n31039), .X(n24443) );
  nand_x1_sg U52266 ( .A(reg_www_6[18]), .B(n32354), .X(n24448) );
  nand_x1_sg U52267 ( .A(reg_ww_6[18]), .B(n35320), .X(n24449) );
  nand_x1_sg U52268 ( .A(reg_www_8[0]), .B(n32406), .X(n24562) );
  nand_x1_sg U52269 ( .A(reg_ww_8[0]), .B(n32724), .X(n24563) );
  nand_x1_sg U52270 ( .A(reg_www_8[3]), .B(n32777), .X(n24568) );
  nand_x1_sg U52271 ( .A(reg_ww_8[3]), .B(n32736), .X(n24569) );
  nand_x1_sg U52272 ( .A(reg_www_8[6]), .B(n31925), .X(n24574) );
  nand_x1_sg U52273 ( .A(reg_ww_8[6]), .B(n32761), .X(n24575) );
  nand_x1_sg U52274 ( .A(reg_www_8[9]), .B(n32451), .X(n24580) );
  nand_x1_sg U52275 ( .A(reg_ww_8[9]), .B(n32730), .X(n24581) );
  nand_x1_sg U52276 ( .A(reg_www_8[12]), .B(n32035), .X(n24586) );
  nand_x1_sg U52277 ( .A(reg_ww_8[12]), .B(n32726), .X(n24587) );
  nand_x1_sg U52278 ( .A(reg_www_8[15]), .B(n32280), .X(n24592) );
  nand_x1_sg U52279 ( .A(reg_ww_8[15]), .B(n30713), .X(n24593) );
  nand_x1_sg U52280 ( .A(reg_www_9[2]), .B(n31637), .X(n23860) );
  nand_x1_sg U52281 ( .A(reg_ww_9[2]), .B(n30899), .X(n23861) );
  nand_x1_sg U52282 ( .A(reg_www_9[5]), .B(n31896), .X(n23866) );
  nand_x1_sg U52283 ( .A(reg_ww_9[5]), .B(n30889), .X(n23867) );
  nand_x1_sg U52284 ( .A(reg_www_9[8]), .B(n32030), .X(n23872) );
  nand_x1_sg U52285 ( .A(reg_ww_9[8]), .B(n32738), .X(n23873) );
  nand_x1_sg U52286 ( .A(reg_www_9[11]), .B(n31904), .X(n23878) );
  nand_x1_sg U52287 ( .A(reg_ww_9[11]), .B(n31056), .X(n23879) );
  nand_x1_sg U52288 ( .A(reg_www_9[14]), .B(n32290), .X(n23884) );
  nand_x1_sg U52289 ( .A(reg_ww_9[14]), .B(n32754), .X(n23885) );
  nand_x1_sg U52290 ( .A(reg_www_10[10]), .B(n35077), .X(n23956) );
  nand_x1_sg U52291 ( .A(reg_ww_10[10]), .B(n35193), .X(n23957) );
  nand_x1_sg U52292 ( .A(reg_www_10[13]), .B(n32429), .X(n23962) );
  nand_x1_sg U52293 ( .A(reg_ww_10[13]), .B(n30724), .X(n23963) );
  nand_x1_sg U52294 ( .A(reg_www_10[16]), .B(n32325), .X(n23968) );
  nand_x1_sg U52295 ( .A(reg_ww_10[16]), .B(n34042), .X(n23969) );
  nand_x1_sg U52296 ( .A(reg_www_10[19]), .B(n32345), .X(n23974) );
  nand_x1_sg U52297 ( .A(reg_ww_10[19]), .B(n30594), .X(n23975) );
  nand_x1_sg U52298 ( .A(reg_www_11[0]), .B(n32366), .X(n24016) );
  nand_x1_sg U52299 ( .A(reg_ww_11[0]), .B(n30881), .X(n24017) );
  nand_x1_sg U52300 ( .A(reg_www_14[6]), .B(n29756), .X(n23698) );
  nand_x1_sg U52301 ( .A(reg_ww_14[6]), .B(n35351), .X(n23699) );
  nand_x1_sg U52302 ( .A(reg_www_14[9]), .B(n32349), .X(n23704) );
  nand_x1_sg U52303 ( .A(reg_ww_14[9]), .B(n34043), .X(n23705) );
  nand_x1_sg U52304 ( .A(reg_www_14[12]), .B(n30599), .X(n23710) );
  nand_x1_sg U52305 ( .A(reg_ww_14[12]), .B(n31206), .X(n23711) );
  nand_x1_sg U52306 ( .A(reg_www_14[15]), .B(n31642), .X(n23716) );
  nand_x1_sg U52307 ( .A(reg_ww_14[15]), .B(n32735), .X(n23717) );
  nand_x1_sg U52308 ( .A(reg_www_14[18]), .B(n31501), .X(n23722) );
  nand_x1_sg U52309 ( .A(reg_ww_14[18]), .B(n31035), .X(n23723) );
  nand_x1_sg U52310 ( .A(reg_ii_3[0]), .B(n32338), .X(n26036) );
  nand_x1_sg U52311 ( .A(n34718), .B(reg_i_3[0]), .X(n26037) );
  nand_x1_sg U52312 ( .A(reg_ii_3[2]), .B(n32215), .X(n26040) );
  nand_x1_sg U52313 ( .A(n32726), .B(reg_i_3[2]), .X(n26041) );
  nand_x1_sg U52314 ( .A(reg_ii_3[3]), .B(n33945), .X(n26042) );
  nand_x1_sg U52315 ( .A(n32755), .B(reg_i_3[3]), .X(n26043) );
  nand_x1_sg U52316 ( .A(reg_ii_3[5]), .B(n34577), .X(n26046) );
  nand_x1_sg U52317 ( .A(n35193), .B(reg_i_3[5]), .X(n26047) );
  nand_x1_sg U52318 ( .A(reg_ii_3[6]), .B(n32295), .X(n26048) );
  nand_x1_sg U52319 ( .A(n35221), .B(reg_i_3[6]), .X(n26049) );
  nand_x1_sg U52320 ( .A(reg_ii_3[8]), .B(n34567), .X(n26052) );
  nand_x1_sg U52321 ( .A(n35332), .B(reg_i_3[8]), .X(n26053) );
  nand_x1_sg U52322 ( .A(reg_ii_3[9]), .B(n31640), .X(n26054) );
  nand_x1_sg U52323 ( .A(n35199), .B(reg_i_3[9]), .X(n26055) );
  nand_x1_sg U52324 ( .A(reg_ii_3[11]), .B(n30170), .X(n26058) );
  nand_x1_sg U52325 ( .A(n34073), .B(reg_i_3[11]), .X(n26059) );
  nand_x1_sg U52326 ( .A(reg_ii_3[12]), .B(n32498), .X(n26060) );
  nand_x1_sg U52327 ( .A(n35164), .B(reg_i_3[12]), .X(n26061) );
  nand_x1_sg U52328 ( .A(reg_ii_3[14]), .B(n32216), .X(n26064) );
  nand_x1_sg U52329 ( .A(n34077), .B(reg_i_3[14]), .X(n26065) );
  nand_x1_sg U52330 ( .A(reg_ii_4[7]), .B(n32026), .X(n26130) );
  nand_x1_sg U52331 ( .A(n34724), .B(reg_i_4[7]), .X(n26131) );
  nand_x1_sg U52332 ( .A(reg_ii_4[8]), .B(n32243), .X(n26132) );
  nand_x1_sg U52333 ( .A(n35358), .B(reg_i_4[8]), .X(n26133) );
  nand_x1_sg U52334 ( .A(reg_ii_4[10]), .B(n32020), .X(n26136) );
  nand_x1_sg U52335 ( .A(n32846), .B(reg_i_4[10]), .X(n26137) );
  nand_x1_sg U52336 ( .A(reg_ii_4[11]), .B(n32287), .X(n26138) );
  nand_x1_sg U52337 ( .A(n35377), .B(reg_i_4[11]), .X(n26139) );
  nand_x1_sg U52338 ( .A(reg_ii_4[13]), .B(n32214), .X(n26142) );
  nand_x1_sg U52339 ( .A(n34095), .B(reg_i_4[13]), .X(n26143) );
  nand_x1_sg U52340 ( .A(reg_ii_4[14]), .B(n32048), .X(n26144) );
  nand_x1_sg U52341 ( .A(n35181), .B(reg_i_4[14]), .X(n26145) );
  nand_x1_sg U52342 ( .A(reg_ii_4[16]), .B(n32407), .X(n26148) );
  nand_x1_sg U52343 ( .A(n32750), .B(reg_i_4[16]), .X(n26149) );
  nand_x1_sg U52344 ( .A(reg_ii_4[17]), .B(n32312), .X(n26150) );
  nand_x1_sg U52345 ( .A(n32732), .B(reg_i_4[17]), .X(n26151) );
  nand_x1_sg U52346 ( .A(reg_ii_5[14]), .B(n32300), .X(n25428) );
  nand_x1_sg U52347 ( .A(n35321), .B(reg_i_5[14]), .X(n25429) );
  nand_x1_sg U52348 ( .A(reg_ii_5[15]), .B(n31505), .X(n25430) );
  nand_x1_sg U52349 ( .A(n35345), .B(reg_i_5[15]), .X(n25431) );
  nand_x1_sg U52350 ( .A(reg_ii_5[17]), .B(n32400), .X(n25434) );
  nand_x1_sg U52351 ( .A(n32831), .B(reg_i_5[17]), .X(n25435) );
  nand_x1_sg U52352 ( .A(reg_ii_5[18]), .B(n32214), .X(n25436) );
  nand_x1_sg U52353 ( .A(n35225), .B(reg_i_5[18]), .X(n25437) );
  nand_x1_sg U52354 ( .A(reg_ii_6[1]), .B(n32026), .X(n25482) );
  nand_x1_sg U52355 ( .A(n35189), .B(reg_i_6[1]), .X(n25483) );
  nand_x1_sg U52356 ( .A(reg_ii_6[2]), .B(n31889), .X(n25484) );
  nand_x1_sg U52357 ( .A(n31873), .B(reg_i_6[2]), .X(n25485) );
  nand_x1_sg U52358 ( .A(reg_ii_6[4]), .B(n31729), .X(n25488) );
  nand_x1_sg U52359 ( .A(n30179), .B(reg_i_6[4]), .X(n25489) );
  nand_x1_sg U52360 ( .A(reg_ii_7[0]), .B(n31743), .X(n25560) );
  nand_x1_sg U52361 ( .A(n30906), .B(reg_i_7[0]), .X(n25561) );
  nand_x1_sg U52362 ( .A(reg_ii_7[1]), .B(n35079), .X(n25562) );
  nand_x1_sg U52363 ( .A(n35231), .B(reg_i_7[1]), .X(n25563) );
  nand_x1_sg U52364 ( .A(reg_ii_7[3]), .B(n32041), .X(n25566) );
  nand_x1_sg U52365 ( .A(n32841), .B(reg_i_7[3]), .X(n25567) );
  nand_x1_sg U52366 ( .A(reg_ii_7[4]), .B(n32012), .X(n25568) );
  nand_x1_sg U52367 ( .A(n32836), .B(reg_i_7[4]), .X(n25569) );
  nand_x1_sg U52368 ( .A(reg_ii_7[6]), .B(n32456), .X(n25572) );
  nand_x1_sg U52369 ( .A(n35093), .B(reg_i_7[6]), .X(n25573) );
  nand_x1_sg U52370 ( .A(reg_ii_7[7]), .B(n32855), .X(n25574) );
  nand_x1_sg U52371 ( .A(n32711), .B(reg_i_7[7]), .X(n25575) );
  nand_x1_sg U52372 ( .A(reg_ii_7[9]), .B(n32321), .X(n25578) );
  nand_x1_sg U52373 ( .A(n35092), .B(reg_i_7[9]), .X(n25579) );
  nand_x1_sg U52374 ( .A(reg_ii_7[10]), .B(n32772), .X(n25580) );
  nand_x1_sg U52375 ( .A(n31672), .B(reg_i_7[10]), .X(n25581) );
  nand_x1_sg U52376 ( .A(reg_ii_7[12]), .B(n31729), .X(n25584) );
  nand_x1_sg U52377 ( .A(n35232), .B(reg_i_7[12]), .X(n25585) );
  nand_x1_sg U52378 ( .A(reg_ii_7[13]), .B(n32156), .X(n25586) );
  nand_x1_sg U52379 ( .A(n32442), .B(reg_i_7[13]), .X(n25587) );
  nand_x1_sg U52380 ( .A(reg_ii_7[15]), .B(n32234), .X(n25590) );
  nand_x1_sg U52381 ( .A(n32835), .B(reg_i_7[15]), .X(n25591) );
  nand_x1_sg U52382 ( .A(reg_ii_7[16]), .B(n32777), .X(n25592) );
  nand_x1_sg U52383 ( .A(n34096), .B(reg_i_7[16]), .X(n25593) );
  nand_x1_sg U52384 ( .A(reg_ii_7[18]), .B(n33946), .X(n25596) );
  nand_x1_sg U52385 ( .A(n34702), .B(reg_i_7[18]), .X(n25597) );
  nand_x1_sg U52386 ( .A(reg_ii_7[19]), .B(n32315), .X(n25598) );
  nand_x1_sg U52387 ( .A(n34091), .B(reg_i_7[19]), .X(n25599) );
  nand_x1_sg U52388 ( .A(reg_ii_9[1]), .B(n35277), .X(n25722) );
  nand_x1_sg U52389 ( .A(n31675), .B(reg_i_9[1]), .X(n25723) );
  nand_x1_sg U52390 ( .A(reg_ii_9[2]), .B(n31896), .X(n25724) );
  nand_x1_sg U52391 ( .A(n34077), .B(reg_i_9[2]), .X(n25725) );
  nand_x1_sg U52392 ( .A(reg_ii_9[4]), .B(n32322), .X(n25728) );
  nand_x1_sg U52393 ( .A(n32723), .B(reg_i_9[4]), .X(n25729) );
  nand_x1_sg U52394 ( .A(reg_ii_9[5]), .B(n34896), .X(n25730) );
  nand_x1_sg U52395 ( .A(n32717), .B(reg_i_9[5]), .X(n25731) );
  nand_x1_sg U52396 ( .A(reg_ii_9[7]), .B(n32401), .X(n25734) );
  nand_x1_sg U52397 ( .A(n34053), .B(reg_i_9[7]), .X(n25735) );
  nand_x1_sg U52398 ( .A(reg_ii_9[8]), .B(n32349), .X(n25736) );
  nand_x1_sg U52399 ( .A(n32847), .B(reg_i_9[8]), .X(n25737) );
  nand_x1_sg U52400 ( .A(reg_ii_9[10]), .B(n32160), .X(n25740) );
  nand_x1_sg U52401 ( .A(n35371), .B(reg_i_9[10]), .X(n25741) );
  nand_x1_sg U52402 ( .A(reg_ii_9[11]), .B(n31630), .X(n25742) );
  nand_x1_sg U52403 ( .A(n35206), .B(reg_i_9[11]), .X(n25743) );
  nand_x1_sg U52404 ( .A(reg_ii_9[19]), .B(n32493), .X(n25002) );
  nand_x1_sg U52405 ( .A(n35350), .B(reg_i_9[19]), .X(n25003) );
  nand_x1_sg U52406 ( .A(reg_ii_10[0]), .B(n32326), .X(n25004) );
  nand_x1_sg U52407 ( .A(n31671), .B(reg_i_10[0]), .X(n25005) );
  nand_x1_sg U52408 ( .A(reg_ii_10[2]), .B(n30599), .X(n25008) );
  nand_x1_sg U52409 ( .A(n34056), .B(reg_i_10[2]), .X(n25009) );
  nand_x1_sg U52410 ( .A(reg_ii_10[3]), .B(n32282), .X(n25010) );
  nand_x1_sg U52411 ( .A(n32840), .B(reg_i_10[3]), .X(n25011) );
  nand_x1_sg U52412 ( .A(reg_ii_10[5]), .B(n30623), .X(n25014) );
  nand_x1_sg U52413 ( .A(n35351), .B(reg_i_10[5]), .X(n25015) );
  nand_x1_sg U52414 ( .A(reg_ii_10[6]), .B(n30596), .X(n25016) );
  nand_x1_sg U52415 ( .A(n35209), .B(reg_i_10[6]), .X(n25017) );
  nand_x1_sg U52416 ( .A(reg_ii_10[8]), .B(n32138), .X(n25020) );
  nand_x1_sg U52417 ( .A(n35398), .B(reg_i_10[8]), .X(n25021) );
  nand_x1_sg U52418 ( .A(reg_ii_10[9]), .B(n32292), .X(n25022) );
  nand_x1_sg U52419 ( .A(n34047), .B(reg_i_10[9]), .X(n25023) );
  nand_x1_sg U52420 ( .A(reg_ii_10[11]), .B(n32318), .X(n25026) );
  nand_x1_sg U52421 ( .A(n34721), .B(reg_i_10[11]), .X(n25027) );
  nand_x1_sg U52422 ( .A(reg_ii_10[12]), .B(n30149), .X(n25028) );
  nand_x1_sg U52423 ( .A(n34050), .B(reg_i_10[12]), .X(n25029) );
  nand_x1_sg U52424 ( .A(reg_ii_10[14]), .B(n32315), .X(n25032) );
  nand_x1_sg U52425 ( .A(n35367), .B(reg_i_10[14]), .X(n25033) );
  nand_x1_sg U52426 ( .A(reg_ii_10[15]), .B(n31896), .X(n25034) );
  nand_x1_sg U52427 ( .A(n33996), .B(reg_i_10[15]), .X(n25035) );
  nand_x1_sg U52428 ( .A(reg_ii_10[17]), .B(n33953), .X(n25038) );
  nand_x1_sg U52429 ( .A(n32832), .B(reg_i_10[17]), .X(n25039) );
  nand_x1_sg U52430 ( .A(reg_ii_10[18]), .B(n32045), .X(n25040) );
  nand_x1_sg U52431 ( .A(n31865), .B(reg_i_10[18]), .X(n25041) );
  nand_x1_sg U52432 ( .A(reg_ii_11[11]), .B(n32280), .X(n25106) );
  nand_x1_sg U52433 ( .A(n31868), .B(reg_i_11[11]), .X(n25107) );
  nand_x1_sg U52434 ( .A(reg_ii_11[13]), .B(n32330), .X(n25110) );
  nand_x1_sg U52435 ( .A(n35233), .B(reg_i_11[13]), .X(n25111) );
  nand_x1_sg U52436 ( .A(reg_ii_11[14]), .B(n34652), .X(n25112) );
  nand_x1_sg U52437 ( .A(n30593), .B(reg_i_11[14]), .X(n25113) );
  nand_x1_sg U52438 ( .A(reg_ii_11[16]), .B(n32232), .X(n25116) );
  nand_x1_sg U52439 ( .A(n30593), .B(reg_i_11[16]), .X(n25117) );
  nand_x1_sg U52440 ( .A(reg_ii_11[17]), .B(n32400), .X(n25118) );
  nand_x1_sg U52441 ( .A(n34076), .B(reg_i_11[17]), .X(n25119) );
  nand_x1_sg U52442 ( .A(reg_ii_11[19]), .B(n31646), .X(n25122) );
  nand_x1_sg U52443 ( .A(n35084), .B(reg_i_11[19]), .X(n25123) );
  nand_x1_sg U52444 ( .A(reg_ii_12[0]), .B(n32493), .X(n25164) );
  nand_x1_sg U52445 ( .A(n32726), .B(reg_i_12[0]), .X(n25165) );
  nand_x1_sg U52446 ( .A(reg_ii_12[1]), .B(n34846), .X(n25166) );
  nand_x1_sg U52447 ( .A(n35362), .B(reg_i_12[1]), .X(n25167) );
  nand_x1_sg U52448 ( .A(reg_ww_2[2]), .B(n34851), .X(n24852) );
  nand_x1_sg U52449 ( .A(n35205), .B(reg_w_2[2]), .X(n24853) );
  nand_x1_sg U52450 ( .A(reg_ww_2[3]), .B(n30145), .X(n24854) );
  nand_x1_sg U52451 ( .A(n34668), .B(reg_w_2[3]), .X(n24855) );
  nand_x1_sg U52452 ( .A(reg_ww_2[5]), .B(n31892), .X(n24858) );
  nand_x1_sg U52453 ( .A(n34094), .B(reg_w_2[5]), .X(n24859) );
  nand_x1_sg U52454 ( .A(reg_ww_2[6]), .B(n32381), .X(n24860) );
  nand_x1_sg U52455 ( .A(n32766), .B(reg_w_2[6]), .X(n24861) );
  nand_x1_sg U52456 ( .A(reg_ww_2[8]), .B(n33972), .X(n24864) );
  nand_x1_sg U52457 ( .A(n34072), .B(reg_w_2[8]), .X(n24865) );
  nand_x1_sg U52458 ( .A(reg_ww_2[9]), .B(n32248), .X(n24866) );
  nand_x1_sg U52459 ( .A(n34713), .B(reg_w_2[9]), .X(n24867) );
  nand_x1_sg U52460 ( .A(reg_ww_2[11]), .B(n32145), .X(n24870) );
  nand_x1_sg U52461 ( .A(n32713), .B(reg_w_2[11]), .X(n24871) );
  nand_x1_sg U52462 ( .A(reg_ww_2[12]), .B(n31889), .X(n24872) );
  nand_x1_sg U52463 ( .A(n34719), .B(reg_w_2[12]), .X(n24873) );
  nand_x1_sg U52464 ( .A(reg_ww_2[14]), .B(n32328), .X(n24876) );
  nand_x1_sg U52465 ( .A(n32741), .B(reg_w_2[14]), .X(n24877) );
  nand_x1_sg U52466 ( .A(reg_ww_2[15]), .B(n32336), .X(n24878) );
  nand_x1_sg U52467 ( .A(n35211), .B(reg_w_2[15]), .X(n24879) );
  nand_x1_sg U52468 ( .A(reg_ww_2[17]), .B(n32367), .X(n24882) );
  nand_x1_sg U52469 ( .A(n35371), .B(reg_w_2[17]), .X(n24883) );
  nand_x1_sg U52470 ( .A(reg_ww_2[18]), .B(n30611), .X(n24884) );
  nand_x1_sg U52471 ( .A(n35353), .B(reg_w_2[18]), .X(n24885) );
  nand_x1_sg U52472 ( .A(reg_ww_5[1]), .B(n33945), .X(n24294) );
  nand_x1_sg U52473 ( .A(n34055), .B(reg_w_5[1]), .X(n24295) );
  nand_x1_sg U52474 ( .A(reg_ww_5[2]), .B(n32348), .X(n24296) );
  nand_x1_sg U52475 ( .A(n35335), .B(reg_w_5[2]), .X(n24297) );
  nand_x1_sg U52476 ( .A(reg_ww_5[4]), .B(n32337), .X(n24300) );
  nand_x1_sg U52477 ( .A(n31692), .B(reg_w_5[4]), .X(n24301) );
  nand_x1_sg U52478 ( .A(reg_ww_5[5]), .B(n31509), .X(n24302) );
  nand_x1_sg U52479 ( .A(n35183), .B(reg_w_5[5]), .X(n24303) );
  nand_x1_sg U52480 ( .A(reg_ww_5[7]), .B(n32356), .X(n24306) );
  nand_x1_sg U52481 ( .A(n35209), .B(reg_w_5[7]), .X(n24307) );
  nand_x1_sg U52482 ( .A(reg_ww_5[8]), .B(n34937), .X(n24308) );
  nand_x1_sg U52483 ( .A(n34668), .B(reg_w_5[8]), .X(n24309) );
  nand_x1_sg U52484 ( .A(reg_ww_5[10]), .B(n32429), .X(n24312) );
  nand_x1_sg U52485 ( .A(n35185), .B(reg_w_5[10]), .X(n24313) );
  nand_x1_sg U52486 ( .A(reg_ww_5[11]), .B(n34583), .X(n24314) );
  nand_x1_sg U52487 ( .A(n35342), .B(reg_w_5[11]), .X(n24315) );
  nand_x1_sg U52488 ( .A(reg_ww_5[13]), .B(n32363), .X(n24318) );
  nand_x1_sg U52489 ( .A(n34081), .B(reg_w_5[13]), .X(n24319) );
  nand_x1_sg U52490 ( .A(reg_ww_5[14]), .B(n32016), .X(n24320) );
  nand_x1_sg U52491 ( .A(n32724), .B(reg_w_5[14]), .X(n24321) );
  nand_x1_sg U52492 ( .A(reg_ww_5[16]), .B(n32359), .X(n24324) );
  nand_x1_sg U52493 ( .A(n35320), .B(reg_w_5[16]), .X(n24325) );
  nand_x1_sg U52494 ( .A(reg_ww_5[17]), .B(n34847), .X(n24326) );
  nand_x1_sg U52495 ( .A(n34055), .B(reg_w_5[17]), .X(n24327) );
  nand_x1_sg U52496 ( .A(reg_ww_5[19]), .B(n31645), .X(n24330) );
  nand_x1_sg U52497 ( .A(n34094), .B(reg_w_5[19]), .X(n24331) );
  nand_x1_sg U52498 ( .A(reg_ww_6[15]), .B(n32455), .X(n24402) );
  nand_x1_sg U52499 ( .A(n31690), .B(reg_w_6[15]), .X(n24403) );
  nand_x1_sg U52500 ( .A(reg_ww_6[16]), .B(n30014), .X(n24404) );
  nand_x1_sg U52501 ( .A(n35210), .B(reg_w_6[16]), .X(n24405) );
  nand_x1_sg U52502 ( .A(reg_ww_6[18]), .B(n32380), .X(n24408) );
  nand_x1_sg U52503 ( .A(n32844), .B(reg_w_6[18]), .X(n24409) );
  nand_x1_sg U52504 ( .A(reg_ww_6[19]), .B(n31643), .X(n24410) );
  nand_x1_sg U52505 ( .A(n32837), .B(reg_w_6[19]), .X(n24411) );
  nand_x1_sg U52506 ( .A(reg_ww_7[0]), .B(n31513), .X(n24452) );
  nand_x1_sg U52507 ( .A(n35379), .B(reg_w_7[0]), .X(n24453) );
  nand_x1_sg U52508 ( .A(reg_ww_7[2]), .B(n32368), .X(n24456) );
  nand_x1_sg U52509 ( .A(n34723), .B(reg_w_7[2]), .X(n24457) );
  nand_x1_sg U52510 ( .A(reg_ww_7[3]), .B(n32151), .X(n24458) );
  nand_x1_sg U52511 ( .A(n35347), .B(reg_w_7[3]), .X(n24459) );
  nand_x1_sg U52512 ( .A(reg_ww_7[5]), .B(n33947), .X(n24462) );
  nand_x1_sg U52513 ( .A(n35341), .B(reg_w_7[5]), .X(n24463) );
  nand_x1_sg U52514 ( .A(reg_ww_7[6]), .B(n32242), .X(n24464) );
  nand_x1_sg U52515 ( .A(n34005), .B(reg_w_7[6]), .X(n24465) );
  nand_x1_sg U52516 ( .A(reg_ww_8[1]), .B(n32232), .X(n24534) );
  nand_x1_sg U52517 ( .A(n35177), .B(reg_w_8[1]), .X(n24535) );
  nand_x1_sg U52518 ( .A(reg_ww_8[2]), .B(n32228), .X(n24536) );
  nand_x1_sg U52519 ( .A(n32735), .B(reg_w_8[2]), .X(n24537) );
  nand_x1_sg U52520 ( .A(reg_ww_8[4]), .B(n31739), .X(n24540) );
  nand_x1_sg U52521 ( .A(n34707), .B(reg_w_8[4]), .X(n24541) );
  nand_x1_sg U52522 ( .A(reg_ww_8[5]), .B(n32338), .X(n24542) );
  nand_x1_sg U52523 ( .A(n35330), .B(reg_w_8[5]), .X(n24543) );
  nand_x1_sg U52524 ( .A(reg_ww_8[7]), .B(n31890), .X(n24546) );
  nand_x1_sg U52525 ( .A(n35359), .B(reg_w_8[7]), .X(n24547) );
  nand_x1_sg U52526 ( .A(reg_ww_8[8]), .B(n32322), .X(n24548) );
  nand_x1_sg U52527 ( .A(n35367), .B(reg_w_8[8]), .X(n24549) );
  nand_x1_sg U52528 ( .A(reg_ww_8[10]), .B(n32311), .X(n24552) );
  nand_x1_sg U52529 ( .A(n35211), .B(reg_w_8[10]), .X(n24553) );
  nand_x1_sg U52530 ( .A(reg_ww_8[11]), .B(n32229), .X(n24554) );
  nand_x1_sg U52531 ( .A(n35361), .B(reg_w_8[11]), .X(n24555) );
  nand_x1_sg U52532 ( .A(reg_ww_8[13]), .B(n31633), .X(n24558) );
  nand_x1_sg U52533 ( .A(n35239), .B(reg_w_8[13]), .X(n24559) );
  nand_x1_sg U52534 ( .A(reg_ww_8[14]), .B(n32141), .X(n24560) );
  nand_x1_sg U52535 ( .A(n34719), .B(reg_w_8[14]), .X(n24561) );
  nand_x1_sg U52536 ( .A(reg_ww_9[5]), .B(n32339), .X(n23826) );
  nand_x1_sg U52537 ( .A(n34718), .B(reg_w_9[5]), .X(n23827) );
  nand_x1_sg U52538 ( .A(reg_ww_9[6]), .B(n31743), .X(n23828) );
  nand_x1_sg U52539 ( .A(n35195), .B(reg_w_9[6]), .X(n23829) );
  nand_x1_sg U52540 ( .A(reg_ww_9[8]), .B(n32012), .X(n23832) );
  nand_x1_sg U52541 ( .A(n29763), .B(reg_w_9[8]), .X(n23833) );
  nand_x1_sg U52542 ( .A(reg_ww_9[9]), .B(n31908), .X(n23834) );
  nand_x1_sg U52543 ( .A(n32829), .B(reg_w_9[9]), .X(n23835) );
  nand_x1_sg U52544 ( .A(reg_ww_9[11]), .B(n32149), .X(n23838) );
  nand_x1_sg U52545 ( .A(n35094), .B(reg_w_9[11]), .X(n23839) );
  nand_x1_sg U52546 ( .A(reg_ww_9[12]), .B(n32286), .X(n23840) );
  nand_x1_sg U52547 ( .A(n34662), .B(reg_w_9[12]), .X(n23841) );
  nand_x1_sg U52548 ( .A(reg_ww_9[14]), .B(n32252), .X(n23844) );
  nand_x1_sg U52549 ( .A(n35214), .B(reg_w_9[14]), .X(n23845) );
  nand_x1_sg U52550 ( .A(reg_ww_9[15]), .B(n32311), .X(n23846) );
  nand_x1_sg U52551 ( .A(n30178), .B(reg_w_9[15]), .X(n23847) );
  nand_x1_sg U52552 ( .A(reg_ww_9[17]), .B(n30195), .X(n23850) );
  nand_x1_sg U52553 ( .A(n34092), .B(reg_w_9[17]), .X(n23851) );
  nand_x1_sg U52554 ( .A(reg_ww_9[18]), .B(n32336), .X(n23852) );
  nand_x1_sg U52555 ( .A(n32760), .B(reg_w_9[18]), .X(n23853) );
  nand_x1_sg U52556 ( .A(reg_ww_11[0]), .B(n32150), .X(n23976) );
  nand_x1_sg U52557 ( .A(n32829), .B(reg_w_11[0]), .X(n23977) );
  nand_x1_sg U52558 ( .A(reg_ww_11[1]), .B(n32298), .X(n23978) );
  nand_x1_sg U52559 ( .A(n35361), .B(reg_w_11[1]), .X(n23979) );
  nand_x1_sg U52560 ( .A(reg_ww_11[3]), .B(n33943), .X(n23982) );
  nand_x1_sg U52561 ( .A(n35088), .B(reg_w_11[3]), .X(n23983) );
  nand_x1_sg U52562 ( .A(reg_ww_11[4]), .B(n32369), .X(n23984) );
  nand_x1_sg U52563 ( .A(n35179), .B(reg_w_11[4]), .X(n23985) );
  nand_x1_sg U52564 ( .A(reg_ww_11[6]), .B(n31515), .X(n23988) );
  nand_x1_sg U52565 ( .A(n35344), .B(reg_w_11[6]), .X(n23989) );
  nand_x1_sg U52566 ( .A(reg_ww_11[7]), .B(n34651), .X(n23990) );
  nand_x1_sg U52567 ( .A(n35210), .B(reg_w_11[7]), .X(n23991) );
  nand_x1_sg U52568 ( .A(reg_ww_11[9]), .B(n30208), .X(n23994) );
  nand_x1_sg U52569 ( .A(n34707), .B(reg_w_11[9]), .X(n23995) );
  nand_x1_sg U52570 ( .A(reg_ww_11[10]), .B(n32336), .X(n23996) );
  nand_x1_sg U52571 ( .A(n35377), .B(reg_w_11[10]), .X(n23997) );
  nand_x1_sg U52572 ( .A(reg_ww_11[12]), .B(n32037), .X(n24000) );
  nand_x1_sg U52573 ( .A(n34709), .B(reg_w_11[12]), .X(n24001) );
  nand_x1_sg U52574 ( .A(reg_ww_11[13]), .B(n32405), .X(n24002) );
  nand_x1_sg U52575 ( .A(n34094), .B(reg_w_11[13]), .X(n24003) );
  nand_x1_sg U52576 ( .A(reg_ww_11[15]), .B(n32372), .X(n24006) );
  nand_x1_sg U52577 ( .A(n31865), .B(reg_w_11[15]), .X(n24007) );
  nand_x1_sg U52578 ( .A(reg_ww_11[16]), .B(n34898), .X(n24008) );
  nand_x1_sg U52579 ( .A(n34703), .B(reg_w_11[16]), .X(n24009) );
  nand_x1_sg U52580 ( .A(reg_ww_11[18]), .B(n34896), .X(n24012) );
  nand_x1_sg U52581 ( .A(n35208), .B(reg_w_11[18]), .X(n24013) );
  nand_x1_sg U52582 ( .A(reg_ww_11[19]), .B(n30147), .X(n24014) );
  nand_x1_sg U52583 ( .A(n34712), .B(reg_w_11[19]), .X(n24015) );
  nand_x1_sg U52584 ( .A(reg_ww_15[0]), .B(n32026), .X(n23726) );
  nand_x1_sg U52585 ( .A(n34074), .B(reg_w_15[0]), .X(n23727) );
  nand_x1_sg U52586 ( .A(reg_ww_15[2]), .B(n32355), .X(n23730) );
  nand_x1_sg U52587 ( .A(n35228), .B(reg_w_15[2]), .X(n23731) );
  nand_x1_sg U52588 ( .A(reg_ww_15[3]), .B(n32454), .X(n23732) );
  nand_x1_sg U52589 ( .A(n35209), .B(reg_w_15[3]), .X(n23733) );
  nand_x1_sg U52590 ( .A(reg_ww_15[5]), .B(n32342), .X(n23736) );
  nand_x1_sg U52591 ( .A(n32717), .B(reg_w_15[5]), .X(n23737) );
  nand_x1_sg U52592 ( .A(reg_ww_15[6]), .B(n33948), .X(n23738) );
  nand_x1_sg U52593 ( .A(n34074), .B(reg_w_15[6]), .X(n23739) );
  nand_x1_sg U52594 ( .A(reg_ww_15[8]), .B(n31719), .X(n23742) );
  nand_x1_sg U52595 ( .A(n31871), .B(reg_w_15[8]), .X(n23743) );
  nand_x1_sg U52596 ( .A(reg_ww_15[9]), .B(n32302), .X(n23744) );
  nand_x1_sg U52597 ( .A(n35228), .B(reg_w_15[9]), .X(n23745) );
  nand_x1_sg U52598 ( .A(reg_ww_15[11]), .B(n31636), .X(n23748) );
  nand_x1_sg U52599 ( .A(n34722), .B(reg_w_15[11]), .X(n23749) );
  nand_x1_sg U52600 ( .A(reg_ww_15[12]), .B(n32428), .X(n23750) );
  nand_x1_sg U52601 ( .A(n31692), .B(reg_w_15[12]), .X(n23751) );
  nand_x1_sg U52602 ( .A(reg_ww_15[14]), .B(n32340), .X(n23754) );
  nand_x1_sg U52603 ( .A(n31690), .B(reg_w_15[14]), .X(n23755) );
  nand_x1_sg U52604 ( .A(reg_ww_15[15]), .B(n32362), .X(n23756) );
  nand_x1_sg U52605 ( .A(n31671), .B(reg_w_15[15]), .X(n23757) );
  nand_x1_sg U52606 ( .A(reg_ww_15[17]), .B(n32280), .X(n23760) );
  nand_x1_sg U52607 ( .A(n32835), .B(reg_w_15[17]), .X(n23761) );
  nand_x1_sg U52608 ( .A(reg_ii_3[1]), .B(n32036), .X(n26038) );
  nand_x1_sg U52609 ( .A(n32714), .B(reg_i_3[1]), .X(n26039) );
  nand_x1_sg U52610 ( .A(reg_ii_3[4]), .B(n32034), .X(n26044) );
  nand_x1_sg U52611 ( .A(n35162), .B(reg_i_3[4]), .X(n26045) );
  nand_x1_sg U52612 ( .A(reg_ii_3[7]), .B(n32288), .X(n26050) );
  nand_x1_sg U52613 ( .A(n32738), .B(reg_i_3[7]), .X(n26051) );
  nand_x1_sg U52614 ( .A(reg_ii_3[10]), .B(n34936), .X(n26056) );
  nand_x1_sg U52615 ( .A(n34048), .B(reg_i_3[10]), .X(n26057) );
  nand_x1_sg U52616 ( .A(reg_ii_3[13]), .B(n32295), .X(n26062) );
  nand_x1_sg U52617 ( .A(n35194), .B(reg_i_3[13]), .X(n26063) );
  nand_x1_sg U52618 ( .A(reg_ii_4[9]), .B(n32300), .X(n26134) );
  nand_x1_sg U52619 ( .A(n34002), .B(reg_i_4[9]), .X(n26135) );
  nand_x1_sg U52620 ( .A(reg_ii_4[12]), .B(n32856), .X(n26140) );
  nand_x1_sg U52621 ( .A(n34666), .B(reg_i_4[12]), .X(n26141) );
  nand_x1_sg U52622 ( .A(reg_ii_4[15]), .B(n30622), .X(n26146) );
  nand_x1_sg U52623 ( .A(n32761), .B(reg_i_4[15]), .X(n26147) );
  nand_x1_sg U52624 ( .A(reg_ii_4[18]), .B(n32401), .X(n26152) );
  nand_x1_sg U52625 ( .A(n35173), .B(reg_i_4[18]), .X(n26153) );
  nand_x1_sg U52626 ( .A(reg_ii_5[13]), .B(n32145), .X(n25426) );
  nand_x1_sg U52627 ( .A(n30023), .B(reg_i_5[13]), .X(n25427) );
  nand_x1_sg U52628 ( .A(reg_ii_5[16]), .B(n32308), .X(n25432) );
  nand_x1_sg U52629 ( .A(n32839), .B(reg_i_5[16]), .X(n25433) );
  nand_x1_sg U52630 ( .A(reg_ii_5[19]), .B(n32362), .X(n25438) );
  nand_x1_sg U52631 ( .A(n35355), .B(reg_i_5[19]), .X(n25439) );
  nand_x1_sg U52632 ( .A(reg_ii_6[0]), .B(n32331), .X(n25480) );
  nand_x1_sg U52633 ( .A(n35240), .B(reg_i_6[0]), .X(n25481) );
  nand_x1_sg U52634 ( .A(reg_ii_6[3]), .B(n32402), .X(n25486) );
  nand_x1_sg U52635 ( .A(n35326), .B(reg_i_6[3]), .X(n25487) );
  nand_x1_sg U52636 ( .A(reg_ii_7[2]), .B(n32292), .X(n25564) );
  nand_x1_sg U52637 ( .A(n35399), .B(reg_i_7[2]), .X(n25565) );
  nand_x1_sg U52638 ( .A(reg_ii_7[5]), .B(n34552), .X(n25570) );
  nand_x1_sg U52639 ( .A(n35336), .B(reg_i_7[5]), .X(n25571) );
  nand_x1_sg U52640 ( .A(reg_ii_7[8]), .B(n32855), .X(n25576) );
  nand_x1_sg U52641 ( .A(n34057), .B(reg_i_7[8]), .X(n25577) );
  nand_x1_sg U52642 ( .A(reg_ii_7[11]), .B(n32144), .X(n25582) );
  nand_x1_sg U52643 ( .A(n35222), .B(reg_i_7[11]), .X(n25583) );
  nand_x1_sg U52644 ( .A(reg_ii_7[14]), .B(n31631), .X(n25588) );
  nand_x1_sg U52645 ( .A(n35396), .B(reg_i_7[14]), .X(n25589) );
  nand_x1_sg U52646 ( .A(reg_ii_7[17]), .B(n32049), .X(n25594) );
  nand_x1_sg U52647 ( .A(n31862), .B(reg_i_7[17]), .X(n25595) );
  nand_x1_sg U52648 ( .A(reg_ii_9[0]), .B(n31719), .X(n25720) );
  nand_x1_sg U52649 ( .A(n35184), .B(reg_i_9[0]), .X(n25721) );
  nand_x1_sg U52650 ( .A(reg_ii_9[3]), .B(n32215), .X(n25726) );
  nand_x1_sg U52651 ( .A(n34073), .B(reg_i_9[3]), .X(n25727) );
  nand_x1_sg U52652 ( .A(reg_ii_9[6]), .B(n31737), .X(n25732) );
  nand_x1_sg U52653 ( .A(n32830), .B(reg_i_9[6]), .X(n25733) );
  nand_x1_sg U52654 ( .A(reg_ii_9[9]), .B(n29755), .X(n25738) );
  nand_x1_sg U52655 ( .A(n32440), .B(reg_i_9[9]), .X(n25739) );
  nand_x1_sg U52656 ( .A(reg_ii_9[12]), .B(n34582), .X(n25744) );
  nand_x1_sg U52657 ( .A(n35218), .B(reg_i_9[12]), .X(n25745) );
  nand_x1_sg U52658 ( .A(reg_ii_9[18]), .B(n32493), .X(n25000) );
  nand_x1_sg U52659 ( .A(n34076), .B(reg_i_9[18]), .X(n25001) );
  nand_x1_sg U52660 ( .A(reg_ii_10[1]), .B(n33942), .X(n25006) );
  nand_x1_sg U52661 ( .A(n35090), .B(reg_i_10[1]), .X(n25007) );
  nand_x1_sg U52662 ( .A(reg_ii_10[4]), .B(n34940), .X(n25012) );
  nand_x1_sg U52663 ( .A(n34665), .B(reg_i_10[4]), .X(n25013) );
  nand_x1_sg U52664 ( .A(reg_ii_10[7]), .B(n33972), .X(n25018) );
  nand_x1_sg U52665 ( .A(n34047), .B(reg_i_10[7]), .X(n25019) );
  nand_x1_sg U52666 ( .A(reg_ii_10[10]), .B(n31889), .X(n25024) );
  nand_x1_sg U52667 ( .A(n32731), .B(reg_i_10[10]), .X(n25025) );
  nand_x1_sg U52668 ( .A(reg_ii_10[13]), .B(n32357), .X(n25030) );
  nand_x1_sg U52669 ( .A(n34052), .B(reg_i_10[13]), .X(n25031) );
  nand_x1_sg U52670 ( .A(reg_ii_10[16]), .B(n32369), .X(n25036) );
  nand_x1_sg U52671 ( .A(n32842), .B(reg_i_10[16]), .X(n25037) );
  nand_x1_sg U52672 ( .A(reg_ii_11[12]), .B(n32297), .X(n25108) );
  nand_x1_sg U52673 ( .A(n35186), .B(reg_i_11[12]), .X(n25109) );
  nand_x1_sg U52674 ( .A(reg_ii_11[15]), .B(n32321), .X(n25114) );
  nand_x1_sg U52675 ( .A(n34042), .B(reg_i_11[15]), .X(n25115) );
  nand_x1_sg U52676 ( .A(reg_ii_11[18]), .B(n31897), .X(n25120) );
  nand_x1_sg U52677 ( .A(n34046), .B(reg_i_11[18]), .X(n25121) );
  nand_x1_sg U52678 ( .A(reg_ii_12[2]), .B(n31713), .X(n25168) );
  nand_x1_sg U52679 ( .A(n35219), .B(reg_i_12[2]), .X(n25169) );
  nand_x1_sg U52680 ( .A(reg_ww_2[1]), .B(n32301), .X(n24850) );
  nand_x1_sg U52681 ( .A(n34663), .B(reg_w_2[1]), .X(n24851) );
  nand_x1_sg U52682 ( .A(reg_ww_2[4]), .B(n30207), .X(n24856) );
  nand_x1_sg U52683 ( .A(n35089), .B(reg_w_2[4]), .X(n24857) );
  nand_x1_sg U52684 ( .A(reg_ww_2[7]), .B(n29755), .X(n24862) );
  nand_x1_sg U52685 ( .A(n31868), .B(reg_w_2[7]), .X(n24863) );
  nand_x1_sg U52686 ( .A(reg_ww_2[10]), .B(n30176), .X(n24868) );
  nand_x1_sg U52687 ( .A(n32731), .B(reg_w_2[10]), .X(n24869) );
  nand_x1_sg U52688 ( .A(reg_ww_2[13]), .B(n32014), .X(n24874) );
  nand_x1_sg U52689 ( .A(n34705), .B(reg_w_2[13]), .X(n24875) );
  nand_x1_sg U52690 ( .A(reg_ww_2[16]), .B(n32217), .X(n24880) );
  nand_x1_sg U52691 ( .A(n31873), .B(reg_w_2[16]), .X(n24881) );
  nand_x1_sg U52692 ( .A(reg_ww_2[19]), .B(n32241), .X(n24886) );
  nand_x1_sg U52693 ( .A(n31869), .B(reg_w_2[19]), .X(n24887) );
  nand_x1_sg U52694 ( .A(reg_ww_5[0]), .B(n32311), .X(n24292) );
  nand_x1_sg U52695 ( .A(n32711), .B(reg_w_5[0]), .X(n24293) );
  nand_x1_sg U52696 ( .A(reg_ww_5[3]), .B(n32040), .X(n24298) );
  nand_x1_sg U52697 ( .A(n34052), .B(reg_w_5[3]), .X(n24299) );
  nand_x1_sg U52698 ( .A(reg_ww_5[6]), .B(n32165), .X(n24304) );
  nand_x1_sg U52699 ( .A(n32841), .B(reg_w_5[6]), .X(n24305) );
  nand_x1_sg U52700 ( .A(reg_ww_5[9]), .B(n32027), .X(n24310) );
  nand_x1_sg U52701 ( .A(n31872), .B(reg_w_5[9]), .X(n24311) );
  nand_x1_sg U52702 ( .A(reg_ww_5[12]), .B(n34697), .X(n24316) );
  nand_x1_sg U52703 ( .A(n35339), .B(reg_w_5[12]), .X(n24317) );
  nand_x1_sg U52704 ( .A(reg_ww_5[15]), .B(n32378), .X(n24322) );
  nand_x1_sg U52705 ( .A(n32708), .B(reg_w_5[15]), .X(n24323) );
  nand_x1_sg U52706 ( .A(reg_ww_5[18]), .B(n32378), .X(n24328) );
  nand_x1_sg U52707 ( .A(n35216), .B(reg_w_5[18]), .X(n24329) );
  nand_x1_sg U52708 ( .A(reg_ww_6[17]), .B(n33951), .X(n24406) );
  nand_x1_sg U52709 ( .A(n34007), .B(reg_w_6[17]), .X(n24407) );
  nand_x1_sg U52710 ( .A(reg_ww_7[1]), .B(n30754), .X(n24454) );
  nand_x1_sg U52711 ( .A(n31673), .B(reg_w_7[1]), .X(n24455) );
  nand_x1_sg U52712 ( .A(reg_ww_7[4]), .B(n32233), .X(n24460) );
  nand_x1_sg U52713 ( .A(n34052), .B(reg_w_7[4]), .X(n24461) );
  nand_x1_sg U52714 ( .A(reg_ww_8[0]), .B(n32770), .X(n24532) );
  nand_x1_sg U52715 ( .A(n35239), .B(reg_w_8[0]), .X(n24533) );
  nand_x1_sg U52716 ( .A(reg_ww_8[3]), .B(n32231), .X(n24538) );
  nand_x1_sg U52717 ( .A(n32840), .B(reg_w_8[3]), .X(n24539) );
  nand_x1_sg U52718 ( .A(reg_ww_8[6]), .B(n32239), .X(n24544) );
  nand_x1_sg U52719 ( .A(n32733), .B(reg_w_8[6]), .X(n24545) );
  nand_x1_sg U52720 ( .A(reg_ww_8[9]), .B(n32303), .X(n24550) );
  nand_x1_sg U52721 ( .A(n34043), .B(reg_w_8[9]), .X(n24551) );
  nand_x1_sg U52722 ( .A(reg_ww_8[12]), .B(n32158), .X(n24556) );
  nand_x1_sg U52723 ( .A(n35228), .B(reg_w_8[12]), .X(n24557) );
  nand_x1_sg U52724 ( .A(reg_ww_9[7]), .B(n32343), .X(n23830) );
  nand_x1_sg U52725 ( .A(n35318), .B(reg_w_9[7]), .X(n23831) );
  nand_x1_sg U52726 ( .A(reg_ww_9[10]), .B(n32155), .X(n23836) );
  nand_x1_sg U52727 ( .A(n35336), .B(reg_w_9[10]), .X(n23837) );
  nand_x1_sg U52728 ( .A(reg_ww_9[13]), .B(n32325), .X(n23842) );
  nand_x1_sg U52729 ( .A(n35395), .B(reg_w_9[13]), .X(n23843) );
  nand_x1_sg U52730 ( .A(reg_ww_9[16]), .B(n32291), .X(n23848) );
  nand_x1_sg U52731 ( .A(n31863), .B(reg_w_9[16]), .X(n23849) );
  nand_x1_sg U52732 ( .A(reg_ww_9[19]), .B(n31900), .X(n23854) );
  nand_x1_sg U52733 ( .A(n32753), .B(reg_w_9[19]), .X(n23855) );
  nand_x1_sg U52734 ( .A(reg_ww_11[2]), .B(n32232), .X(n23980) );
  nand_x1_sg U52735 ( .A(n34096), .B(reg_w_11[2]), .X(n23981) );
  nand_x1_sg U52736 ( .A(reg_ww_11[5]), .B(n31740), .X(n23986) );
  nand_x1_sg U52737 ( .A(n35344), .B(reg_w_11[5]), .X(n23987) );
  nand_x1_sg U52738 ( .A(reg_ww_11[8]), .B(n31645), .X(n23992) );
  nand_x1_sg U52739 ( .A(n34703), .B(reg_w_11[8]), .X(n23993) );
  nand_x1_sg U52740 ( .A(reg_ww_11[11]), .B(n32385), .X(n23998) );
  nand_x1_sg U52741 ( .A(n35165), .B(reg_w_11[11]), .X(n23999) );
  nand_x1_sg U52742 ( .A(reg_ww_11[14]), .B(n32044), .X(n24004) );
  nand_x1_sg U52743 ( .A(n34097), .B(reg_w_11[14]), .X(n24005) );
  nand_x1_sg U52744 ( .A(reg_ww_11[17]), .B(n32368), .X(n24010) );
  nand_x1_sg U52745 ( .A(n34708), .B(reg_w_11[17]), .X(n24011) );
  nand_x1_sg U52746 ( .A(reg_ww_15[1]), .B(n34572), .X(n23728) );
  nand_x1_sg U52747 ( .A(n34081), .B(reg_w_15[1]), .X(n23729) );
  nand_x1_sg U52748 ( .A(reg_ww_15[4]), .B(n34570), .X(n23734) );
  nand_x1_sg U52749 ( .A(n30592), .B(reg_w_15[4]), .X(n23735) );
  nand_x1_sg U52750 ( .A(reg_ww_15[7]), .B(n32339), .X(n23740) );
  nand_x1_sg U52751 ( .A(n34076), .B(reg_w_15[7]), .X(n23741) );
  nand_x1_sg U52752 ( .A(reg_ww_15[10]), .B(n31631), .X(n23746) );
  nand_x1_sg U52753 ( .A(n34717), .B(reg_w_15[10]), .X(n23747) );
  nand_x1_sg U52754 ( .A(reg_ww_15[13]), .B(n32494), .X(n23752) );
  nand_x1_sg U52755 ( .A(n35198), .B(reg_w_15[13]), .X(n23753) );
  nand_x1_sg U52756 ( .A(reg_ww_15[16]), .B(n32010), .X(n23758) );
  nand_x1_sg U52757 ( .A(n32442), .B(reg_w_15[16]), .X(n23759) );
  nand_x1_sg U52758 ( .A(reg_iii_0[19]), .B(n31727), .X(n25874) );
  nand_x1_sg U52759 ( .A(reg_ii_0[19]), .B(n30882), .X(n25875) );
  nand_x1_sg U52760 ( .A(reg_iii_1[0]), .B(n32320), .X(n25916) );
  nand_x1_sg U52761 ( .A(reg_ii_1[0]), .B(n35223), .X(n25917) );
  nand_x1_sg U52762 ( .A(reg_ii_1[1]), .B(n32310), .X(n25878) );
  nand_x1_sg U52763 ( .A(n31862), .B(reg_i_1[1]), .X(n25879) );
  nand_x1_sg U52764 ( .A(reg_iii_1[2]), .B(n32302), .X(n25920) );
  nand_x1_sg U52765 ( .A(reg_ii_1[2]), .B(n32708), .X(n25921) );
  nand_x1_sg U52766 ( .A(reg_ii_1[2]), .B(n32386), .X(n25880) );
  nand_x1_sg U52767 ( .A(n35239), .B(reg_i_1[2]), .X(n25881) );
  nand_x1_sg U52768 ( .A(reg_iii_1[3]), .B(n32345), .X(n25922) );
  nand_x1_sg U52769 ( .A(reg_ii_1[3]), .B(n32847), .X(n25923) );
  nand_x1_sg U52770 ( .A(reg_ii_1[4]), .B(n31509), .X(n25884) );
  nand_x1_sg U52771 ( .A(n34705), .B(reg_i_1[4]), .X(n25885) );
  nand_x1_sg U52772 ( .A(reg_iii_1[5]), .B(n33967), .X(n25926) );
  nand_x1_sg U52773 ( .A(reg_ii_1[5]), .B(n32759), .X(n25927) );
  nand_x1_sg U52774 ( .A(reg_ii_1[5]), .B(n32383), .X(n25886) );
  nand_x1_sg U52775 ( .A(n35220), .B(reg_i_1[5]), .X(n25887) );
  nand_x1_sg U52776 ( .A(reg_iii_1[6]), .B(n32027), .X(n25928) );
  nand_x1_sg U52777 ( .A(reg_ii_1[6]), .B(n31491), .X(n25929) );
  nand_x1_sg U52778 ( .A(reg_ii_1[7]), .B(n32028), .X(n25890) );
  nand_x1_sg U52779 ( .A(n35379), .B(reg_i_1[7]), .X(n25891) );
  nand_x1_sg U52780 ( .A(reg_iii_1[8]), .B(n32313), .X(n25932) );
  nand_x1_sg U52781 ( .A(reg_ii_1[8]), .B(n35164), .X(n25933) );
  nand_x1_sg U52782 ( .A(reg_ii_1[8]), .B(n30914), .X(n25892) );
  nand_x1_sg U52783 ( .A(n35329), .B(reg_i_1[8]), .X(n25893) );
  nand_x1_sg U52784 ( .A(reg_iii_1[9]), .B(n32374), .X(n25934) );
  nand_x1_sg U52785 ( .A(reg_ii_1[9]), .B(n32765), .X(n25935) );
  nand_x1_sg U52786 ( .A(reg_ii_1[10]), .B(n33976), .X(n25896) );
  nand_x1_sg U52787 ( .A(n35184), .B(reg_i_1[10]), .X(n25897) );
  nand_x1_sg U52788 ( .A(reg_iii_1[11]), .B(n32348), .X(n25938) );
  nand_x1_sg U52789 ( .A(reg_ii_1[11]), .B(n30902), .X(n25939) );
  nand_x1_sg U52790 ( .A(reg_ii_1[11]), .B(n32406), .X(n25898) );
  nand_x1_sg U52791 ( .A(n31870), .B(reg_i_1[11]), .X(n25899) );
  nand_x1_sg U52792 ( .A(reg_iii_1[12]), .B(n31721), .X(n25940) );
  nand_x1_sg U52793 ( .A(reg_ii_1[12]), .B(n35189), .X(n25941) );
  nand_x1_sg U52794 ( .A(reg_ii_1[13]), .B(n32287), .X(n25902) );
  nand_x1_sg U52795 ( .A(n32730), .B(reg_i_1[13]), .X(n25903) );
  nand_x1_sg U52796 ( .A(reg_iii_1[14]), .B(n32326), .X(n25944) );
  nand_x1_sg U52797 ( .A(reg_ii_1[14]), .B(n30865), .X(n25945) );
  nand_x1_sg U52798 ( .A(reg_ii_1[14]), .B(n32325), .X(n25904) );
  nand_x1_sg U52799 ( .A(n31862), .B(reg_i_1[14]), .X(n25905) );
  nand_x1_sg U52800 ( .A(reg_iii_1[15]), .B(n32149), .X(n25946) );
  nand_x1_sg U52801 ( .A(reg_ii_1[15]), .B(n30867), .X(n25947) );
  nand_x1_sg U52802 ( .A(reg_ii_1[16]), .B(n31725), .X(n25908) );
  nand_x1_sg U52803 ( .A(n32767), .B(reg_i_1[16]), .X(n25909) );
  nand_x1_sg U52804 ( .A(reg_iii_1[17]), .B(n31901), .X(n25950) );
  nand_x1_sg U52805 ( .A(reg_ii_1[17]), .B(n35214), .X(n25951) );
  nand_x1_sg U52806 ( .A(reg_ii_1[17]), .B(n32326), .X(n25910) );
  nand_x1_sg U52807 ( .A(n35317), .B(reg_i_1[17]), .X(n25911) );
  nand_x1_sg U52808 ( .A(reg_iii_1[18]), .B(n32158), .X(n25952) );
  nand_x1_sg U52809 ( .A(reg_ii_1[18]), .B(n35212), .X(n25953) );
  nand_x1_sg U52810 ( .A(reg_ii_1[19]), .B(n32362), .X(n25914) );
  nand_x1_sg U52811 ( .A(n32743), .B(reg_i_1[19]), .X(n25915) );
  nand_x1_sg U52812 ( .A(reg_ii_2[0]), .B(n32361), .X(n25956) );
  nand_x1_sg U52813 ( .A(n34077), .B(reg_i_2[0]), .X(n25957) );
  nand_x1_sg U52814 ( .A(reg_iii_2[1]), .B(n32020), .X(n25998) );
  nand_x1_sg U52815 ( .A(reg_ii_2[1]), .B(n30872), .X(n25999) );
  nand_x1_sg U52816 ( .A(reg_ii_2[1]), .B(n30621), .X(n25958) );
  nand_x1_sg U52817 ( .A(n35350), .B(reg_i_2[1]), .X(n25959) );
  nand_x1_sg U52818 ( .A(reg_iii_2[2]), .B(n31906), .X(n26000) );
  nand_x1_sg U52819 ( .A(reg_ii_2[2]), .B(n35183), .X(n26001) );
  nand_x1_sg U52820 ( .A(reg_ii_2[3]), .B(n32317), .X(n25962) );
  nand_x1_sg U52821 ( .A(n31691), .B(reg_i_2[3]), .X(n25963) );
  nand_x1_sg U52822 ( .A(reg_ii_2[4]), .B(n32238), .X(n25964) );
  nand_x1_sg U52823 ( .A(n35217), .B(reg_i_2[4]), .X(n25965) );
  nand_x1_sg U52824 ( .A(reg_ii_2[6]), .B(n32769), .X(n25968) );
  nand_x1_sg U52825 ( .A(n31674), .B(reg_i_2[6]), .X(n25969) );
  nand_x1_sg U52826 ( .A(reg_ii_2[7]), .B(n30755), .X(n25970) );
  nand_x1_sg U52827 ( .A(n31691), .B(reg_i_2[7]), .X(n25971) );
  nand_x1_sg U52828 ( .A(reg_ii_2[9]), .B(n31723), .X(n25974) );
  nand_x1_sg U52829 ( .A(n34667), .B(reg_i_2[9]), .X(n25975) );
  nand_x1_sg U52830 ( .A(reg_ii_2[10]), .B(n31898), .X(n25976) );
  nand_x1_sg U52831 ( .A(n35214), .B(reg_i_2[10]), .X(n25977) );
  nand_x1_sg U52832 ( .A(reg_ii_2[12]), .B(n32283), .X(n25980) );
  nand_x1_sg U52833 ( .A(n35320), .B(reg_i_2[12]), .X(n25981) );
  nand_x1_sg U52834 ( .A(reg_ii_2[13]), .B(n31731), .X(n25982) );
  nand_x1_sg U52835 ( .A(n34097), .B(reg_i_2[13]), .X(n25983) );
  nand_x1_sg U52836 ( .A(reg_ii_2[15]), .B(n32351), .X(n25986) );
  nand_x1_sg U52837 ( .A(n34072), .B(reg_i_2[15]), .X(n25987) );
  nand_x1_sg U52838 ( .A(reg_ii_2[16]), .B(n32501), .X(n25988) );
  nand_x1_sg U52839 ( .A(n35326), .B(reg_i_2[16]), .X(n25989) );
  nand_x1_sg U52840 ( .A(reg_ii_2[18]), .B(n33968), .X(n25992) );
  nand_x1_sg U52841 ( .A(n35379), .B(reg_i_2[18]), .X(n25993) );
  nand_x1_sg U52842 ( .A(reg_ii_2[19]), .B(n31630), .X(n25994) );
  nand_x1_sg U52843 ( .A(n34045), .B(reg_i_2[19]), .X(n25995) );
  nand_x1_sg U52844 ( .A(reg_ii_4[19]), .B(n32231), .X(n25398) );
  nand_x1_sg U52845 ( .A(n34074), .B(reg_i_4[19]), .X(n25399) );
  nand_x1_sg U52846 ( .A(reg_ii_5[0]), .B(n32237), .X(n25400) );
  nand_x1_sg U52847 ( .A(n34094), .B(reg_i_5[0]), .X(n25401) );
  nand_x1_sg U52848 ( .A(reg_ii_5[2]), .B(n32352), .X(n25404) );
  nand_x1_sg U52849 ( .A(n32760), .B(reg_i_5[2]), .X(n25405) );
  nand_x1_sg U52850 ( .A(reg_ii_5[3]), .B(n31715), .X(n25406) );
  nand_x1_sg U52851 ( .A(n34707), .B(reg_i_5[3]), .X(n25407) );
  nand_x1_sg U52852 ( .A(reg_ii_5[5]), .B(n32281), .X(n25410) );
  nand_x1_sg U52853 ( .A(n34057), .B(reg_i_5[5]), .X(n25411) );
  nand_x1_sg U52854 ( .A(reg_ii_5[6]), .B(n34697), .X(n25412) );
  nand_x1_sg U52855 ( .A(n31871), .B(reg_i_5[6]), .X(n25413) );
  nand_x1_sg U52856 ( .A(reg_ii_5[8]), .B(n30916), .X(n25416) );
  nand_x1_sg U52857 ( .A(n34716), .B(reg_i_5[8]), .X(n25417) );
  nand_x1_sg U52858 ( .A(reg_ii_5[9]), .B(n32500), .X(n25418) );
  nand_x1_sg U52859 ( .A(n32719), .B(reg_i_5[9]), .X(n25419) );
  nand_x1_sg U52860 ( .A(reg_ii_5[11]), .B(n34898), .X(n25422) );
  nand_x1_sg U52861 ( .A(n35404), .B(reg_i_5[11]), .X(n25423) );
  nand_x1_sg U52862 ( .A(reg_ii_5[12]), .B(n31898), .X(n25424) );
  nand_x1_sg U52863 ( .A(n34050), .B(reg_i_5[12]), .X(n25425) );
  nand_x1_sg U52864 ( .A(reg_iii_7[10]), .B(n32239), .X(n25620) );
  nand_x1_sg U52865 ( .A(reg_ii_7[10]), .B(n32741), .X(n25621) );
  nand_x1_sg U52866 ( .A(reg_iii_7[11]), .B(n31639), .X(n25622) );
  nand_x1_sg U52867 ( .A(reg_ii_7[11]), .B(n31490), .X(n25623) );
  nand_x1_sg U52868 ( .A(reg_iii_7[13]), .B(n32401), .X(n25626) );
  nand_x1_sg U52869 ( .A(reg_ii_7[13]), .B(n31041), .X(n25627) );
  nand_x1_sg U52870 ( .A(reg_iii_7[14]), .B(n32287), .X(n25628) );
  nand_x1_sg U52871 ( .A(reg_ii_7[14]), .B(n30868), .X(n25629) );
  nand_x1_sg U52872 ( .A(reg_iii_7[16]), .B(n34696), .X(n25632) );
  nand_x1_sg U52873 ( .A(reg_ii_7[16]), .B(n34043), .X(n25633) );
  nand_x1_sg U52874 ( .A(reg_iii_7[17]), .B(n32028), .X(n25634) );
  nand_x1_sg U52875 ( .A(reg_ii_7[17]), .B(n30586), .X(n25635) );
  nand_x1_sg U52876 ( .A(reg_iii_7[19]), .B(n32281), .X(n25638) );
  nand_x1_sg U52877 ( .A(reg_ii_7[19]), .B(n30720), .X(n25639) );
  nand_x1_sg U52878 ( .A(reg_iii_8[0]), .B(n34575), .X(n25680) );
  nand_x1_sg U52879 ( .A(reg_ii_8[0]), .B(n31093), .X(n25681) );
  nand_x1_sg U52880 ( .A(reg_ii_8[0]), .B(n32138), .X(n25640) );
  nand_x1_sg U52881 ( .A(n31863), .B(reg_i_8[0]), .X(n25641) );
  nand_x1_sg U52882 ( .A(reg_ii_8[2]), .B(n32045), .X(n25644) );
  nand_x1_sg U52883 ( .A(n35198), .B(reg_i_8[2]), .X(n25645) );
  nand_x1_sg U52884 ( .A(reg_ii_8[3]), .B(n32216), .X(n25646) );
  nand_x1_sg U52885 ( .A(n35321), .B(reg_i_8[3]), .X(n25647) );
  nand_x1_sg U52886 ( .A(reg_ii_8[5]), .B(n32328), .X(n25650) );
  nand_x1_sg U52887 ( .A(n35197), .B(reg_i_8[5]), .X(n25651) );
  nand_x1_sg U52888 ( .A(reg_ii_8[6]), .B(n31744), .X(n25652) );
  nand_x1_sg U52889 ( .A(n34708), .B(reg_i_8[6]), .X(n25653) );
  nand_x1_sg U52890 ( .A(reg_ii_8[8]), .B(n34698), .X(n25656) );
  nand_x1_sg U52891 ( .A(n31097), .B(reg_i_8[8]), .X(n25657) );
  nand_x1_sg U52892 ( .A(reg_ii_8[9]), .B(n30198), .X(n25658) );
  nand_x1_sg U52893 ( .A(n34706), .B(reg_i_8[9]), .X(n25659) );
  nand_x1_sg U52894 ( .A(reg_ii_8[11]), .B(n32144), .X(n25662) );
  nand_x1_sg U52895 ( .A(n35081), .B(reg_i_8[11]), .X(n25663) );
  nand_x1_sg U52896 ( .A(reg_ii_8[12]), .B(n32034), .X(n25664) );
  nand_x1_sg U52897 ( .A(n30892), .B(reg_i_8[12]), .X(n25665) );
  nand_x1_sg U52898 ( .A(reg_ii_8[14]), .B(n31736), .X(n25668) );
  nand_x1_sg U52899 ( .A(n34081), .B(reg_i_8[14]), .X(n25669) );
  nand_x1_sg U52900 ( .A(reg_ii_8[15]), .B(n32402), .X(n25670) );
  nand_x1_sg U52901 ( .A(n32725), .B(reg_i_8[15]), .X(n25671) );
  nand_x1_sg U52902 ( .A(reg_ii_8[17]), .B(n31735), .X(n25674) );
  nand_x1_sg U52903 ( .A(n31674), .B(reg_i_8[17]), .X(n25675) );
  nand_x1_sg U52904 ( .A(reg_ii_8[18]), .B(n34898), .X(n25676) );
  nand_x1_sg U52905 ( .A(n35207), .B(reg_i_8[18]), .X(n25677) );
  nand_x1_sg U52906 ( .A(reg_iii_10[0]), .B(n32500), .X(n25044) );
  nand_x1_sg U52907 ( .A(reg_ii_10[0]), .B(n30883), .X(n25045) );
  nand_x1_sg U52908 ( .A(reg_iii_10[1]), .B(n31648), .X(n25046) );
  nand_x1_sg U52909 ( .A(reg_ii_10[1]), .B(n35380), .X(n25047) );
  nand_x1_sg U52910 ( .A(reg_iii_10[3]), .B(n32855), .X(n25050) );
  nand_x1_sg U52911 ( .A(reg_ii_10[3]), .B(n32756), .X(n25051) );
  nand_x1_sg U52912 ( .A(reg_iii_10[4]), .B(n32855), .X(n25052) );
  nand_x1_sg U52913 ( .A(reg_ii_10[4]), .B(n35179), .X(n25053) );
  nand_x1_sg U52914 ( .A(reg_iii_10[6]), .B(n32164), .X(n25056) );
  nand_x1_sg U52915 ( .A(reg_ii_10[6]), .B(n35206), .X(n25057) );
  nand_x1_sg U52916 ( .A(reg_iii_10[7]), .B(n34572), .X(n25058) );
  nand_x1_sg U52917 ( .A(reg_ii_10[7]), .B(n35348), .X(n25059) );
  nand_x1_sg U52918 ( .A(reg_iii_10[9]), .B(n31499), .X(n25062) );
  nand_x1_sg U52919 ( .A(reg_ii_10[9]), .B(n30876), .X(n25063) );
  nand_x1_sg U52920 ( .A(reg_iii_10[10]), .B(n31904), .X(n25064) );
  nand_x1_sg U52921 ( .A(reg_ii_10[10]), .B(n30174), .X(n25065) );
  nand_x1_sg U52922 ( .A(reg_iii_10[12]), .B(n34568), .X(n25068) );
  nand_x1_sg U52923 ( .A(reg_ii_10[12]), .B(n35318), .X(n25069) );
  nand_x1_sg U52924 ( .A(reg_iii_10[13]), .B(n30175), .X(n25070) );
  nand_x1_sg U52925 ( .A(reg_ii_10[13]), .B(n32757), .X(n25071) );
  nand_x1_sg U52926 ( .A(reg_iii_10[15]), .B(n30755), .X(n25074) );
  nand_x1_sg U52927 ( .A(reg_ii_10[15]), .B(n32441), .X(n25075) );
  nand_x1_sg U52928 ( .A(reg_iii_10[16]), .B(n31733), .X(n25076) );
  nand_x1_sg U52929 ( .A(reg_ii_10[16]), .B(n32713), .X(n25077) );
  nand_x1_sg U52930 ( .A(reg_iii_10[18]), .B(n32031), .X(n25080) );
  nand_x1_sg U52931 ( .A(reg_ii_10[18]), .B(n35175), .X(n25081) );
  nand_x1_sg U52932 ( .A(reg_iii_10[19]), .B(n32015), .X(n25082) );
  nand_x1_sg U52933 ( .A(reg_ii_10[19]), .B(n30591), .X(n25083) );
  nand_x1_sg U52934 ( .A(reg_ii_11[1]), .B(n34573), .X(n25086) );
  nand_x1_sg U52935 ( .A(n32749), .B(reg_i_11[1]), .X(n25087) );
  nand_x1_sg U52936 ( .A(reg_ii_11[2]), .B(n33971), .X(n25088) );
  nand_x1_sg U52937 ( .A(n30718), .B(reg_i_11[2]), .X(n25089) );
  nand_x1_sg U52938 ( .A(reg_ii_11[4]), .B(n32360), .X(n25092) );
  nand_x1_sg U52939 ( .A(n35088), .B(reg_i_11[4]), .X(n25093) );
  nand_x1_sg U52940 ( .A(reg_ii_11[5]), .B(n32148), .X(n25094) );
  nand_x1_sg U52941 ( .A(n35089), .B(reg_i_11[5]), .X(n25095) );
  nand_x1_sg U52942 ( .A(reg_ii_11[7]), .B(n32371), .X(n25098) );
  nand_x1_sg U52943 ( .A(n35167), .B(reg_i_11[7]), .X(n25099) );
  nand_x1_sg U52944 ( .A(reg_ii_11[8]), .B(n32252), .X(n25100) );
  nand_x1_sg U52945 ( .A(n32747), .B(reg_i_11[8]), .X(n25101) );
  nand_x1_sg U52946 ( .A(reg_ii_11[10]), .B(n32044), .X(n25104) );
  nand_x1_sg U52947 ( .A(n35333), .B(reg_i_11[10]), .X(n25105) );
  nand_x1_sg U52948 ( .A(reg_iii_13[7]), .B(n34577), .X(n25298) );
  nand_x1_sg U52949 ( .A(reg_ii_13[7]), .B(n30725), .X(n25299) );
  nand_x1_sg U52950 ( .A(reg_iii_13[9]), .B(n32428), .X(n25302) );
  nand_x1_sg U52951 ( .A(reg_ii_13[9]), .B(n30878), .X(n25303) );
  nand_x1_sg U52952 ( .A(reg_iii_13[10]), .B(n34581), .X(n25304) );
  nand_x1_sg U52953 ( .A(reg_ii_13[10]), .B(n30593), .X(n25305) );
  nand_x1_sg U52954 ( .A(reg_iii_13[12]), .B(n32034), .X(n25308) );
  nand_x1_sg U52955 ( .A(reg_ii_13[12]), .B(n34045), .X(n25309) );
  nand_x1_sg U52956 ( .A(reg_iii_13[13]), .B(n32312), .X(n25310) );
  nand_x1_sg U52957 ( .A(reg_ii_13[13]), .B(n32720), .X(n25311) );
  nand_x1_sg U52958 ( .A(reg_iii_13[15]), .B(n31901), .X(n25314) );
  nand_x1_sg U52959 ( .A(reg_ii_13[15]), .B(n30593), .X(n25315) );
  nand_x1_sg U52960 ( .A(reg_iii_13[16]), .B(n32494), .X(n25316) );
  nand_x1_sg U52961 ( .A(reg_ii_13[16]), .B(n30709), .X(n25317) );
  nand_x1_sg U52962 ( .A(reg_iii_13[18]), .B(n32769), .X(n25320) );
  nand_x1_sg U52963 ( .A(reg_ii_13[18]), .B(n35164), .X(n25321) );
  nand_x1_sg U52964 ( .A(reg_iii_13[19]), .B(n30622), .X(n25322) );
  nand_x1_sg U52965 ( .A(reg_ii_13[19]), .B(n35207), .X(n25323) );
  nand_x1_sg U52966 ( .A(reg_iii_14[0]), .B(n31720), .X(n25358) );
  nand_x1_sg U52967 ( .A(reg_ii_14[0]), .B(n32831), .X(n25359) );
  nand_x1_sg U52968 ( .A(reg_ii_14[1]), .B(n32342), .X(n25326) );
  nand_x1_sg U52969 ( .A(n35224), .B(reg_i_14[1]), .X(n25327) );
  nand_x1_sg U52970 ( .A(reg_iii_14[2]), .B(n32044), .X(n25362) );
  nand_x1_sg U52971 ( .A(reg_ii_14[2]), .B(n35333), .X(n25363) );
  nand_x1_sg U52972 ( .A(reg_ii_14[2]), .B(n32776), .X(n25328) );
  nand_x1_sg U52973 ( .A(n32762), .B(reg_i_14[2]), .X(n25329) );
  nand_x1_sg U52974 ( .A(reg_iii_14[3]), .B(n34937), .X(n25364) );
  nand_x1_sg U52975 ( .A(reg_ii_14[3]), .B(n35219), .X(n25365) );
  nand_x1_sg U52976 ( .A(reg_ii_14[4]), .B(n32769), .X(n25332) );
  nand_x1_sg U52977 ( .A(n32737), .B(reg_i_14[4]), .X(n25333) );
  nand_x1_sg U52978 ( .A(reg_iii_14[5]), .B(n35077), .X(n25368) );
  nand_x1_sg U52979 ( .A(reg_ii_14[5]), .B(n32831), .X(n25369) );
  nand_x1_sg U52980 ( .A(reg_ii_14[5]), .B(n32498), .X(n25334) );
  nand_x1_sg U52981 ( .A(n32741), .B(reg_i_14[5]), .X(n25335) );
  nand_x1_sg U52982 ( .A(reg_iii_14[6]), .B(n32405), .X(n25370) );
  nand_x1_sg U52983 ( .A(reg_ii_14[6]), .B(n30865), .X(n25371) );
  nand_x1_sg U52984 ( .A(reg_ii_14[7]), .B(n31497), .X(n25338) );
  nand_x1_sg U52985 ( .A(n35380), .B(reg_i_14[7]), .X(n25339) );
  nand_x1_sg U52986 ( .A(reg_iii_14[8]), .B(n31900), .X(n25374) );
  nand_x1_sg U52987 ( .A(reg_ii_14[8]), .B(n30906), .X(n25375) );
  nand_x1_sg U52988 ( .A(reg_ii_14[8]), .B(n32499), .X(n25340) );
  nand_x1_sg U52989 ( .A(n34056), .B(reg_i_14[8]), .X(n25341) );
  nand_x1_sg U52990 ( .A(reg_iii_14[9]), .B(n32496), .X(n25376) );
  nand_x1_sg U52991 ( .A(reg_ii_14[9]), .B(n32735), .X(n25377) );
  nand_x1_sg U52992 ( .A(reg_ii_14[10]), .B(n31639), .X(n25344) );
  nand_x1_sg U52993 ( .A(n29758), .B(reg_i_14[10]), .X(n25345) );
  nand_x1_sg U52994 ( .A(reg_iii_14[11]), .B(n34581), .X(n25380) );
  nand_x1_sg U52995 ( .A(reg_ii_14[11]), .B(n35222), .X(n25381) );
  nand_x1_sg U52996 ( .A(reg_ii_14[11]), .B(n32498), .X(n25346) );
  nand_x1_sg U52997 ( .A(n35208), .B(reg_i_14[11]), .X(n25347) );
  nand_x1_sg U52998 ( .A(reg_iii_14[12]), .B(n35079), .X(n25382) );
  nand_x1_sg U52999 ( .A(reg_ii_14[12]), .B(n32841), .X(n25383) );
  nand_x1_sg U53000 ( .A(reg_ii_14[13]), .B(n32226), .X(n25350) );
  nand_x1_sg U53001 ( .A(n32766), .B(reg_i_14[13]), .X(n25351) );
  nand_x1_sg U53002 ( .A(reg_iii_14[14]), .B(n31739), .X(n25386) );
  nand_x1_sg U53003 ( .A(reg_ii_14[14]), .B(n30171), .X(n25387) );
  nand_x1_sg U53004 ( .A(reg_ii_14[14]), .B(n32254), .X(n25352) );
  nand_x1_sg U53005 ( .A(n32744), .B(reg_i_14[14]), .X(n25353) );
  nand_x1_sg U53006 ( .A(reg_iii_14[15]), .B(n31910), .X(n25388) );
  nand_x1_sg U53007 ( .A(reg_ii_14[15]), .B(n35165), .X(n25389) );
  nand_x1_sg U53008 ( .A(reg_ii_14[16]), .B(n31637), .X(n25356) );
  nand_x1_sg U53009 ( .A(n31873), .B(reg_i_14[16]), .X(n25357) );
  nand_x1_sg U53010 ( .A(reg_iii_14[17]), .B(n30597), .X(n25392) );
  nand_x1_sg U53011 ( .A(reg_ii_14[17]), .B(n31039), .X(n25393) );
  nand_x1_sg U53012 ( .A(reg_iii_14[18]), .B(n31744), .X(n25394) );
  nand_x1_sg U53013 ( .A(reg_ii_14[18]), .B(n32732), .X(n25395) );
  nand_x1_sg U53014 ( .A(reg_www_0[0]), .B(n34652), .X(n24728) );
  nand_x1_sg U53015 ( .A(reg_ww_0[0]), .B(n30875), .X(n24729) );
  nand_x1_sg U53016 ( .A(reg_www_0[2]), .B(n32450), .X(n24732) );
  nand_x1_sg U53017 ( .A(reg_ww_0[2]), .B(n35321), .X(n24733) );
  nand_x1_sg U53018 ( .A(reg_www_0[3]), .B(n32354), .X(n24734) );
  nand_x1_sg U53019 ( .A(reg_ww_0[3]), .B(n32725), .X(n24735) );
  nand_x1_sg U53020 ( .A(reg_www_0[5]), .B(n34936), .X(n24738) );
  nand_x1_sg U53021 ( .A(reg_ww_0[5]), .B(n35236), .X(n24739) );
  nand_x1_sg U53022 ( .A(reg_www_0[6]), .B(n32237), .X(n24740) );
  nand_x1_sg U53023 ( .A(reg_ww_0[6]), .B(n32716), .X(n24741) );
  nand_x1_sg U53024 ( .A(reg_www_0[8]), .B(n30140), .X(n24744) );
  nand_x1_sg U53025 ( .A(reg_ww_0[8]), .B(n30748), .X(n24745) );
  nand_x1_sg U53026 ( .A(reg_www_0[9]), .B(n32359), .X(n24746) );
  nand_x1_sg U53027 ( .A(reg_ww_0[9]), .B(n30707), .X(n24747) );
  nand_x1_sg U53028 ( .A(reg_www_0[11]), .B(n32012), .X(n24750) );
  nand_x1_sg U53029 ( .A(reg_ww_0[11]), .B(n35208), .X(n24751) );
  nand_x1_sg U53030 ( .A(reg_www_0[12]), .B(n32030), .X(n24752) );
  nand_x1_sg U53031 ( .A(reg_ww_0[12]), .B(n35355), .X(n24753) );
  nand_x1_sg U53032 ( .A(reg_www_0[14]), .B(n31503), .X(n24756) );
  nand_x1_sg U53033 ( .A(reg_ww_0[14]), .B(n35202), .X(n24757) );
  nand_x1_sg U53034 ( .A(reg_www_0[15]), .B(n30198), .X(n24758) );
  nand_x1_sg U53035 ( .A(reg_ww_0[15]), .B(n34713), .X(n24759) );
  nand_x1_sg U53036 ( .A(reg_www_0[17]), .B(n31908), .X(n24762) );
  nand_x1_sg U53037 ( .A(reg_ww_0[17]), .B(n30870), .X(n24763) );
  nand_x1_sg U53038 ( .A(reg_ww_0[17]), .B(n30197), .X(n24722) );
  nand_x1_sg U53039 ( .A(n35207), .B(reg_w_0[17]), .X(n24723) );
  nand_x1_sg U53040 ( .A(reg_www_0[18]), .B(n32770), .X(n24764) );
  nand_x1_sg U53041 ( .A(reg_ww_0[18]), .B(n31206), .X(n24765) );
  nand_x1_sg U53042 ( .A(reg_ww_0[19]), .B(n31900), .X(n24726) );
  nand_x1_sg U53043 ( .A(n34078), .B(reg_w_0[19]), .X(n24727) );
  nand_x1_sg U53044 ( .A(reg_ww_1[0]), .B(n32339), .X(n24768) );
  nand_x1_sg U53045 ( .A(n35236), .B(reg_w_1[0]), .X(n24769) );
  nand_x1_sg U53046 ( .A(reg_www_1[1]), .B(n32454), .X(n24810) );
  nand_x1_sg U53047 ( .A(reg_ww_1[1]), .B(n32764), .X(n24811) );
  nand_x1_sg U53048 ( .A(reg_ww_1[1]), .B(n31729), .X(n24770) );
  nand_x1_sg U53049 ( .A(n32725), .B(reg_w_1[1]), .X(n24771) );
  nand_x1_sg U53050 ( .A(reg_www_1[2]), .B(n32364), .X(n24812) );
  nand_x1_sg U53051 ( .A(reg_ww_1[2]), .B(n30713), .X(n24813) );
  nand_x1_sg U53052 ( .A(reg_ww_1[3]), .B(n32280), .X(n24774) );
  nand_x1_sg U53053 ( .A(n35200), .B(reg_w_1[3]), .X(n24775) );
  nand_x1_sg U53054 ( .A(reg_www_1[4]), .B(n33977), .X(n24816) );
  nand_x1_sg U53055 ( .A(reg_ww_1[4]), .B(n30716), .X(n24817) );
  nand_x1_sg U53056 ( .A(reg_ww_1[4]), .B(n31717), .X(n24776) );
  nand_x1_sg U53057 ( .A(n35169), .B(reg_w_1[4]), .X(n24777) );
  nand_x1_sg U53058 ( .A(reg_www_1[5]), .B(n32143), .X(n24818) );
  nand_x1_sg U53059 ( .A(reg_ww_1[5]), .B(n30729), .X(n24819) );
  nand_x1_sg U53060 ( .A(reg_ww_1[6]), .B(n32352), .X(n24780) );
  nand_x1_sg U53061 ( .A(n34091), .B(reg_w_1[6]), .X(n24781) );
  nand_x1_sg U53062 ( .A(reg_www_1[7]), .B(n30014), .X(n24822) );
  nand_x1_sg U53063 ( .A(reg_ww_1[7]), .B(n35232), .X(n24823) );
  nand_x1_sg U53064 ( .A(reg_ww_1[7]), .B(n32148), .X(n24782) );
  nand_x1_sg U53065 ( .A(n32756), .B(reg_w_1[7]), .X(n24783) );
  nand_x1_sg U53066 ( .A(reg_www_1[8]), .B(n32016), .X(n24824) );
  nand_x1_sg U53067 ( .A(reg_ww_1[8]), .B(n34710), .X(n24825) );
  nand_x1_sg U53068 ( .A(reg_ww_1[9]), .B(n32301), .X(n24786) );
  nand_x1_sg U53069 ( .A(n35368), .B(reg_w_1[9]), .X(n24787) );
  nand_x1_sg U53070 ( .A(reg_www_1[10]), .B(n32501), .X(n24828) );
  nand_x1_sg U53071 ( .A(reg_ww_1[10]), .B(n31056), .X(n24829) );
  nand_x1_sg U53072 ( .A(reg_ww_1[10]), .B(n32379), .X(n24788) );
  nand_x1_sg U53073 ( .A(n29764), .B(reg_w_1[10]), .X(n24789) );
  nand_x1_sg U53074 ( .A(reg_www_1[11]), .B(n32301), .X(n24830) );
  nand_x1_sg U53075 ( .A(reg_ww_1[11]), .B(n35240), .X(n24831) );
  nand_x1_sg U53076 ( .A(reg_ww_1[12]), .B(n31713), .X(n24792) );
  nand_x1_sg U53077 ( .A(n35399), .B(reg_w_1[12]), .X(n24793) );
  nand_x1_sg U53078 ( .A(reg_www_1[13]), .B(n31744), .X(n24834) );
  nand_x1_sg U53079 ( .A(reg_ww_1[13]), .B(n32720), .X(n24835) );
  nand_x1_sg U53080 ( .A(reg_ww_1[13]), .B(n34580), .X(n24794) );
  nand_x1_sg U53081 ( .A(n32716), .B(reg_w_1[13]), .X(n24795) );
  nand_x1_sg U53082 ( .A(reg_www_1[14]), .B(n32032), .X(n24836) );
  nand_x1_sg U53083 ( .A(reg_ww_1[14]), .B(n35239), .X(n24837) );
  nand_x1_sg U53084 ( .A(reg_ww_1[15]), .B(n35080), .X(n24798) );
  nand_x1_sg U53085 ( .A(n35403), .B(reg_w_1[15]), .X(n24799) );
  nand_x1_sg U53086 ( .A(reg_www_1[16]), .B(n32501), .X(n24840) );
  nand_x1_sg U53087 ( .A(reg_ww_1[16]), .B(n32736), .X(n24841) );
  nand_x1_sg U53088 ( .A(reg_ww_1[16]), .B(n32774), .X(n24800) );
  nand_x1_sg U53089 ( .A(n35229), .B(reg_w_1[16]), .X(n24801) );
  nand_x1_sg U53090 ( .A(reg_www_1[17]), .B(n33968), .X(n24842) );
  nand_x1_sg U53091 ( .A(reg_ww_1[17]), .B(n32712), .X(n24843) );
  nand_x1_sg U53092 ( .A(reg_ww_1[18]), .B(n31646), .X(n24804) );
  nand_x1_sg U53093 ( .A(n35230), .B(reg_w_1[18]), .X(n24805) );
  nand_x1_sg U53094 ( .A(reg_www_1[19]), .B(n32363), .X(n24846) );
  nand_x1_sg U53095 ( .A(reg_ww_1[19]), .B(n30722), .X(n24847) );
  nand_x1_sg U53096 ( .A(reg_ww_1[19]), .B(n32020), .X(n24806) );
  nand_x1_sg U53097 ( .A(n31672), .B(reg_w_1[19]), .X(n24807) );
  nand_x1_sg U53098 ( .A(reg_ww_2[0]), .B(n32306), .X(n24848) );
  nand_x1_sg U53099 ( .A(n35355), .B(reg_w_2[0]), .X(n24849) );
  nand_x1_sg U53100 ( .A(reg_ww_3[16]), .B(n32854), .X(n24204) );
  nand_x1_sg U53101 ( .A(n31673), .B(reg_w_3[16]), .X(n24205) );
  nand_x1_sg U53102 ( .A(reg_ww_3[17]), .B(n34583), .X(n24206) );
  nand_x1_sg U53103 ( .A(n32846), .B(reg_w_3[17]), .X(n24207) );
  nand_x1_sg U53104 ( .A(reg_ww_3[19]), .B(n32364), .X(n24210) );
  nand_x1_sg U53105 ( .A(n34097), .B(reg_w_3[19]), .X(n24211) );
  nand_x1_sg U53106 ( .A(reg_www_4[0]), .B(n32345), .X(n24252) );
  nand_x1_sg U53107 ( .A(reg_ww_4[0]), .B(n35081), .X(n24253) );
  nand_x1_sg U53108 ( .A(reg_ww_4[0]), .B(n32030), .X(n24212) );
  nand_x1_sg U53109 ( .A(n35171), .B(reg_w_4[0]), .X(n24213) );
  nand_x1_sg U53110 ( .A(reg_www_4[1]), .B(n32145), .X(n24254) );
  nand_x1_sg U53111 ( .A(reg_ww_4[1]), .B(n35342), .X(n24255) );
  nand_x1_sg U53112 ( .A(reg_ww_4[2]), .B(n29756), .X(n24216) );
  nand_x1_sg U53113 ( .A(n32761), .B(reg_w_4[2]), .X(n24217) );
  nand_x1_sg U53114 ( .A(reg_www_4[3]), .B(n31724), .X(n24258) );
  nand_x1_sg U53115 ( .A(reg_ww_4[3]), .B(n31093), .X(n24259) );
  nand_x1_sg U53116 ( .A(reg_ww_4[3]), .B(n34846), .X(n24218) );
  nand_x1_sg U53117 ( .A(n29765), .B(reg_w_4[3]), .X(n24219) );
  nand_x1_sg U53118 ( .A(reg_www_4[4]), .B(n30149), .X(n24260) );
  nand_x1_sg U53119 ( .A(reg_ww_4[4]), .B(n35183), .X(n24261) );
  nand_x1_sg U53120 ( .A(reg_ww_4[5]), .B(n32285), .X(n24222) );
  nand_x1_sg U53121 ( .A(n35193), .B(reg_w_4[5]), .X(n24223) );
  nand_x1_sg U53122 ( .A(reg_www_4[6]), .B(n32011), .X(n24264) );
  nand_x1_sg U53123 ( .A(reg_ww_4[6]), .B(n35230), .X(n24265) );
  nand_x1_sg U53124 ( .A(reg_ww_4[6]), .B(n32323), .X(n24224) );
  nand_x1_sg U53125 ( .A(n32736), .B(reg_w_4[6]), .X(n24225) );
  nand_x1_sg U53126 ( .A(reg_www_4[7]), .B(n30213), .X(n24266) );
  nand_x1_sg U53127 ( .A(reg_ww_4[7]), .B(n35165), .X(n24267) );
  nand_x1_sg U53128 ( .A(reg_ww_4[8]), .B(n32159), .X(n24228) );
  nand_x1_sg U53129 ( .A(n35182), .B(reg_w_4[8]), .X(n24229) );
  nand_x1_sg U53130 ( .A(reg_www_4[9]), .B(n32310), .X(n24270) );
  nand_x1_sg U53131 ( .A(reg_ww_4[9]), .B(n30892), .X(n24271) );
  nand_x1_sg U53132 ( .A(reg_ww_4[9]), .B(n32360), .X(n24230) );
  nand_x1_sg U53133 ( .A(n35175), .B(reg_w_4[9]), .X(n24231) );
  nand_x1_sg U53134 ( .A(reg_www_4[10]), .B(n32500), .X(n24272) );
  nand_x1_sg U53135 ( .A(reg_ww_4[10]), .B(n32725), .X(n24273) );
  nand_x1_sg U53136 ( .A(reg_ww_4[11]), .B(n32032), .X(n24234) );
  nand_x1_sg U53137 ( .A(n35368), .B(reg_w_4[11]), .X(n24235) );
  nand_x1_sg U53138 ( .A(reg_ww_4[12]), .B(n34847), .X(n24236) );
  nand_x1_sg U53139 ( .A(n34704), .B(reg_w_4[12]), .X(n24237) );
  nand_x1_sg U53140 ( .A(reg_ww_4[14]), .B(n29755), .X(n24240) );
  nand_x1_sg U53141 ( .A(n34711), .B(reg_w_4[14]), .X(n24241) );
  nand_x1_sg U53142 ( .A(reg_ww_4[15]), .B(n31739), .X(n24242) );
  nand_x1_sg U53143 ( .A(n30898), .B(reg_w_4[15]), .X(n24243) );
  nand_x1_sg U53144 ( .A(reg_ww_4[17]), .B(n32290), .X(n24246) );
  nand_x1_sg U53145 ( .A(n35403), .B(reg_w_4[17]), .X(n24247) );
  nand_x1_sg U53146 ( .A(reg_ww_4[18]), .B(n32333), .X(n24248) );
  nand_x1_sg U53147 ( .A(n30179), .B(reg_w_4[18]), .X(n24249) );
  nand_x1_sg U53148 ( .A(reg_www_7[0]), .B(n32306), .X(n24492) );
  nand_x1_sg U53149 ( .A(reg_ww_7[0]), .B(n32441), .X(n24493) );
  nand_x1_sg U53150 ( .A(reg_www_7[1]), .B(n32335), .X(n24494) );
  nand_x1_sg U53151 ( .A(reg_ww_7[1]), .B(n35234), .X(n24495) );
  nand_x1_sg U53152 ( .A(reg_www_7[3]), .B(n31645), .X(n24498) );
  nand_x1_sg U53153 ( .A(reg_ww_7[3]), .B(n32752), .X(n24499) );
  nand_x1_sg U53154 ( .A(reg_www_7[4]), .B(n32014), .X(n24500) );
  nand_x1_sg U53155 ( .A(reg_ww_7[4]), .B(n32719), .X(n24501) );
  nand_x1_sg U53156 ( .A(reg_www_7[6]), .B(n32499), .X(n24504) );
  nand_x1_sg U53157 ( .A(reg_ww_7[6]), .B(n30716), .X(n24505) );
  nand_x1_sg U53158 ( .A(reg_www_7[7]), .B(n34696), .X(n24506) );
  nand_x1_sg U53159 ( .A(reg_ww_7[7]), .B(n30881), .X(n24507) );
  nand_x1_sg U53160 ( .A(reg_ww_7[8]), .B(n31503), .X(n24468) );
  nand_x1_sg U53161 ( .A(n34662), .B(reg_w_7[8]), .X(n24469) );
  nand_x1_sg U53162 ( .A(reg_www_7[9]), .B(n32286), .X(n24510) );
  nand_x1_sg U53163 ( .A(reg_ww_7[9]), .B(n31490), .X(n24511) );
  nand_x1_sg U53164 ( .A(reg_ww_7[9]), .B(n34852), .X(n24470) );
  nand_x1_sg U53165 ( .A(n35162), .B(reg_w_7[9]), .X(n24471) );
  nand_x1_sg U53166 ( .A(reg_www_7[10]), .B(n32229), .X(n24512) );
  nand_x1_sg U53167 ( .A(reg_ww_7[10]), .B(n30172), .X(n24513) );
  nand_x1_sg U53168 ( .A(reg_ww_7[11]), .B(n32253), .X(n24474) );
  nand_x1_sg U53169 ( .A(n35085), .B(reg_w_7[11]), .X(n24475) );
  nand_x1_sg U53170 ( .A(reg_www_7[12]), .B(n32330), .X(n24516) );
  nand_x1_sg U53171 ( .A(reg_ww_7[12]), .B(n35333), .X(n24517) );
  nand_x1_sg U53172 ( .A(reg_ww_7[12]), .B(n30144), .X(n24476) );
  nand_x1_sg U53173 ( .A(n35181), .B(reg_w_7[12]), .X(n24477) );
  nand_x1_sg U53174 ( .A(reg_www_7[13]), .B(n32227), .X(n24518) );
  nand_x1_sg U53175 ( .A(reg_ww_7[13]), .B(n31025), .X(n24519) );
  nand_x1_sg U53176 ( .A(reg_ww_7[14]), .B(n31728), .X(n24480) );
  nand_x1_sg U53177 ( .A(n34703), .B(reg_w_7[14]), .X(n24481) );
  nand_x1_sg U53178 ( .A(reg_www_7[15]), .B(n32403), .X(n24522) );
  nand_x1_sg U53179 ( .A(reg_ww_7[15]), .B(n35204), .X(n24523) );
  nand_x1_sg U53180 ( .A(reg_ww_7[15]), .B(n34653), .X(n24482) );
  nand_x1_sg U53181 ( .A(n34083), .B(reg_w_7[15]), .X(n24483) );
  nand_x1_sg U53182 ( .A(reg_www_7[16]), .B(n31925), .X(n24524) );
  nand_x1_sg U53183 ( .A(reg_ww_7[16]), .B(n30720), .X(n24525) );
  nand_x1_sg U53184 ( .A(reg_ww_7[17]), .B(n30918), .X(n24486) );
  nand_x1_sg U53185 ( .A(n35161), .B(reg_w_7[17]), .X(n24487) );
  nand_x1_sg U53186 ( .A(reg_www_7[18]), .B(n29756), .X(n24528) );
  nand_x1_sg U53187 ( .A(reg_ww_7[18]), .B(n31058), .X(n24529) );
  nand_x1_sg U53188 ( .A(reg_ww_7[18]), .B(n32281), .X(n24488) );
  nand_x1_sg U53189 ( .A(n32765), .B(reg_w_7[18]), .X(n24489) );
  nand_x1_sg U53190 ( .A(reg_www_9[18]), .B(n32297), .X(n23892) );
  nand_x1_sg U53191 ( .A(reg_ww_9[18]), .B(n31207), .X(n23893) );
  nand_x1_sg U53192 ( .A(reg_www_9[19]), .B(n32347), .X(n23894) );
  nand_x1_sg U53193 ( .A(reg_ww_9[19]), .B(n35338), .X(n23895) );
  nand_x1_sg U53194 ( .A(reg_www_10[0]), .B(n32285), .X(n23936) );
  nand_x1_sg U53195 ( .A(reg_ww_10[0]), .B(n30712), .X(n23937) );
  nand_x1_sg U53196 ( .A(reg_ww_10[1]), .B(n32160), .X(n23898) );
  nand_x1_sg U53197 ( .A(n31869), .B(reg_w_10[1]), .X(n23899) );
  nand_x1_sg U53198 ( .A(reg_www_10[2]), .B(n32371), .X(n23940) );
  nand_x1_sg U53199 ( .A(reg_ww_10[2]), .B(n30705), .X(n23941) );
  nand_x1_sg U53200 ( .A(reg_ww_10[2]), .B(n32331), .X(n23900) );
  nand_x1_sg U53201 ( .A(n30906), .B(reg_w_10[2]), .X(n23901) );
  nand_x1_sg U53202 ( .A(reg_www_10[3]), .B(n32156), .X(n23942) );
  nand_x1_sg U53203 ( .A(reg_ww_10[3]), .B(n35329), .X(n23943) );
  nand_x1_sg U53204 ( .A(reg_ww_10[4]), .B(n32046), .X(n23904) );
  nand_x1_sg U53205 ( .A(n33997), .B(reg_w_10[4]), .X(n23905) );
  nand_x1_sg U53206 ( .A(reg_www_10[5]), .B(n31642), .X(n23946) );
  nand_x1_sg U53207 ( .A(reg_ww_10[5]), .B(n35200), .X(n23947) );
  nand_x1_sg U53208 ( .A(reg_ww_10[5]), .B(n32356), .X(n23906) );
  nand_x1_sg U53209 ( .A(n30899), .B(reg_w_10[5]), .X(n23907) );
  nand_x1_sg U53210 ( .A(reg_www_10[6]), .B(n34578), .X(n23948) );
  nand_x1_sg U53211 ( .A(reg_ww_10[6]), .B(n35229), .X(n23949) );
  nand_x1_sg U53212 ( .A(reg_ww_10[7]), .B(n32139), .X(n23910) );
  nand_x1_sg U53213 ( .A(n32839), .B(reg_w_10[7]), .X(n23911) );
  nand_x1_sg U53214 ( .A(reg_www_10[8]), .B(n33953), .X(n23952) );
  nand_x1_sg U53215 ( .A(reg_ww_10[8]), .B(n32839), .X(n23953) );
  nand_x1_sg U53216 ( .A(reg_ww_10[8]), .B(n32327), .X(n23912) );
  nand_x1_sg U53217 ( .A(n32836), .B(reg_w_10[8]), .X(n23913) );
  nand_x1_sg U53218 ( .A(reg_ww_10[10]), .B(n32228), .X(n23916) );
  nand_x1_sg U53219 ( .A(n30729), .B(reg_w_10[10]), .X(n23917) );
  nand_x1_sg U53220 ( .A(reg_ww_10[11]), .B(n32236), .X(n23918) );
  nand_x1_sg U53221 ( .A(n34080), .B(reg_w_10[11]), .X(n23919) );
  nand_x1_sg U53222 ( .A(reg_ww_10[13]), .B(n34568), .X(n23922) );
  nand_x1_sg U53223 ( .A(n32729), .B(reg_w_10[13]), .X(n23923) );
  nand_x1_sg U53224 ( .A(reg_ww_10[14]), .B(n34553), .X(n23924) );
  nand_x1_sg U53225 ( .A(n32708), .B(reg_w_10[14]), .X(n23925) );
  nand_x1_sg U53226 ( .A(reg_ww_10[16]), .B(n34573), .X(n23928) );
  nand_x1_sg U53227 ( .A(n34051), .B(reg_w_10[16]), .X(n23929) );
  nand_x1_sg U53228 ( .A(reg_ww_10[17]), .B(n31732), .X(n23930) );
  nand_x1_sg U53229 ( .A(n35362), .B(reg_w_10[17]), .X(n23931) );
  nand_x1_sg U53230 ( .A(reg_ww_10[19]), .B(n32046), .X(n23934) );
  nand_x1_sg U53231 ( .A(n35164), .B(reg_w_10[19]), .X(n23935) );
  nand_x1_sg U53232 ( .A(reg_www_13[0]), .B(n32298), .X(n24164) );
  nand_x1_sg U53233 ( .A(reg_ww_13[0]), .B(n35195), .X(n24165) );
  nand_x1_sg U53234 ( .A(reg_www_13[2]), .B(n30145), .X(n24168) );
  nand_x1_sg U53235 ( .A(reg_ww_13[2]), .B(n35353), .X(n24169) );
  nand_x1_sg U53236 ( .A(reg_www_13[3]), .B(n32138), .X(n24170) );
  nand_x1_sg U53237 ( .A(reg_ww_13[3]), .B(n35086), .X(n24171) );
  nand_x1_sg U53238 ( .A(reg_www_13[5]), .B(n31735), .X(n24174) );
  nand_x1_sg U53239 ( .A(reg_ww_13[5]), .B(n31060), .X(n24175) );
  nand_x1_sg U53240 ( .A(reg_ww_13[5]), .B(n34565), .X(n24146) );
  nand_x1_sg U53241 ( .A(n35317), .B(reg_w_13[5]), .X(n24147) );
  nand_x1_sg U53242 ( .A(reg_www_13[6]), .B(n32337), .X(n24176) );
  nand_x1_sg U53243 ( .A(reg_ww_13[6]), .B(n35169), .X(n24177) );
  nand_x1_sg U53244 ( .A(reg_ww_13[7]), .B(n32226), .X(n24150) );
  nand_x1_sg U53245 ( .A(n30587), .B(reg_w_13[7]), .X(n24151) );
  nand_x1_sg U53246 ( .A(reg_www_13[8]), .B(n33952), .X(n24180) );
  nand_x1_sg U53247 ( .A(reg_ww_13[8]), .B(n30864), .X(n24181) );
  nand_x1_sg U53248 ( .A(reg_ww_13[8]), .B(n32253), .X(n24152) );
  nand_x1_sg U53249 ( .A(n30037), .B(reg_w_13[8]), .X(n24153) );
  nand_x1_sg U53250 ( .A(reg_www_13[9]), .B(n32161), .X(n24182) );
  nand_x1_sg U53251 ( .A(reg_ww_13[9]), .B(n32748), .X(n24183) );
  nand_x1_sg U53252 ( .A(reg_ww_13[10]), .B(n32146), .X(n24156) );
  nand_x1_sg U53253 ( .A(n34667), .B(reg_w_13[10]), .X(n24157) );
  nand_x1_sg U53254 ( .A(reg_www_13[11]), .B(n34650), .X(n24186) );
  nand_x1_sg U53255 ( .A(reg_ww_13[11]), .B(n30869), .X(n24187) );
  nand_x1_sg U53256 ( .A(reg_ww_13[11]), .B(n32037), .X(n24158) );
  nand_x1_sg U53257 ( .A(n35398), .B(reg_w_13[11]), .X(n24159) );
  nand_x1_sg U53258 ( .A(reg_www_13[12]), .B(n32405), .X(n24188) );
  nand_x1_sg U53259 ( .A(reg_ww_13[12]), .B(n35209), .X(n24189) );
  nand_x1_sg U53260 ( .A(reg_ww_13[13]), .B(n32244), .X(n24162) );
  nand_x1_sg U53261 ( .A(n32745), .B(reg_w_13[13]), .X(n24163) );
  nand_x1_sg U53262 ( .A(reg_www_13[14]), .B(n34898), .X(n24192) );
  nand_x1_sg U53263 ( .A(reg_ww_13[14]), .B(n31054), .X(n24193) );
  nand_x1_sg U53264 ( .A(reg_ww_13[14]), .B(n31926), .X(n23633) );
  nand_x1_sg U53265 ( .A(n34711), .B(reg_w_13[14]), .X(n23634) );
  nand_x1_sg U53266 ( .A(reg_www_13[15]), .B(n32251), .X(n24194) );
  nand_x1_sg U53267 ( .A(reg_ww_13[15]), .B(n35179), .X(n24195) );
  nand_x1_sg U53268 ( .A(reg_ww_13[15]), .B(n31639), .X(n23636) );
  nand_x1_sg U53269 ( .A(n31869), .B(reg_w_13[15]), .X(n23637) );
  nand_x1_sg U53270 ( .A(reg_www_13[17]), .B(n32139), .X(n24198) );
  nand_x1_sg U53271 ( .A(reg_ww_13[17]), .B(n35194), .X(n24199) );
  nand_x1_sg U53272 ( .A(reg_ww_13[17]), .B(n32049), .X(n23640) );
  nand_x1_sg U53273 ( .A(n34046), .B(reg_w_13[17]), .X(n23641) );
  nand_x1_sg U53274 ( .A(reg_www_13[18]), .B(n31897), .X(n24200) );
  nand_x1_sg U53275 ( .A(reg_ww_13[18]), .B(n30725), .X(n24201) );
  nand_x1_sg U53276 ( .A(reg_ww_13[18]), .B(n32143), .X(n23642) );
  nand_x1_sg U53277 ( .A(n31870), .B(reg_w_13[18]), .X(n23643) );
  nand_x1_sg U53278 ( .A(reg_ww_14[0]), .B(n32241), .X(n23646) );
  nand_x1_sg U53279 ( .A(n34723), .B(reg_w_14[0]), .X(n23647) );
  nand_x1_sg U53280 ( .A(reg_www_14[1]), .B(n32143), .X(n23688) );
  nand_x1_sg U53281 ( .A(reg_ww_14[1]), .B(n30883), .X(n23689) );
  nand_x1_sg U53282 ( .A(reg_ww_14[1]), .B(n32031), .X(n23648) );
  nand_x1_sg U53283 ( .A(n33999), .B(reg_w_14[1]), .X(n23649) );
  nand_x1_sg U53284 ( .A(reg_www_14[2]), .B(n31909), .X(n23690) );
  nand_x1_sg U53285 ( .A(reg_ww_14[2]), .B(n32767), .X(n23691) );
  nand_x1_sg U53286 ( .A(reg_ww_14[3]), .B(n31717), .X(n23652) );
  nand_x1_sg U53287 ( .A(n34092), .B(reg_w_14[3]), .X(n23653) );
  nand_x1_sg U53288 ( .A(reg_www_14[4]), .B(n33952), .X(n23694) );
  nand_x1_sg U53289 ( .A(reg_ww_14[4]), .B(n30711), .X(n23695) );
  nand_x1_sg U53290 ( .A(reg_ww_14[4]), .B(n32018), .X(n23654) );
  nand_x1_sg U53291 ( .A(n35187), .B(reg_w_14[4]), .X(n23655) );
  nand_x1_sg U53292 ( .A(reg_www_14[5]), .B(n32238), .X(n23696) );
  nand_x1_sg U53293 ( .A(reg_ww_14[5]), .B(n30716), .X(n23697) );
  nand_x1_sg U53294 ( .A(reg_ww_14[6]), .B(n31731), .X(n23658) );
  nand_x1_sg U53295 ( .A(n35202), .B(reg_w_14[6]), .X(n23659) );
  nand_x1_sg U53296 ( .A(reg_ww_14[7]), .B(n31511), .X(n23660) );
  nand_x1_sg U53297 ( .A(n32754), .B(reg_w_14[7]), .X(n23661) );
  nand_x1_sg U53298 ( .A(reg_ww_14[9]), .B(n32237), .X(n23664) );
  nand_x1_sg U53299 ( .A(n32740), .B(reg_w_14[9]), .X(n23665) );
  nand_x1_sg U53300 ( .A(reg_ww_14[10]), .B(n32217), .X(n23666) );
  nand_x1_sg U53301 ( .A(n35201), .B(reg_w_14[10]), .X(n23667) );
  nand_x1_sg U53302 ( .A(reg_ww_14[12]), .B(n32322), .X(n23670) );
  nand_x1_sg U53303 ( .A(n34665), .B(reg_w_14[12]), .X(n23671) );
  nand_x1_sg U53304 ( .A(reg_ww_14[13]), .B(n34849), .X(n23672) );
  nand_x1_sg U53305 ( .A(n35171), .B(reg_w_14[13]), .X(n23673) );
  nand_x1_sg U53306 ( .A(reg_ww_14[15]), .B(n32301), .X(n23676) );
  nand_x1_sg U53307 ( .A(n34699), .B(reg_w_14[15]), .X(n23677) );
  nand_x1_sg U53308 ( .A(reg_ww_14[16]), .B(n32249), .X(n23678) );
  nand_x1_sg U53309 ( .A(n34699), .B(reg_w_14[16]), .X(n23679) );
  nand_x1_sg U53310 ( .A(reg_ww_14[18]), .B(n32331), .X(n23682) );
  nand_x1_sg U53311 ( .A(n32747), .B(reg_w_14[18]), .X(n23683) );
  nand_x1_sg U53312 ( .A(reg_ww_14[19]), .B(n32285), .X(n23684) );
  nand_x1_sg U53313 ( .A(n32735), .B(reg_w_14[19]), .X(n23685) );
  nand_x1_sg U53314 ( .A(reg_ii_1[0]), .B(n35080), .X(n25876) );
  nand_x1_sg U53315 ( .A(n35086), .B(reg_i_1[0]), .X(n25877) );
  nand_x1_sg U53316 ( .A(reg_iii_1[1]), .B(n30920), .X(n25918) );
  nand_x1_sg U53317 ( .A(reg_ii_1[1]), .B(n35186), .X(n25919) );
  nand_x1_sg U53318 ( .A(reg_ii_1[3]), .B(n32292), .X(n25882) );
  nand_x1_sg U53319 ( .A(n32765), .B(reg_i_1[3]), .X(n25883) );
  nand_x1_sg U53320 ( .A(reg_iii_1[4]), .B(n34651), .X(n25924) );
  nand_x1_sg U53321 ( .A(reg_ii_1[4]), .B(n35330), .X(n25925) );
  nand_x1_sg U53322 ( .A(reg_ii_1[6]), .B(n32247), .X(n25888) );
  nand_x1_sg U53323 ( .A(n30717), .B(reg_i_1[6]), .X(n25889) );
  nand_x1_sg U53324 ( .A(reg_iii_1[7]), .B(n31511), .X(n25930) );
  nand_x1_sg U53325 ( .A(reg_ii_1[7]), .B(n35345), .X(n25931) );
  nand_x1_sg U53326 ( .A(reg_ii_1[9]), .B(n32150), .X(n25894) );
  nand_x1_sg U53327 ( .A(n35348), .B(reg_i_1[9]), .X(n25895) );
  nand_x1_sg U53328 ( .A(reg_iii_1[10]), .B(n34846), .X(n25936) );
  nand_x1_sg U53329 ( .A(reg_ii_1[10]), .B(n31033), .X(n25937) );
  nand_x1_sg U53330 ( .A(reg_ii_1[12]), .B(n30153), .X(n25900) );
  nand_x1_sg U53331 ( .A(n31872), .B(reg_i_1[12]), .X(n25901) );
  nand_x1_sg U53332 ( .A(reg_iii_1[13]), .B(n33946), .X(n25942) );
  nand_x1_sg U53333 ( .A(reg_ii_1[13]), .B(n32844), .X(n25943) );
  nand_x1_sg U53334 ( .A(reg_ii_1[15]), .B(n30169), .X(n25906) );
  nand_x1_sg U53335 ( .A(n34091), .B(reg_i_1[15]), .X(n25907) );
  nand_x1_sg U53336 ( .A(reg_iii_1[16]), .B(n32361), .X(n25948) );
  nand_x1_sg U53337 ( .A(reg_ii_1[16]), .B(n35205), .X(n25949) );
  nand_x1_sg U53338 ( .A(reg_ii_1[18]), .B(n31719), .X(n25912) );
  nand_x1_sg U53339 ( .A(n32750), .B(reg_i_1[18]), .X(n25913) );
  nand_x1_sg U53340 ( .A(reg_iii_1[19]), .B(n30754), .X(n25954) );
  nand_x1_sg U53341 ( .A(reg_ii_1[19]), .B(n31039), .X(n25955) );
  nand_x1_sg U53342 ( .A(reg_iii_2[0]), .B(n32772), .X(n25996) );
  nand_x1_sg U53343 ( .A(reg_ii_2[0]), .B(n30864), .X(n25997) );
  nand_x1_sg U53344 ( .A(reg_ii_2[2]), .B(n31905), .X(n25960) );
  nand_x1_sg U53345 ( .A(n32718), .B(reg_i_2[2]), .X(n25961) );
  nand_x1_sg U53346 ( .A(reg_ii_2[5]), .B(n32350), .X(n25966) );
  nand_x1_sg U53347 ( .A(n35338), .B(reg_i_2[5]), .X(n25967) );
  nand_x1_sg U53348 ( .A(reg_ii_2[8]), .B(n32777), .X(n25972) );
  nand_x1_sg U53349 ( .A(n32847), .B(reg_i_2[8]), .X(n25973) );
  nand_x1_sg U53350 ( .A(reg_ii_2[11]), .B(n32351), .X(n25978) );
  nand_x1_sg U53351 ( .A(n31865), .B(reg_i_2[11]), .X(n25979) );
  nand_x1_sg U53352 ( .A(reg_ii_2[14]), .B(n31910), .X(n25984) );
  nand_x1_sg U53353 ( .A(n32762), .B(reg_i_2[14]), .X(n25985) );
  nand_x1_sg U53354 ( .A(reg_ii_2[17]), .B(n32153), .X(n25990) );
  nand_x1_sg U53355 ( .A(n31870), .B(reg_i_2[17]), .X(n25991) );
  nand_x1_sg U53356 ( .A(reg_ii_5[1]), .B(n32402), .X(n25402) );
  nand_x1_sg U53357 ( .A(n30592), .B(reg_i_5[1]), .X(n25403) );
  nand_x1_sg U53358 ( .A(reg_ii_5[4]), .B(n32041), .X(n25408) );
  nand_x1_sg U53359 ( .A(n32743), .B(reg_i_5[4]), .X(n25409) );
  nand_x1_sg U53360 ( .A(reg_ii_5[7]), .B(n31723), .X(n25414) );
  nand_x1_sg U53361 ( .A(n31675), .B(reg_i_5[7]), .X(n25415) );
  nand_x1_sg U53362 ( .A(reg_ii_5[10]), .B(n32246), .X(n25420) );
  nand_x1_sg U53363 ( .A(n30172), .B(reg_i_5[10]), .X(n25421) );
  nand_x1_sg U53364 ( .A(reg_iii_7[9]), .B(n33967), .X(n25618) );
  nand_x1_sg U53365 ( .A(reg_ii_7[9]), .B(n32829), .X(n25619) );
  nand_x1_sg U53366 ( .A(reg_iii_7[12]), .B(n32253), .X(n25624) );
  nand_x1_sg U53367 ( .A(reg_ii_7[12]), .B(n35167), .X(n25625) );
  nand_x1_sg U53368 ( .A(reg_iii_7[15]), .B(n34893), .X(n25630) );
  nand_x1_sg U53369 ( .A(reg_ii_7[15]), .B(n35216), .X(n25631) );
  nand_x1_sg U53370 ( .A(reg_iii_7[18]), .B(n32317), .X(n25636) );
  nand_x1_sg U53371 ( .A(reg_ii_7[18]), .B(n35212), .X(n25637) );
  nand_x1_sg U53372 ( .A(reg_ii_8[1]), .B(n32143), .X(n25642) );
  nand_x1_sg U53373 ( .A(n35175), .B(reg_i_8[1]), .X(n25643) );
  nand_x1_sg U53374 ( .A(reg_ii_8[4]), .B(n31499), .X(n25648) );
  nand_x1_sg U53375 ( .A(n34702), .B(reg_i_8[4]), .X(n25649) );
  nand_x1_sg U53376 ( .A(reg_ii_8[7]), .B(n32291), .X(n25654) );
  nand_x1_sg U53377 ( .A(n32742), .B(reg_i_8[7]), .X(n25655) );
  nand_x1_sg U53378 ( .A(reg_ii_8[10]), .B(n31640), .X(n25660) );
  nand_x1_sg U53379 ( .A(n32736), .B(reg_i_8[10]), .X(n25661) );
  nand_x1_sg U53380 ( .A(reg_ii_8[13]), .B(n32355), .X(n25666) );
  nand_x1_sg U53381 ( .A(n35353), .B(reg_i_8[13]), .X(n25667) );
  nand_x1_sg U53382 ( .A(reg_ii_8[16]), .B(n32350), .X(n25672) );
  nand_x1_sg U53383 ( .A(n30180), .B(reg_i_8[16]), .X(n25673) );
  nand_x1_sg U53384 ( .A(reg_ii_8[19]), .B(n32286), .X(n25678) );
  nand_x1_sg U53385 ( .A(n34057), .B(reg_i_8[19]), .X(n25679) );
  nand_x1_sg U53386 ( .A(reg_iii_10[2]), .B(n30599), .X(n25048) );
  nand_x1_sg U53387 ( .A(reg_ii_10[2]), .B(n30720), .X(n25049) );
  nand_x1_sg U53388 ( .A(reg_iii_10[5]), .B(n31634), .X(n25054) );
  nand_x1_sg U53389 ( .A(reg_ii_10[5]), .B(n31206), .X(n25055) );
  nand_x1_sg U53390 ( .A(reg_iii_10[8]), .B(n32338), .X(n25060) );
  nand_x1_sg U53391 ( .A(reg_ii_10[8]), .B(n35379), .X(n25061) );
  nand_x1_sg U53392 ( .A(reg_iii_10[11]), .B(n31925), .X(n25066) );
  nand_x1_sg U53393 ( .A(reg_ii_10[11]), .B(n30895), .X(n25067) );
  nand_x1_sg U53394 ( .A(reg_iii_10[14]), .B(n34698), .X(n25072) );
  nand_x1_sg U53395 ( .A(reg_ii_10[14]), .B(n35361), .X(n25073) );
  nand_x1_sg U53396 ( .A(reg_iii_10[17]), .B(n32384), .X(n25078) );
  nand_x1_sg U53397 ( .A(reg_ii_10[17]), .B(n35399), .X(n25079) );
  nand_x1_sg U53398 ( .A(reg_ii_10[19]), .B(n32453), .X(n25042) );
  nand_x1_sg U53399 ( .A(n31864), .B(reg_i_10[19]), .X(n25043) );
  nand_x1_sg U53400 ( .A(reg_ii_11[0]), .B(n32146), .X(n25084) );
  nand_x1_sg U53401 ( .A(n32759), .B(reg_i_11[0]), .X(n25085) );
  nand_x1_sg U53402 ( .A(reg_ii_11[3]), .B(n32028), .X(n25090) );
  nand_x1_sg U53403 ( .A(n34084), .B(reg_i_11[3]), .X(n25091) );
  nand_x1_sg U53404 ( .A(reg_ii_11[6]), .B(n34565), .X(n25096) );
  nand_x1_sg U53405 ( .A(n32757), .B(reg_i_11[6]), .X(n25097) );
  nand_x1_sg U53406 ( .A(reg_ii_11[9]), .B(n31893), .X(n25102) );
  nand_x1_sg U53407 ( .A(n32738), .B(reg_i_11[9]), .X(n25103) );
  nand_x1_sg U53408 ( .A(reg_iii_13[8]), .B(n34578), .X(n25300) );
  nand_x1_sg U53409 ( .A(reg_ii_13[8]), .B(n30589), .X(n25301) );
  nand_x1_sg U53410 ( .A(reg_iii_13[11]), .B(n32293), .X(n25306) );
  nand_x1_sg U53411 ( .A(reg_ii_13[11]), .B(n32766), .X(n25307) );
  nand_x1_sg U53412 ( .A(reg_iii_13[14]), .B(n34846), .X(n25312) );
  nand_x1_sg U53413 ( .A(reg_ii_13[14]), .B(n35203), .X(n25313) );
  nand_x1_sg U53414 ( .A(reg_iii_13[17]), .B(n32144), .X(n25318) );
  nand_x1_sg U53415 ( .A(reg_ii_13[17]), .B(n30876), .X(n25319) );
  nand_x1_sg U53416 ( .A(reg_ii_14[0]), .B(n32373), .X(n25324) );
  nand_x1_sg U53417 ( .A(n35358), .B(reg_i_14[0]), .X(n25325) );
  nand_x1_sg U53418 ( .A(reg_iii_14[1]), .B(n31716), .X(n25360) );
  nand_x1_sg U53419 ( .A(reg_ii_14[1]), .B(n32841), .X(n25361) );
  nand_x1_sg U53420 ( .A(reg_ii_14[3]), .B(n31509), .X(n25330) );
  nand_x1_sg U53421 ( .A(n32745), .B(reg_i_14[3]), .X(n25331) );
  nand_x1_sg U53422 ( .A(reg_iii_14[4]), .B(n32351), .X(n25366) );
  nand_x1_sg U53423 ( .A(reg_ii_14[4]), .B(n30591), .X(n25367) );
  nand_x1_sg U53424 ( .A(reg_ii_14[6]), .B(n34894), .X(n25336) );
  nand_x1_sg U53425 ( .A(n35225), .B(reg_i_14[6]), .X(n25337) );
  nand_x1_sg U53426 ( .A(reg_iii_14[7]), .B(n32343), .X(n25372) );
  nand_x1_sg U53427 ( .A(reg_ii_14[7]), .B(n29763), .X(n25373) );
  nand_x1_sg U53428 ( .A(reg_ii_14[9]), .B(n31890), .X(n25342) );
  nand_x1_sg U53429 ( .A(n32842), .B(reg_i_14[9]), .X(n25343) );
  nand_x1_sg U53430 ( .A(reg_iii_14[10]), .B(n34896), .X(n25378) );
  nand_x1_sg U53431 ( .A(reg_ii_14[10]), .B(n30861), .X(n25379) );
  nand_x1_sg U53432 ( .A(reg_ii_14[12]), .B(n32163), .X(n25348) );
  nand_x1_sg U53433 ( .A(n35086), .B(reg_i_14[12]), .X(n25349) );
  nand_x1_sg U53434 ( .A(reg_iii_14[13]), .B(n32493), .X(n25384) );
  nand_x1_sg U53435 ( .A(reg_ii_14[13]), .B(n32836), .X(n25385) );
  nand_x1_sg U53436 ( .A(reg_ii_14[15]), .B(n32153), .X(n25354) );
  nand_x1_sg U53437 ( .A(n30178), .B(reg_i_14[15]), .X(n25355) );
  nand_x1_sg U53438 ( .A(reg_iii_14[16]), .B(n32217), .X(n25390) );
  nand_x1_sg U53439 ( .A(reg_ii_14[16]), .B(n31033), .X(n25391) );
  nand_x1_sg U53440 ( .A(reg_iii_14[19]), .B(n32774), .X(n25396) );
  nand_x1_sg U53441 ( .A(reg_ii_14[19]), .B(n32836), .X(n25397) );
  nand_x1_sg U53442 ( .A(reg_www_0[1]), .B(n31741), .X(n24730) );
  nand_x1_sg U53443 ( .A(reg_ww_0[1]), .B(n30883), .X(n24731) );
  nand_x1_sg U53444 ( .A(reg_www_0[4]), .B(n31712), .X(n24736) );
  nand_x1_sg U53445 ( .A(reg_ww_0[4]), .B(n35358), .X(n24737) );
  nand_x1_sg U53446 ( .A(reg_www_0[7]), .B(n31640), .X(n24742) );
  nand_x1_sg U53447 ( .A(reg_ww_0[7]), .B(n32744), .X(n24743) );
  nand_x1_sg U53448 ( .A(reg_www_0[10]), .B(n32160), .X(n24748) );
  nand_x1_sg U53449 ( .A(reg_ww_0[10]), .B(n31492), .X(n24749) );
  nand_x1_sg U53450 ( .A(reg_www_0[13]), .B(n34580), .X(n24754) );
  nand_x1_sg U53451 ( .A(reg_ww_0[13]), .B(n35220), .X(n24755) );
  nand_x1_sg U53452 ( .A(reg_www_0[16]), .B(n31648), .X(n24760) );
  nand_x1_sg U53453 ( .A(reg_ww_0[16]), .B(n31207), .X(n24761) );
  nand_x1_sg U53454 ( .A(reg_ww_0[18]), .B(n31715), .X(n24724) );
  nand_x1_sg U53455 ( .A(n34082), .B(reg_w_0[18]), .X(n24725) );
  nand_x1_sg U53456 ( .A(reg_www_0[19]), .B(n35277), .X(n24766) );
  nand_x1_sg U53457 ( .A(reg_ww_0[19]), .B(n35348), .X(n24767) );
  nand_x1_sg U53458 ( .A(reg_www_1[0]), .B(n34572), .X(n24808) );
  nand_x1_sg U53459 ( .A(reg_ww_1[0]), .B(n30705), .X(n24809) );
  nand_x1_sg U53460 ( .A(reg_ww_1[2]), .B(n32298), .X(n24772) );
  nand_x1_sg U53461 ( .A(n34084), .B(reg_w_1[2]), .X(n24773) );
  nand_x1_sg U53462 ( .A(reg_www_1[3]), .B(n30920), .X(n24814) );
  nand_x1_sg U53463 ( .A(reg_ww_1[3]), .B(n30592), .X(n24815) );
  nand_x1_sg U53464 ( .A(reg_ww_1[5]), .B(n32372), .X(n24778) );
  nand_x1_sg U53465 ( .A(n35181), .B(reg_w_1[5]), .X(n24779) );
  nand_x1_sg U53466 ( .A(reg_www_1[6]), .B(n34895), .X(n24820) );
  nand_x1_sg U53467 ( .A(reg_ww_1[6]), .B(n34719), .X(n24821) );
  nand_x1_sg U53468 ( .A(reg_ww_1[8]), .B(n31892), .X(n24784) );
  nand_x1_sg U53469 ( .A(n32749), .B(reg_w_1[8]), .X(n24785) );
  nand_x1_sg U53470 ( .A(reg_www_1[9]), .B(n30151), .X(n24826) );
  nand_x1_sg U53471 ( .A(reg_ww_1[9]), .B(n32830), .X(n24827) );
  nand_x1_sg U53472 ( .A(reg_ww_1[11]), .B(n34897), .X(n24790) );
  nand_x1_sg U53473 ( .A(n34046), .B(reg_w_1[11]), .X(n24791) );
  nand_x1_sg U53474 ( .A(reg_www_1[12]), .B(n31513), .X(n24832) );
  nand_x1_sg U53475 ( .A(reg_ww_1[12]), .B(n35204), .X(n24833) );
  nand_x1_sg U53476 ( .A(reg_ww_1[14]), .B(n32238), .X(n24796) );
  nand_x1_sg U53477 ( .A(n34058), .B(reg_w_1[14]), .X(n24797) );
  nand_x1_sg U53478 ( .A(reg_www_1[15]), .B(n32154), .X(n24838) );
  nand_x1_sg U53479 ( .A(reg_ww_1[15]), .B(n30903), .X(n24839) );
  nand_x1_sg U53480 ( .A(reg_ww_1[17]), .B(n30597), .X(n24802) );
  nand_x1_sg U53481 ( .A(n30024), .B(reg_w_1[17]), .X(n24803) );
  nand_x1_sg U53482 ( .A(reg_www_1[18]), .B(n32050), .X(n24844) );
  nand_x1_sg U53483 ( .A(reg_ww_1[18]), .B(n32830), .X(n24845) );
  nand_x1_sg U53484 ( .A(reg_ww_3[18]), .B(n32140), .X(n24208) );
  nand_x1_sg U53485 ( .A(n32830), .B(reg_w_3[18]), .X(n24209) );
  nand_x1_sg U53486 ( .A(reg_ww_4[1]), .B(n34573), .X(n24214) );
  nand_x1_sg U53487 ( .A(n35173), .B(reg_w_4[1]), .X(n24215) );
  nand_x1_sg U53488 ( .A(reg_www_4[2]), .B(n32037), .X(n24256) );
  nand_x1_sg U53489 ( .A(reg_ww_4[2]), .B(n31094), .X(n24257) );
  nand_x1_sg U53490 ( .A(reg_ww_4[4]), .B(n32428), .X(n24220) );
  nand_x1_sg U53491 ( .A(n35404), .B(reg_w_4[4]), .X(n24221) );
  nand_x1_sg U53492 ( .A(reg_www_4[5]), .B(n32291), .X(n24262) );
  nand_x1_sg U53493 ( .A(reg_ww_4[5]), .B(n35335), .X(n24263) );
  nand_x1_sg U53494 ( .A(reg_ww_4[7]), .B(n32296), .X(n24226) );
  nand_x1_sg U53495 ( .A(n34048), .B(reg_w_4[7]), .X(n24227) );
  nand_x1_sg U53496 ( .A(reg_www_4[8]), .B(n31736), .X(n24268) );
  nand_x1_sg U53497 ( .A(reg_ww_4[8]), .B(n30727), .X(n24269) );
  nand_x1_sg U53498 ( .A(reg_ww_4[10]), .B(n31894), .X(n24232) );
  nand_x1_sg U53499 ( .A(n34083), .B(reg_w_4[10]), .X(n24233) );
  nand_x1_sg U53500 ( .A(reg_ww_4[13]), .B(n33968), .X(n24238) );
  nand_x1_sg U53501 ( .A(n34706), .B(reg_w_4[13]), .X(n24239) );
  nand_x1_sg U53502 ( .A(reg_ww_4[16]), .B(n32500), .X(n24244) );
  nand_x1_sg U53503 ( .A(n34714), .B(reg_w_4[16]), .X(n24245) );
  nand_x1_sg U53504 ( .A(reg_ww_4[19]), .B(n32011), .X(n24250) );
  nand_x1_sg U53505 ( .A(n34717), .B(reg_w_4[19]), .X(n24251) );
  nand_x1_sg U53506 ( .A(reg_www_7[2]), .B(n31636), .X(n24496) );
  nand_x1_sg U53507 ( .A(reg_ww_7[2]), .B(n35194), .X(n24497) );
  nand_x1_sg U53508 ( .A(reg_www_7[5]), .B(n32380), .X(n24502) );
  nand_x1_sg U53509 ( .A(reg_ww_7[5]), .B(n35347), .X(n24503) );
  nand_x1_sg U53510 ( .A(reg_ww_7[7]), .B(n31648), .X(n24466) );
  nand_x1_sg U53511 ( .A(n35091), .B(reg_w_7[7]), .X(n24467) );
  nand_x1_sg U53512 ( .A(reg_www_7[8]), .B(n32027), .X(n24508) );
  nand_x1_sg U53513 ( .A(reg_ww_7[8]), .B(n32743), .X(n24509) );
  nand_x1_sg U53514 ( .A(reg_ww_7[10]), .B(n33950), .X(n24472) );
  nand_x1_sg U53515 ( .A(n32831), .B(reg_w_7[10]), .X(n24473) );
  nand_x1_sg U53516 ( .A(reg_www_7[11]), .B(n34651), .X(n24514) );
  nand_x1_sg U53517 ( .A(reg_ww_7[11]), .B(n30898), .X(n24515) );
  nand_x1_sg U53518 ( .A(reg_ww_7[13]), .B(n30730), .X(n24478) );
  nand_x1_sg U53519 ( .A(n31863), .B(reg_w_7[13]), .X(n24479) );
  nand_x1_sg U53520 ( .A(reg_www_7[14]), .B(n32771), .X(n24520) );
  nand_x1_sg U53521 ( .A(reg_ww_7[14]), .B(n35342), .X(n24521) );
  nand_x1_sg U53522 ( .A(reg_ww_7[16]), .B(n31727), .X(n24484) );
  nand_x1_sg U53523 ( .A(n34096), .B(reg_w_7[16]), .X(n24485) );
  nand_x1_sg U53524 ( .A(reg_www_7[17]), .B(n32038), .X(n24526) );
  nand_x1_sg U53525 ( .A(reg_ww_7[17]), .B(n30588), .X(n24527) );
  nand_x1_sg U53526 ( .A(reg_ww_7[19]), .B(n32347), .X(n24490) );
  nand_x1_sg U53527 ( .A(n32748), .B(reg_w_7[19]), .X(n24491) );
  nand_x1_sg U53528 ( .A(reg_www_9[17]), .B(n32214), .X(n23890) );
  nand_x1_sg U53529 ( .A(reg_ww_9[17]), .B(n30875), .X(n23891) );
  nand_x1_sg U53530 ( .A(reg_ww_10[0]), .B(n31888), .X(n23896) );
  nand_x1_sg U53531 ( .A(n32737), .B(reg_w_10[0]), .X(n23897) );
  nand_x1_sg U53532 ( .A(reg_www_10[1]), .B(n32243), .X(n23938) );
  nand_x1_sg U53533 ( .A(reg_ww_10[1]), .B(n32766), .X(n23939) );
  nand_x1_sg U53534 ( .A(reg_ww_10[3]), .B(n32499), .X(n23902) );
  nand_x1_sg U53535 ( .A(n35318), .B(reg_w_10[3]), .X(n23903) );
  nand_x1_sg U53536 ( .A(reg_www_10[4]), .B(n34852), .X(n23944) );
  nand_x1_sg U53537 ( .A(reg_ww_10[4]), .B(n35201), .X(n23945) );
  nand_x1_sg U53538 ( .A(reg_ww_10[6]), .B(n32326), .X(n23908) );
  nand_x1_sg U53539 ( .A(n35223), .B(reg_w_10[6]), .X(n23909) );
  nand_x1_sg U53540 ( .A(reg_www_10[7]), .B(n32383), .X(n23950) );
  nand_x1_sg U53541 ( .A(reg_ww_10[7]), .B(n31041), .X(n23951) );
  nand_x1_sg U53542 ( .A(reg_ww_10[9]), .B(n32228), .X(n23914) );
  nand_x1_sg U53543 ( .A(n35224), .B(reg_w_10[9]), .X(n23915) );
  nand_x1_sg U53544 ( .A(reg_ww_10[12]), .B(n31725), .X(n23920) );
  nand_x1_sg U53545 ( .A(n30037), .B(reg_w_10[12]), .X(n23921) );
  nand_x1_sg U53546 ( .A(reg_ww_10[15]), .B(n32343), .X(n23926) );
  nand_x1_sg U53547 ( .A(n34051), .B(reg_w_10[15]), .X(n23927) );
  nand_x1_sg U53548 ( .A(reg_ww_10[18]), .B(n32037), .X(n23932) );
  nand_x1_sg U53549 ( .A(n30899), .B(reg_w_10[18]), .X(n23933) );
  nand_x1_sg U53550 ( .A(reg_www_13[1]), .B(n32336), .X(n24166) );
  nand_x1_sg U53551 ( .A(reg_ww_13[1]), .B(n35332), .X(n24167) );
  nand_x1_sg U53552 ( .A(reg_www_13[4]), .B(n32231), .X(n24172) );
  nand_x1_sg U53553 ( .A(reg_ww_13[4]), .B(n32740), .X(n24173) );
  nand_x1_sg U53554 ( .A(reg_ww_13[6]), .B(n31636), .X(n24148) );
  nand_x1_sg U53555 ( .A(n34004), .B(reg_w_13[6]), .X(n24149) );
  nand_x1_sg U53556 ( .A(reg_www_13[7]), .B(n32456), .X(n24178) );
  nand_x1_sg U53557 ( .A(reg_ww_13[7]), .B(n35184), .X(n24179) );
  nand_x1_sg U53558 ( .A(reg_ww_13[9]), .B(n32018), .X(n24154) );
  nand_x1_sg U53559 ( .A(n35237), .B(reg_w_13[9]), .X(n24155) );
  nand_x1_sg U53560 ( .A(reg_www_13[10]), .B(n31646), .X(n24184) );
  nand_x1_sg U53561 ( .A(reg_ww_13[10]), .B(n32741), .X(n24185) );
  nand_x1_sg U53562 ( .A(reg_ww_13[12]), .B(n31642), .X(n24160) );
  nand_x1_sg U53563 ( .A(n32752), .B(reg_w_13[12]), .X(n24161) );
  nand_x1_sg U53564 ( .A(reg_www_13[13]), .B(n32295), .X(n24190) );
  nand_x1_sg U53565 ( .A(reg_ww_13[13]), .B(n32731), .X(n24191) );
  nand_x1_sg U53566 ( .A(reg_www_13[16]), .B(n32307), .X(n24196) );
  nand_x1_sg U53567 ( .A(reg_ww_13[16]), .B(n35353), .X(n24197) );
  nand_x1_sg U53568 ( .A(reg_ww_13[16]), .B(n32321), .X(n23638) );
  nand_x1_sg U53569 ( .A(n35191), .B(reg_w_13[16]), .X(n23639) );
  nand_x1_sg U53570 ( .A(reg_www_13[19]), .B(n34893), .X(n24202) );
  nand_x1_sg U53571 ( .A(reg_ww_13[19]), .B(n32723), .X(n24203) );
  nand_x1_sg U53572 ( .A(reg_ww_13[19]), .B(n32386), .X(n23644) );
  nand_x1_sg U53573 ( .A(n32724), .B(reg_w_13[19]), .X(n23645) );
  nand_x1_sg U53574 ( .A(reg_www_14[0]), .B(n32363), .X(n23686) );
  nand_x1_sg U53575 ( .A(reg_ww_14[0]), .B(n30875), .X(n23687) );
  nand_x1_sg U53576 ( .A(reg_ww_14[2]), .B(n32495), .X(n23650) );
  nand_x1_sg U53577 ( .A(n34001), .B(reg_w_14[2]), .X(n23651) );
  nand_x1_sg U53578 ( .A(reg_www_14[3]), .B(n32293), .X(n23692) );
  nand_x1_sg U53579 ( .A(reg_ww_14[3]), .B(n30595), .X(n23693) );
  nand_x1_sg U53580 ( .A(reg_ww_14[5]), .B(n32408), .X(n23656) );
  nand_x1_sg U53581 ( .A(n32764), .B(reg_w_14[5]), .X(n23657) );
  nand_x1_sg U53582 ( .A(reg_ww_14[8]), .B(n32343), .X(n23662) );
  nand_x1_sg U53583 ( .A(n32740), .B(reg_w_14[8]), .X(n23663) );
  nand_x1_sg U53584 ( .A(reg_ww_14[11]), .B(n32163), .X(n23668) );
  nand_x1_sg U53585 ( .A(n34662), .B(reg_w_14[11]), .X(n23669) );
  nand_x1_sg U53586 ( .A(reg_ww_14[14]), .B(n32296), .X(n23674) );
  nand_x1_sg U53587 ( .A(n35376), .B(reg_w_14[14]), .X(n23675) );
  nand_x1_sg U53588 ( .A(reg_ww_14[17]), .B(n32303), .X(n23680) );
  nand_x1_sg U53589 ( .A(n32759), .B(reg_w_14[17]), .X(n23681) );
  nand_x1_sg U53590 ( .A(reg_iii_0[0]), .B(n34937), .X(n25836) );
  nand_x1_sg U53591 ( .A(reg_ii_0[0]), .B(n31492), .X(n25837) );
  nand_x1_sg U53592 ( .A(reg_iii_0[1]), .B(n33943), .X(n25838) );
  nand_x1_sg U53593 ( .A(reg_ii_0[1]), .B(n35395), .X(n25839) );
  nand_x1_sg U53594 ( .A(reg_iii_0[2]), .B(n30153), .X(n25840) );
  nand_x1_sg U53595 ( .A(reg_ii_0[2]), .B(n29762), .X(n25841) );
  nand_x1_sg U53596 ( .A(reg_iii_0[3]), .B(n32305), .X(n25842) );
  nand_x1_sg U53597 ( .A(reg_ii_0[3]), .B(n32443), .X(n25843) );
  nand_x1_sg U53598 ( .A(reg_iii_0[4]), .B(n31509), .X(n25844) );
  nand_x1_sg U53599 ( .A(reg_ii_0[4]), .B(n30747), .X(n25845) );
  nand_x1_sg U53600 ( .A(reg_iii_0[5]), .B(n32308), .X(n25846) );
  nand_x1_sg U53601 ( .A(reg_ii_0[5]), .B(n30729), .X(n25847) );
  nand_x1_sg U53602 ( .A(reg_iii_0[6]), .B(n32320), .X(n25848) );
  nand_x1_sg U53603 ( .A(reg_ii_0[6]), .B(n35092), .X(n25849) );
  nand_x1_sg U53604 ( .A(reg_iii_0[7]), .B(n32332), .X(n25850) );
  nand_x1_sg U53605 ( .A(reg_ii_0[7]), .B(n32713), .X(n25851) );
  nand_x1_sg U53606 ( .A(reg_iii_0[8]), .B(n32291), .X(n25852) );
  nand_x1_sg U53607 ( .A(reg_ii_0[8]), .B(n30889), .X(n25853) );
  nand_x1_sg U53608 ( .A(reg_iii_0[9]), .B(n32854), .X(n25854) );
  nand_x1_sg U53609 ( .A(reg_ii_0[9]), .B(n35167), .X(n25855) );
  nand_x1_sg U53610 ( .A(reg_iii_0[10]), .B(n32455), .X(n25856) );
  nand_x1_sg U53611 ( .A(reg_ii_0[10]), .B(n35198), .X(n25857) );
  nand_x1_sg U53612 ( .A(reg_iii_0[11]), .B(n32328), .X(n25858) );
  nand_x1_sg U53613 ( .A(reg_ii_0[11]), .B(n30748), .X(n25859) );
  nand_x1_sg U53614 ( .A(reg_iii_0[12]), .B(n32019), .X(n25860) );
  nand_x1_sg U53615 ( .A(reg_ii_0[12]), .B(n30589), .X(n25861) );
  nand_x1_sg U53616 ( .A(reg_iii_0[13]), .B(n32317), .X(n25862) );
  nand_x1_sg U53617 ( .A(reg_ii_0[13]), .B(n31489), .X(n25863) );
  nand_x1_sg U53618 ( .A(reg_iii_0[14]), .B(n32355), .X(n25864) );
  nand_x1_sg U53619 ( .A(reg_ii_0[14]), .B(n30725), .X(n25865) );
  nand_x1_sg U53620 ( .A(reg_iii_0[15]), .B(n30208), .X(n25866) );
  nand_x1_sg U53621 ( .A(reg_ii_0[15]), .B(n31097), .X(n25867) );
  nand_x1_sg U53622 ( .A(reg_iii_0[16]), .B(n31904), .X(n25868) );
  nand_x1_sg U53623 ( .A(reg_ii_0[16]), .B(n35187), .X(n25869) );
  nand_x1_sg U53624 ( .A(reg_iii_0[17]), .B(n34571), .X(n25870) );
  nand_x1_sg U53625 ( .A(reg_ii_0[17]), .B(n30718), .X(n25871) );
  nand_x1_sg U53626 ( .A(reg_iii_0[18]), .B(n31499), .X(n25872) );
  nand_x1_sg U53627 ( .A(reg_ii_0[18]), .B(n31095), .X(n25873) );
  nand_x1_sg U53628 ( .A(reg_iii_3[0]), .B(n32348), .X(n26076) );
  nand_x1_sg U53629 ( .A(reg_ii_3[0]), .B(n30869), .X(n26077) );
  nand_x1_sg U53630 ( .A(reg_iii_3[1]), .B(n32282), .X(n26078) );
  nand_x1_sg U53631 ( .A(reg_ii_3[1]), .B(n32755), .X(n26079) );
  nand_x1_sg U53632 ( .A(reg_iii_3[2]), .B(n31745), .X(n26080) );
  nand_x1_sg U53633 ( .A(reg_ii_3[2]), .B(n30173), .X(n26081) );
  nand_x1_sg U53634 ( .A(reg_iii_3[3]), .B(n31515), .X(n26082) );
  nand_x1_sg U53635 ( .A(reg_ii_3[3]), .B(n30712), .X(n26083) );
  nand_x1_sg U53636 ( .A(reg_iii_3[4]), .B(n32776), .X(n26084) );
  nand_x1_sg U53637 ( .A(reg_ii_3[4]), .B(n32712), .X(n26085) );
  nand_x1_sg U53638 ( .A(reg_iii_3[5]), .B(n32015), .X(n26086) );
  nand_x1_sg U53639 ( .A(reg_ii_3[5]), .B(n30586), .X(n26087) );
  nand_x1_sg U53640 ( .A(reg_iii_3[6]), .B(n32495), .X(n26088) );
  nand_x1_sg U53641 ( .A(reg_ii_3[6]), .B(n33999), .X(n26089) );
  nand_x1_sg U53642 ( .A(reg_iii_3[7]), .B(n35078), .X(n26090) );
  nand_x1_sg U53643 ( .A(reg_ii_3[7]), .B(n31029), .X(n26091) );
  nand_x1_sg U53644 ( .A(reg_iii_3[8]), .B(n32349), .X(n26092) );
  nand_x1_sg U53645 ( .A(reg_ii_3[8]), .B(n32842), .X(n26093) );
  nand_x1_sg U53646 ( .A(reg_iii_3[9]), .B(n32159), .X(n26094) );
  nand_x1_sg U53647 ( .A(reg_ii_3[9]), .B(n31095), .X(n26095) );
  nand_x1_sg U53648 ( .A(reg_iii_3[10]), .B(n32408), .X(n26096) );
  nand_x1_sg U53649 ( .A(reg_ii_3[10]), .B(n34714), .X(n26097) );
  nand_x1_sg U53650 ( .A(reg_iii_3[11]), .B(n32288), .X(n26098) );
  nand_x1_sg U53651 ( .A(reg_ii_3[11]), .B(n32721), .X(n26099) );
  nand_x1_sg U53652 ( .A(reg_iii_3[12]), .B(n31905), .X(n26100) );
  nand_x1_sg U53653 ( .A(reg_ii_3[12]), .B(n32834), .X(n26101) );
  nand_x1_sg U53654 ( .A(reg_iii_3[13]), .B(n31497), .X(n26102) );
  nand_x1_sg U53655 ( .A(reg_ii_3[13]), .B(n35162), .X(n26103) );
  nand_x1_sg U53656 ( .A(reg_iii_3[14]), .B(n32166), .X(n26104) );
  nand_x1_sg U53657 ( .A(reg_ii_3[14]), .B(n30724), .X(n26105) );
  nand_x1_sg U53658 ( .A(reg_iii_3[15]), .B(n32040), .X(n26106) );
  nand_x1_sg U53659 ( .A(reg_ii_3[15]), .B(n31031), .X(n26107) );
  nand_x1_sg U53660 ( .A(reg_iii_3[16]), .B(n35077), .X(n26108) );
  nand_x1_sg U53661 ( .A(reg_ii_3[16]), .B(n35197), .X(n26109) );
  nand_x1_sg U53662 ( .A(reg_iii_3[17]), .B(n32305), .X(n26110) );
  nand_x1_sg U53663 ( .A(reg_ii_3[17]), .B(n35160), .X(n26111) );
  nand_x1_sg U53664 ( .A(reg_iii_3[18]), .B(n31896), .X(n26112) );
  nand_x1_sg U53665 ( .A(reg_ii_3[18]), .B(n31054), .X(n26113) );
  nand_x1_sg U53666 ( .A(reg_iii_3[19]), .B(n30623), .X(n26114) );
  nand_x1_sg U53667 ( .A(reg_ii_3[19]), .B(n31489), .X(n26115) );
  nand_x1_sg U53668 ( .A(reg_iii_6[0]), .B(n30169), .X(n25520) );
  nand_x1_sg U53669 ( .A(reg_ii_6[0]), .B(n30887), .X(n25521) );
  nand_x1_sg U53670 ( .A(reg_iii_6[1]), .B(n34571), .X(n25522) );
  nand_x1_sg U53671 ( .A(reg_ii_6[1]), .B(n35177), .X(n25523) );
  nand_x1_sg U53672 ( .A(reg_iii_6[2]), .B(n32360), .X(n25524) );
  nand_x1_sg U53673 ( .A(reg_ii_6[2]), .B(n32723), .X(n25525) );
  nand_x1_sg U53674 ( .A(reg_iii_6[3]), .B(n31902), .X(n25526) );
  nand_x1_sg U53675 ( .A(reg_ii_6[3]), .B(n30869), .X(n25527) );
  nand_x1_sg U53676 ( .A(reg_iii_6[4]), .B(n32769), .X(n25528) );
  nand_x1_sg U53677 ( .A(reg_ii_6[4]), .B(n30870), .X(n25529) );
  nand_x1_sg U53678 ( .A(reg_iii_6[5]), .B(n31910), .X(n25530) );
  nand_x1_sg U53679 ( .A(reg_ii_6[5]), .B(n30887), .X(n25531) );
  nand_x1_sg U53680 ( .A(reg_iii_6[6]), .B(n32499), .X(n25532) );
  nand_x1_sg U53681 ( .A(reg_ii_6[6]), .B(n34091), .X(n25533) );
  nand_x1_sg U53682 ( .A(reg_iii_6[7]), .B(n31719), .X(n25534) );
  nand_x1_sg U53683 ( .A(reg_ii_6[7]), .B(n35167), .X(n25535) );
  nand_x1_sg U53684 ( .A(reg_iii_6[8]), .B(n31925), .X(n25536) );
  nand_x1_sg U53685 ( .A(reg_ii_6[8]), .B(n35225), .X(n25537) );
  nand_x1_sg U53686 ( .A(reg_iii_6[9]), .B(n31499), .X(n25538) );
  nand_x1_sg U53687 ( .A(reg_ii_6[9]), .B(n35222), .X(n25539) );
  nand_x1_sg U53688 ( .A(reg_iii_6[10]), .B(n32244), .X(n25540) );
  nand_x1_sg U53689 ( .A(reg_ii_6[10]), .B(n31671), .X(n25541) );
  nand_x1_sg U53690 ( .A(reg_iii_6[11]), .B(n32429), .X(n25542) );
  nand_x1_sg U53691 ( .A(reg_ii_6[11]), .B(n31054), .X(n25543) );
  nand_x1_sg U53692 ( .A(reg_iii_6[12]), .B(n32229), .X(n25544) );
  nand_x1_sg U53693 ( .A(reg_ii_6[12]), .B(n30712), .X(n25545) );
  nand_x1_sg U53694 ( .A(reg_iii_6[13]), .B(n31909), .X(n25546) );
  nand_x1_sg U53695 ( .A(reg_ii_6[13]), .B(n30867), .X(n25547) );
  nand_x1_sg U53696 ( .A(reg_iii_6[14]), .B(n31736), .X(n25548) );
  nand_x1_sg U53697 ( .A(reg_ii_6[14]), .B(n33997), .X(n25549) );
  nand_x1_sg U53698 ( .A(reg_iii_6[15]), .B(n32776), .X(n25550) );
  nand_x1_sg U53699 ( .A(reg_ii_6[15]), .B(n30588), .X(n25551) );
  nand_x1_sg U53700 ( .A(reg_iii_6[16]), .B(n32347), .X(n25552) );
  nand_x1_sg U53701 ( .A(reg_ii_6[16]), .B(n32845), .X(n25553) );
  nand_x1_sg U53702 ( .A(reg_iii_9[0]), .B(n32153), .X(n25756) );
  nand_x1_sg U53703 ( .A(reg_ii_9[0]), .B(n32762), .X(n25757) );
  nand_x1_sg U53704 ( .A(reg_iii_9[1]), .B(n32335), .X(n25758) );
  nand_x1_sg U53705 ( .A(reg_ii_9[1]), .B(n34083), .X(n25759) );
  nand_x1_sg U53706 ( .A(reg_iii_9[2]), .B(n32151), .X(n25760) );
  nand_x1_sg U53707 ( .A(reg_ii_9[2]), .B(n30874), .X(n25761) );
  nand_x1_sg U53708 ( .A(reg_iii_9[3]), .B(n32032), .X(n25762) );
  nand_x1_sg U53709 ( .A(reg_ii_9[3]), .B(n30877), .X(n25763) );
  nand_x1_sg U53710 ( .A(reg_iii_9[4]), .B(n32313), .X(n25764) );
  nand_x1_sg U53711 ( .A(reg_ii_9[4]), .B(n31031), .X(n25765) );
  nand_x1_sg U53712 ( .A(reg_iii_9[5]), .B(n32232), .X(n25766) );
  nand_x1_sg U53713 ( .A(reg_ii_9[5]), .B(n34699), .X(n25767) );
  nand_x1_sg U53714 ( .A(reg_iii_9[6]), .B(n32308), .X(n25768) );
  nand_x1_sg U53715 ( .A(reg_ii_9[6]), .B(n32759), .X(n25769) );
  nand_x1_sg U53716 ( .A(reg_iii_9[7]), .B(n32154), .X(n25770) );
  nand_x1_sg U53717 ( .A(reg_ii_9[7]), .B(n32443), .X(n25771) );
  nand_x1_sg U53718 ( .A(reg_iii_9[8]), .B(n34850), .X(n25772) );
  nand_x1_sg U53719 ( .A(reg_ii_9[8]), .B(n35351), .X(n25773) );
  nand_x1_sg U53720 ( .A(reg_iii_9[9]), .B(n32381), .X(n25774) );
  nand_x1_sg U53721 ( .A(reg_ii_9[9]), .B(n35182), .X(n25775) );
  nand_x1_sg U53722 ( .A(reg_iii_9[10]), .B(n32771), .X(n25776) );
  nand_x1_sg U53723 ( .A(reg_ii_9[10]), .B(n31491), .X(n25777) );
  nand_x1_sg U53724 ( .A(reg_iii_9[11]), .B(n32166), .X(n25778) );
  nand_x1_sg U53725 ( .A(reg_ii_9[11]), .B(n35082), .X(n25779) );
  nand_x1_sg U53726 ( .A(reg_iii_9[12]), .B(n32450), .X(n25780) );
  nand_x1_sg U53727 ( .A(reg_ii_9[12]), .B(n31673), .X(n25781) );
  nand_x1_sg U53728 ( .A(reg_iii_9[13]), .B(n31741), .X(n25782) );
  nand_x1_sg U53729 ( .A(reg_ii_9[13]), .B(n35320), .X(n25783) );
  nand_x1_sg U53730 ( .A(reg_iii_9[14]), .B(n31505), .X(n25784) );
  nand_x1_sg U53731 ( .A(reg_ii_9[14]), .B(n35093), .X(n25785) );
  nand_x1_sg U53732 ( .A(reg_iii_9[15]), .B(n30140), .X(n25786) );
  nand_x1_sg U53733 ( .A(reg_ii_9[15]), .B(n35229), .X(n25787) );
  nand_x1_sg U53734 ( .A(reg_iii_9[16]), .B(n32316), .X(n25788) );
  nand_x1_sg U53735 ( .A(reg_ii_9[16]), .B(n35332), .X(n25789) );
  nand_x1_sg U53736 ( .A(reg_iii_9[17]), .B(n30916), .X(n25790) );
  nand_x1_sg U53737 ( .A(reg_ii_9[17]), .B(n35355), .X(n25791) );
  nand_x1_sg U53738 ( .A(reg_iii_9[18]), .B(n32249), .X(n25792) );
  nand_x1_sg U53739 ( .A(reg_ii_9[18]), .B(n34709), .X(n25793) );
  nand_x1_sg U53740 ( .A(reg_iii_9[19]), .B(n32300), .X(n25794) );
  nand_x1_sg U53741 ( .A(reg_ii_9[19]), .B(n34714), .X(n25795) );
  nand_x1_sg U53742 ( .A(reg_iii_12[0]), .B(n32296), .X(n25204) );
  nand_x1_sg U53743 ( .A(reg_ii_12[0]), .B(n31491), .X(n25205) );
  nand_x1_sg U53744 ( .A(reg_iii_12[1]), .B(n32400), .X(n25206) );
  nand_x1_sg U53745 ( .A(reg_ii_12[1]), .B(n35326), .X(n25207) );
  nand_x1_sg U53746 ( .A(reg_iii_12[2]), .B(n32495), .X(n25208) );
  nand_x1_sg U53747 ( .A(reg_ii_12[2]), .B(n35317), .X(n25209) );
  nand_x1_sg U53748 ( .A(reg_iii_12[3]), .B(n32236), .X(n25210) );
  nand_x1_sg U53749 ( .A(reg_ii_12[3]), .B(n35087), .X(n25211) );
  nand_x1_sg U53750 ( .A(reg_iii_12[4]), .B(n31728), .X(n25212) );
  nand_x1_sg U53751 ( .A(reg_ii_12[4]), .B(n30898), .X(n25213) );
  nand_x1_sg U53752 ( .A(reg_iii_12[5]), .B(n30151), .X(n25214) );
  nand_x1_sg U53753 ( .A(reg_ii_12[5]), .B(n32743), .X(n25215) );
  nand_x1_sg U53754 ( .A(reg_iii_12[6]), .B(n32048), .X(n25216) );
  nand_x1_sg U53755 ( .A(reg_ii_12[6]), .B(n34712), .X(n25217) );
  nand_x1_sg U53756 ( .A(reg_iii_12[7]), .B(n32166), .X(n25218) );
  nand_x1_sg U53757 ( .A(reg_ii_12[7]), .B(n31206), .X(n25219) );
  nand_x1_sg U53758 ( .A(reg_iii_12[8]), .B(n34552), .X(n25220) );
  nand_x1_sg U53759 ( .A(reg_ii_12[8]), .B(n30861), .X(n25221) );
  nand_x1_sg U53760 ( .A(reg_iii_12[9]), .B(n32016), .X(n25222) );
  nand_x1_sg U53761 ( .A(reg_ii_12[9]), .B(n30587), .X(n25223) );
  nand_x1_sg U53762 ( .A(reg_iii_12[10]), .B(n32453), .X(n25224) );
  nand_x1_sg U53763 ( .A(reg_ii_12[10]), .B(n32846), .X(n25225) );
  nand_x1_sg U53764 ( .A(reg_iii_12[11]), .B(n32282), .X(n25226) );
  nand_x1_sg U53765 ( .A(reg_ii_12[11]), .B(n31060), .X(n25227) );
  nand_x1_sg U53766 ( .A(reg_iii_12[12]), .B(n32035), .X(n25228) );
  nand_x1_sg U53767 ( .A(reg_ii_12[12]), .B(n31489), .X(n25229) );
  nand_x1_sg U53768 ( .A(reg_iii_12[13]), .B(n32320), .X(n25230) );
  nand_x1_sg U53769 ( .A(reg_ii_12[13]), .B(n34704), .X(n25231) );
  nand_x1_sg U53770 ( .A(reg_iii_12[14]), .B(n32369), .X(n25232) );
  nand_x1_sg U53771 ( .A(reg_ii_12[14]), .B(n32737), .X(n25233) );
  nand_x1_sg U53772 ( .A(reg_iii_12[15]), .B(n32012), .X(n25234) );
  nand_x1_sg U53773 ( .A(reg_ii_12[15]), .B(n32718), .X(n25235) );
  nand_x1_sg U53774 ( .A(reg_iii_12[16]), .B(n32241), .X(n25236) );
  nand_x1_sg U53775 ( .A(reg_ii_12[16]), .B(n30884), .X(n25237) );
  nand_x1_sg U53776 ( .A(reg_iii_12[17]), .B(n32496), .X(n25238) );
  nand_x1_sg U53777 ( .A(reg_ii_12[17]), .B(n35321), .X(n25239) );
  nand_x1_sg U53778 ( .A(reg_iii_12[18]), .B(n34566), .X(n25240) );
  nand_x1_sg U53779 ( .A(reg_ii_12[18]), .B(n35185), .X(n25241) );
  nand_x1_sg U53780 ( .A(reg_iii_12[19]), .B(n30920), .X(n25242) );
  nand_x1_sg U53781 ( .A(reg_ii_12[19]), .B(n35186), .X(n25243) );
  nand_x1_sg U53782 ( .A(reg_iii_13[0]), .B(n32042), .X(n25284) );
  nand_x1_sg U53783 ( .A(reg_ii_13[0]), .B(n31056), .X(n25285) );
  nand_x1_sg U53784 ( .A(reg_iii_13[1]), .B(n32375), .X(n25286) );
  nand_x1_sg U53785 ( .A(reg_ii_13[1]), .B(n35093), .X(n25287) );
  nand_x1_sg U53786 ( .A(reg_iii_13[2]), .B(n32408), .X(n25288) );
  nand_x1_sg U53787 ( .A(reg_ii_13[2]), .B(n32730), .X(n25289) );
  nand_x1_sg U53788 ( .A(reg_iii_13[3]), .B(n32316), .X(n25290) );
  nand_x1_sg U53789 ( .A(reg_ii_13[3]), .B(n35396), .X(n25291) );
  nand_x1_sg U53790 ( .A(reg_iii_13[4]), .B(n31894), .X(n25292) );
  nand_x1_sg U53791 ( .A(reg_ii_13[4]), .B(n35376), .X(n25293) );
  nand_x1_sg U53792 ( .A(reg_iii_13[5]), .B(n33943), .X(n25294) );
  nand_x1_sg U53793 ( .A(reg_ii_13[5]), .B(n35399), .X(n25295) );
  nand_x1_sg U53794 ( .A(reg_iii_13[6]), .B(n34553), .X(n25296) );
  nand_x1_sg U53795 ( .A(reg_ii_13[6]), .B(n30726), .X(n25297) );
  nand_x1_sg U53796 ( .A(reg_iii_15[0]), .B(n32018), .X(n24648) );
  nand_x1_sg U53797 ( .A(reg_ii_15[0]), .B(n32732), .X(n24649) );
  nand_x1_sg U53798 ( .A(reg_iii_15[1]), .B(n32041), .X(n24650) );
  nand_x1_sg U53799 ( .A(reg_ii_15[1]), .B(n35205), .X(n24651) );
  nand_x1_sg U53800 ( .A(reg_iii_15[2]), .B(n33947), .X(n24652) );
  nand_x1_sg U53801 ( .A(reg_ii_15[2]), .B(n32764), .X(n24653) );
  nand_x1_sg U53802 ( .A(reg_iii_15[3]), .B(n32237), .X(n24654) );
  nand_x1_sg U53803 ( .A(reg_ii_15[3]), .B(n35403), .X(n24655) );
  nand_x1_sg U53804 ( .A(reg_iii_15[4]), .B(n34936), .X(n24656) );
  nand_x1_sg U53805 ( .A(reg_ii_15[4]), .B(n34724), .X(n24657) );
  nand_x1_sg U53806 ( .A(reg_iii_15[5]), .B(n31717), .X(n24658) );
  nand_x1_sg U53807 ( .A(reg_ii_15[5]), .B(n30707), .X(n24659) );
  nand_x1_sg U53808 ( .A(reg_iii_15[6]), .B(n32161), .X(n24660) );
  nand_x1_sg U53809 ( .A(reg_ii_15[6]), .B(n35213), .X(n24661) );
  nand_x1_sg U53810 ( .A(reg_iii_15[7]), .B(n31630), .X(n24662) );
  nand_x1_sg U53811 ( .A(reg_ii_15[7]), .B(n35227), .X(n24663) );
  nand_x1_sg U53812 ( .A(reg_iii_15[8]), .B(n33976), .X(n24664) );
  nand_x1_sg U53813 ( .A(reg_ii_15[8]), .B(n32747), .X(n24665) );
  nand_x1_sg U53814 ( .A(reg_iii_15[9]), .B(n31897), .X(n24666) );
  nand_x1_sg U53815 ( .A(reg_ii_15[9]), .B(n31035), .X(n24667) );
  nand_x1_sg U53816 ( .A(reg_iii_15[10]), .B(n32406), .X(n24668) );
  nand_x1_sg U53817 ( .A(reg_ii_15[10]), .B(n35087), .X(n24669) );
  nand_x1_sg U53818 ( .A(reg_iii_15[11]), .B(n31743), .X(n24670) );
  nand_x1_sg U53819 ( .A(reg_ii_15[11]), .B(n34708), .X(n24671) );
  nand_x1_sg U53820 ( .A(reg_iii_15[12]), .B(n32328), .X(n24672) );
  nand_x1_sg U53821 ( .A(reg_ii_15[12]), .B(n32839), .X(n24673) );
  nand_x1_sg U53822 ( .A(reg_iii_15[13]), .B(n33942), .X(n24674) );
  nand_x1_sg U53823 ( .A(reg_ii_15[13]), .B(n32845), .X(n24675) );
  nand_x1_sg U53824 ( .A(reg_iii_15[14]), .B(n31503), .X(n24676) );
  nand_x1_sg U53825 ( .A(reg_ii_15[14]), .B(n30727), .X(n24677) );
  nand_x1_sg U53826 ( .A(reg_iii_15[15]), .B(n32454), .X(n24678) );
  nand_x1_sg U53827 ( .A(reg_ii_15[15]), .B(n35395), .X(n24679) );
  nand_x1_sg U53828 ( .A(reg_iii_15[16]), .B(n32015), .X(n24680) );
  nand_x1_sg U53829 ( .A(reg_ii_15[16]), .B(n32847), .X(n24681) );
  nand_x1_sg U53830 ( .A(reg_iii_15[17]), .B(n32234), .X(n24682) );
  nand_x1_sg U53831 ( .A(reg_ii_15[17]), .B(n32829), .X(n24683) );
  nand_x1_sg U53832 ( .A(reg_iii_15[18]), .B(n32287), .X(n24684) );
  nand_x1_sg U53833 ( .A(reg_ii_15[18]), .B(n32844), .X(n24685) );
  nand_x1_sg U53834 ( .A(reg_iii_15[19]), .B(n34578), .X(n24686) );
  nand_x1_sg U53835 ( .A(reg_ii_15[19]), .B(n35184), .X(n24687) );
  nand_x1_sg U53836 ( .A(reg_www_2[13]), .B(n34570), .X(n24914) );
  nand_x1_sg U53837 ( .A(reg_ww_2[13]), .B(n31043), .X(n24915) );
  nand_x1_sg U53838 ( .A(reg_www_2[14]), .B(n30144), .X(n24916) );
  nand_x1_sg U53839 ( .A(reg_ww_2[14]), .B(n30727), .X(n24917) );
  nand_x1_sg U53840 ( .A(reg_www_2[15]), .B(n31745), .X(n24918) );
  nand_x1_sg U53841 ( .A(reg_ww_2[15]), .B(n31492), .X(n24919) );
  nand_x1_sg U53842 ( .A(reg_www_2[16]), .B(n31712), .X(n24920) );
  nand_x1_sg U53843 ( .A(reg_ww_2[16]), .B(n35358), .X(n24921) );
  nand_x1_sg U53844 ( .A(reg_www_2[17]), .B(n34580), .X(n24922) );
  nand_x1_sg U53845 ( .A(reg_ww_2[17]), .B(n32846), .X(n24923) );
  nand_x1_sg U53846 ( .A(reg_www_2[18]), .B(n32384), .X(n24924) );
  nand_x1_sg U53847 ( .A(reg_ww_2[18]), .B(n35183), .X(n24925) );
  nand_x1_sg U53848 ( .A(reg_www_2[19]), .B(n33942), .X(n24926) );
  nand_x1_sg U53849 ( .A(reg_ww_2[19]), .B(n35233), .X(n24927) );
  nand_x1_sg U53850 ( .A(reg_www_3[0]), .B(n32226), .X(n24960) );
  nand_x1_sg U53851 ( .A(reg_ww_3[0]), .B(n32749), .X(n24961) );
  nand_x1_sg U53852 ( .A(reg_www_3[1]), .B(n33977), .X(n24962) );
  nand_x1_sg U53853 ( .A(reg_ww_3[1]), .B(n32834), .X(n24963) );
  nand_x1_sg U53854 ( .A(reg_www_3[2]), .B(n32231), .X(n24964) );
  nand_x1_sg U53855 ( .A(reg_ww_3[2]), .B(n35370), .X(n24965) );
  nand_x1_sg U53856 ( .A(reg_www_3[3]), .B(n31731), .X(n24966) );
  nand_x1_sg U53857 ( .A(reg_ww_3[3]), .B(n34704), .X(n24967) );
  nand_x1_sg U53858 ( .A(reg_www_3[4]), .B(n32036), .X(n24968) );
  nand_x1_sg U53859 ( .A(reg_ww_3[4]), .B(n35376), .X(n24969) );
  nand_x1_sg U53860 ( .A(reg_www_3[5]), .B(n31902), .X(n24970) );
  nand_x1_sg U53861 ( .A(reg_ww_3[5]), .B(n34668), .X(n24971) );
  nand_x1_sg U53862 ( .A(reg_www_3[6]), .B(n32376), .X(n24972) );
  nand_x1_sg U53863 ( .A(reg_ww_3[6]), .B(n32733), .X(n24973) );
  nand_x1_sg U53864 ( .A(reg_www_3[7]), .B(n32148), .X(n24974) );
  nand_x1_sg U53865 ( .A(reg_ww_3[7]), .B(n35231), .X(n24975) );
  nand_x1_sg U53866 ( .A(reg_www_3[8]), .B(n32351), .X(n24976) );
  nand_x1_sg U53867 ( .A(reg_ww_3[8]), .B(n35220), .X(n24977) );
  nand_x1_sg U53868 ( .A(reg_www_5[3]), .B(n32405), .X(n24338) );
  nand_x1_sg U53869 ( .A(reg_ww_5[3]), .B(n30722), .X(n24339) );
  nand_x1_sg U53870 ( .A(reg_www_5[4]), .B(n32242), .X(n24340) );
  nand_x1_sg U53871 ( .A(reg_ww_5[4]), .B(n34042), .X(n24341) );
  nand_x1_sg U53872 ( .A(reg_www_5[5]), .B(n31649), .X(n24342) );
  nand_x1_sg U53873 ( .A(reg_ww_5[5]), .B(n30881), .X(n24343) );
  nand_x1_sg U53874 ( .A(reg_www_5[6]), .B(n32366), .X(n24344) );
  nand_x1_sg U53875 ( .A(reg_ww_5[6]), .B(n30711), .X(n24345) );
  nand_x1_sg U53876 ( .A(reg_www_5[7]), .B(n34576), .X(n24346) );
  nand_x1_sg U53877 ( .A(reg_ww_5[7]), .B(n35211), .X(n24347) );
  nand_x1_sg U53878 ( .A(reg_www_5[8]), .B(n32048), .X(n24348) );
  nand_x1_sg U53879 ( .A(reg_ww_5[8]), .B(n32717), .X(n24349) );
  nand_x1_sg U53880 ( .A(reg_www_5[9]), .B(n32318), .X(n24350) );
  nand_x1_sg U53881 ( .A(reg_ww_5[9]), .B(n30879), .X(n24351) );
  nand_x1_sg U53882 ( .A(reg_www_5[10]), .B(n34695), .X(n24352) );
  nand_x1_sg U53883 ( .A(reg_ww_5[10]), .B(n30876), .X(n24353) );
  nand_x1_sg U53884 ( .A(reg_www_5[11]), .B(n31643), .X(n24354) );
  nand_x1_sg U53885 ( .A(reg_ww_5[11]), .B(n35212), .X(n24355) );
  nand_x1_sg U53886 ( .A(reg_www_5[12]), .B(n34582), .X(n24356) );
  nand_x1_sg U53887 ( .A(reg_ww_5[12]), .B(n35089), .X(n24357) );
  nand_x1_sg U53888 ( .A(reg_www_5[13]), .B(n32360), .X(n24358) );
  nand_x1_sg U53889 ( .A(reg_ww_5[13]), .B(n30884), .X(n24359) );
  nand_x1_sg U53890 ( .A(reg_www_5[14]), .B(n31731), .X(n24360) );
  nand_x1_sg U53891 ( .A(reg_ww_5[14]), .B(n33996), .X(n24361) );
  nand_x1_sg U53892 ( .A(reg_www_5[15]), .B(n32155), .X(n24362) );
  nand_x1_sg U53893 ( .A(reg_ww_5[15]), .B(n34667), .X(n24363) );
  nand_x1_sg U53894 ( .A(reg_www_5[16]), .B(n31711), .X(n24364) );
  nand_x1_sg U53895 ( .A(reg_ww_5[16]), .B(n35367), .X(n24365) );
  nand_x1_sg U53896 ( .A(reg_www_5[17]), .B(n30918), .X(n24366) );
  nand_x1_sg U53897 ( .A(reg_ww_5[17]), .B(n30891), .X(n24367) );
  nand_x1_sg U53898 ( .A(reg_www_5[18]), .B(n32214), .X(n24368) );
  nand_x1_sg U53899 ( .A(reg_ww_5[18]), .B(n33997), .X(n24369) );
  nand_x1_sg U53900 ( .A(reg_www_5[19]), .B(n31892), .X(n24370) );
  nand_x1_sg U53901 ( .A(reg_ww_5[19]), .B(n35347), .X(n24371) );
  nand_x1_sg U53902 ( .A(reg_www_8[16]), .B(n32140), .X(n24594) );
  nand_x1_sg U53903 ( .A(reg_ww_8[16]), .B(n31096), .X(n24595) );
  nand_x1_sg U53904 ( .A(reg_www_8[17]), .B(n32251), .X(n24596) );
  nand_x1_sg U53905 ( .A(reg_ww_8[17]), .B(n35350), .X(n24597) );
  nand_x1_sg U53906 ( .A(reg_www_8[18]), .B(n31501), .X(n24598) );
  nand_x1_sg U53907 ( .A(reg_ww_8[18]), .B(n31027), .X(n24599) );
  nand_x1_sg U53908 ( .A(reg_www_8[19]), .B(n32359), .X(n24600) );
  nand_x1_sg U53909 ( .A(reg_ww_8[19]), .B(n30905), .X(n24601) );
  nand_x1_sg U53910 ( .A(reg_www_11[1]), .B(n32384), .X(n24018) );
  nand_x1_sg U53911 ( .A(reg_ww_11[1]), .B(n31037), .X(n24019) );
  nand_x1_sg U53912 ( .A(reg_www_11[2]), .B(n32318), .X(n24020) );
  nand_x1_sg U53913 ( .A(reg_ww_11[2]), .B(n34043), .X(n24021) );
  nand_x1_sg U53914 ( .A(reg_www_11[3]), .B(n32227), .X(n24022) );
  nand_x1_sg U53915 ( .A(reg_ww_11[3]), .B(n35356), .X(n24023) );
  nand_x1_sg U53916 ( .A(reg_www_11[4]), .B(n30596), .X(n24024) );
  nand_x1_sg U53917 ( .A(reg_ww_11[4]), .B(n29767), .X(n24025) );
  nand_x1_sg U53918 ( .A(reg_www_11[5]), .B(n34936), .X(n24026) );
  nand_x1_sg U53919 ( .A(reg_ww_11[5]), .B(n32832), .X(n24027) );
  nand_x1_sg U53920 ( .A(reg_www_11[6]), .B(n32401), .X(n24028) );
  nand_x1_sg U53921 ( .A(reg_ww_11[6]), .B(n30882), .X(n24029) );
  nand_x1_sg U53922 ( .A(reg_www_11[7]), .B(n31511), .X(n24030) );
  nand_x1_sg U53923 ( .A(reg_ww_11[7]), .B(n35218), .X(n24031) );
  nand_x1_sg U53924 ( .A(reg_www_11[8]), .B(n31740), .X(n24032) );
  nand_x1_sg U53925 ( .A(reg_ww_11[8]), .B(n35368), .X(n24033) );
  nand_x1_sg U53926 ( .A(reg_www_11[9]), .B(n30730), .X(n24034) );
  nand_x1_sg U53927 ( .A(reg_ww_11[9]), .B(n30707), .X(n24035) );
  nand_x1_sg U53928 ( .A(reg_www_11[10]), .B(n33982), .X(n24036) );
  nand_x1_sg U53929 ( .A(reg_ww_11[10]), .B(n32765), .X(n24037) );
  nand_x1_sg U53930 ( .A(reg_www_11[11]), .B(n31643), .X(n24038) );
  nand_x1_sg U53931 ( .A(reg_ww_11[11]), .B(n30173), .X(n24039) );
  nand_x1_sg U53932 ( .A(reg_www_11[12]), .B(n32247), .X(n24040) );
  nand_x1_sg U53933 ( .A(reg_ww_11[12]), .B(n35338), .X(n24041) );
  nand_x1_sg U53934 ( .A(reg_www_11[13]), .B(n32045), .X(n24042) );
  nand_x1_sg U53935 ( .A(reg_ww_11[13]), .B(n30859), .X(n24043) );
  nand_x1_sg U53936 ( .A(reg_www_11[14]), .B(n32140), .X(n24044) );
  nand_x1_sg U53937 ( .A(reg_ww_11[14]), .B(n30878), .X(n24045) );
  nand_x1_sg U53938 ( .A(reg_www_11[15]), .B(n32011), .X(n24046) );
  nand_x1_sg U53939 ( .A(reg_ww_11[15]), .B(n30902), .X(n24047) );
  nand_x1_sg U53940 ( .A(reg_www_11[16]), .B(n32020), .X(n24048) );
  nand_x1_sg U53941 ( .A(reg_ww_11[16]), .B(n35344), .X(n24049) );
  nand_x1_sg U53942 ( .A(reg_www_11[17]), .B(n32049), .X(n24050) );
  nand_x1_sg U53943 ( .A(reg_ww_11[17]), .B(n30866), .X(n24051) );
  nand_x1_sg U53944 ( .A(reg_www_11[18]), .B(n31720), .X(n24052) );
  nand_x1_sg U53945 ( .A(reg_ww_11[18]), .B(n31043), .X(n24053) );
  nand_x1_sg U53946 ( .A(reg_www_11[19]), .B(n32148), .X(n24054) );
  nand_x1_sg U53947 ( .A(reg_ww_11[19]), .B(n31041), .X(n24055) );
  nand_x1_sg U53948 ( .A(reg_www_12[0]), .B(n31633), .X(n24096) );
  nand_x1_sg U53949 ( .A(reg_ww_12[0]), .B(n35330), .X(n24097) );
  nand_x1_sg U53950 ( .A(reg_www_12[1]), .B(n32375), .X(n24098) );
  nand_x1_sg U53951 ( .A(reg_ww_12[1]), .B(n32747), .X(n24099) );
  nand_x1_sg U53952 ( .A(reg_www_12[2]), .B(n34567), .X(n24100) );
  nand_x1_sg U53953 ( .A(reg_ww_12[2]), .B(n30895), .X(n24101) );
  nand_x1_sg U53954 ( .A(reg_www_12[3]), .B(n30157), .X(n24102) );
  nand_x1_sg U53955 ( .A(reg_ww_12[3]), .B(n32729), .X(n24103) );
  nand_x1_sg U53956 ( .A(reg_www_12[4]), .B(n32376), .X(n24104) );
  nand_x1_sg U53957 ( .A(reg_ww_12[4]), .B(n31029), .X(n24105) );
  nand_x1_sg U53958 ( .A(reg_www_12[5]), .B(n33950), .X(n24106) );
  nand_x1_sg U53959 ( .A(reg_ww_12[5]), .B(n32443), .X(n24107) );
  nand_x1_sg U53960 ( .A(reg_www_12[6]), .B(n34897), .X(n24108) );
  nand_x1_sg U53961 ( .A(reg_ww_12[6]), .B(n35175), .X(n24109) );
  nand_x1_sg U53962 ( .A(reg_www_12[7]), .B(n32350), .X(n24110) );
  nand_x1_sg U53963 ( .A(reg_ww_12[7]), .B(n32717), .X(n24111) );
  nand_x1_sg U53964 ( .A(reg_www_12[8]), .B(n32254), .X(n24112) );
  nand_x1_sg U53965 ( .A(reg_ww_12[8]), .B(n29768), .X(n24113) );
  nand_x1_sg U53966 ( .A(reg_www_12[9]), .B(n31649), .X(n24114) );
  nand_x1_sg U53967 ( .A(reg_ww_12[9]), .B(n30905), .X(n24115) );
  nand_x1_sg U53968 ( .A(reg_www_12[10]), .B(n32386), .X(n24116) );
  nand_x1_sg U53969 ( .A(reg_ww_12[10]), .B(n32719), .X(n24117) );
  nand_x1_sg U53970 ( .A(reg_www_12[11]), .B(n32307), .X(n24118) );
  nand_x1_sg U53971 ( .A(reg_ww_12[11]), .B(n35083), .X(n24119) );
  nand_x1_sg U53972 ( .A(reg_www_12[12]), .B(n32367), .X(n24120) );
  nand_x1_sg U53973 ( .A(reg_ww_12[12]), .B(n31675), .X(n24121) );
  nand_x1_sg U53974 ( .A(reg_www_12[13]), .B(n32161), .X(n24122) );
  nand_x1_sg U53975 ( .A(reg_ww_12[13]), .B(n31043), .X(n24123) );
  nand_x1_sg U53976 ( .A(reg_www_12[14]), .B(n30157), .X(n24124) );
  nand_x1_sg U53977 ( .A(reg_ww_12[14]), .B(n30747), .X(n24125) );
  nand_x1_sg U53978 ( .A(reg_www_12[15]), .B(n31902), .X(n24126) );
  nand_x1_sg U53979 ( .A(reg_ww_12[15]), .B(n30594), .X(n24127) );
  nand_x1_sg U53980 ( .A(reg_www_12[16]), .B(n32247), .X(n24128) );
  nand_x1_sg U53981 ( .A(reg_ww_12[16]), .B(n34714), .X(n24129) );
  nand_x1_sg U53982 ( .A(reg_www_12[17]), .B(n32313), .X(n24130) );
  nand_x1_sg U53983 ( .A(reg_ww_12[17]), .B(n32761), .X(n24131) );
  nand_x1_sg U53984 ( .A(reg_www_12[18]), .B(n31713), .X(n24132) );
  nand_x1_sg U53985 ( .A(reg_ww_12[18]), .B(n32755), .X(n24133) );
  nand_x1_sg U53986 ( .A(reg_www_12[19]), .B(n31905), .X(n24134) );
  nand_x1_sg U53987 ( .A(reg_ww_12[19]), .B(n31037), .X(n24135) );
  nand_x1_sg U53988 ( .A(reg_www_15[0]), .B(n30196), .X(n23766) );
  nand_x1_sg U53989 ( .A(reg_ww_15[0]), .B(n32441), .X(n23767) );
  nand_x1_sg U53990 ( .A(reg_www_15[1]), .B(n32050), .X(n23768) );
  nand_x1_sg U53991 ( .A(reg_ww_15[1]), .B(n30905), .X(n23769) );
  nand_x1_sg U53992 ( .A(reg_www_15[2]), .B(n32026), .X(n23770) );
  nand_x1_sg U53993 ( .A(reg_ww_15[2]), .B(n32750), .X(n23771) );
  nand_x1_sg U53994 ( .A(reg_www_15[3]), .B(n32368), .X(n23772) );
  nand_x1_sg U53995 ( .A(reg_ww_15[3]), .B(n30859), .X(n23773) );
  nand_x1_sg U53996 ( .A(reg_www_15[4]), .B(n31893), .X(n23774) );
  nand_x1_sg U53997 ( .A(reg_ww_15[4]), .B(n32714), .X(n23775) );
  nand_x1_sg U53998 ( .A(reg_www_15[5]), .B(n34575), .X(n23776) );
  nand_x1_sg U53999 ( .A(reg_ww_15[5]), .B(n35199), .X(n23777) );
  nand_x1_sg U54000 ( .A(reg_www_15[6]), .B(n32159), .X(n23778) );
  nand_x1_sg U54001 ( .A(reg_ww_15[6]), .B(n35336), .X(n23779) );
  nand_x1_sg U54002 ( .A(reg_www_15[7]), .B(n32381), .X(n23780) );
  nand_x1_sg U54003 ( .A(reg_ww_15[7]), .B(n30711), .X(n23781) );
  nand_x1_sg U54004 ( .A(reg_www_15[8]), .B(n32248), .X(n23782) );
  nand_x1_sg U54005 ( .A(reg_ww_15[8]), .B(n35368), .X(n23783) );
  nand_x1_sg U54006 ( .A(reg_www_15[9]), .B(n31631), .X(n23784) );
  nand_x1_sg U54007 ( .A(reg_ww_15[9]), .B(n35371), .X(n23785) );
  nand_x1_sg U54008 ( .A(reg_www_15[10]), .B(n31889), .X(n23786) );
  nand_x1_sg U54009 ( .A(reg_ww_15[10]), .B(n35350), .X(n23787) );
  nand_x1_sg U54010 ( .A(reg_www_15[11]), .B(n32040), .X(n23788) );
  nand_x1_sg U54011 ( .A(reg_ww_15[11]), .B(n35210), .X(n23789) );
  nand_x1_sg U54012 ( .A(reg_www_15[12]), .B(n30599), .X(n23790) );
  nand_x1_sg U54013 ( .A(reg_ww_15[12]), .B(n31058), .X(n23791) );
  nand_x1_sg U54014 ( .A(reg_www_15[13]), .B(n32045), .X(n23792) );
  nand_x1_sg U54015 ( .A(reg_ww_15[13]), .B(n32754), .X(n23793) );
  nand_x1_sg U54016 ( .A(reg_www_15[14]), .B(n32283), .X(n23794) );
  nand_x1_sg U54017 ( .A(reg_ww_15[14]), .B(n32718), .X(n23795) );
  nand_x1_sg U54018 ( .A(reg_www_15[15]), .B(n33948), .X(n23796) );
  nand_x1_sg U54019 ( .A(reg_ww_15[15]), .B(n30705), .X(n23797) );
  nand_x1_sg U54020 ( .A(reg_www_15[16]), .B(n31723), .X(n23798) );
  nand_x1_sg U54021 ( .A(reg_ww_15[16]), .B(n31094), .X(n23799) );
  nand_x1_sg U54022 ( .A(reg_www_15[17]), .B(n32352), .X(n23800) );
  nand_x1_sg U54023 ( .A(reg_ww_15[17]), .B(n31674), .X(n23801) );
  nand_x1_sg U54024 ( .A(reg_www_15[18]), .B(n32312), .X(n23802) );
  nand_x1_sg U54025 ( .A(reg_ww_15[18]), .B(n31037), .X(n23803) );
  nand_x1_sg U54026 ( .A(reg_www_15[19]), .B(n32339), .X(n23804) );
  nand_x1_sg U54027 ( .A(reg_ww_15[19]), .B(n30592), .X(n23805) );
  nand_x1_sg U54028 ( .A(reg_ii_0[0]), .B(n32321), .X(n25796) );
  nand_x1_sg U54029 ( .A(n30179), .B(reg_i_0[0]), .X(n25797) );
  nand_x1_sg U54030 ( .A(reg_ii_0[2]), .B(n31732), .X(n25800) );
  nand_x1_sg U54031 ( .A(n32719), .B(reg_i_0[2]), .X(n25801) );
  nand_x1_sg U54032 ( .A(reg_ii_0[3]), .B(n31511), .X(n25802) );
  nand_x1_sg U54033 ( .A(n31207), .B(reg_i_0[3]), .X(n25803) );
  nand_x1_sg U54034 ( .A(reg_ii_0[5]), .B(n33971), .X(n25806) );
  nand_x1_sg U54035 ( .A(n35185), .B(reg_i_0[5]), .X(n25807) );
  nand_x1_sg U54036 ( .A(reg_ii_0[6]), .B(n32454), .X(n25808) );
  nand_x1_sg U54037 ( .A(n32728), .B(reg_i_0[6]), .X(n25809) );
  nand_x1_sg U54038 ( .A(reg_ii_0[8]), .B(n31631), .X(n25812) );
  nand_x1_sg U54039 ( .A(n33999), .B(reg_i_0[8]), .X(n25813) );
  nand_x1_sg U54040 ( .A(reg_ii_0[9]), .B(n34571), .X(n25814) );
  nand_x1_sg U54041 ( .A(n35376), .B(reg_i_0[9]), .X(n25815) );
  nand_x1_sg U54042 ( .A(reg_ii_0[11]), .B(n31888), .X(n25818) );
  nand_x1_sg U54043 ( .A(n34004), .B(reg_i_0[11]), .X(n25819) );
  nand_x1_sg U54044 ( .A(reg_ii_0[12]), .B(n31721), .X(n25820) );
  nand_x1_sg U54045 ( .A(n30863), .B(reg_i_0[12]), .X(n25821) );
  nand_x1_sg U54046 ( .A(reg_ii_0[14]), .B(n32016), .X(n25824) );
  nand_x1_sg U54047 ( .A(n30171), .B(reg_i_0[14]), .X(n25825) );
  nand_x1_sg U54048 ( .A(reg_ii_0[15]), .B(n31711), .X(n25826) );
  nand_x1_sg U54049 ( .A(n31671), .B(reg_i_0[15]), .X(n25827) );
  nand_x1_sg U54050 ( .A(reg_ii_0[17]), .B(n34571), .X(n25830) );
  nand_x1_sg U54051 ( .A(n32845), .B(reg_i_0[17]), .X(n25831) );
  nand_x1_sg U54052 ( .A(reg_ii_0[18]), .B(n34583), .X(n25832) );
  nand_x1_sg U54053 ( .A(n29757), .B(reg_i_0[18]), .X(n25833) );
  nand_x1_sg U54054 ( .A(reg_ii_3[15]), .B(n31711), .X(n26066) );
  nand_x1_sg U54055 ( .A(n35395), .B(reg_i_3[15]), .X(n26067) );
  nand_x1_sg U54056 ( .A(reg_ii_3[17]), .B(n32330), .X(n26070) );
  nand_x1_sg U54057 ( .A(n32712), .B(reg_i_3[17]), .X(n26071) );
  nand_x1_sg U54058 ( .A(reg_ii_3[18]), .B(n32295), .X(n26072) );
  nand_x1_sg U54059 ( .A(n35090), .B(reg_i_3[18]), .X(n26073) );
  nand_x1_sg U54060 ( .A(reg_ii_4[1]), .B(n32772), .X(n26118) );
  nand_x1_sg U54061 ( .A(n35227), .B(reg_i_4[1]), .X(n26119) );
  nand_x1_sg U54062 ( .A(reg_ii_4[2]), .B(n30140), .X(n26120) );
  nand_x1_sg U54063 ( .A(n34001), .B(reg_i_4[2]), .X(n26121) );
  nand_x1_sg U54064 ( .A(reg_ii_4[4]), .B(n32252), .X(n26124) );
  nand_x1_sg U54065 ( .A(n34006), .B(reg_i_4[4]), .X(n26125) );
  nand_x1_sg U54066 ( .A(reg_ii_4[5]), .B(n31909), .X(n26126) );
  nand_x1_sg U54067 ( .A(n32845), .B(reg_i_4[5]), .X(n26127) );
  nand_x1_sg U54068 ( .A(reg_ii_6[5]), .B(n32335), .X(n25490) );
  nand_x1_sg U54069 ( .A(n32728), .B(reg_i_6[5]), .X(n25491) );
  nand_x1_sg U54070 ( .A(reg_ii_6[7]), .B(n30176), .X(n25494) );
  nand_x1_sg U54071 ( .A(n31689), .B(reg_i_6[7]), .X(n25495) );
  nand_x1_sg U54072 ( .A(reg_ii_6[8]), .B(n32771), .X(n25496) );
  nand_x1_sg U54073 ( .A(n35087), .B(reg_i_6[8]), .X(n25497) );
  nand_x1_sg U54074 ( .A(reg_ii_6[10]), .B(n31733), .X(n25500) );
  nand_x1_sg U54075 ( .A(n35208), .B(reg_i_6[10]), .X(n25501) );
  nand_x1_sg U54076 ( .A(reg_ii_6[11]), .B(n32155), .X(n25502) );
  nand_x1_sg U54077 ( .A(n34701), .B(reg_i_6[11]), .X(n25503) );
  nand_x1_sg U54078 ( .A(reg_ii_6[13]), .B(n32453), .X(n25506) );
  nand_x1_sg U54079 ( .A(n31491), .B(reg_i_6[13]), .X(n25507) );
  nand_x1_sg U54080 ( .A(reg_ii_6[14]), .B(n31715), .X(n25508) );
  nand_x1_sg U54081 ( .A(n30594), .B(reg_i_6[14]), .X(n25509) );
  nand_x1_sg U54082 ( .A(reg_ii_6[16]), .B(n32251), .X(n25512) );
  nand_x1_sg U54083 ( .A(n31676), .B(reg_i_6[16]), .X(n25513) );
  nand_x1_sg U54084 ( .A(reg_ii_6[17]), .B(n32031), .X(n25514) );
  nand_x1_sg U54085 ( .A(n34716), .B(reg_i_6[17]), .X(n25515) );
  nand_x1_sg U54086 ( .A(reg_ii_6[19]), .B(n32352), .X(n25518) );
  nand_x1_sg U54087 ( .A(n31692), .B(reg_i_6[19]), .X(n25519) );
  nand_x1_sg U54088 ( .A(reg_ii_9[13]), .B(n32014), .X(n25746) );
  nand_x1_sg U54089 ( .A(n34092), .B(reg_i_9[13]), .X(n25747) );
  nand_x1_sg U54090 ( .A(reg_ii_9[14]), .B(n32770), .X(n25748) );
  nand_x1_sg U54091 ( .A(n32764), .B(reg_i_9[14]), .X(n25749) );
  nand_x1_sg U54092 ( .A(reg_ii_9[16]), .B(n32357), .X(n25752) );
  nand_x1_sg U54093 ( .A(n32753), .B(reg_i_9[16]), .X(n25753) );
  nand_x1_sg U54094 ( .A(reg_ii_9[17]), .B(n31501), .X(n25754) );
  nand_x1_sg U54095 ( .A(n34710), .B(reg_i_9[17]), .X(n25755) );
  nand_x1_sg U54096 ( .A(reg_ii_12[3]), .B(n32297), .X(n25170) );
  nand_x1_sg U54097 ( .A(n34722), .B(reg_i_12[3]), .X(n25171) );
  nand_x1_sg U54098 ( .A(reg_ii_12[4]), .B(n34573), .X(n25172) );
  nand_x1_sg U54099 ( .A(n29769), .B(reg_i_12[4]), .X(n25173) );
  nand_x1_sg U54100 ( .A(reg_ii_12[6]), .B(n32385), .X(n25176) );
  nand_x1_sg U54101 ( .A(n34007), .B(reg_i_12[6]), .X(n25177) );
  nand_x1_sg U54102 ( .A(reg_ii_12[7]), .B(n34570), .X(n25178) );
  nand_x1_sg U54103 ( .A(n35206), .B(reg_i_12[7]), .X(n25179) );
  nand_x1_sg U54104 ( .A(reg_ii_12[9]), .B(n33946), .X(n25182) );
  nand_x1_sg U54105 ( .A(n34000), .B(reg_i_12[9]), .X(n25183) );
  nand_x1_sg U54106 ( .A(reg_ii_12[10]), .B(n32158), .X(n25184) );
  nand_x1_sg U54107 ( .A(n34663), .B(reg_i_12[10]), .X(n25185) );
  nand_x1_sg U54108 ( .A(reg_ii_12[12]), .B(n32375), .X(n25188) );
  nand_x1_sg U54109 ( .A(n35351), .B(reg_i_12[12]), .X(n25189) );
  nand_x1_sg U54110 ( .A(reg_ii_12[13]), .B(n32028), .X(n25190) );
  nand_x1_sg U54111 ( .A(n32440), .B(reg_i_12[13]), .X(n25191) );
  nand_x1_sg U54112 ( .A(reg_ii_12[15]), .B(n32296), .X(n25194) );
  nand_x1_sg U54113 ( .A(n35189), .B(reg_i_12[15]), .X(n25195) );
  nand_x1_sg U54114 ( .A(reg_ii_12[16]), .B(n32330), .X(n25196) );
  nand_x1_sg U54115 ( .A(n34096), .B(reg_i_12[16]), .X(n25197) );
  nand_x1_sg U54116 ( .A(reg_ii_12[18]), .B(n32048), .X(n25200) );
  nand_x1_sg U54117 ( .A(n34058), .B(reg_i_12[18]), .X(n25201) );
  nand_x1_sg U54118 ( .A(reg_ii_12[19]), .B(n32138), .X(n25202) );
  nand_x1_sg U54119 ( .A(n35380), .B(reg_i_12[19]), .X(n25203) );
  nand_x1_sg U54120 ( .A(reg_ii_13[0]), .B(n33951), .X(n25244) );
  nand_x1_sg U54121 ( .A(n34056), .B(reg_i_13[0]), .X(n25245) );
  nand_x1_sg U54122 ( .A(reg_ii_13[2]), .B(n32286), .X(n25248) );
  nand_x1_sg U54123 ( .A(n35317), .B(reg_i_13[2]), .X(n25249) );
  nand_x1_sg U54124 ( .A(reg_ii_13[3]), .B(n34695), .X(n25250) );
  nand_x1_sg U54125 ( .A(n34663), .B(reg_i_13[3]), .X(n25251) );
  nand_x1_sg U54126 ( .A(reg_ii_13[5]), .B(n31715), .X(n25254) );
  nand_x1_sg U54127 ( .A(n32755), .B(reg_i_13[5]), .X(n25255) );
  nand_x1_sg U54128 ( .A(reg_ii_13[6]), .B(n35277), .X(n25256) );
  nand_x1_sg U54129 ( .A(n32754), .B(reg_i_13[6]), .X(n25257) );
  nand_x1_sg U54130 ( .A(reg_ii_13[8]), .B(n31745), .X(n25260) );
  nand_x1_sg U54131 ( .A(n34711), .B(reg_i_13[8]), .X(n25261) );
  nand_x1_sg U54132 ( .A(reg_ii_13[9]), .B(n32366), .X(n25262) );
  nand_x1_sg U54133 ( .A(n35213), .B(reg_i_13[9]), .X(n25263) );
  nand_x1_sg U54134 ( .A(reg_ii_13[11]), .B(n32285), .X(n25266) );
  nand_x1_sg U54135 ( .A(n31868), .B(reg_i_13[11]), .X(n25267) );
  nand_x1_sg U54136 ( .A(reg_ii_13[12]), .B(n31637), .X(n25268) );
  nand_x1_sg U54137 ( .A(n32721), .B(reg_i_13[12]), .X(n25269) );
  nand_x1_sg U54138 ( .A(reg_ii_13[14]), .B(n30621), .X(n25272) );
  nand_x1_sg U54139 ( .A(n30172), .B(reg_i_13[14]), .X(n25273) );
  nand_x1_sg U54140 ( .A(reg_ii_13[15]), .B(n34575), .X(n25274) );
  nand_x1_sg U54141 ( .A(n34000), .B(reg_i_13[15]), .X(n25275) );
  nand_x1_sg U54142 ( .A(reg_ii_13[17]), .B(n32140), .X(n25278) );
  nand_x1_sg U54143 ( .A(n35398), .B(reg_i_13[17]), .X(n25279) );
  nand_x1_sg U54144 ( .A(reg_ii_13[18]), .B(n30147), .X(n25280) );
  nand_x1_sg U54145 ( .A(n31864), .B(reg_i_13[18]), .X(n25281) );
  nand_x1_sg U54146 ( .A(reg_ii_14[17]), .B(n32015), .X(n24602) );
  nand_x1_sg U54147 ( .A(n30595), .B(reg_i_14[17]), .X(n24603) );
  nand_x1_sg U54148 ( .A(reg_ii_14[19]), .B(n32384), .X(n24606) );
  nand_x1_sg U54149 ( .A(n31872), .B(reg_i_14[19]), .X(n24607) );
  nand_x1_sg U54150 ( .A(reg_ii_15[0]), .B(n30623), .X(n24608) );
  nand_x1_sg U54151 ( .A(n32720), .B(reg_i_15[0]), .X(n24609) );
  nand_x1_sg U54152 ( .A(reg_ii_15[2]), .B(n32290), .X(n24612) );
  nand_x1_sg U54153 ( .A(n32718), .B(reg_i_15[2]), .X(n24613) );
  nand_x1_sg U54154 ( .A(reg_ii_15[3]), .B(n32857), .X(n24614) );
  nand_x1_sg U54155 ( .A(n34082), .B(reg_i_15[3]), .X(n24615) );
  nand_x1_sg U54156 ( .A(reg_ii_15[5]), .B(n32139), .X(n24618) );
  nand_x1_sg U54157 ( .A(n34078), .B(reg_i_15[5]), .X(n24619) );
  nand_x1_sg U54158 ( .A(reg_ii_15[6]), .B(n31926), .X(n24620) );
  nand_x1_sg U54159 ( .A(n32730), .B(reg_i_15[6]), .X(n24621) );
  nand_x1_sg U54160 ( .A(reg_ii_15[8]), .B(n32233), .X(n24624) );
  nand_x1_sg U54161 ( .A(n32714), .B(reg_i_15[8]), .X(n24625) );
  nand_x1_sg U54162 ( .A(reg_ii_15[9]), .B(n31637), .X(n24626) );
  nand_x1_sg U54163 ( .A(n35327), .B(reg_i_15[9]), .X(n24627) );
  nand_x1_sg U54164 ( .A(reg_ii_15[11]), .B(n32019), .X(n24630) );
  nand_x1_sg U54165 ( .A(n31690), .B(reg_i_15[11]), .X(n24631) );
  nand_x1_sg U54166 ( .A(reg_ii_15[12]), .B(n32378), .X(n24632) );
  nand_x1_sg U54167 ( .A(n34006), .B(reg_i_15[12]), .X(n24633) );
  nand_x1_sg U54168 ( .A(reg_ii_15[14]), .B(n32153), .X(n24636) );
  nand_x1_sg U54169 ( .A(n35370), .B(reg_i_15[14]), .X(n24637) );
  nand_x1_sg U54170 ( .A(reg_ii_15[15]), .B(n32241), .X(n24638) );
  nand_x1_sg U54171 ( .A(n35182), .B(reg_i_15[15]), .X(n24639) );
  nand_x1_sg U54172 ( .A(reg_ii_15[17]), .B(n32342), .X(n24642) );
  nand_x1_sg U54173 ( .A(n35206), .B(reg_i_15[17]), .X(n24643) );
  nand_x1_sg U54174 ( .A(reg_ii_15[18]), .B(n32451), .X(n24644) );
  nand_x1_sg U54175 ( .A(n32834), .B(reg_i_15[18]), .X(n24645) );
  nand_x1_sg U54176 ( .A(reg_ww_0[1]), .B(n34568), .X(n24690) );
  nand_x1_sg U54177 ( .A(n35362), .B(reg_w_0[1]), .X(n24691) );
  nand_x1_sg U54178 ( .A(reg_ww_0[2]), .B(n32450), .X(n24692) );
  nand_x1_sg U54179 ( .A(n34002), .B(reg_w_0[2]), .X(n24693) );
  nand_x1_sg U54180 ( .A(reg_ww_0[4]), .B(n31893), .X(n24696) );
  nand_x1_sg U54181 ( .A(n31672), .B(reg_w_0[4]), .X(n24697) );
  nand_x1_sg U54182 ( .A(reg_ww_0[5]), .B(n32154), .X(n24698) );
  nand_x1_sg U54183 ( .A(n35333), .B(reg_w_0[5]), .X(n24699) );
  nand_x1_sg U54184 ( .A(reg_ww_0[7]), .B(n32366), .X(n24702) );
  nand_x1_sg U54185 ( .A(n35356), .B(reg_w_0[7]), .X(n24703) );
  nand_x1_sg U54186 ( .A(reg_ww_0[8]), .B(n32254), .X(n24704) );
  nand_x1_sg U54187 ( .A(n32832), .B(reg_w_0[8]), .X(n24705) );
  nand_x1_sg U54188 ( .A(reg_ww_0[10]), .B(n32770), .X(n24708) );
  nand_x1_sg U54189 ( .A(n35083), .B(reg_w_0[10]), .X(n24709) );
  nand_x1_sg U54190 ( .A(reg_ww_0[11]), .B(n32035), .X(n24710) );
  nand_x1_sg U54191 ( .A(n30864), .B(reg_w_0[11]), .X(n24711) );
  nand_x1_sg U54192 ( .A(reg_ww_0[13]), .B(n32375), .X(n24714) );
  nand_x1_sg U54193 ( .A(n34095), .B(reg_w_0[13]), .X(n24715) );
  nand_x1_sg U54194 ( .A(reg_ww_0[14]), .B(n32367), .X(n24716) );
  nand_x1_sg U54195 ( .A(n29768), .B(reg_w_0[14]), .X(n24717) );
  nand_x1_sg U54196 ( .A(reg_ww_0[16]), .B(n32038), .X(n24720) );
  nand_x1_sg U54197 ( .A(n34712), .B(reg_w_0[16]), .X(n24721) );
  nand_x1_sg U54198 ( .A(reg_ww_3[1]), .B(n32331), .X(n24930) );
  nand_x1_sg U54199 ( .A(n35318), .B(reg_w_3[1]), .X(n24931) );
  nand_x1_sg U54200 ( .A(reg_ww_3[2]), .B(n30175), .X(n24932) );
  nand_x1_sg U54201 ( .A(n34721), .B(reg_w_3[2]), .X(n24933) );
  nand_x1_sg U54202 ( .A(reg_ww_3[4]), .B(n35277), .X(n24936) );
  nand_x1_sg U54203 ( .A(n35092), .B(reg_w_3[4]), .X(n24937) );
  nand_x1_sg U54204 ( .A(reg_ww_3[5]), .B(n32042), .X(n24938) );
  nand_x1_sg U54205 ( .A(n35231), .B(reg_w_3[5]), .X(n24939) );
  nand_x1_sg U54206 ( .A(reg_ww_3[7]), .B(n32050), .X(n24942) );
  nand_x1_sg U54207 ( .A(n35338), .B(reg_w_3[7]), .X(n24943) );
  nand_x1_sg U54208 ( .A(reg_ww_3[8]), .B(n31888), .X(n24944) );
  nand_x1_sg U54209 ( .A(n35163), .B(reg_w_3[8]), .X(n24945) );
  nand_x1_sg U54210 ( .A(reg_ww_3[10]), .B(n32494), .X(n24948) );
  nand_x1_sg U54211 ( .A(n34000), .B(reg_w_3[10]), .X(n24949) );
  nand_x1_sg U54212 ( .A(reg_ww_3[11]), .B(n32049), .X(n24950) );
  nand_x1_sg U54213 ( .A(n35215), .B(reg_w_3[11]), .X(n24951) );
  nand_x1_sg U54214 ( .A(reg_ww_3[13]), .B(n34576), .X(n24954) );
  nand_x1_sg U54215 ( .A(n35356), .B(reg_w_3[13]), .X(n24955) );
  nand_x1_sg U54216 ( .A(reg_ww_3[14]), .B(n35079), .X(n24956) );
  nand_x1_sg U54217 ( .A(n32837), .B(reg_w_3[14]), .X(n24957) );
  nand_x1_sg U54218 ( .A(reg_ww_6[0]), .B(n32233), .X(n24372) );
  nand_x1_sg U54219 ( .A(n35396), .B(reg_w_6[0]), .X(n24373) );
  nand_x1_sg U54220 ( .A(reg_ww_6[1]), .B(n30914), .X(n24374) );
  nand_x1_sg U54221 ( .A(n35087), .B(reg_w_6[1]), .X(n24375) );
  nand_x1_sg U54222 ( .A(reg_ww_6[3]), .B(n31735), .X(n24378) );
  nand_x1_sg U54223 ( .A(n35359), .B(reg_w_6[3]), .X(n24379) );
  nand_x1_sg U54224 ( .A(reg_ww_6[4]), .B(n32315), .X(n24380) );
  nand_x1_sg U54225 ( .A(n32752), .B(reg_w_6[4]), .X(n24381) );
  nand_x1_sg U54226 ( .A(reg_ww_6[6]), .B(n30197), .X(n24384) );
  nand_x1_sg U54227 ( .A(n34048), .B(reg_w_6[6]), .X(n24385) );
  nand_x1_sg U54228 ( .A(reg_ww_6[7]), .B(n34695), .X(n24386) );
  nand_x1_sg U54229 ( .A(n35171), .B(reg_w_6[7]), .X(n24387) );
  nand_x1_sg U54230 ( .A(reg_ww_6[9]), .B(n32155), .X(n24390) );
  nand_x1_sg U54231 ( .A(n34082), .B(reg_w_6[9]), .X(n24391) );
  nand_x1_sg U54232 ( .A(reg_ww_6[10]), .B(n31716), .X(n24392) );
  nand_x1_sg U54233 ( .A(n34047), .B(reg_w_6[10]), .X(n24393) );
  nand_x1_sg U54234 ( .A(reg_ww_6[12]), .B(n34897), .X(n24396) );
  nand_x1_sg U54235 ( .A(n34006), .B(reg_w_6[12]), .X(n24397) );
  nand_x1_sg U54236 ( .A(reg_ww_6[13]), .B(n32857), .X(n24398) );
  nand_x1_sg U54237 ( .A(n35202), .B(reg_w_6[13]), .X(n24399) );
  nand_x1_sg U54238 ( .A(reg_ww_8[16]), .B(n34567), .X(n23808) );
  nand_x1_sg U54239 ( .A(n35332), .B(reg_w_8[16]), .X(n23809) );
  nand_x1_sg U54240 ( .A(reg_ww_8[17]), .B(n32154), .X(n23810) );
  nand_x1_sg U54241 ( .A(n34058), .B(reg_w_8[17]), .X(n23811) );
  nand_x1_sg U54242 ( .A(reg_ww_8[19]), .B(n31720), .X(n23814) );
  nand_x1_sg U54243 ( .A(n35227), .B(reg_w_8[19]), .X(n23815) );
  nand_x1_sg U54244 ( .A(reg_ww_9[0]), .B(n32354), .X(n23816) );
  nand_x1_sg U54245 ( .A(n31676), .B(reg_w_9[0]), .X(n23817) );
  nand_x1_sg U54246 ( .A(reg_ww_9[2]), .B(n32158), .X(n23820) );
  nand_x1_sg U54247 ( .A(n35339), .B(reg_w_9[2]), .X(n23821) );
  nand_x1_sg U54248 ( .A(reg_ww_9[3]), .B(n32234), .X(n23822) );
  nand_x1_sg U54249 ( .A(n35160), .B(reg_w_9[3]), .X(n23823) );
  nand_x1_sg U54250 ( .A(reg_ww_12[0]), .B(n30622), .X(n24056) );
  nand_x1_sg U54251 ( .A(n35083), .B(reg_w_12[0]), .X(n24057) );
  nand_x1_sg U54252 ( .A(reg_ww_12[2]), .B(n33982), .X(n24060) );
  nand_x1_sg U54253 ( .A(n35240), .B(reg_w_12[2]), .X(n24061) );
  nand_x1_sg U54254 ( .A(reg_ww_12[3]), .B(n30621), .X(n24062) );
  nand_x1_sg U54255 ( .A(n32723), .B(reg_w_12[3]), .X(n24063) );
  nand_x1_sg U54256 ( .A(reg_ww_12[5]), .B(n31501), .X(n24066) );
  nand_x1_sg U54257 ( .A(n31871), .B(reg_w_12[5]), .X(n24067) );
  nand_x1_sg U54258 ( .A(reg_ww_12[6]), .B(n32372), .X(n24068) );
  nand_x1_sg U54259 ( .A(n35224), .B(reg_w_12[6]), .X(n24069) );
  nand_x1_sg U54260 ( .A(reg_ww_12[8]), .B(n31888), .X(n24072) );
  nand_x1_sg U54261 ( .A(n34718), .B(reg_w_12[8]), .X(n24073) );
  nand_x1_sg U54262 ( .A(reg_ww_12[9]), .B(n35078), .X(n24074) );
  nand_x1_sg U54263 ( .A(n32709), .B(reg_w_12[9]), .X(n24075) );
  nand_x1_sg U54264 ( .A(reg_ww_12[11]), .B(n32226), .X(n24078) );
  nand_x1_sg U54265 ( .A(n35347), .B(reg_w_12[11]), .X(n24079) );
  nand_x1_sg U54266 ( .A(reg_ww_12[12]), .B(n33947), .X(n24080) );
  nand_x1_sg U54267 ( .A(n32712), .B(reg_w_12[12]), .X(n24081) );
  nand_x1_sg U54268 ( .A(reg_ww_12[14]), .B(n34894), .X(n24084) );
  nand_x1_sg U54269 ( .A(n34050), .B(reg_w_12[14]), .X(n24085) );
  nand_x1_sg U54270 ( .A(reg_ww_12[15]), .B(n34577), .X(n24086) );
  nand_x1_sg U54271 ( .A(n35187), .B(reg_w_12[15]), .X(n24087) );
  nand_x1_sg U54272 ( .A(reg_ww_12[17]), .B(n32337), .X(n24090) );
  nand_x1_sg U54273 ( .A(n35370), .B(reg_w_12[17]), .X(n24091) );
  nand_x1_sg U54274 ( .A(reg_ww_12[18]), .B(n32236), .X(n24092) );
  nand_x1_sg U54275 ( .A(n32443), .B(reg_w_12[18]), .X(n24093) );
  nand_x1_sg U54276 ( .A(reg_ww_13[1]), .B(n30195), .X(n24138) );
  nand_x1_sg U54277 ( .A(n34084), .B(reg_w_13[1]), .X(n24139) );
  nand_x1_sg U54278 ( .A(reg_ww_13[2]), .B(n32306), .X(n24140) );
  nand_x1_sg U54279 ( .A(n35201), .B(reg_w_13[2]), .X(n24141) );
  nand_x1_sg U54280 ( .A(reg_ww_13[4]), .B(n32165), .X(n24144) );
  nand_x1_sg U54281 ( .A(n35094), .B(reg_w_13[4]), .X(n24145) );
  nand_x1_sg U54282 ( .A(reg_ww_15[18]), .B(n32403), .X(n23762) );
  nand_x1_sg U54283 ( .A(n35213), .B(reg_w_15[18]), .X(n23763) );
  nand_x1_sg U54284 ( .A(reg_ii_0[1]), .B(n32379), .X(n25798) );
  nand_x1_sg U54285 ( .A(n35335), .B(reg_i_0[1]), .X(n25799) );
  nand_x1_sg U54286 ( .A(reg_ii_0[4]), .B(n32164), .X(n25804) );
  nand_x1_sg U54287 ( .A(n34073), .B(reg_i_0[4]), .X(n25805) );
  nand_x1_sg U54288 ( .A(reg_ii_0[7]), .B(n31513), .X(n25810) );
  nand_x1_sg U54289 ( .A(n34723), .B(reg_i_0[7]), .X(n25811) );
  nand_x1_sg U54290 ( .A(reg_ii_0[10]), .B(n30196), .X(n25816) );
  nand_x1_sg U54291 ( .A(n34053), .B(reg_i_0[10]), .X(n25817) );
  nand_x1_sg U54292 ( .A(reg_ii_0[13]), .B(n32344), .X(n25822) );
  nand_x1_sg U54293 ( .A(n32441), .B(reg_i_0[13]), .X(n25823) );
  nand_x1_sg U54294 ( .A(reg_ii_0[16]), .B(n32050), .X(n25828) );
  nand_x1_sg U54295 ( .A(n31689), .B(reg_i_0[16]), .X(n25829) );
  nand_x1_sg U54296 ( .A(reg_ii_0[19]), .B(n31904), .X(n25834) );
  nand_x1_sg U54297 ( .A(n34080), .B(reg_i_0[19]), .X(n25835) );
  nand_x1_sg U54298 ( .A(reg_ii_3[16]), .B(n32775), .X(n26068) );
  nand_x1_sg U54299 ( .A(n32721), .B(reg_i_3[16]), .X(n26069) );
  nand_x1_sg U54300 ( .A(reg_ii_3[19]), .B(n33976), .X(n26074) );
  nand_x1_sg U54301 ( .A(n34005), .B(reg_i_3[19]), .X(n26075) );
  nand_x1_sg U54302 ( .A(reg_ii_4[0]), .B(n32407), .X(n26116) );
  nand_x1_sg U54303 ( .A(n35093), .B(reg_i_4[0]), .X(n26117) );
  nand_x1_sg U54304 ( .A(reg_ii_4[3]), .B(n32776), .X(n26122) );
  nand_x1_sg U54305 ( .A(n35204), .B(reg_i_4[3]), .X(n26123) );
  nand_x1_sg U54306 ( .A(reg_ii_4[6]), .B(n32371), .X(n26128) );
  nand_x1_sg U54307 ( .A(n32834), .B(reg_i_4[6]), .X(n26129) );
  nand_x1_sg U54308 ( .A(reg_ii_6[6]), .B(n32242), .X(n25492) );
  nand_x1_sg U54309 ( .A(n34724), .B(reg_i_6[6]), .X(n25493) );
  nand_x1_sg U54310 ( .A(reg_ii_6[9]), .B(n32010), .X(n25498) );
  nand_x1_sg U54311 ( .A(n35088), .B(reg_i_6[9]), .X(n25499) );
  nand_x1_sg U54312 ( .A(reg_ii_6[12]), .B(n32302), .X(n25504) );
  nand_x1_sg U54313 ( .A(n30177), .B(reg_i_6[12]), .X(n25505) );
  nand_x1_sg U54314 ( .A(reg_ii_6[15]), .B(n30155), .X(n25510) );
  nand_x1_sg U54315 ( .A(n31676), .B(reg_i_6[15]), .X(n25511) );
  nand_x1_sg U54316 ( .A(reg_ii_6[18]), .B(n34852), .X(n25516) );
  nand_x1_sg U54317 ( .A(n34053), .B(reg_i_6[18]), .X(n25517) );
  nand_x1_sg U54318 ( .A(reg_ii_9[15]), .B(n32407), .X(n25750) );
  nand_x1_sg U54319 ( .A(n35185), .B(reg_i_9[15]), .X(n25751) );
  nand_x1_sg U54320 ( .A(reg_ii_12[5]), .B(n31634), .X(n25174) );
  nand_x1_sg U54321 ( .A(n29762), .B(reg_i_12[5]), .X(n25175) );
  nand_x1_sg U54322 ( .A(reg_ii_12[8]), .B(n32311), .X(n25180) );
  nand_x1_sg U54323 ( .A(n34007), .B(reg_i_12[8]), .X(n25181) );
  nand_x1_sg U54324 ( .A(reg_ii_12[11]), .B(n31515), .X(n25186) );
  nand_x1_sg U54325 ( .A(n35204), .B(reg_i_12[11]), .X(n25187) );
  nand_x1_sg U54326 ( .A(reg_ii_12[14]), .B(n32306), .X(n25192) );
  nand_x1_sg U54327 ( .A(n34095), .B(reg_i_12[14]), .X(n25193) );
  nand_x1_sg U54328 ( .A(reg_ii_12[17]), .B(n32383), .X(n25198) );
  nand_x1_sg U54329 ( .A(n32767), .B(reg_i_12[17]), .X(n25199) );
  nand_x1_sg U54330 ( .A(reg_ii_13[1]), .B(n32376), .X(n25246) );
  nand_x1_sg U54331 ( .A(n31673), .B(reg_i_13[1]), .X(n25247) );
  nand_x1_sg U54332 ( .A(reg_ii_13[4]), .B(n33945), .X(n25252) );
  nand_x1_sg U54333 ( .A(n30178), .B(reg_i_13[4]), .X(n25253) );
  nand_x1_sg U54334 ( .A(reg_ii_13[7]), .B(n32363), .X(n25258) );
  nand_x1_sg U54335 ( .A(n35236), .B(reg_i_13[7]), .X(n25259) );
  nand_x1_sg U54336 ( .A(reg_ii_13[10]), .B(n32227), .X(n25264) );
  nand_x1_sg U54337 ( .A(n31675), .B(reg_i_13[10]), .X(n25265) );
  nand_x1_sg U54338 ( .A(reg_ii_13[13]), .B(n33982), .X(n25270) );
  nand_x1_sg U54339 ( .A(n32716), .B(reg_i_13[13]), .X(n25271) );
  nand_x1_sg U54340 ( .A(reg_ii_13[16]), .B(n32288), .X(n25276) );
  nand_x1_sg U54341 ( .A(n35179), .B(reg_i_13[16]), .X(n25277) );
  nand_x1_sg U54342 ( .A(reg_ii_13[19]), .B(n32310), .X(n25282) );
  nand_x1_sg U54343 ( .A(n35218), .B(reg_i_13[19]), .X(n25283) );
  nand_x1_sg U54344 ( .A(reg_ii_14[18]), .B(n32316), .X(n24604) );
  nand_x1_sg U54345 ( .A(n34045), .B(reg_i_14[18]), .X(n24605) );
  nand_x1_sg U54346 ( .A(reg_ii_15[1]), .B(n30918), .X(n24610) );
  nand_x1_sg U54347 ( .A(n35177), .B(reg_i_15[1]), .X(n24611) );
  nand_x1_sg U54348 ( .A(reg_ii_15[4]), .B(n32373), .X(n24616) );
  nand_x1_sg U54349 ( .A(n34713), .B(reg_i_15[4]), .X(n24617) );
  nand_x1_sg U54350 ( .A(reg_ii_15[7]), .B(n30611), .X(n24622) );
  nand_x1_sg U54351 ( .A(n35341), .B(reg_i_15[7]), .X(n24623) );
  nand_x1_sg U54352 ( .A(reg_ii_15[10]), .B(n32293), .X(n24628) );
  nand_x1_sg U54353 ( .A(n34002), .B(reg_i_15[10]), .X(n24629) );
  nand_x1_sg U54354 ( .A(reg_ii_15[13]), .B(n32494), .X(n24634) );
  nand_x1_sg U54355 ( .A(n32844), .B(reg_i_15[13]), .X(n24635) );
  nand_x1_sg U54356 ( .A(reg_ii_15[16]), .B(n32332), .X(n24640) );
  nand_x1_sg U54357 ( .A(n35361), .B(reg_i_15[16]), .X(n24641) );
  nand_x1_sg U54358 ( .A(reg_ii_15[19]), .B(n31737), .X(n24646) );
  nand_x1_sg U54359 ( .A(n31674), .B(reg_i_15[19]), .X(n24647) );
  nand_x1_sg U54360 ( .A(reg_ww_0[0]), .B(n32027), .X(n24688) );
  nand_x1_sg U54361 ( .A(n35181), .B(reg_w_0[0]), .X(n24689) );
  nand_x1_sg U54362 ( .A(reg_ww_0[3]), .B(n31649), .X(n24694) );
  nand_x1_sg U54363 ( .A(n35234), .B(reg_w_0[3]), .X(n24695) );
  nand_x1_sg U54364 ( .A(reg_ww_0[6]), .B(n32041), .X(n24700) );
  nand_x1_sg U54365 ( .A(n35165), .B(reg_w_0[6]), .X(n24701) );
  nand_x1_sg U54366 ( .A(reg_ww_0[9]), .B(n30207), .X(n24706) );
  nand_x1_sg U54367 ( .A(n35367), .B(reg_w_0[9]), .X(n24707) );
  nand_x1_sg U54368 ( .A(reg_ww_0[12]), .B(n32355), .X(n24712) );
  nand_x1_sg U54369 ( .A(n35212), .B(reg_w_0[12]), .X(n24713) );
  nand_x1_sg U54370 ( .A(reg_ww_0[15]), .B(n33967), .X(n24718) );
  nand_x1_sg U54371 ( .A(n32748), .B(reg_w_0[15]), .X(n24719) );
  nand_x1_sg U54372 ( .A(reg_ww_3[0]), .B(n34847), .X(n24928) );
  nand_x1_sg U54373 ( .A(n32720), .B(reg_w_3[0]), .X(n24929) );
  nand_x1_sg U54374 ( .A(reg_ww_3[3]), .B(n32367), .X(n24934) );
  nand_x1_sg U54375 ( .A(n30171), .B(reg_w_3[3]), .X(n24935) );
  nand_x1_sg U54376 ( .A(reg_ww_3[6]), .B(n30140), .X(n24940) );
  nand_x1_sg U54377 ( .A(n34051), .B(reg_w_3[6]), .X(n24941) );
  nand_x1_sg U54378 ( .A(reg_ww_3[9]), .B(n31735), .X(n24946) );
  nand_x1_sg U54379 ( .A(n34055), .B(reg_w_3[9]), .X(n24947) );
  nand_x1_sg U54380 ( .A(reg_ww_3[12]), .B(n34575), .X(n24952) );
  nand_x1_sg U54381 ( .A(n34083), .B(reg_w_3[12]), .X(n24953) );
  nand_x1_sg U54382 ( .A(reg_ww_3[15]), .B(n31649), .X(n24958) );
  nand_x1_sg U54383 ( .A(n32713), .B(reg_w_3[15]), .X(n24959) );
  nand_x1_sg U54384 ( .A(reg_ww_6[2]), .B(n33948), .X(n24376) );
  nand_x1_sg U54385 ( .A(n34701), .B(reg_w_6[2]), .X(n24377) );
  nand_x1_sg U54386 ( .A(reg_ww_6[5]), .B(n32014), .X(n24382) );
  nand_x1_sg U54387 ( .A(n32742), .B(reg_w_6[5]), .X(n24383) );
  nand_x1_sg U54388 ( .A(reg_ww_6[8]), .B(n34696), .X(n24388) );
  nand_x1_sg U54389 ( .A(n35216), .B(reg_w_6[8]), .X(n24389) );
  nand_x1_sg U54390 ( .A(reg_ww_6[11]), .B(n31633), .X(n24394) );
  nand_x1_sg U54391 ( .A(n32729), .B(reg_w_6[11]), .X(n24395) );
  nand_x1_sg U54392 ( .A(reg_ww_6[14]), .B(n34652), .X(n24400) );
  nand_x1_sg U54393 ( .A(n35191), .B(reg_w_6[14]), .X(n24401) );
  nand_x1_sg U54394 ( .A(reg_ww_8[15]), .B(n32243), .X(n23806) );
  nand_x1_sg U54395 ( .A(n32709), .B(reg_w_8[15]), .X(n23807) );
  nand_x1_sg U54396 ( .A(reg_ww_8[18]), .B(n32038), .X(n23812) );
  nand_x1_sg U54397 ( .A(n31691), .B(reg_w_8[18]), .X(n23813) );
  nand_x1_sg U54398 ( .A(reg_ww_9[1]), .B(n32307), .X(n23818) );
  nand_x1_sg U54399 ( .A(n35082), .B(reg_w_9[1]), .X(n23819) );
  nand_x1_sg U54400 ( .A(reg_ww_9[4]), .B(n30213), .X(n23824) );
  nand_x1_sg U54401 ( .A(n34072), .B(reg_w_9[4]), .X(n23825) );
  nand_x1_sg U54402 ( .A(reg_ww_12[1]), .B(n31732), .X(n24058) );
  nand_x1_sg U54403 ( .A(n34078), .B(reg_w_12[1]), .X(n24059) );
  nand_x1_sg U54404 ( .A(reg_ww_12[4]), .B(n32380), .X(n24064) );
  nand_x1_sg U54405 ( .A(n35201), .B(reg_w_12[4]), .X(n24065) );
  nand_x1_sg U54406 ( .A(reg_ww_12[7]), .B(n31740), .X(n24070) );
  nand_x1_sg U54407 ( .A(n34080), .B(reg_w_12[7]), .X(n24071) );
  nand_x1_sg U54408 ( .A(reg_ww_12[10]), .B(n31893), .X(n24076) );
  nand_x1_sg U54409 ( .A(n34704), .B(reg_w_12[10]), .X(n24077) );
  nand_x1_sg U54410 ( .A(reg_ww_12[13]), .B(n32379), .X(n24082) );
  nand_x1_sg U54411 ( .A(n31689), .B(reg_w_12[13]), .X(n24083) );
  nand_x1_sg U54412 ( .A(reg_ww_12[16]), .B(n32451), .X(n24088) );
  nand_x1_sg U54413 ( .A(n30903), .B(reg_w_12[16]), .X(n24089) );
  nand_x1_sg U54414 ( .A(reg_ww_12[19]), .B(n31741), .X(n24094) );
  nand_x1_sg U54415 ( .A(n34666), .B(reg_w_12[19]), .X(n24095) );
  nand_x1_sg U54416 ( .A(reg_ww_13[0]), .B(n32348), .X(n24136) );
  nand_x1_sg U54417 ( .A(n31864), .B(reg_w_13[0]), .X(n24137) );
  nand_x1_sg U54418 ( .A(reg_ww_13[3]), .B(n32305), .X(n24142) );
  nand_x1_sg U54419 ( .A(n30179), .B(reg_w_13[3]), .X(n24143) );
  nand_x1_sg U54420 ( .A(reg_ww_15[19]), .B(n32293), .X(n23764) );
  nand_x1_sg U54421 ( .A(n35203), .B(reg_w_15[19]), .X(n23765) );
  nor_x1_sg U54422 ( .A(n30511), .B(n21320), .X(n21319) );
  nor_x1_sg U54423 ( .A(n30507), .B(n34992), .X(n21318) );
  nand_x1_sg U54424 ( .A(n42772), .B(n42773), .X(n21320) );
  nand_x1_sg U54425 ( .A(n31707), .B(n30540), .X(n20903) );
  nand_x1_sg U54426 ( .A(n20905), .B(n20906), .X(n20902) );
  nor_x1_sg U54427 ( .A(n20907), .B(n20908), .X(n20905) );
  nand_x1_sg U54428 ( .A(n31659), .B(n30540), .X(n20933) );
  nand_x1_sg U54429 ( .A(n20906), .B(n20935), .X(n20934) );
  nand_x1_sg U54430 ( .A(n20936), .B(n20937), .X(n20935) );
  nand_x1_sg U54431 ( .A(n31597), .B(n21326), .X(n21346) );
  nand_x1_sg U54432 ( .A(n21327), .B(n21347), .X(n21345) );
  nand_x1_sg U54433 ( .A(n21348), .B(n21349), .X(n21347) );
  nand_x1_sg U54434 ( .A(n31595), .B(n21326), .X(n21369) );
  nand_x1_sg U54435 ( .A(n21327), .B(n21371), .X(n21368) );
  nor_x1_sg U54436 ( .A(n30449), .B(n21740), .X(n21739) );
  nor_x1_sg U54437 ( .A(n30445), .B(n35248), .X(n21738) );
  nand_x1_sg U54438 ( .A(n42655), .B(n42656), .X(n21740) );
  nand_x1_sg U54439 ( .A(n35457), .B(state[0]), .X(n22220) );
  nand_x1_sg U54440 ( .A(filter_output_shifter_input_taken), .B(n20894), .X(
        n29668) );
  nor_x1_sg U54441 ( .A(filter_state[0]), .B(n42531), .X(n20894) );
  nor_x1_sg U54442 ( .A(filter_state[1]), .B(filter_state[0]), .X(n28256) );
  nor_x1_sg U54443 ( .A(n42413), .B(n26584), .X(n28255) );
  inv_x1_sg U54444 ( .A(filter_state[1]), .X(n42531) );
  nand_x1_sg U54445 ( .A(n32007), .B(n26589), .X(\filter_0/n9633 ) );
  nand_x1_sg U54446 ( .A(n32784), .B(mask_output_filter_input_taken), .X(
        n26589) );
  nand_x1_sg U54447 ( .A(n33924), .B(n28147), .X(n28146) );
  nand_x1_sg U54448 ( .A(\filter_0/reg_xor_w_mask[10] ), .B(n32826), .X(n28145) );
  nand_x1_sg U54449 ( .A(n28148), .B(n42457), .X(n28147) );
  nand_x1_sg U54450 ( .A(n34019), .B(n28132), .X(n28131) );
  nand_x1_sg U54451 ( .A(\filter_0/reg_xor_w_mask[7] ), .B(n31915), .X(n28130)
         );
  nand_x1_sg U54452 ( .A(n28133), .B(n42454), .X(n28132) );
  nand_x1_sg U54453 ( .A(n34886), .B(n28117), .X(n28116) );
  nand_x1_sg U54454 ( .A(\filter_0/reg_xor_w_mask[4] ), .B(n32782), .X(n28115)
         );
  nand_x1_sg U54455 ( .A(n28118), .B(n42451), .X(n28117) );
  nand_x1_sg U54456 ( .A(n34912), .B(n28102), .X(n28101) );
  nand_x1_sg U54457 ( .A(\filter_0/reg_xor_w_mask[1] ), .B(n32807), .X(n28100)
         );
  nand_x1_sg U54458 ( .A(n28103), .B(n42448), .X(n28102) );
  nand_x1_sg U54459 ( .A(n30030), .B(n28087), .X(n28086) );
  nand_x1_sg U54460 ( .A(\filter_0/reg_xor_i_mask[30] ), .B(n32871), .X(n28085) );
  nand_x1_sg U54461 ( .A(n28088), .B(n42445), .X(n28087) );
  nand_x1_sg U54462 ( .A(n32258), .B(n28072), .X(n28071) );
  nand_x1_sg U54463 ( .A(\filter_0/reg_xor_i_mask[27] ), .B(n32483), .X(n28070) );
  nand_x1_sg U54464 ( .A(n28073), .B(n42442), .X(n28072) );
  nand_x1_sg U54465 ( .A(n32270), .B(n28057), .X(n28056) );
  nand_x1_sg U54466 ( .A(\filter_0/reg_xor_i_mask[24] ), .B(n32876), .X(n28055) );
  nand_x1_sg U54467 ( .A(n28058), .B(n42439), .X(n28057) );
  nand_x1_sg U54468 ( .A(n33906), .B(n28027), .X(n28026) );
  nand_x1_sg U54469 ( .A(\filter_0/reg_xor_i_mask[18] ), .B(n34677), .X(n28025) );
  nand_x1_sg U54470 ( .A(n28028), .B(n42433), .X(n28027) );
  nand_x1_sg U54471 ( .A(n31678), .B(n28012), .X(n28011) );
  nand_x1_sg U54472 ( .A(\filter_0/reg_xor_i_mask[15] ), .B(n34646), .X(n28010) );
  nand_x1_sg U54473 ( .A(n28013), .B(n42430), .X(n28012) );
  nand_x1_sg U54474 ( .A(n34906), .B(n27997), .X(n27996) );
  nand_x1_sg U54475 ( .A(\filter_0/reg_xor_i_mask[12] ), .B(n32801), .X(n27995) );
  nand_x1_sg U54476 ( .A(n27998), .B(n42427), .X(n27997) );
  nand_x1_sg U54477 ( .A(n33926), .B(n27982), .X(n27981) );
  nand_x1_sg U54478 ( .A(\filter_0/reg_xor_i_mask[9] ), .B(n32436), .X(n27980)
         );
  nand_x1_sg U54479 ( .A(n27983), .B(n42424), .X(n27982) );
  nand_x1_sg U54480 ( .A(n31681), .B(n27967), .X(n27966) );
  nand_x1_sg U54481 ( .A(\filter_0/reg_xor_i_mask[6] ), .B(n30166), .X(n27965)
         );
  nand_x1_sg U54482 ( .A(n27968), .B(n42421), .X(n27967) );
  nand_x1_sg U54483 ( .A(n31680), .B(n27952), .X(n27951) );
  nand_x1_sg U54484 ( .A(\filter_0/reg_xor_i_mask[3] ), .B(n32861), .X(n27950)
         );
  nand_x1_sg U54485 ( .A(n27953), .B(n42418), .X(n27952) );
  nand_x1_sg U54486 ( .A(n33938), .B(n28142), .X(n28141) );
  nand_x1_sg U54487 ( .A(\filter_0/reg_xor_w_mask[9] ), .B(n34687), .X(n28140)
         );
  nand_x1_sg U54488 ( .A(n28143), .B(n42456), .X(n28142) );
  nand_x1_sg U54489 ( .A(n33928), .B(n28137), .X(n28136) );
  nand_x1_sg U54490 ( .A(\filter_0/reg_xor_w_mask[8] ), .B(n34670), .X(n28135)
         );
  nand_x1_sg U54491 ( .A(n28138), .B(n42455), .X(n28137) );
  nand_x1_sg U54492 ( .A(n31677), .B(n28127), .X(n28126) );
  nand_x1_sg U54493 ( .A(\filter_0/reg_xor_w_mask[6] ), .B(n32434), .X(n28125)
         );
  nand_x1_sg U54494 ( .A(n28128), .B(n42453), .X(n28127) );
  nand_x1_sg U54495 ( .A(n34013), .B(n28122), .X(n28121) );
  nand_x1_sg U54496 ( .A(\filter_0/reg_xor_w_mask[5] ), .B(n30758), .X(n28120)
         );
  nand_x1_sg U54497 ( .A(n28123), .B(n42452), .X(n28122) );
  nand_x1_sg U54498 ( .A(n34014), .B(n28112), .X(n28111) );
  nand_x1_sg U54499 ( .A(\filter_0/reg_xor_w_mask[3] ), .B(n35070), .X(n28110)
         );
  nand_x1_sg U54500 ( .A(n28113), .B(n42450), .X(n28112) );
  nand_x1_sg U54501 ( .A(n33901), .B(n28107), .X(n28106) );
  nand_x1_sg U54502 ( .A(\filter_0/reg_xor_w_mask[2] ), .B(n30773), .X(n28105)
         );
  nand_x1_sg U54503 ( .A(n28108), .B(n42449), .X(n28107) );
  nand_x1_sg U54504 ( .A(n31686), .B(n28097), .X(n28096) );
  nand_x1_sg U54505 ( .A(\filter_0/reg_xor_w_mask[0] ), .B(n30765), .X(n28095)
         );
  nand_x1_sg U54506 ( .A(n28098), .B(n42447), .X(n28097) );
  nand_x1_sg U54507 ( .A(n33892), .B(n28092), .X(n28091) );
  nand_x1_sg U54508 ( .A(\filter_0/reg_xor_i_mask[31] ), .B(n30247), .X(n28090) );
  nand_x1_sg U54509 ( .A(n28093), .B(n42446), .X(n28092) );
  nand_x1_sg U54510 ( .A(n30033), .B(n28082), .X(n28081) );
  nand_x1_sg U54511 ( .A(\filter_0/reg_xor_i_mask[29] ), .B(n32866), .X(n28080) );
  nand_x1_sg U54512 ( .A(n28083), .B(n42444), .X(n28082) );
  nand_x1_sg U54513 ( .A(n32267), .B(n28077), .X(n28076) );
  nand_x1_sg U54514 ( .A(\filter_0/reg_xor_i_mask[28] ), .B(n30772), .X(n28075) );
  nand_x1_sg U54515 ( .A(n28078), .B(n42443), .X(n28077) );
  nand_x1_sg U54516 ( .A(n33921), .B(n28067), .X(n28066) );
  nand_x1_sg U54517 ( .A(\filter_0/reg_xor_i_mask[26] ), .B(n34682), .X(n28065) );
  nand_x1_sg U54518 ( .A(n28068), .B(n42441), .X(n28067) );
  nand_x1_sg U54519 ( .A(n33896), .B(n28062), .X(n28061) );
  nand_x1_sg U54520 ( .A(\filter_0/reg_xor_i_mask[25] ), .B(n32462), .X(n28060) );
  nand_x1_sg U54521 ( .A(n28063), .B(n42440), .X(n28062) );
  nand_x1_sg U54522 ( .A(n33894), .B(n28052), .X(n28051) );
  nand_x1_sg U54523 ( .A(\filter_0/reg_xor_i_mask[23] ), .B(n32490), .X(n28050) );
  nand_x1_sg U54524 ( .A(n28053), .B(n42438), .X(n28052) );
  nand_x1_sg U54525 ( .A(n31688), .B(n28047), .X(n28046) );
  nand_x1_sg U54526 ( .A(\filter_0/reg_xor_i_mask[22] ), .B(n32797), .X(n28045) );
  nand_x1_sg U54527 ( .A(n28048), .B(n42437), .X(n28047) );
  nand_x1_sg U54528 ( .A(n30034), .B(n28032), .X(n28031) );
  nand_x1_sg U54529 ( .A(\filter_0/reg_xor_i_mask[19] ), .B(n34634), .X(n28030) );
  nand_x1_sg U54530 ( .A(n28033), .B(n42434), .X(n28032) );
  nand_x1_sg U54531 ( .A(n33911), .B(n28022), .X(n28021) );
  nand_x1_sg U54532 ( .A(\filter_0/reg_xor_i_mask[17] ), .B(n34629), .X(n28020) );
  nand_x1_sg U54533 ( .A(n28023), .B(n42432), .X(n28022) );
  nand_x1_sg U54534 ( .A(n33918), .B(n28017), .X(n28016) );
  nand_x1_sg U54535 ( .A(\filter_0/reg_xor_i_mask[16] ), .B(n32469), .X(n28015) );
  nand_x1_sg U54536 ( .A(n28018), .B(n42431), .X(n28017) );
  nand_x1_sg U54537 ( .A(n35411), .B(n28007), .X(n28006) );
  nand_x1_sg U54538 ( .A(\filter_0/reg_xor_i_mask[14] ), .B(n30745), .X(n28005) );
  nand_x1_sg U54539 ( .A(n28008), .B(n42429), .X(n28007) );
  nand_x1_sg U54540 ( .A(n30205), .B(n28002), .X(n28001) );
  nand_x1_sg U54541 ( .A(\filter_0/reg_xor_i_mask[13] ), .B(n32430), .X(n28000) );
  nand_x1_sg U54542 ( .A(n28003), .B(n42428), .X(n28002) );
  nand_x1_sg U54543 ( .A(n33902), .B(n27992), .X(n27991) );
  nand_x1_sg U54544 ( .A(\filter_0/reg_xor_i_mask[11] ), .B(n32811), .X(n27990) );
  nand_x1_sg U54545 ( .A(n27993), .B(n42426), .X(n27992) );
  nand_x1_sg U54546 ( .A(n30036), .B(n27987), .X(n27986) );
  nand_x1_sg U54547 ( .A(\filter_0/reg_xor_i_mask[10] ), .B(n32476), .X(n27985) );
  nand_x1_sg U54548 ( .A(n27988), .B(n42425), .X(n27987) );
  nand_x1_sg U54549 ( .A(n34604), .B(n27977), .X(n27976) );
  nand_x1_sg U54550 ( .A(\filter_0/reg_xor_i_mask[8] ), .B(n32877), .X(n27975)
         );
  nand_x1_sg U54551 ( .A(n27978), .B(n42423), .X(n27977) );
  nand_x1_sg U54552 ( .A(n31683), .B(n27972), .X(n27971) );
  nand_x1_sg U54553 ( .A(\filter_0/reg_xor_i_mask[7] ), .B(n30762), .X(n27970)
         );
  nand_x1_sg U54554 ( .A(n27973), .B(n42422), .X(n27972) );
  nand_x1_sg U54555 ( .A(n34018), .B(n27962), .X(n27961) );
  nand_x1_sg U54556 ( .A(\filter_0/reg_xor_i_mask[5] ), .B(n32881), .X(n27960)
         );
  nand_x1_sg U54557 ( .A(n27963), .B(n42420), .X(n27962) );
  nand_x1_sg U54558 ( .A(n33929), .B(n27957), .X(n27956) );
  nand_x1_sg U54559 ( .A(\filter_0/reg_xor_i_mask[4] ), .B(n34692), .X(n27955)
         );
  nand_x1_sg U54560 ( .A(n27958), .B(n42419), .X(n27957) );
  nand_x1_sg U54561 ( .A(n34911), .B(n27947), .X(n27946) );
  nand_x1_sg U54562 ( .A(\filter_0/reg_xor_i_mask[2] ), .B(n32821), .X(n27945)
         );
  nand_x1_sg U54563 ( .A(n27948), .B(n42417), .X(n27947) );
  nand_x1_sg U54564 ( .A(n29692), .B(reg_www_15[19]), .X(n27869) );
  nand_x1_sg U54565 ( .A(\filter_0/reg_w_15[19] ), .B(n32438), .X(n27870) );
  nand_x1_sg U54566 ( .A(n30935), .B(reg_www_15[18]), .X(n27867) );
  nand_x1_sg U54567 ( .A(\filter_0/reg_w_15[18] ), .B(n32483), .X(n27868) );
  nand_x1_sg U54568 ( .A(n30923), .B(reg_www_15[17]), .X(n27865) );
  nand_x1_sg U54569 ( .A(\filter_0/reg_w_15[17] ), .B(n32800), .X(n27866) );
  nand_x1_sg U54570 ( .A(n34602), .B(reg_www_15[16]), .X(n27863) );
  nand_x1_sg U54571 ( .A(\filter_0/reg_w_15[16] ), .B(n32489), .X(n27864) );
  nand_x1_sg U54572 ( .A(n29694), .B(reg_www_15[15]), .X(n27861) );
  nand_x1_sg U54573 ( .A(\filter_0/reg_w_15[15] ), .B(n32874), .X(n27862) );
  nand_x1_sg U54574 ( .A(n34039), .B(reg_www_15[14]), .X(n27859) );
  nand_x1_sg U54575 ( .A(\filter_0/reg_w_15[14] ), .B(n32458), .X(n27860) );
  nand_x1_sg U54576 ( .A(n34024), .B(reg_www_15[13]), .X(n27857) );
  nand_x1_sg U54577 ( .A(\filter_0/reg_w_15[13] ), .B(n34670), .X(n27858) );
  nand_x1_sg U54578 ( .A(n31530), .B(reg_www_15[12]), .X(n27855) );
  nand_x1_sg U54579 ( .A(\filter_0/reg_w_15[12] ), .B(n32457), .X(n27856) );
  nand_x1_sg U54580 ( .A(n35264), .B(reg_www_15[11]), .X(n27853) );
  nand_x1_sg U54581 ( .A(\filter_0/reg_w_15[11] ), .B(n32864), .X(n27854) );
  nand_x1_sg U54582 ( .A(n33919), .B(reg_www_15[10]), .X(n27851) );
  nand_x1_sg U54583 ( .A(\filter_0/reg_w_15[10] ), .B(n31208), .X(n27852) );
  nand_x1_sg U54584 ( .A(n34031), .B(reg_www_15[9]), .X(n27849) );
  nand_x1_sg U54585 ( .A(\filter_0/reg_w_15[9] ), .B(n30248), .X(n27850) );
  nand_x1_sg U54586 ( .A(n31523), .B(reg_www_15[8]), .X(n27847) );
  nand_x1_sg U54587 ( .A(\filter_0/reg_w_15[8] ), .B(n32779), .X(n27848) );
  nand_x1_sg U54588 ( .A(n34030), .B(reg_www_14[9]), .X(n27809) );
  nand_x1_sg U54589 ( .A(\filter_0/reg_w_14[9] ), .B(n34636), .X(n27810) );
  nand_x1_sg U54590 ( .A(n31681), .B(reg_www_14[8]), .X(n27807) );
  nand_x1_sg U54591 ( .A(\filter_0/reg_w_14[8] ), .B(n32790), .X(n27808) );
  nand_x1_sg U54592 ( .A(n33941), .B(reg_www_14[7]), .X(n27805) );
  nand_x1_sg U54593 ( .A(\filter_0/reg_w_14[7] ), .B(n32876), .X(n27806) );
  nand_x1_sg U54594 ( .A(n31686), .B(reg_www_14[6]), .X(n27803) );
  nand_x1_sg U54595 ( .A(\filter_0/reg_w_14[6] ), .B(n32811), .X(n27804) );
  nand_x1_sg U54596 ( .A(n31531), .B(reg_www_14[5]), .X(n27801) );
  nand_x1_sg U54597 ( .A(\filter_0/reg_w_14[5] ), .B(n32791), .X(n27802) );
  nand_x1_sg U54598 ( .A(n34029), .B(reg_www_14[4]), .X(n27799) );
  nand_x1_sg U54599 ( .A(\filter_0/reg_w_14[4] ), .B(n32864), .X(n27800) );
  nand_x1_sg U54600 ( .A(n30209), .B(reg_www_14[3]), .X(n27797) );
  nand_x1_sg U54601 ( .A(\filter_0/reg_w_14[3] ), .B(n32826), .X(n27798) );
  nand_x1_sg U54602 ( .A(n31522), .B(reg_www_14[2]), .X(n27795) );
  nand_x1_sg U54603 ( .A(\filter_0/reg_w_14[2] ), .B(n30247), .X(n27796) );
  nand_x1_sg U54604 ( .A(n34883), .B(reg_www_14[1]), .X(n27793) );
  nand_x1_sg U54605 ( .A(\filter_0/reg_w_14[1] ), .B(n31292), .X(n27794) );
  nand_x1_sg U54606 ( .A(n30158), .B(reg_www_14[0]), .X(n27791) );
  nand_x1_sg U54607 ( .A(\filter_0/reg_w_14[0] ), .B(n34642), .X(n27792) );
  nand_x1_sg U54608 ( .A(n33930), .B(reg_www_13[19]), .X(n27789) );
  nand_x1_sg U54609 ( .A(\filter_0/reg_w_13[19] ), .B(n30739), .X(n27790) );
  nand_x1_sg U54610 ( .A(n34912), .B(reg_www_13[18]), .X(n27787) );
  nand_x1_sg U54611 ( .A(\filter_0/reg_w_13[18] ), .B(n32877), .X(n27788) );
  nand_x1_sg U54612 ( .A(n34038), .B(reg_www_13[17]), .X(n27785) );
  nand_x1_sg U54613 ( .A(\filter_0/reg_w_13[17] ), .B(n30164), .X(n27786) );
  nand_x1_sg U54614 ( .A(n34031), .B(reg_www_13[16]), .X(n27783) );
  nand_x1_sg U54615 ( .A(\filter_0/reg_w_13[16] ), .B(n31921), .X(n27784) );
  nand_x1_sg U54616 ( .A(n31084), .B(reg_www_13[15]), .X(n27781) );
  nand_x1_sg U54617 ( .A(\filter_0/reg_w_13[15] ), .B(n32431), .X(n27782) );
  nand_x1_sg U54618 ( .A(n32223), .B(reg_www_13[14]), .X(n27779) );
  nand_x1_sg U54619 ( .A(\filter_0/reg_w_13[14] ), .B(n32879), .X(n27780) );
  nand_x1_sg U54620 ( .A(n31070), .B(reg_www_13[13]), .X(n27777) );
  nand_x1_sg U54621 ( .A(\filter_0/reg_w_13[13] ), .B(n34638), .X(n27778) );
  nand_x1_sg U54622 ( .A(n30627), .B(reg_www_13[12]), .X(n27775) );
  nand_x1_sg U54623 ( .A(\filter_0/reg_w_13[12] ), .B(n32865), .X(n27776) );
  nand_x1_sg U54624 ( .A(n35412), .B(reg_www_13[11]), .X(n27773) );
  nand_x1_sg U54625 ( .A(\filter_0/reg_w_13[11] ), .B(n32432), .X(n27774) );
  nand_x1_sg U54626 ( .A(n34601), .B(reg_www_12[11]), .X(n27733) );
  nand_x1_sg U54627 ( .A(\filter_0/reg_w_12[11] ), .B(n34688), .X(n27734) );
  nand_x1_sg U54628 ( .A(n33931), .B(reg_www_12[10]), .X(n27731) );
  nand_x1_sg U54629 ( .A(\filter_0/reg_w_12[10] ), .B(n34677), .X(n27732) );
  nand_x1_sg U54630 ( .A(n31526), .B(reg_www_12[9]), .X(n27729) );
  nand_x1_sg U54631 ( .A(\filter_0/reg_w_12[9] ), .B(n32465), .X(n27730) );
  nand_x1_sg U54632 ( .A(n33941), .B(reg_www_12[8]), .X(n27727) );
  nand_x1_sg U54633 ( .A(\filter_0/reg_w_12[8] ), .B(n32787), .X(n27728) );
  nand_x1_sg U54634 ( .A(n29696), .B(reg_www_12[7]), .X(n27725) );
  nand_x1_sg U54635 ( .A(\filter_0/reg_w_12[7] ), .B(n31920), .X(n27726) );
  nand_x1_sg U54636 ( .A(n34031), .B(reg_www_12[6]), .X(n27723) );
  nand_x1_sg U54637 ( .A(\filter_0/reg_w_12[6] ), .B(n32468), .X(n27724) );
  nand_x1_sg U54638 ( .A(n33901), .B(reg_www_12[4]), .X(n27719) );
  nand_x1_sg U54639 ( .A(\filter_0/reg_w_12[4] ), .B(n32790), .X(n27720) );
  nand_x1_sg U54640 ( .A(n33924), .B(reg_www_12[3]), .X(n27717) );
  nand_x1_sg U54641 ( .A(\filter_0/reg_w_12[3] ), .B(n32490), .X(n27718) );
  nand_x1_sg U54642 ( .A(n32259), .B(reg_www_12[2]), .X(n27715) );
  nand_x1_sg U54643 ( .A(\filter_0/reg_w_12[2] ), .B(n32469), .X(n27716) );
  nand_x1_sg U54644 ( .A(n30921), .B(reg_www_12[1]), .X(n27713) );
  nand_x1_sg U54645 ( .A(\filter_0/reg_w_12[1] ), .B(n32461), .X(n27714) );
  nand_x1_sg U54646 ( .A(n34033), .B(reg_www_12[0]), .X(n27711) );
  nand_x1_sg U54647 ( .A(\filter_0/reg_w_12[0] ), .B(n34673), .X(n27712) );
  nand_x1_sg U54648 ( .A(n34888), .B(reg_www_11[19]), .X(n27709) );
  nand_x1_sg U54649 ( .A(\filter_0/reg_w_11[19] ), .B(n30168), .X(n27710) );
  nand_x1_sg U54650 ( .A(n32275), .B(reg_www_11[18]), .X(n27707) );
  nand_x1_sg U54651 ( .A(\filter_0/reg_w_11[18] ), .B(n32779), .X(n27708) );
  nand_x1_sg U54652 ( .A(n31085), .B(reg_www_11[17]), .X(n27705) );
  nand_x1_sg U54653 ( .A(\filter_0/reg_w_11[17] ), .B(n30745), .X(n27706) );
  nand_x1_sg U54654 ( .A(n33900), .B(reg_www_11[16]), .X(n27703) );
  nand_x1_sg U54655 ( .A(\filter_0/reg_w_11[16] ), .B(n35074), .X(n27704) );
  nand_x1_sg U54656 ( .A(n30386), .B(reg_www_11[15]), .X(n27701) );
  nand_x1_sg U54657 ( .A(\filter_0/reg_w_11[15] ), .B(n32792), .X(n27702) );
  nand_x1_sg U54658 ( .A(n30775), .B(reg_www_11[14]), .X(n27699) );
  nand_x1_sg U54659 ( .A(\filter_0/reg_w_11[14] ), .B(n32465), .X(n27700) );
  nand_x1_sg U54660 ( .A(n33889), .B(reg_www_11[13]), .X(n27697) );
  nand_x1_sg U54661 ( .A(\filter_0/reg_w_11[13] ), .B(n32482), .X(n27698) );
  nand_x1_sg U54662 ( .A(n32267), .B(reg_www_11[12]), .X(n27695) );
  nand_x1_sg U54663 ( .A(\filter_0/reg_w_11[12] ), .B(n34692), .X(n27696) );
  nand_x1_sg U54664 ( .A(n34019), .B(reg_www_11[11]), .X(n27693) );
  nand_x1_sg U54665 ( .A(\filter_0/reg_w_11[11] ), .B(n32479), .X(n27694) );
  nand_x1_sg U54666 ( .A(n34891), .B(reg_www_11[10]), .X(n27691) );
  nand_x1_sg U54667 ( .A(\filter_0/reg_w_11[10] ), .B(n32477), .X(n27692) );
  nand_x1_sg U54668 ( .A(n29702), .B(reg_www_11[9]), .X(n27689) );
  nand_x1_sg U54669 ( .A(\filter_0/reg_w_11[9] ), .B(n32780), .X(n27690) );
  nand_x1_sg U54670 ( .A(n30159), .B(reg_www_11[8]), .X(n27687) );
  nand_x1_sg U54671 ( .A(\filter_0/reg_w_11[8] ), .B(n32806), .X(n27688) );
  nand_x1_sg U54672 ( .A(n33926), .B(reg_www_11[7]), .X(n27685) );
  nand_x1_sg U54673 ( .A(\filter_0/reg_w_11[7] ), .B(n32802), .X(n27686) );
  nand_x1_sg U54674 ( .A(n31529), .B(reg_www_11[6]), .X(n27683) );
  nand_x1_sg U54675 ( .A(\filter_0/reg_w_11[6] ), .B(n34685), .X(n27684) );
  nand_x1_sg U54676 ( .A(n30927), .B(reg_www_11[5]), .X(n27681) );
  nand_x1_sg U54677 ( .A(\filter_0/reg_w_11[5] ), .B(n32486), .X(n27682) );
  nand_x1_sg U54678 ( .A(n33912), .B(reg_www_11[4]), .X(n27679) );
  nand_x1_sg U54679 ( .A(\filter_0/reg_w_11[4] ), .B(n32786), .X(n27680) );
  nand_x1_sg U54680 ( .A(n30933), .B(reg_www_11[3]), .X(n27677) );
  nand_x1_sg U54681 ( .A(\filter_0/reg_w_11[3] ), .B(n31914), .X(n27678) );
  nand_x1_sg U54682 ( .A(n34026), .B(reg_www_11[2]), .X(n27675) );
  nand_x1_sg U54683 ( .A(\filter_0/reg_w_11[2] ), .B(n32799), .X(n27676) );
  nand_x1_sg U54684 ( .A(n30026), .B(reg_www_11[1]), .X(n27673) );
  nand_x1_sg U54685 ( .A(\filter_0/reg_w_11[1] ), .B(n34676), .X(n27674) );
  nand_x1_sg U54686 ( .A(n31524), .B(reg_www_11[0]), .X(n27671) );
  nand_x1_sg U54687 ( .A(\filter_0/reg_w_11[0] ), .B(n30767), .X(n27672) );
  nand_x1_sg U54688 ( .A(n33935), .B(reg_www_10[19]), .X(n27669) );
  nand_x1_sg U54689 ( .A(\filter_0/reg_w_10[19] ), .B(n32463), .X(n27670) );
  nand_x1_sg U54690 ( .A(n31529), .B(reg_www_10[18]), .X(n27667) );
  nand_x1_sg U54691 ( .A(\filter_0/reg_w_10[18] ), .B(n32432), .X(n27668) );
  nand_x1_sg U54692 ( .A(n33934), .B(reg_www_10[17]), .X(n27665) );
  nand_x1_sg U54693 ( .A(\filter_0/reg_w_10[17] ), .B(n32432), .X(n27666) );
  nand_x1_sg U54694 ( .A(n30027), .B(reg_www_10[16]), .X(n27663) );
  nand_x1_sg U54695 ( .A(\filter_0/reg_w_10[16] ), .B(n32460), .X(n27664) );
  nand_x1_sg U54696 ( .A(n35265), .B(reg_www_10[15]), .X(n27661) );
  nand_x1_sg U54697 ( .A(\filter_0/reg_w_10[15] ), .B(n30249), .X(n27662) );
  nand_x1_sg U54698 ( .A(n30927), .B(reg_www_10[14]), .X(n27659) );
  nand_x1_sg U54699 ( .A(\filter_0/reg_w_10[14] ), .B(n32475), .X(n27660) );
  nand_x1_sg U54700 ( .A(n33914), .B(reg_www_10[13]), .X(n27657) );
  nand_x1_sg U54701 ( .A(\filter_0/reg_w_10[13] ), .B(n30742), .X(n27658) );
  nand_x1_sg U54702 ( .A(n31243), .B(reg_www_10[12]), .X(n27655) );
  nand_x1_sg U54703 ( .A(\filter_0/reg_w_10[12] ), .B(n32812), .X(n27656) );
  nand_x1_sg U54704 ( .A(n32277), .B(reg_www_10[11]), .X(n27653) );
  nand_x1_sg U54705 ( .A(\filter_0/reg_w_10[11] ), .B(n32787), .X(n27654) );
  nand_x1_sg U54706 ( .A(n34019), .B(reg_www_10[10]), .X(n27651) );
  nand_x1_sg U54707 ( .A(\filter_0/reg_w_10[10] ), .B(n32815), .X(n27652) );
  nand_x1_sg U54708 ( .A(n30210), .B(reg_www_10[9]), .X(n27649) );
  nand_x1_sg U54709 ( .A(\filter_0/reg_w_10[9] ), .B(n30764), .X(n27650) );
  nand_x1_sg U54710 ( .A(n30929), .B(reg_www_10[8]), .X(n27647) );
  nand_x1_sg U54711 ( .A(\filter_0/reg_w_10[8] ), .B(n32790), .X(n27648) );
  nand_x1_sg U54712 ( .A(n31522), .B(reg_www_10[7]), .X(n27645) );
  nand_x1_sg U54713 ( .A(\filter_0/reg_w_10[7] ), .B(n32879), .X(n27646) );
  nand_x1_sg U54714 ( .A(n30627), .B(reg_www_10[6]), .X(n27643) );
  nand_x1_sg U54715 ( .A(\filter_0/reg_w_10[6] ), .B(n32875), .X(n27644) );
  nand_x1_sg U54716 ( .A(n34885), .B(reg_www_10[5]), .X(n27641) );
  nand_x1_sg U54717 ( .A(\filter_0/reg_w_10[5] ), .B(n32460), .X(n27642) );
  nand_x1_sg U54718 ( .A(n30256), .B(reg_www_10[4]), .X(n27639) );
  nand_x1_sg U54719 ( .A(\filter_0/reg_w_10[4] ), .B(n30764), .X(n27640) );
  nand_x1_sg U54720 ( .A(n31075), .B(reg_www_10[3]), .X(n27637) );
  nand_x1_sg U54721 ( .A(\filter_0/reg_w_10[3] ), .B(n32787), .X(n27638) );
  nand_x1_sg U54722 ( .A(n30777), .B(reg_www_10[2]), .X(n27635) );
  nand_x1_sg U54723 ( .A(\filter_0/reg_w_10[2] ), .B(n32791), .X(n27636) );
  nand_x1_sg U54724 ( .A(n32255), .B(reg_www_10[1]), .X(n27633) );
  nand_x1_sg U54725 ( .A(\filter_0/reg_w_10[1] ), .B(n31912), .X(n27634) );
  nand_x1_sg U54726 ( .A(n34040), .B(reg_www_10[0]), .X(n27631) );
  nand_x1_sg U54727 ( .A(\filter_0/reg_w_10[0] ), .B(n34671), .X(n27632) );
  nand_x1_sg U54728 ( .A(n34913), .B(reg_www_9[19]), .X(n27629) );
  nand_x1_sg U54729 ( .A(\filter_0/reg_w_9[19] ), .B(n32785), .X(n27630) );
  nand_x1_sg U54730 ( .A(n34883), .B(reg_www_9[18]), .X(n27627) );
  nand_x1_sg U54731 ( .A(\filter_0/reg_w_9[18] ), .B(n31912), .X(n27628) );
  nand_x1_sg U54732 ( .A(n32266), .B(reg_www_9[17]), .X(n27625) );
  nand_x1_sg U54733 ( .A(\filter_0/reg_w_9[17] ), .B(n32431), .X(n27626) );
  nand_x1_sg U54734 ( .A(n34041), .B(reg_www_9[16]), .X(n27623) );
  nand_x1_sg U54735 ( .A(\filter_0/reg_w_9[16] ), .B(n31295), .X(n27624) );
  nand_x1_sg U54736 ( .A(n32275), .B(reg_www_9[15]), .X(n27621) );
  nand_x1_sg U54737 ( .A(\filter_0/reg_w_9[15] ), .B(n32464), .X(n27622) );
  nand_x1_sg U54738 ( .A(n33903), .B(reg_www_9[14]), .X(n27619) );
  nand_x1_sg U54739 ( .A(\filter_0/reg_w_9[14] ), .B(n32805), .X(n27620) );
  nand_x1_sg U54740 ( .A(n34911), .B(reg_www_9[13]), .X(n27617) );
  nand_x1_sg U54741 ( .A(\filter_0/reg_w_9[13] ), .B(n32877), .X(n27618) );
  nand_x1_sg U54742 ( .A(n32271), .B(reg_www_9[12]), .X(n27615) );
  nand_x1_sg U54743 ( .A(\filter_0/reg_w_9[12] ), .B(n31912), .X(n27616) );
  nand_x1_sg U54744 ( .A(n32268), .B(reg_www_9[11]), .X(n27613) );
  nand_x1_sg U54745 ( .A(\filter_0/reg_w_9[11] ), .B(n32867), .X(n27614) );
  nand_x1_sg U54746 ( .A(n34884), .B(reg_www_9[10]), .X(n27611) );
  nand_x1_sg U54747 ( .A(\filter_0/reg_w_9[10] ), .B(n30248), .X(n27612) );
  nand_x1_sg U54748 ( .A(n31524), .B(reg_www_9[9]), .X(n27609) );
  nand_x1_sg U54749 ( .A(\filter_0/reg_w_9[9] ), .B(n30168), .X(n27610) );
  nand_x1_sg U54750 ( .A(n30025), .B(reg_www_9[2]), .X(n27595) );
  nand_x1_sg U54751 ( .A(\filter_0/reg_w_9[2] ), .B(n34692), .X(n27596) );
  nand_x1_sg U54752 ( .A(n31529), .B(reg_www_9[1]), .X(n27593) );
  nand_x1_sg U54753 ( .A(\filter_0/reg_w_9[1] ), .B(n31294), .X(n27594) );
  nand_x1_sg U54754 ( .A(n30209), .B(reg_www_9[0]), .X(n27591) );
  nand_x1_sg U54755 ( .A(\filter_0/reg_w_9[0] ), .B(n34677), .X(n27592) );
  nand_x1_sg U54756 ( .A(n34906), .B(reg_www_8[19]), .X(n27589) );
  nand_x1_sg U54757 ( .A(\filter_0/reg_w_8[19] ), .B(n34682), .X(n27590) );
  nand_x1_sg U54758 ( .A(n34914), .B(reg_www_8[18]), .X(n27587) );
  nand_x1_sg U54759 ( .A(\filter_0/reg_w_8[18] ), .B(n34675), .X(n27588) );
  nand_x1_sg U54760 ( .A(n33895), .B(reg_www_8[17]), .X(n27585) );
  nand_x1_sg U54761 ( .A(\filter_0/reg_w_8[17] ), .B(n32434), .X(n27586) );
  nand_x1_sg U54762 ( .A(n33894), .B(reg_www_8[16]), .X(n27583) );
  nand_x1_sg U54763 ( .A(\filter_0/reg_w_8[16] ), .B(n34680), .X(n27584) );
  nand_x1_sg U54764 ( .A(n34880), .B(reg_www_8[15]), .X(n27581) );
  nand_x1_sg U54765 ( .A(\filter_0/reg_w_8[15] ), .B(n31912), .X(n27582) );
  nand_x1_sg U54766 ( .A(n34039), .B(reg_www_8[14]), .X(n27579) );
  nand_x1_sg U54767 ( .A(\filter_0/reg_w_8[14] ), .B(n32871), .X(n27580) );
  nand_x1_sg U54768 ( .A(n32263), .B(reg_www_8[13]), .X(n27577) );
  nand_x1_sg U54769 ( .A(\filter_0/reg_w_8[13] ), .B(n32820), .X(n27578) );
  nand_x1_sg U54770 ( .A(n34914), .B(reg_www_8[12]), .X(n27575) );
  nand_x1_sg U54771 ( .A(\filter_0/reg_w_8[12] ), .B(n34670), .X(n27576) );
  nand_x1_sg U54772 ( .A(n34028), .B(reg_www_8[11]), .X(n27573) );
  nand_x1_sg U54773 ( .A(\filter_0/reg_w_8[11] ), .B(n32486), .X(n27574) );
  nand_x1_sg U54774 ( .A(n34038), .B(reg_www_8[10]), .X(n27571) );
  nand_x1_sg U54775 ( .A(\filter_0/reg_w_8[10] ), .B(n30166), .X(n27572) );
  nand_x1_sg U54776 ( .A(n33893), .B(reg_www_8[9]), .X(n27569) );
  nand_x1_sg U54777 ( .A(\filter_0/reg_w_8[9] ), .B(n30736), .X(n27570) );
  nand_x1_sg U54778 ( .A(n34889), .B(reg_www_8[8]), .X(n27567) );
  nand_x1_sg U54779 ( .A(\filter_0/reg_w_8[8] ), .B(n32865), .X(n27568) );
  nand_x1_sg U54780 ( .A(n33892), .B(reg_www_8[7]), .X(n27565) );
  nand_x1_sg U54781 ( .A(\filter_0/reg_w_8[7] ), .B(n32485), .X(n27566) );
  nand_x1_sg U54782 ( .A(n33897), .B(reg_www_8[6]), .X(n27563) );
  nand_x1_sg U54783 ( .A(\filter_0/reg_w_8[6] ), .B(n32801), .X(n27564) );
  nand_x1_sg U54784 ( .A(n29694), .B(reg_www_8[5]), .X(n27561) );
  nand_x1_sg U54785 ( .A(\filter_0/reg_w_8[5] ), .B(n34648), .X(n27562) );
  nand_x1_sg U54786 ( .A(n31679), .B(reg_www_8[4]), .X(n27559) );
  nand_x1_sg U54787 ( .A(\filter_0/reg_w_8[4] ), .B(n32865), .X(n27560) );
  nand_x1_sg U54788 ( .A(n30256), .B(reg_www_7[10]), .X(n27531) );
  nand_x1_sg U54789 ( .A(\filter_0/reg_w_7[10] ), .B(n32862), .X(n27532) );
  nand_x1_sg U54790 ( .A(n33892), .B(reg_www_7[9]), .X(n27529) );
  nand_x1_sg U54791 ( .A(\filter_0/reg_w_7[9] ), .B(n32877), .X(n27530) );
  nand_x1_sg U54792 ( .A(n34036), .B(reg_www_7[8]), .X(n27527) );
  nand_x1_sg U54793 ( .A(\filter_0/reg_w_7[8] ), .B(n32817), .X(n27528) );
  nand_x1_sg U54794 ( .A(n33941), .B(reg_www_7[7]), .X(n27525) );
  nand_x1_sg U54795 ( .A(\filter_0/reg_w_7[7] ), .B(n32810), .X(n27526) );
  nand_x1_sg U54796 ( .A(n31522), .B(reg_www_7[6]), .X(n27523) );
  nand_x1_sg U54797 ( .A(\filter_0/reg_w_7[6] ), .B(n30768), .X(n27524) );
  nand_x1_sg U54798 ( .A(n33934), .B(reg_www_7[5]), .X(n27521) );
  nand_x1_sg U54799 ( .A(\filter_0/reg_w_7[5] ), .B(n32464), .X(n27522) );
  nand_x1_sg U54800 ( .A(n34021), .B(reg_www_7[4]), .X(n27519) );
  nand_x1_sg U54801 ( .A(\filter_0/reg_w_7[4] ), .B(n32807), .X(n27520) );
  nand_x1_sg U54802 ( .A(n34603), .B(reg_www_7[3]), .X(n27517) );
  nand_x1_sg U54803 ( .A(\filter_0/reg_w_7[3] ), .B(n34631), .X(n27518) );
  nand_x1_sg U54804 ( .A(n33904), .B(reg_www_7[2]), .X(n27515) );
  nand_x1_sg U54805 ( .A(\filter_0/reg_w_7[2] ), .B(n34631), .X(n27516) );
  nand_x1_sg U54806 ( .A(n31518), .B(reg_www_7[1]), .X(n27513) );
  nand_x1_sg U54807 ( .A(\filter_0/reg_w_7[1] ), .B(n32794), .X(n27514) );
  nand_x1_sg U54808 ( .A(n32278), .B(reg_www_7[0]), .X(n27511) );
  nand_x1_sg U54809 ( .A(\filter_0/reg_w_7[0] ), .B(n34683), .X(n27512) );
  nand_x1_sg U54810 ( .A(n32263), .B(reg_www_6[19]), .X(n27509) );
  nand_x1_sg U54811 ( .A(\filter_0/reg_w_6[19] ), .B(n35070), .X(n27510) );
  nand_x1_sg U54812 ( .A(n33908), .B(reg_www_6[18]), .X(n27507) );
  nand_x1_sg U54813 ( .A(\filter_0/reg_w_6[18] ), .B(n31920), .X(n27508) );
  nand_x1_sg U54814 ( .A(n31089), .B(reg_www_6[17]), .X(n27505) );
  nand_x1_sg U54815 ( .A(\filter_0/reg_w_6[17] ), .B(n32779), .X(n27506) );
  nand_x1_sg U54816 ( .A(n31069), .B(reg_www_6[16]), .X(n27503) );
  nand_x1_sg U54817 ( .A(\filter_0/reg_w_6[16] ), .B(n30735), .X(n27504) );
  nand_x1_sg U54818 ( .A(n33896), .B(reg_www_6[15]), .X(n27501) );
  nand_x1_sg U54819 ( .A(\filter_0/reg_w_6[15] ), .B(n30761), .X(n27502) );
  nand_x1_sg U54820 ( .A(n33901), .B(reg_www_6[14]), .X(n27499) );
  nand_x1_sg U54821 ( .A(\filter_0/reg_w_6[14] ), .B(n32467), .X(n27500) );
  nand_x1_sg U54822 ( .A(n29700), .B(reg_www_6[13]), .X(n27497) );
  nand_x1_sg U54823 ( .A(\filter_0/reg_w_6[13] ), .B(n34686), .X(n27498) );
  nand_x1_sg U54824 ( .A(n31242), .B(reg_www_6[12]), .X(n27495) );
  nand_x1_sg U54825 ( .A(\filter_0/reg_w_6[12] ), .B(n34683), .X(n27496) );
  nand_x1_sg U54826 ( .A(n31686), .B(reg_www_6[11]), .X(n27493) );
  nand_x1_sg U54827 ( .A(\filter_0/reg_w_6[11] ), .B(n32458), .X(n27494) );
  nand_x1_sg U54828 ( .A(n35159), .B(reg_www_6[10]), .X(n27491) );
  nand_x1_sg U54829 ( .A(\filter_0/reg_w_6[10] ), .B(n32804), .X(n27492) );
  nand_x1_sg U54830 ( .A(n34009), .B(reg_www_6[9]), .X(n27489) );
  nand_x1_sg U54831 ( .A(\filter_0/reg_w_6[9] ), .B(n34624), .X(n27490) );
  nand_x1_sg U54832 ( .A(n34886), .B(reg_www_6[8]), .X(n27487) );
  nand_x1_sg U54833 ( .A(\filter_0/reg_w_6[8] ), .B(n30735), .X(n27488) );
  nand_x1_sg U54834 ( .A(n35411), .B(reg_www_6[7]), .X(n27485) );
  nand_x1_sg U54835 ( .A(\filter_0/reg_w_6[7] ), .B(n34641), .X(n27486) );
  nand_x1_sg U54836 ( .A(n30937), .B(reg_www_6[6]), .X(n27483) );
  nand_x1_sg U54837 ( .A(\filter_0/reg_w_6[6] ), .B(n34671), .X(n27484) );
  nand_x1_sg U54838 ( .A(n34907), .B(reg_www_6[5]), .X(n27481) );
  nand_x1_sg U54839 ( .A(\filter_0/reg_w_6[5] ), .B(n34672), .X(n27482) );
  nand_x1_sg U54840 ( .A(n30026), .B(reg_www_6[4]), .X(n27479) );
  nand_x1_sg U54841 ( .A(\filter_0/reg_w_6[4] ), .B(n34690), .X(n27480) );
  nand_x1_sg U54842 ( .A(n32224), .B(reg_www_6[3]), .X(n27477) );
  nand_x1_sg U54843 ( .A(\filter_0/reg_w_6[3] ), .B(n34672), .X(n27478) );
  nand_x1_sg U54844 ( .A(n31080), .B(reg_www_6[2]), .X(n27475) );
  nand_x1_sg U54845 ( .A(\filter_0/reg_w_6[2] ), .B(n34631), .X(n27476) );
  nand_x1_sg U54846 ( .A(n33935), .B(reg_www_6[1]), .X(n27473) );
  nand_x1_sg U54847 ( .A(\filter_0/reg_w_6[1] ), .B(n32822), .X(n27474) );
  nand_x1_sg U54848 ( .A(n34908), .B(reg_www_6[0]), .X(n27471) );
  nand_x1_sg U54849 ( .A(\filter_0/reg_w_6[0] ), .B(n31917), .X(n27472) );
  nand_x1_sg U54850 ( .A(n33934), .B(reg_www_5[19]), .X(n27469) );
  nand_x1_sg U54851 ( .A(\filter_0/reg_w_5[19] ), .B(n34621), .X(n27470) );
  nand_x1_sg U54852 ( .A(n31084), .B(reg_www_5[18]), .X(n27467) );
  nand_x1_sg U54853 ( .A(\filter_0/reg_w_5[18] ), .B(n34630), .X(n27468) );
  nand_x1_sg U54854 ( .A(n32271), .B(reg_www_5[17]), .X(n27465) );
  nand_x1_sg U54855 ( .A(\filter_0/reg_w_5[17] ), .B(n30732), .X(n27466) );
  nand_x1_sg U54856 ( .A(n34025), .B(reg_www_5[16]), .X(n27463) );
  nand_x1_sg U54857 ( .A(\filter_0/reg_w_5[16] ), .B(n32816), .X(n27464) );
  nand_x1_sg U54858 ( .A(n31075), .B(reg_www_5[15]), .X(n27461) );
  nand_x1_sg U54859 ( .A(\filter_0/reg_w_5[15] ), .B(n34642), .X(n27462) );
  nand_x1_sg U54860 ( .A(n34903), .B(reg_www_5[14]), .X(n27459) );
  nand_x1_sg U54861 ( .A(\filter_0/reg_w_5[14] ), .B(n34693), .X(n27460) );
  nand_x1_sg U54862 ( .A(n34879), .B(reg_www_5[13]), .X(n27457) );
  nand_x1_sg U54863 ( .A(\filter_0/reg_w_5[13] ), .B(n32430), .X(n27458) );
  nand_x1_sg U54864 ( .A(n33930), .B(reg_www_5[0]), .X(n27431) );
  nand_x1_sg U54865 ( .A(\filter_0/reg_w_5[0] ), .B(n32814), .X(n27432) );
  nand_x1_sg U54866 ( .A(n31516), .B(reg_www_4[19]), .X(n27429) );
  nand_x1_sg U54867 ( .A(\filter_0/reg_w_4[19] ), .B(n30762), .X(n27430) );
  nand_x1_sg U54868 ( .A(n34604), .B(reg_www_4[18]), .X(n27427) );
  nand_x1_sg U54869 ( .A(\filter_0/reg_w_4[18] ), .B(n35068), .X(n27428) );
  nand_x1_sg U54870 ( .A(n34601), .B(reg_www_4[17]), .X(n27425) );
  nand_x1_sg U54871 ( .A(\filter_0/reg_w_4[17] ), .B(n32468), .X(n27426) );
  nand_x1_sg U54872 ( .A(n34013), .B(reg_www_4[16]), .X(n27423) );
  nand_x1_sg U54873 ( .A(\filter_0/reg_w_4[16] ), .B(n32478), .X(n27424) );
  nand_x1_sg U54874 ( .A(n32261), .B(reg_www_4[15]), .X(n27421) );
  nand_x1_sg U54875 ( .A(\filter_0/reg_w_4[15] ), .B(n34633), .X(n27422) );
  nand_x1_sg U54876 ( .A(n31079), .B(reg_www_4[14]), .X(n27419) );
  nand_x1_sg U54877 ( .A(\filter_0/reg_w_4[14] ), .B(n34688), .X(n27420) );
  nand_x1_sg U54878 ( .A(n33924), .B(reg_www_4[13]), .X(n27417) );
  nand_x1_sg U54879 ( .A(\filter_0/reg_w_4[13] ), .B(n30742), .X(n27418) );
  nand_x1_sg U54880 ( .A(n31528), .B(reg_www_4[12]), .X(n27415) );
  nand_x1_sg U54881 ( .A(\filter_0/reg_w_4[12] ), .B(n34635), .X(n27416) );
  nand_x1_sg U54882 ( .A(n32260), .B(reg_www_4[11]), .X(n27413) );
  nand_x1_sg U54883 ( .A(\filter_0/reg_w_4[11] ), .B(n32825), .X(n27414) );
  nand_x1_sg U54884 ( .A(n31519), .B(reg_www_4[10]), .X(n27411) );
  nand_x1_sg U54885 ( .A(\filter_0/reg_w_4[10] ), .B(n31297), .X(n27412) );
  nand_x1_sg U54886 ( .A(n32272), .B(reg_www_4[9]), .X(n27409) );
  nand_x1_sg U54887 ( .A(\filter_0/reg_w_4[9] ), .B(n30164), .X(n27410) );
  nand_x1_sg U54888 ( .A(n31688), .B(reg_www_4[8]), .X(n27407) );
  nand_x1_sg U54889 ( .A(\filter_0/reg_w_4[8] ), .B(n35067), .X(n27408) );
  nand_x1_sg U54890 ( .A(n31516), .B(reg_www_3[8]), .X(n27367) );
  nand_x1_sg U54891 ( .A(\filter_0/reg_w_3[8] ), .B(n30764), .X(n27368) );
  nand_x1_sg U54892 ( .A(n31070), .B(reg_www_3[7]), .X(n27365) );
  nand_x1_sg U54893 ( .A(\filter_0/reg_w_3[7] ), .B(n34642), .X(n27366) );
  nand_x1_sg U54894 ( .A(n31065), .B(reg_www_3[6]), .X(n27363) );
  nand_x1_sg U54895 ( .A(\filter_0/reg_w_3[6] ), .B(n32870), .X(n27364) );
  nand_x1_sg U54896 ( .A(n31529), .B(reg_www_3[5]), .X(n27361) );
  nand_x1_sg U54897 ( .A(\filter_0/reg_w_3[5] ), .B(n34626), .X(n27362) );
  nand_x1_sg U54898 ( .A(n34884), .B(reg_www_3[4]), .X(n27359) );
  nand_x1_sg U54899 ( .A(\filter_0/reg_w_3[4] ), .B(n34647), .X(n27360) );
  nand_x1_sg U54900 ( .A(n32256), .B(reg_www_3[3]), .X(n27357) );
  nand_x1_sg U54901 ( .A(\filter_0/reg_w_3[3] ), .B(n34624), .X(n27358) );
  nand_x1_sg U54902 ( .A(n30775), .B(reg_www_3[2]), .X(n27355) );
  nand_x1_sg U54903 ( .A(\filter_0/reg_w_3[2] ), .B(n32869), .X(n27356) );
  nand_x1_sg U54904 ( .A(n31247), .B(reg_www_3[1]), .X(n27353) );
  nand_x1_sg U54905 ( .A(\filter_0/reg_w_3[1] ), .B(n32457), .X(n27354) );
  nand_x1_sg U54906 ( .A(n34609), .B(reg_www_3[0]), .X(n27351) );
  nand_x1_sg U54907 ( .A(\filter_0/reg_w_3[0] ), .B(n32782), .X(n27352) );
  nand_x1_sg U54908 ( .A(n34904), .B(reg_www_2[19]), .X(n27349) );
  nand_x1_sg U54909 ( .A(\filter_0/reg_w_2[19] ), .B(n32819), .X(n27350) );
  nand_x1_sg U54910 ( .A(n31533), .B(reg_www_2[18]), .X(n27347) );
  nand_x1_sg U54911 ( .A(\filter_0/reg_w_2[18] ), .B(n34620), .X(n27348) );
  nand_x1_sg U54912 ( .A(n29690), .B(reg_www_2[17]), .X(n27345) );
  nand_x1_sg U54913 ( .A(\filter_0/reg_w_2[17] ), .B(n34625), .X(n27346) );
  nand_x1_sg U54914 ( .A(n33893), .B(reg_www_2[9]), .X(n27329) );
  nand_x1_sg U54915 ( .A(\filter_0/reg_w_2[9] ), .B(n35070), .X(n27330) );
  nand_x1_sg U54916 ( .A(n33930), .B(reg_www_2[8]), .X(n27327) );
  nand_x1_sg U54917 ( .A(\filter_0/reg_w_2[8] ), .B(n30742), .X(n27328) );
  nand_x1_sg U54918 ( .A(n31248), .B(reg_www_2[7]), .X(n27325) );
  nand_x1_sg U54919 ( .A(\filter_0/reg_w_2[7] ), .B(n30164), .X(n27326) );
  nand_x1_sg U54920 ( .A(n32270), .B(reg_www_2[6]), .X(n27323) );
  nand_x1_sg U54921 ( .A(\filter_0/reg_w_2[6] ), .B(n31911), .X(n27324) );
  nand_x1_sg U54922 ( .A(n29700), .B(reg_www_2[5]), .X(n27321) );
  nand_x1_sg U54923 ( .A(\filter_0/reg_w_2[5] ), .B(n34646), .X(n27322) );
  nand_x1_sg U54924 ( .A(n31079), .B(reg_www_2[4]), .X(n27319) );
  nand_x1_sg U54925 ( .A(\filter_0/reg_w_2[4] ), .B(n34629), .X(n27320) );
  nand_x1_sg U54926 ( .A(n33900), .B(reg_www_2[3]), .X(n27317) );
  nand_x1_sg U54927 ( .A(\filter_0/reg_w_2[3] ), .B(n32817), .X(n27318) );
  nand_x1_sg U54928 ( .A(n34011), .B(reg_www_2[2]), .X(n27315) );
  nand_x1_sg U54929 ( .A(\filter_0/reg_w_2[2] ), .B(n34628), .X(n27316) );
  nand_x1_sg U54930 ( .A(n34881), .B(reg_www_2[1]), .X(n27313) );
  nand_x1_sg U54931 ( .A(\filter_0/reg_w_2[1] ), .B(n35067), .X(n27314) );
  nand_x1_sg U54932 ( .A(n34878), .B(reg_www_2[0]), .X(n27311) );
  nand_x1_sg U54933 ( .A(\filter_0/reg_w_2[0] ), .B(n35067), .X(n27312) );
  nand_x1_sg U54934 ( .A(n34889), .B(reg_www_1[19]), .X(n27309) );
  nand_x1_sg U54935 ( .A(\filter_0/reg_w_1[19] ), .B(n34683), .X(n27310) );
  nand_x1_sg U54936 ( .A(n34031), .B(reg_www_1[18]), .X(n27307) );
  nand_x1_sg U54937 ( .A(\filter_0/reg_w_1[18] ), .B(n35069), .X(n27308) );
  nand_x1_sg U54938 ( .A(n34878), .B(reg_www_1[17]), .X(n27305) );
  nand_x1_sg U54939 ( .A(\filter_0/reg_w_1[17] ), .B(n34681), .X(n27306) );
  nand_x1_sg U54940 ( .A(n32261), .B(reg_www_1[16]), .X(n27303) );
  nand_x1_sg U54941 ( .A(\filter_0/reg_w_1[16] ), .B(n32430), .X(n27304) );
  nand_x1_sg U54942 ( .A(n31084), .B(reg_www_1[15]), .X(n27301) );
  nand_x1_sg U54943 ( .A(\filter_0/reg_w_1[15] ), .B(n34634), .X(n27302) );
  nand_x1_sg U54944 ( .A(n30935), .B(reg_www_1[14]), .X(n27299) );
  nand_x1_sg U54945 ( .A(\filter_0/reg_w_1[14] ), .B(n32439), .X(n27300) );
  nand_x1_sg U54946 ( .A(n33890), .B(reg_www_1[13]), .X(n27297) );
  nand_x1_sg U54947 ( .A(\filter_0/reg_w_1[13] ), .B(n32795), .X(n27298) );
  nand_x1_sg U54948 ( .A(n32272), .B(reg_www_1[12]), .X(n27295) );
  nand_x1_sg U54949 ( .A(\filter_0/reg_w_1[12] ), .B(n32785), .X(n27296) );
  nand_x1_sg U54950 ( .A(n31525), .B(reg_www_1[11]), .X(n27293) );
  nand_x1_sg U54951 ( .A(\filter_0/reg_w_1[11] ), .B(n32782), .X(n27294) );
  nand_x1_sg U54952 ( .A(n32265), .B(reg_www_1[10]), .X(n27291) );
  nand_x1_sg U54953 ( .A(\filter_0/reg_w_1[10] ), .B(n32481), .X(n27292) );
  nand_x1_sg U54954 ( .A(n31085), .B(reg_www_1[9]), .X(n27289) );
  nand_x1_sg U54955 ( .A(\filter_0/reg_w_1[9] ), .B(n32490), .X(n27290) );
  nand_x1_sg U54956 ( .A(n31687), .B(reg_www_1[8]), .X(n27287) );
  nand_x1_sg U54957 ( .A(\filter_0/reg_w_1[8] ), .B(n30761), .X(n27288) );
  nand_x1_sg U54958 ( .A(n31678), .B(reg_www_1[7]), .X(n27285) );
  nand_x1_sg U54959 ( .A(\filter_0/reg_w_1[7] ), .B(n34683), .X(n27286) );
  nand_x1_sg U54960 ( .A(n33913), .B(reg_www_1[6]), .X(n27283) );
  nand_x1_sg U54961 ( .A(\filter_0/reg_w_1[6] ), .B(n30741), .X(n27284) );
  nand_x1_sg U54962 ( .A(n34041), .B(reg_www_1[5]), .X(n27281) );
  nand_x1_sg U54963 ( .A(\filter_0/reg_w_1[5] ), .B(n30250), .X(n27282) );
  nand_x1_sg U54964 ( .A(n33928), .B(reg_www_1[4]), .X(n27279) );
  nand_x1_sg U54965 ( .A(\filter_0/reg_w_1[4] ), .B(n31297), .X(n27280) );
  nand_x1_sg U54966 ( .A(n30158), .B(reg_www_1[3]), .X(n27277) );
  nand_x1_sg U54967 ( .A(\filter_0/reg_w_1[3] ), .B(n31918), .X(n27278) );
  nand_x1_sg U54968 ( .A(n34903), .B(reg_www_1[2]), .X(n27275) );
  nand_x1_sg U54969 ( .A(\filter_0/reg_w_1[2] ), .B(n32864), .X(n27276) );
  nand_x1_sg U54970 ( .A(n34014), .B(reg_www_1[1]), .X(n27273) );
  nand_x1_sg U54971 ( .A(\filter_0/reg_w_1[1] ), .B(n34675), .X(n27274) );
  nand_x1_sg U54972 ( .A(n34604), .B(reg_www_1[0]), .X(n27271) );
  nand_x1_sg U54973 ( .A(\filter_0/reg_w_1[0] ), .B(n31917), .X(n27272) );
  nand_x1_sg U54974 ( .A(n33911), .B(reg_www_0[19]), .X(n27269) );
  nand_x1_sg U54975 ( .A(\filter_0/reg_w_0[19] ), .B(n35074), .X(n27270) );
  nand_x1_sg U54976 ( .A(n31247), .B(reg_www_0[18]), .X(n27267) );
  nand_x1_sg U54977 ( .A(\filter_0/reg_w_0[18] ), .B(n32866), .X(n27268) );
  nand_x1_sg U54978 ( .A(n33906), .B(reg_www_0[17]), .X(n27265) );
  nand_x1_sg U54979 ( .A(\filter_0/reg_w_0[17] ), .B(n34681), .X(n27266) );
  nand_x1_sg U54980 ( .A(n32278), .B(reg_www_0[16]), .X(n27263) );
  nand_x1_sg U54981 ( .A(\filter_0/reg_w_0[16] ), .B(n32865), .X(n27264) );
  nand_x1_sg U54982 ( .A(n30927), .B(reg_www_0[15]), .X(n27261) );
  nand_x1_sg U54983 ( .A(\filter_0/reg_w_0[15] ), .B(n32435), .X(n27262) );
  nand_x1_sg U54984 ( .A(n31686), .B(reg_www_0[14]), .X(n27259) );
  nand_x1_sg U54985 ( .A(\filter_0/reg_w_0[14] ), .B(n34636), .X(n27260) );
  nand_x1_sg U54986 ( .A(n34883), .B(reg_www_0[13]), .X(n27257) );
  nand_x1_sg U54987 ( .A(\filter_0/reg_w_0[13] ), .B(n34642), .X(n27258) );
  nand_x1_sg U54988 ( .A(n34881), .B(reg_www_0[12]), .X(n27255) );
  nand_x1_sg U54989 ( .A(\filter_0/reg_w_0[12] ), .B(n30741), .X(n27256) );
  nand_x1_sg U54990 ( .A(n34912), .B(reg_www_0[11]), .X(n27253) );
  nand_x1_sg U54991 ( .A(\filter_0/reg_w_0[11] ), .B(n32792), .X(n27254) );
  nand_x1_sg U54992 ( .A(n30027), .B(reg_www_0[10]), .X(n27251) );
  nand_x1_sg U54993 ( .A(\filter_0/reg_w_0[10] ), .B(n32815), .X(n27252) );
  nand_x1_sg U54994 ( .A(n33938), .B(reg_www_0[9]), .X(n27249) );
  nand_x1_sg U54995 ( .A(\filter_0/reg_w_0[9] ), .B(n32468), .X(n27250) );
  nand_x1_sg U54996 ( .A(n31090), .B(reg_www_0[8]), .X(n27247) );
  nand_x1_sg U54997 ( .A(\filter_0/reg_w_0[8] ), .B(n31294), .X(n27248) );
  nand_x1_sg U54998 ( .A(n32259), .B(reg_www_0[7]), .X(n27245) );
  nand_x1_sg U54999 ( .A(\filter_0/reg_w_0[7] ), .B(n32474), .X(n27246) );
  nand_x1_sg U55000 ( .A(n32264), .B(reg_www_0[6]), .X(n27243) );
  nand_x1_sg U55001 ( .A(\filter_0/reg_w_0[6] ), .B(n31922), .X(n27244) );
  nand_x1_sg U55002 ( .A(n31523), .B(reg_iii_15[13]), .X(n27217) );
  nand_x1_sg U55003 ( .A(\filter_0/reg_i_15[13] ), .B(n32821), .X(n27218) );
  nand_x1_sg U55004 ( .A(n34025), .B(reg_iii_15[12]), .X(n27215) );
  nand_x1_sg U55005 ( .A(\filter_0/reg_i_15[12] ), .B(n32817), .X(n27216) );
  nand_x1_sg U55006 ( .A(n35466), .B(reg_iii_15[11]), .X(n27213) );
  nand_x1_sg U55007 ( .A(\filter_0/reg_i_15[11] ), .B(n32460), .X(n27214) );
  nand_x1_sg U55008 ( .A(n31247), .B(reg_iii_15[10]), .X(n27211) );
  nand_x1_sg U55009 ( .A(\filter_0/reg_i_15[10] ), .B(n32809), .X(n27212) );
  nand_x1_sg U55010 ( .A(n33933), .B(reg_iii_15[9]), .X(n27209) );
  nand_x1_sg U55011 ( .A(\filter_0/reg_i_15[9] ), .B(n30758), .X(n27210) );
  nand_x1_sg U55012 ( .A(n30627), .B(reg_iii_15[8]), .X(n27207) );
  nand_x1_sg U55013 ( .A(\filter_0/reg_i_15[8] ), .B(n31921), .X(n27208) );
  nand_x1_sg U55014 ( .A(n34035), .B(reg_iii_15[7]), .X(n27205) );
  nand_x1_sg U55015 ( .A(\filter_0/reg_i_15[7] ), .B(n34681), .X(n27206) );
  nand_x1_sg U55016 ( .A(n31520), .B(reg_iii_15[6]), .X(n27203) );
  nand_x1_sg U55017 ( .A(\filter_0/reg_i_15[6] ), .B(n30738), .X(n27204) );
  nand_x1_sg U55018 ( .A(n33936), .B(reg_iii_15[5]), .X(n27201) );
  nand_x1_sg U55019 ( .A(\filter_0/reg_i_15[5] ), .B(n34631), .X(n27202) );
  nand_x1_sg U55020 ( .A(n31243), .B(reg_iii_15[4]), .X(n27199) );
  nand_x1_sg U55021 ( .A(\filter_0/reg_i_15[4] ), .B(n32457), .X(n27200) );
  nand_x1_sg U55022 ( .A(n31248), .B(reg_iii_15[3]), .X(n27197) );
  nand_x1_sg U55023 ( .A(\filter_0/reg_i_15[3] ), .B(n31292), .X(n27198) );
  nand_x1_sg U55024 ( .A(n31074), .B(reg_iii_15[2]), .X(n27195) );
  nand_x1_sg U55025 ( .A(\filter_0/reg_i_15[2] ), .B(n32469), .X(n27196) );
  nand_x1_sg U55026 ( .A(n33911), .B(reg_iii_15[1]), .X(n27193) );
  nand_x1_sg U55027 ( .A(\filter_0/reg_i_15[1] ), .B(n32794), .X(n27194) );
  nand_x1_sg U55028 ( .A(n33928), .B(reg_iii_15[0]), .X(n27191) );
  nand_x1_sg U55029 ( .A(\filter_0/reg_i_15[0] ), .B(n34682), .X(n27192) );
  nand_x1_sg U55030 ( .A(n34030), .B(reg_iii_14[19]), .X(n27189) );
  nand_x1_sg U55031 ( .A(\filter_0/reg_i_14[19] ), .B(n32819), .X(n27190) );
  nand_x1_sg U55032 ( .A(n34884), .B(reg_iii_14[18]), .X(n27187) );
  nand_x1_sg U55033 ( .A(\filter_0/reg_i_14[18] ), .B(n32797), .X(n27188) );
  nand_x1_sg U55034 ( .A(n31519), .B(reg_iii_14[17]), .X(n27185) );
  nand_x1_sg U55035 ( .A(\filter_0/reg_i_14[17] ), .B(n32820), .X(n27186) );
  nand_x1_sg U55036 ( .A(n32223), .B(reg_iii_14[16]), .X(n27183) );
  nand_x1_sg U55037 ( .A(\filter_0/reg_i_14[16] ), .B(n32433), .X(n27184) );
  nand_x1_sg U55038 ( .A(n35265), .B(reg_iii_14[15]), .X(n27181) );
  nand_x1_sg U55039 ( .A(\filter_0/reg_i_14[15] ), .B(n30161), .X(n27182) );
  nand_x1_sg U55040 ( .A(n31064), .B(reg_iii_14[7]), .X(n27165) );
  nand_x1_sg U55041 ( .A(\filter_0/reg_i_14[7] ), .B(n32824), .X(n27166) );
  nand_x1_sg U55042 ( .A(n32255), .B(reg_iii_14[6]), .X(n27163) );
  nand_x1_sg U55043 ( .A(\filter_0/reg_i_14[6] ), .B(n34691), .X(n27164) );
  nand_x1_sg U55044 ( .A(n31528), .B(reg_iii_14[5]), .X(n27161) );
  nand_x1_sg U55045 ( .A(\filter_0/reg_i_14[5] ), .B(n35069), .X(n27162) );
  nand_x1_sg U55046 ( .A(n32276), .B(reg_iii_14[4]), .X(n27159) );
  nand_x1_sg U55047 ( .A(\filter_0/reg_i_14[4] ), .B(n32794), .X(n27160) );
  nand_x1_sg U55048 ( .A(n33890), .B(reg_iii_14[3]), .X(n27157) );
  nand_x1_sg U55049 ( .A(\filter_0/reg_i_14[3] ), .B(n34640), .X(n27158) );
  nand_x1_sg U55050 ( .A(n34022), .B(reg_iii_14[2]), .X(n27155) );
  nand_x1_sg U55051 ( .A(\filter_0/reg_i_14[2] ), .B(n34675), .X(n27156) );
  nand_x1_sg U55052 ( .A(n34021), .B(reg_iii_14[1]), .X(n27153) );
  nand_x1_sg U55053 ( .A(\filter_0/reg_i_14[1] ), .B(n32786), .X(n27154) );
  nand_x1_sg U55054 ( .A(n31528), .B(reg_iii_14[0]), .X(n27151) );
  nand_x1_sg U55055 ( .A(\filter_0/reg_i_14[0] ), .B(n32815), .X(n27152) );
  nand_x1_sg U55056 ( .A(n33920), .B(reg_iii_13[19]), .X(n27149) );
  nand_x1_sg U55057 ( .A(\filter_0/reg_i_13[19] ), .B(n34623), .X(n27150) );
  nand_x1_sg U55058 ( .A(n31521), .B(reg_iii_13[18]), .X(n27147) );
  nand_x1_sg U55059 ( .A(\filter_0/reg_i_13[18] ), .B(n32882), .X(n27148) );
  nand_x1_sg U55060 ( .A(n33914), .B(reg_iii_13[17]), .X(n27145) );
  nand_x1_sg U55061 ( .A(\filter_0/reg_i_13[17] ), .B(n32785), .X(n27146) );
  nand_x1_sg U55062 ( .A(n30937), .B(reg_iii_13[16]), .X(n27143) );
  nand_x1_sg U55063 ( .A(\filter_0/reg_i_13[16] ), .B(n32470), .X(n27144) );
  nand_x1_sg U55064 ( .A(n33907), .B(reg_iii_13[15]), .X(n27141) );
  nand_x1_sg U55065 ( .A(\filter_0/reg_i_13[15] ), .B(n32819), .X(n27142) );
  nand_x1_sg U55066 ( .A(n32224), .B(reg_iii_13[14]), .X(n27139) );
  nand_x1_sg U55067 ( .A(\filter_0/reg_i_13[14] ), .B(n34678), .X(n27140) );
  nand_x1_sg U55068 ( .A(n32271), .B(reg_iii_13[13]), .X(n27137) );
  nand_x1_sg U55069 ( .A(\filter_0/reg_i_13[13] ), .B(n32822), .X(n27138) );
  nand_x1_sg U55070 ( .A(n31521), .B(reg_iii_13[12]), .X(n27135) );
  nand_x1_sg U55071 ( .A(\filter_0/reg_i_13[12] ), .B(n32489), .X(n27136) );
  nand_x1_sg U55072 ( .A(n30777), .B(reg_iii_13[11]), .X(n27133) );
  nand_x1_sg U55073 ( .A(\filter_0/reg_i_13[11] ), .B(n32826), .X(n27134) );
  nand_x1_sg U55074 ( .A(n33918), .B(reg_iii_13[10]), .X(n27131) );
  nand_x1_sg U55075 ( .A(\filter_0/reg_i_13[10] ), .B(n30249), .X(n27132) );
  nand_x1_sg U55076 ( .A(n35411), .B(reg_iii_13[9]), .X(n27129) );
  nand_x1_sg U55077 ( .A(\filter_0/reg_i_13[9] ), .B(n32859), .X(n27130) );
  nand_x1_sg U55078 ( .A(n33908), .B(reg_iii_13[8]), .X(n27127) );
  nand_x1_sg U55079 ( .A(\filter_0/reg_i_13[8] ), .B(n32438), .X(n27128) );
  nand_x1_sg U55080 ( .A(n34023), .B(reg_iii_13[7]), .X(n27125) );
  nand_x1_sg U55081 ( .A(\filter_0/reg_i_13[7] ), .B(n34693), .X(n27126) );
  nand_x1_sg U55082 ( .A(n33890), .B(reg_iii_13[6]), .X(n27123) );
  nand_x1_sg U55083 ( .A(\filter_0/reg_i_13[6] ), .B(n32804), .X(n27124) );
  nand_x1_sg U55084 ( .A(n31525), .B(reg_iii_13[5]), .X(n27121) );
  nand_x1_sg U55085 ( .A(\filter_0/reg_i_13[5] ), .B(n32806), .X(n27122) );
  nand_x1_sg U55086 ( .A(n34016), .B(reg_iii_13[4]), .X(n27119) );
  nand_x1_sg U55087 ( .A(\filter_0/reg_i_13[4] ), .B(n34690), .X(n27120) );
  nand_x1_sg U55088 ( .A(n33940), .B(reg_iii_13[3]), .X(n27117) );
  nand_x1_sg U55089 ( .A(\filter_0/reg_i_13[3] ), .B(n32799), .X(n27118) );
  nand_x1_sg U55090 ( .A(n34034), .B(reg_iii_13[2]), .X(n27115) );
  nand_x1_sg U55091 ( .A(\filter_0/reg_i_13[2] ), .B(n35073), .X(n27116) );
  nand_x1_sg U55092 ( .A(n33925), .B(reg_iii_13[1]), .X(n27113) );
  nand_x1_sg U55093 ( .A(\filter_0/reg_i_13[1] ), .B(n34638), .X(n27114) );
  nand_x1_sg U55094 ( .A(n34606), .B(reg_iii_13[0]), .X(n27111) );
  nand_x1_sg U55095 ( .A(\filter_0/reg_i_13[0] ), .B(n30249), .X(n27112) );
  nand_x1_sg U55096 ( .A(n31685), .B(reg_iii_12[19]), .X(n27109) );
  nand_x1_sg U55097 ( .A(\filter_0/reg_i_12[19] ), .B(n32872), .X(n27110) );
  nand_x1_sg U55098 ( .A(n30775), .B(reg_iii_12[18]), .X(n27107) );
  nand_x1_sg U55099 ( .A(\filter_0/reg_i_12[18] ), .B(n32779), .X(n27108) );
  nand_x1_sg U55100 ( .A(n31685), .B(reg_iii_12[17]), .X(n27105) );
  nand_x1_sg U55101 ( .A(\filter_0/reg_i_12[17] ), .B(n34643), .X(n27106) );
  nand_x1_sg U55102 ( .A(n34906), .B(reg_iii_12[16]), .X(n27103) );
  nand_x1_sg U55103 ( .A(\filter_0/reg_i_12[16] ), .B(n31922), .X(n27104) );
  nand_x1_sg U55104 ( .A(n34608), .B(reg_iii_12[15]), .X(n27101) );
  nand_x1_sg U55105 ( .A(\filter_0/reg_i_12[15] ), .B(n32814), .X(n27102) );
  nand_x1_sg U55106 ( .A(n34603), .B(reg_iii_12[14]), .X(n27099) );
  nand_x1_sg U55107 ( .A(\filter_0/reg_i_12[14] ), .B(n32861), .X(n27100) );
  nand_x1_sg U55108 ( .A(n34602), .B(reg_iii_12[13]), .X(n27097) );
  nand_x1_sg U55109 ( .A(\filter_0/reg_i_12[13] ), .B(n32874), .X(n27098) );
  nand_x1_sg U55110 ( .A(n32264), .B(reg_iii_12[12]), .X(n27095) );
  nand_x1_sg U55111 ( .A(\filter_0/reg_i_12[12] ), .B(n32866), .X(n27096) );
  nand_x1_sg U55112 ( .A(n31526), .B(reg_iii_12[11]), .X(n27093) );
  nand_x1_sg U55113 ( .A(\filter_0/reg_i_12[11] ), .B(n32864), .X(n27094) );
  nand_x1_sg U55114 ( .A(n31684), .B(reg_iii_12[10]), .X(n27091) );
  nand_x1_sg U55115 ( .A(\filter_0/reg_i_12[10] ), .B(n32474), .X(n27092) );
  nand_x1_sg U55116 ( .A(n33926), .B(reg_iii_12[9]), .X(n27089) );
  nand_x1_sg U55117 ( .A(\filter_0/reg_i_12[9] ), .B(n32462), .X(n27090) );
  nand_x1_sg U55118 ( .A(n30935), .B(reg_iii_12[8]), .X(n27087) );
  nand_x1_sg U55119 ( .A(\filter_0/reg_i_12[8] ), .B(n32809), .X(n27088) );
  nand_x1_sg U55120 ( .A(n34021), .B(reg_iii_12[7]), .X(n27085) );
  nand_x1_sg U55121 ( .A(\filter_0/reg_i_12[7] ), .B(n32481), .X(n27086) );
  nand_x1_sg U55122 ( .A(n31089), .B(reg_iii_12[6]), .X(n27083) );
  nand_x1_sg U55123 ( .A(\filter_0/reg_i_12[6] ), .B(n32814), .X(n27084) );
  nand_x1_sg U55124 ( .A(n34601), .B(reg_iii_12[5]), .X(n27081) );
  nand_x1_sg U55125 ( .A(\filter_0/reg_i_12[5] ), .B(n32790), .X(n27082) );
  nand_x1_sg U55126 ( .A(n30387), .B(reg_iii_12[4]), .X(n27079) );
  nand_x1_sg U55127 ( .A(\filter_0/reg_i_12[4] ), .B(n34638), .X(n27080) );
  nand_x1_sg U55128 ( .A(n34602), .B(reg_iii_12[3]), .X(n27077) );
  nand_x1_sg U55129 ( .A(\filter_0/reg_i_12[3] ), .B(n32490), .X(n27078) );
  nand_x1_sg U55130 ( .A(n29689), .B(reg_iii_12[2]), .X(n27075) );
  nand_x1_sg U55131 ( .A(\filter_0/reg_i_12[2] ), .B(n32781), .X(n27076) );
  nand_x1_sg U55132 ( .A(n30931), .B(reg_iii_12[1]), .X(n27073) );
  nand_x1_sg U55133 ( .A(\filter_0/reg_i_12[1] ), .B(n32465), .X(n27074) );
  nand_x1_sg U55134 ( .A(n34609), .B(reg_iii_12[0]), .X(n27071) );
  nand_x1_sg U55135 ( .A(\filter_0/reg_i_12[0] ), .B(n31915), .X(n27072) );
  nand_x1_sg U55136 ( .A(n34036), .B(reg_iii_11[19]), .X(n27069) );
  nand_x1_sg U55137 ( .A(\filter_0/reg_i_11[19] ), .B(n31295), .X(n27070) );
  nand_x1_sg U55138 ( .A(n31520), .B(reg_iii_11[18]), .X(n27067) );
  nand_x1_sg U55139 ( .A(\filter_0/reg_i_11[18] ), .B(n31920), .X(n27068) );
  nand_x1_sg U55140 ( .A(n33929), .B(reg_iii_11[11]), .X(n27053) );
  nand_x1_sg U55141 ( .A(\filter_0/reg_i_11[11] ), .B(n34626), .X(n27054) );
  nand_x1_sg U55142 ( .A(n33904), .B(reg_iii_11[10]), .X(n27051) );
  nand_x1_sg U55143 ( .A(\filter_0/reg_i_11[10] ), .B(n32439), .X(n27052) );
  nand_x1_sg U55144 ( .A(n34608), .B(reg_iii_11[9]), .X(n27049) );
  nand_x1_sg U55145 ( .A(\filter_0/reg_i_11[9] ), .B(n34621), .X(n27050) );
  nand_x1_sg U55146 ( .A(n34025), .B(reg_iii_11[8]), .X(n27047) );
  nand_x1_sg U55147 ( .A(\filter_0/reg_i_11[8] ), .B(n30248), .X(n27048) );
  nand_x1_sg U55148 ( .A(n34036), .B(reg_iii_11[7]), .X(n27045) );
  nand_x1_sg U55149 ( .A(\filter_0/reg_i_11[7] ), .B(n31295), .X(n27046) );
  nand_x1_sg U55150 ( .A(n34028), .B(reg_iii_11[6]), .X(n27043) );
  nand_x1_sg U55151 ( .A(\filter_0/reg_i_11[6] ), .B(n34624), .X(n27044) );
  nand_x1_sg U55152 ( .A(n31530), .B(reg_iii_11[5]), .X(n27041) );
  nand_x1_sg U55153 ( .A(\filter_0/reg_i_11[5] ), .B(n30252), .X(n27042) );
  nand_x1_sg U55154 ( .A(n34040), .B(reg_iii_10[5]), .X(n27001) );
  nand_x1_sg U55155 ( .A(\filter_0/reg_i_10[5] ), .B(n31297), .X(n27002) );
  nand_x1_sg U55156 ( .A(n31085), .B(reg_iii_10[4]), .X(n26999) );
  nand_x1_sg U55157 ( .A(\filter_0/reg_i_10[4] ), .B(n31297), .X(n27000) );
  nand_x1_sg U55158 ( .A(n32275), .B(reg_iii_10[3]), .X(n26997) );
  nand_x1_sg U55159 ( .A(\filter_0/reg_i_10[3] ), .B(n32805), .X(n26998) );
  nand_x1_sg U55160 ( .A(n34018), .B(reg_iii_10[2]), .X(n26995) );
  nand_x1_sg U55161 ( .A(\filter_0/reg_i_10[2] ), .B(n30768), .X(n26996) );
  nand_x1_sg U55162 ( .A(n34011), .B(reg_iii_10[1]), .X(n26993) );
  nand_x1_sg U55163 ( .A(\filter_0/reg_i_10[1] ), .B(n32804), .X(n26994) );
  nand_x1_sg U55164 ( .A(n34607), .B(reg_iii_10[0]), .X(n26991) );
  nand_x1_sg U55165 ( .A(\filter_0/reg_i_10[0] ), .B(n30738), .X(n26992) );
  nand_x1_sg U55166 ( .A(n33925), .B(reg_iii_9[19]), .X(n26989) );
  nand_x1_sg U55167 ( .A(\filter_0/reg_i_9[19] ), .B(n32472), .X(n26990) );
  nand_x1_sg U55168 ( .A(n31533), .B(reg_iii_9[18]), .X(n26987) );
  nand_x1_sg U55169 ( .A(\filter_0/reg_i_9[18] ), .B(n31916), .X(n26988) );
  nand_x1_sg U55170 ( .A(n32263), .B(reg_iii_9[17]), .X(n26985) );
  nand_x1_sg U55171 ( .A(\filter_0/reg_i_9[17] ), .B(n32789), .X(n26986) );
  nand_x1_sg U55172 ( .A(n30921), .B(reg_iii_9[16]), .X(n26983) );
  nand_x1_sg U55173 ( .A(\filter_0/reg_i_9[16] ), .B(n31915), .X(n26984) );
  nand_x1_sg U55174 ( .A(n30921), .B(reg_iii_9[15]), .X(n26981) );
  nand_x1_sg U55175 ( .A(\filter_0/reg_i_9[15] ), .B(n34640), .X(n26982) );
  nand_x1_sg U55176 ( .A(n30025), .B(reg_iii_9[14]), .X(n26979) );
  nand_x1_sg U55177 ( .A(\filter_0/reg_i_9[14] ), .B(n32786), .X(n26980) );
  nand_x1_sg U55178 ( .A(n34039), .B(reg_iii_9[13]), .X(n26977) );
  nand_x1_sg U55179 ( .A(\filter_0/reg_i_9[13] ), .B(n32439), .X(n26978) );
  nand_x1_sg U55180 ( .A(n31085), .B(reg_iii_9[12]), .X(n26975) );
  nand_x1_sg U55181 ( .A(\filter_0/reg_i_9[12] ), .B(n31918), .X(n26976) );
  nand_x1_sg U55182 ( .A(n34914), .B(reg_iii_9[11]), .X(n26973) );
  nand_x1_sg U55183 ( .A(\filter_0/reg_i_9[11] ), .B(n32797), .X(n26974) );
  nand_x1_sg U55184 ( .A(n31069), .B(reg_iii_9[10]), .X(n26971) );
  nand_x1_sg U55185 ( .A(\filter_0/reg_i_9[10] ), .B(n32481), .X(n26972) );
  nand_x1_sg U55186 ( .A(n34041), .B(reg_iii_9[9]), .X(n26969) );
  nand_x1_sg U55187 ( .A(\filter_0/reg_i_9[9] ), .B(n31295), .X(n26970) );
  nand_x1_sg U55188 ( .A(n34604), .B(reg_iii_9[8]), .X(n26967) );
  nand_x1_sg U55189 ( .A(\filter_0/reg_i_9[8] ), .B(n34687), .X(n26968) );
  nand_x1_sg U55190 ( .A(n31533), .B(reg_iii_8[14]), .X(n26939) );
  nand_x1_sg U55191 ( .A(\filter_0/reg_i_8[14] ), .B(n31209), .X(n26940) );
  nand_x1_sg U55192 ( .A(n34888), .B(reg_iii_8[13]), .X(n26937) );
  nand_x1_sg U55193 ( .A(\filter_0/reg_i_8[13] ), .B(n34645), .X(n26938) );
  nand_x1_sg U55194 ( .A(n33900), .B(reg_iii_8[12]), .X(n26935) );
  nand_x1_sg U55195 ( .A(\filter_0/reg_i_8[12] ), .B(n35072), .X(n26936) );
  nand_x1_sg U55196 ( .A(n34021), .B(reg_iii_8[11]), .X(n26933) );
  nand_x1_sg U55197 ( .A(\filter_0/reg_i_8[11] ), .B(n34648), .X(n26934) );
  nand_x1_sg U55198 ( .A(n34908), .B(reg_iii_8[10]), .X(n26931) );
  nand_x1_sg U55199 ( .A(\filter_0/reg_i_8[10] ), .B(n30736), .X(n26932) );
  nand_x1_sg U55200 ( .A(n31242), .B(reg_iii_8[9]), .X(n26929) );
  nand_x1_sg U55201 ( .A(\filter_0/reg_i_8[9] ), .B(n31208), .X(n26930) );
  nand_x1_sg U55202 ( .A(n33909), .B(reg_iii_8[8]), .X(n26927) );
  nand_x1_sg U55203 ( .A(\filter_0/reg_i_8[8] ), .B(n32875), .X(n26928) );
  nand_x1_sg U55204 ( .A(n30028), .B(reg_iii_8[7]), .X(n26925) );
  nand_x1_sg U55205 ( .A(\filter_0/reg_i_8[7] ), .B(n34633), .X(n26926) );
  nand_x1_sg U55206 ( .A(n29698), .B(reg_iii_8[6]), .X(n26923) );
  nand_x1_sg U55207 ( .A(\filter_0/reg_i_8[6] ), .B(n32862), .X(n26924) );
  nand_x1_sg U55208 ( .A(n32268), .B(reg_iii_8[5]), .X(n26921) );
  nand_x1_sg U55209 ( .A(\filter_0/reg_i_8[5] ), .B(n30252), .X(n26922) );
  nand_x1_sg U55210 ( .A(n34891), .B(reg_iii_8[4]), .X(n26919) );
  nand_x1_sg U55211 ( .A(\filter_0/reg_i_8[4] ), .B(n32479), .X(n26920) );
  nand_x1_sg U55212 ( .A(n34888), .B(reg_iii_8[3]), .X(n26917) );
  nand_x1_sg U55213 ( .A(\filter_0/reg_i_8[3] ), .B(n31294), .X(n26918) );
  nand_x1_sg U55214 ( .A(n32260), .B(reg_iii_8[2]), .X(n26915) );
  nand_x1_sg U55215 ( .A(\filter_0/reg_i_8[2] ), .B(n31917), .X(n26916) );
  nand_x1_sg U55216 ( .A(n34914), .B(reg_iii_8[1]), .X(n26913) );
  nand_x1_sg U55217 ( .A(\filter_0/reg_i_8[1] ), .B(n34647), .X(n26914) );
  nand_x1_sg U55218 ( .A(n31080), .B(reg_iii_8[0]), .X(n26911) );
  nand_x1_sg U55219 ( .A(\filter_0/reg_i_8[0] ), .B(n32791), .X(n26912) );
  nand_x1_sg U55220 ( .A(n34012), .B(reg_iii_7[19]), .X(n26909) );
  nand_x1_sg U55221 ( .A(\filter_0/reg_i_7[19] ), .B(n34673), .X(n26910) );
  nand_x1_sg U55222 ( .A(n30387), .B(reg_iii_7[18]), .X(n26907) );
  nand_x1_sg U55223 ( .A(\filter_0/reg_i_7[18] ), .B(n32800), .X(n26908) );
  nand_x1_sg U55224 ( .A(n30031), .B(reg_iii_7[17]), .X(n26905) );
  nand_x1_sg U55225 ( .A(\filter_0/reg_i_7[17] ), .B(n31911), .X(n26906) );
  nand_x1_sg U55226 ( .A(n30029), .B(reg_iii_7[16]), .X(n26903) );
  nand_x1_sg U55227 ( .A(\filter_0/reg_i_7[16] ), .B(n32824), .X(n26904) );
  nand_x1_sg U55228 ( .A(n34909), .B(reg_iii_7[15]), .X(n26901) );
  nand_x1_sg U55229 ( .A(\filter_0/reg_i_7[15] ), .B(n32804), .X(n26902) );
  nand_x1_sg U55230 ( .A(n34606), .B(reg_iii_7[14]), .X(n26899) );
  nand_x1_sg U55231 ( .A(\filter_0/reg_i_7[14] ), .B(n32875), .X(n26900) );
  nand_x1_sg U55232 ( .A(n31677), .B(reg_iii_7[13]), .X(n26897) );
  nand_x1_sg U55233 ( .A(\filter_0/reg_i_7[13] ), .B(n31209), .X(n26898) );
  nand_x1_sg U55234 ( .A(n34035), .B(reg_iii_7[12]), .X(n26895) );
  nand_x1_sg U55235 ( .A(\filter_0/reg_i_7[12] ), .B(n32462), .X(n26896) );
  nand_x1_sg U55236 ( .A(n34039), .B(reg_iii_7[11]), .X(n26893) );
  nand_x1_sg U55237 ( .A(\filter_0/reg_i_7[11] ), .B(n32806), .X(n26894) );
  nand_x1_sg U55238 ( .A(n32258), .B(reg_iii_7[10]), .X(n26891) );
  nand_x1_sg U55239 ( .A(\filter_0/reg_i_7[10] ), .B(n32781), .X(n26892) );
  nand_x1_sg U55240 ( .A(n34879), .B(reg_iii_7[9]), .X(n26889) );
  nand_x1_sg U55241 ( .A(\filter_0/reg_i_7[9] ), .B(n34643), .X(n26890) );
  nand_x1_sg U55242 ( .A(n31533), .B(reg_iii_7[8]), .X(n26887) );
  nand_x1_sg U55243 ( .A(\filter_0/reg_i_7[8] ), .B(n34686), .X(n26888) );
  nand_x1_sg U55244 ( .A(n31516), .B(reg_iii_7[7]), .X(n26885) );
  nand_x1_sg U55245 ( .A(\filter_0/reg_i_7[7] ), .B(n30250), .X(n26886) );
  nand_x1_sg U55246 ( .A(n33920), .B(reg_iii_7[6]), .X(n26883) );
  nand_x1_sg U55247 ( .A(\filter_0/reg_i_7[6] ), .B(n30732), .X(n26884) );
  nand_x1_sg U55248 ( .A(n34028), .B(reg_iii_7[5]), .X(n26881) );
  nand_x1_sg U55249 ( .A(\filter_0/reg_i_7[5] ), .B(n32458), .X(n26882) );
  nand_x1_sg U55250 ( .A(n35412), .B(reg_iii_7[4]), .X(n26879) );
  nand_x1_sg U55251 ( .A(\filter_0/reg_i_7[4] ), .B(n34647), .X(n26880) );
  nand_x1_sg U55252 ( .A(n32256), .B(reg_iii_7[3]), .X(n26877) );
  nand_x1_sg U55253 ( .A(\filter_0/reg_i_7[3] ), .B(n34630), .X(n26878) );
  nand_x1_sg U55254 ( .A(n33899), .B(reg_iii_6[4]), .X(n26839) );
  nand_x1_sg U55255 ( .A(\filter_0/reg_i_6[4] ), .B(n32816), .X(n26840) );
  nand_x1_sg U55256 ( .A(n31521), .B(reg_iii_6[3]), .X(n26837) );
  nand_x1_sg U55257 ( .A(\filter_0/reg_i_6[3] ), .B(n32815), .X(n26838) );
  nand_x1_sg U55258 ( .A(n33907), .B(reg_iii_6[2]), .X(n26835) );
  nand_x1_sg U55259 ( .A(\filter_0/reg_i_6[2] ), .B(n32796), .X(n26836) );
  nand_x1_sg U55260 ( .A(n31685), .B(reg_iii_6[1]), .X(n26833) );
  nand_x1_sg U55261 ( .A(\filter_0/reg_i_6[1] ), .B(n32789), .X(n26834) );
  nand_x1_sg U55262 ( .A(n32256), .B(reg_iii_6[0]), .X(n26831) );
  nand_x1_sg U55263 ( .A(\filter_0/reg_i_6[0] ), .B(n32471), .X(n26832) );
  nand_x1_sg U55264 ( .A(n31064), .B(reg_iii_5[19]), .X(n26829) );
  nand_x1_sg U55265 ( .A(\filter_0/reg_i_5[19] ), .B(n34634), .X(n26830) );
  nand_x1_sg U55266 ( .A(n30158), .B(reg_iii_5[18]), .X(n26827) );
  nand_x1_sg U55267 ( .A(\filter_0/reg_i_5[18] ), .B(n30741), .X(n26828) );
  nand_x1_sg U55268 ( .A(n32277), .B(reg_iii_5[17]), .X(n26825) );
  nand_x1_sg U55269 ( .A(\filter_0/reg_i_5[17] ), .B(n30168), .X(n26826) );
  nand_x1_sg U55270 ( .A(n31089), .B(reg_iii_5[16]), .X(n26823) );
  nand_x1_sg U55271 ( .A(\filter_0/reg_i_5[16] ), .B(n34625), .X(n26824) );
  nand_x1_sg U55272 ( .A(n33904), .B(reg_iii_5[15]), .X(n26821) );
  nand_x1_sg U55273 ( .A(\filter_0/reg_i_5[15] ), .B(n30738), .X(n26822) );
  nand_x1_sg U55274 ( .A(n32264), .B(reg_iii_5[14]), .X(n26819) );
  nand_x1_sg U55275 ( .A(\filter_0/reg_i_5[14] ), .B(n32467), .X(n26820) );
  nand_x1_sg U55276 ( .A(n29690), .B(reg_iii_5[13]), .X(n26817) );
  nand_x1_sg U55277 ( .A(\filter_0/reg_i_5[13] ), .B(n32433), .X(n26818) );
  nand_x1_sg U55278 ( .A(n34035), .B(reg_iii_5[12]), .X(n26815) );
  nand_x1_sg U55279 ( .A(\filter_0/reg_i_5[12] ), .B(n34687), .X(n26816) );
  nand_x1_sg U55280 ( .A(n32276), .B(reg_iii_5[11]), .X(n26813) );
  nand_x1_sg U55281 ( .A(\filter_0/reg_i_5[11] ), .B(n30733), .X(n26814) );
  nand_x1_sg U55282 ( .A(n30625), .B(reg_iii_5[10]), .X(n26811) );
  nand_x1_sg U55283 ( .A(\filter_0/reg_i_5[10] ), .B(n32781), .X(n26812) );
  nand_x1_sg U55284 ( .A(n32265), .B(reg_iii_5[9]), .X(n26809) );
  nand_x1_sg U55285 ( .A(\filter_0/reg_i_5[9] ), .B(n30736), .X(n26810) );
  nand_x1_sg U55286 ( .A(n34008), .B(reg_iii_5[8]), .X(n26807) );
  nand_x1_sg U55287 ( .A(\filter_0/reg_i_5[8] ), .B(n32802), .X(n26808) );
  nand_x1_sg U55288 ( .A(n31517), .B(reg_iii_5[7]), .X(n26805) );
  nand_x1_sg U55289 ( .A(\filter_0/reg_i_5[7] ), .B(n34685), .X(n26806) );
  nand_x1_sg U55290 ( .A(n32258), .B(reg_iii_5[6]), .X(n26803) );
  nand_x1_sg U55291 ( .A(\filter_0/reg_i_5[6] ), .B(n34623), .X(n26804) );
  nand_x1_sg U55292 ( .A(n31532), .B(reg_iii_5[4]), .X(n26799) );
  nand_x1_sg U55293 ( .A(\filter_0/reg_i_5[4] ), .B(n32434), .X(n26800) );
  nand_x1_sg U55294 ( .A(n34886), .B(reg_iii_5[3]), .X(n26797) );
  nand_x1_sg U55295 ( .A(\filter_0/reg_i_5[3] ), .B(n32811), .X(n26798) );
  nand_x1_sg U55296 ( .A(n31528), .B(reg_iii_5[2]), .X(n26795) );
  nand_x1_sg U55297 ( .A(\filter_0/reg_i_5[2] ), .B(n31208), .X(n26796) );
  nand_x1_sg U55298 ( .A(n30933), .B(reg_iii_5[1]), .X(n26793) );
  nand_x1_sg U55299 ( .A(\filter_0/reg_i_5[1] ), .B(n32795), .X(n26794) );
  nand_x1_sg U55300 ( .A(n30923), .B(reg_iii_5[0]), .X(n26791) );
  nand_x1_sg U55301 ( .A(\filter_0/reg_i_5[0] ), .B(n32476), .X(n26792) );
  nand_x1_sg U55302 ( .A(n34904), .B(reg_iii_4[19]), .X(n26789) );
  nand_x1_sg U55303 ( .A(\filter_0/reg_i_4[19] ), .B(n32807), .X(n26790) );
  nand_x1_sg U55304 ( .A(n31074), .B(reg_iii_4[18]), .X(n26787) );
  nand_x1_sg U55305 ( .A(\filter_0/reg_i_4[18] ), .B(n32457), .X(n26788) );
  nand_x1_sg U55306 ( .A(n33893), .B(reg_iii_4[17]), .X(n26785) );
  nand_x1_sg U55307 ( .A(\filter_0/reg_i_4[17] ), .B(n30767), .X(n26786) );
  nand_x1_sg U55308 ( .A(n31532), .B(reg_iii_4[16]), .X(n26783) );
  nand_x1_sg U55309 ( .A(\filter_0/reg_i_4[16] ), .B(n32784), .X(n26784) );
  nand_x1_sg U55310 ( .A(n29698), .B(reg_iii_4[15]), .X(n26781) );
  nand_x1_sg U55311 ( .A(\filter_0/reg_i_4[15] ), .B(n32796), .X(n26782) );
  nand_x1_sg U55312 ( .A(n34911), .B(reg_iii_4[14]), .X(n26779) );
  nand_x1_sg U55313 ( .A(\filter_0/reg_i_4[14] ), .B(n32432), .X(n26780) );
  nand_x1_sg U55314 ( .A(n31679), .B(reg_iii_4[13]), .X(n26777) );
  nand_x1_sg U55315 ( .A(\filter_0/reg_i_4[13] ), .B(n32477), .X(n26778) );
  nand_x1_sg U55316 ( .A(n31524), .B(reg_iii_4[12]), .X(n26775) );
  nand_x1_sg U55317 ( .A(\filter_0/reg_i_4[12] ), .B(n32789), .X(n26776) );
  nand_x1_sg U55318 ( .A(n30777), .B(reg_iii_4[11]), .X(n26773) );
  nand_x1_sg U55319 ( .A(\filter_0/reg_i_4[11] ), .B(n32876), .X(n26774) );
  nand_x1_sg U55320 ( .A(n33902), .B(reg_iii_4[10]), .X(n26771) );
  nand_x1_sg U55321 ( .A(\filter_0/reg_i_4[10] ), .B(n32874), .X(n26772) );
  nand_x1_sg U55322 ( .A(n34008), .B(reg_iii_4[9]), .X(n26769) );
  nand_x1_sg U55323 ( .A(\filter_0/reg_i_4[9] ), .B(n32431), .X(n26770) );
  nand_x1_sg U55324 ( .A(n33939), .B(reg_iii_4[8]), .X(n26767) );
  nand_x1_sg U55325 ( .A(\filter_0/reg_i_4[8] ), .B(n32471), .X(n26768) );
  nand_x1_sg U55326 ( .A(n34907), .B(reg_iii_4[7]), .X(n26765) );
  nand_x1_sg U55327 ( .A(\filter_0/reg_i_4[7] ), .B(n32472), .X(n26766) );
  nand_x1_sg U55328 ( .A(n34012), .B(reg_iii_4[6]), .X(n26763) );
  nand_x1_sg U55329 ( .A(\filter_0/reg_i_4[6] ), .B(n32796), .X(n26764) );
  nand_x1_sg U55330 ( .A(n33918), .B(reg_iii_4[5]), .X(n26761) );
  nand_x1_sg U55331 ( .A(\filter_0/reg_i_4[5] ), .B(n30765), .X(n26762) );
  nand_x1_sg U55332 ( .A(n31521), .B(reg_iii_4[4]), .X(n26759) );
  nand_x1_sg U55333 ( .A(\filter_0/reg_i_4[4] ), .B(n32799), .X(n26760) );
  nand_x1_sg U55334 ( .A(n32268), .B(reg_iii_4[3]), .X(n26757) );
  nand_x1_sg U55335 ( .A(\filter_0/reg_i_4[3] ), .B(n32784), .X(n26758) );
  nand_x1_sg U55336 ( .A(n33938), .B(reg_iii_4[2]), .X(n26755) );
  nand_x1_sg U55337 ( .A(\filter_0/reg_i_4[2] ), .B(n32467), .X(n26756) );
  nand_x1_sg U55338 ( .A(n31683), .B(reg_iii_4[1]), .X(n26753) );
  nand_x1_sg U55339 ( .A(\filter_0/reg_i_4[1] ), .B(n34687), .X(n26754) );
  nand_x1_sg U55340 ( .A(n31517), .B(reg_iii_4[0]), .X(n26751) );
  nand_x1_sg U55341 ( .A(\filter_0/reg_i_4[0] ), .B(n32805), .X(n26752) );
  nand_x1_sg U55342 ( .A(n34608), .B(reg_iii_3[19]), .X(n26749) );
  nand_x1_sg U55343 ( .A(\filter_0/reg_i_3[19] ), .B(n32435), .X(n26750) );
  nand_x1_sg U55344 ( .A(n31242), .B(reg_iii_3[18]), .X(n26747) );
  nand_x1_sg U55345 ( .A(\filter_0/reg_i_3[18] ), .B(n32437), .X(n26748) );
  nand_x1_sg U55346 ( .A(n34012), .B(reg_iii_3[17]), .X(n26745) );
  nand_x1_sg U55347 ( .A(\filter_0/reg_i_3[17] ), .B(n34645), .X(n26746) );
  nand_x1_sg U55348 ( .A(n31079), .B(reg_iii_3[16]), .X(n26743) );
  nand_x1_sg U55349 ( .A(\filter_0/reg_i_3[16] ), .B(n31914), .X(n26744) );
  nand_x1_sg U55350 ( .A(n34026), .B(reg_iii_3[15]), .X(n26741) );
  nand_x1_sg U55351 ( .A(\filter_0/reg_i_3[15] ), .B(n32461), .X(n26742) );
  nand_x1_sg U55352 ( .A(n34028), .B(reg_iii_3[14]), .X(n26739) );
  nand_x1_sg U55353 ( .A(\filter_0/reg_i_3[14] ), .B(n32794), .X(n26740) );
  nand_x1_sg U55354 ( .A(n31064), .B(reg_iii_3[13]), .X(n26737) );
  nand_x1_sg U55355 ( .A(\filter_0/reg_i_3[13] ), .B(n32482), .X(n26738) );
  nand_x1_sg U55356 ( .A(n31248), .B(reg_iii_3[12]), .X(n26735) );
  nand_x1_sg U55357 ( .A(\filter_0/reg_i_3[12] ), .B(n34680), .X(n26736) );
  nand_x1_sg U55358 ( .A(n30929), .B(reg_iii_3[11]), .X(n26733) );
  nand_x1_sg U55359 ( .A(\filter_0/reg_i_3[11] ), .B(n32797), .X(n26734) );
  nand_x1_sg U55360 ( .A(n34019), .B(reg_iii_3[10]), .X(n26731) );
  nand_x1_sg U55361 ( .A(\filter_0/reg_i_3[10] ), .B(n32881), .X(n26732) );
  nand_x1_sg U55362 ( .A(n31089), .B(reg_iii_3[9]), .X(n26729) );
  nand_x1_sg U55363 ( .A(\filter_0/reg_i_3[9] ), .B(n34691), .X(n26730) );
  nand_x1_sg U55364 ( .A(n32259), .B(reg_iii_3[8]), .X(n26727) );
  nand_x1_sg U55365 ( .A(\filter_0/reg_i_3[8] ), .B(n32824), .X(n26728) );
  nand_x1_sg U55366 ( .A(n32276), .B(reg_iii_3[7]), .X(n26725) );
  nand_x1_sg U55367 ( .A(\filter_0/reg_i_3[7] ), .B(n30735), .X(n26726) );
  nand_x1_sg U55368 ( .A(n31074), .B(reg_iii_3[6]), .X(n26723) );
  nand_x1_sg U55369 ( .A(\filter_0/reg_i_3[6] ), .B(n32462), .X(n26724) );
  nand_x1_sg U55370 ( .A(n34013), .B(reg_iii_3[5]), .X(n26721) );
  nand_x1_sg U55371 ( .A(\filter_0/reg_i_3[5] ), .B(n32485), .X(n26722) );
  nand_x1_sg U55372 ( .A(n30929), .B(reg_iii_3[4]), .X(n26719) );
  nand_x1_sg U55373 ( .A(\filter_0/reg_i_3[4] ), .B(n32436), .X(n26720) );
  nand_x1_sg U55374 ( .A(n31090), .B(reg_iii_3[3]), .X(n26717) );
  nand_x1_sg U55375 ( .A(\filter_0/reg_i_3[3] ), .B(n32489), .X(n26718) );
  nand_x1_sg U55376 ( .A(n33889), .B(reg_iii_3[2]), .X(n26715) );
  nand_x1_sg U55377 ( .A(\filter_0/reg_i_3[2] ), .B(n32881), .X(n26716) );
  nand_x1_sg U55378 ( .A(n30625), .B(reg_iii_3[1]), .X(n26713) );
  nand_x1_sg U55379 ( .A(\filter_0/reg_i_3[1] ), .B(n34672), .X(n26714) );
  nand_x1_sg U55380 ( .A(n32256), .B(reg_iii_3[0]), .X(n26711) );
  nand_x1_sg U55381 ( .A(\filter_0/reg_i_3[0] ), .B(n32827), .X(n26712) );
  nand_x1_sg U55382 ( .A(n31065), .B(reg_iii_2[19]), .X(n26709) );
  nand_x1_sg U55383 ( .A(\filter_0/reg_i_2[19] ), .B(n34693), .X(n26710) );
  nand_x1_sg U55384 ( .A(n32268), .B(reg_iii_2[18]), .X(n26707) );
  nand_x1_sg U55385 ( .A(\filter_0/reg_i_2[18] ), .B(n32483), .X(n26708) );
  nand_x1_sg U55386 ( .A(n34908), .B(reg_iii_2[17]), .X(n26705) );
  nand_x1_sg U55387 ( .A(\filter_0/reg_i_2[17] ), .B(n35072), .X(n26706) );
  nand_x1_sg U55388 ( .A(n32277), .B(reg_iii_2[16]), .X(n26703) );
  nand_x1_sg U55389 ( .A(\filter_0/reg_i_2[16] ), .B(n32799), .X(n26704) );
  nand_x1_sg U55390 ( .A(n31248), .B(reg_iii_2[15]), .X(n26701) );
  nand_x1_sg U55391 ( .A(\filter_0/reg_i_2[15] ), .B(n32463), .X(n26702) );
  nand_x1_sg U55392 ( .A(n33941), .B(reg_iii_2[14]), .X(n26699) );
  nand_x1_sg U55393 ( .A(\filter_0/reg_i_2[14] ), .B(n30767), .X(n26700) );
  nand_x1_sg U55394 ( .A(n30937), .B(reg_iii_2[13]), .X(n26697) );
  nand_x1_sg U55395 ( .A(\filter_0/reg_i_2[13] ), .B(n34685), .X(n26698) );
  nand_x1_sg U55396 ( .A(n34909), .B(reg_iii_2[12]), .X(n26695) );
  nand_x1_sg U55397 ( .A(\filter_0/reg_i_2[12] ), .B(n31293), .X(n26696) );
  nand_x1_sg U55398 ( .A(n33923), .B(reg_iii_2[11]), .X(n26693) );
  nand_x1_sg U55399 ( .A(\filter_0/reg_i_2[11] ), .B(n34641), .X(n26694) );
  nand_x1_sg U55400 ( .A(n31677), .B(reg_iii_2[10]), .X(n26691) );
  nand_x1_sg U55401 ( .A(\filter_0/reg_i_2[10] ), .B(n32434), .X(n26692) );
  nand_x1_sg U55402 ( .A(n34026), .B(reg_iii_2[9]), .X(n26689) );
  nand_x1_sg U55403 ( .A(\filter_0/reg_i_2[9] ), .B(n34625), .X(n26690) );
  nand_x1_sg U55404 ( .A(n31526), .B(reg_iii_2[8]), .X(n26687) );
  nand_x1_sg U55405 ( .A(\filter_0/reg_i_2[8] ), .B(n34620), .X(n26688) );
  nand_x1_sg U55406 ( .A(n34878), .B(reg_iii_2[7]), .X(n26685) );
  nand_x1_sg U55407 ( .A(\filter_0/reg_i_2[7] ), .B(n32431), .X(n26686) );
  nand_x1_sg U55408 ( .A(n32265), .B(reg_iii_2[6]), .X(n26683) );
  nand_x1_sg U55409 ( .A(\filter_0/reg_i_2[6] ), .B(n32786), .X(n26684) );
  nand_x1_sg U55410 ( .A(n33904), .B(reg_iii_2[5]), .X(n26681) );
  nand_x1_sg U55411 ( .A(\filter_0/reg_i_2[5] ), .B(n32866), .X(n26682) );
  nand_x1_sg U55412 ( .A(n31532), .B(reg_iii_2[4]), .X(n26679) );
  nand_x1_sg U55413 ( .A(\filter_0/reg_i_2[4] ), .B(n34633), .X(n26680) );
  nand_x1_sg U55414 ( .A(n31243), .B(reg_iii_2[3]), .X(n26677) );
  nand_x1_sg U55415 ( .A(\filter_0/reg_i_2[3] ), .B(n35072), .X(n26678) );
  nand_x1_sg U55416 ( .A(n34880), .B(reg_iii_2[2]), .X(n26675) );
  nand_x1_sg U55417 ( .A(\filter_0/reg_i_2[2] ), .B(n34637), .X(n26676) );
  nand_x1_sg U55418 ( .A(n34909), .B(reg_iii_1[2]), .X(n26635) );
  nand_x1_sg U55419 ( .A(\filter_0/reg_i_1[2] ), .B(n31915), .X(n26636) );
  nand_x1_sg U55420 ( .A(n34607), .B(reg_iii_1[1]), .X(n26633) );
  nand_x1_sg U55421 ( .A(\filter_0/reg_i_1[1] ), .B(n32800), .X(n26634) );
  nand_x1_sg U55422 ( .A(n33903), .B(reg_iii_1[0]), .X(n26631) );
  nand_x1_sg U55423 ( .A(\filter_0/reg_i_1[0] ), .B(n32430), .X(n26632) );
  nand_x1_sg U55424 ( .A(n31688), .B(reg_iii_0[19]), .X(n26629) );
  nand_x1_sg U55425 ( .A(\filter_0/reg_i_0[19] ), .B(n35074), .X(n26630) );
  nand_x1_sg U55426 ( .A(n34609), .B(reg_iii_0[18]), .X(n26627) );
  nand_x1_sg U55427 ( .A(\filter_0/reg_i_0[18] ), .B(n32437), .X(n26628) );
  nand_x1_sg U55428 ( .A(n34913), .B(reg_iii_0[17]), .X(n26625) );
  nand_x1_sg U55429 ( .A(\filter_0/reg_i_0[17] ), .B(n35072), .X(n26626) );
  nand_x1_sg U55430 ( .A(n31682), .B(reg_iii_0[16]), .X(n26623) );
  nand_x1_sg U55431 ( .A(\filter_0/reg_i_0[16] ), .B(n32874), .X(n26624) );
  nand_x1_sg U55432 ( .A(n34022), .B(reg_iii_0[15]), .X(n26621) );
  nand_x1_sg U55433 ( .A(\filter_0/reg_i_0[15] ), .B(n30742), .X(n26622) );
  nand_x1_sg U55434 ( .A(n34009), .B(reg_iii_0[14]), .X(n26619) );
  nand_x1_sg U55435 ( .A(\filter_0/reg_i_0[14] ), .B(n32491), .X(n26620) );
  nand_x1_sg U55436 ( .A(n32273), .B(reg_iii_0[13]), .X(n26617) );
  nand_x1_sg U55437 ( .A(\filter_0/reg_i_0[13] ), .B(n32810), .X(n26618) );
  nand_x1_sg U55438 ( .A(n31075), .B(reg_iii_0[12]), .X(n26615) );
  nand_x1_sg U55439 ( .A(\filter_0/reg_i_0[12] ), .B(n32436), .X(n26616) );
  nand_x1_sg U55440 ( .A(n34881), .B(reg_iii_0[11]), .X(n26613) );
  nand_x1_sg U55441 ( .A(\filter_0/reg_i_0[11] ), .B(n32872), .X(n26614) );
  nand_x1_sg U55442 ( .A(n34024), .B(reg_iii_0[10]), .X(n26611) );
  nand_x1_sg U55443 ( .A(\filter_0/reg_i_0[10] ), .B(n32876), .X(n26612) );
  nand_x1_sg U55444 ( .A(n34890), .B(reg_iii_0[9]), .X(n26609) );
  nand_x1_sg U55445 ( .A(\filter_0/reg_i_0[9] ), .B(n32477), .X(n26610) );
  nand_x1_sg U55446 ( .A(n34011), .B(reg_iii_0[8]), .X(n26607) );
  nand_x1_sg U55447 ( .A(\filter_0/reg_i_0[8] ), .B(n32484), .X(n26608) );
  nand_x1_sg U55448 ( .A(n34009), .B(reg_iii_0[7]), .X(n26605) );
  nand_x1_sg U55449 ( .A(\filter_0/reg_i_0[7] ), .B(n30757), .X(n26606) );
  nand_x1_sg U55450 ( .A(n31518), .B(reg_iii_0[6]), .X(n26603) );
  nand_x1_sg U55451 ( .A(\filter_0/reg_i_0[6] ), .B(n34693), .X(n26604) );
  nand_x1_sg U55452 ( .A(n34023), .B(reg_iii_0[5]), .X(n26601) );
  nand_x1_sg U55453 ( .A(\filter_0/reg_i_0[5] ), .B(n32875), .X(n26602) );
  nand_x1_sg U55454 ( .A(n31065), .B(reg_iii_0[4]), .X(n26599) );
  nand_x1_sg U55455 ( .A(\filter_0/reg_i_0[4] ), .B(n32471), .X(n26600) );
  nand_x1_sg U55456 ( .A(n34024), .B(reg_iii_0[3]), .X(n26597) );
  nand_x1_sg U55457 ( .A(\filter_0/reg_i_0[3] ), .B(n32463), .X(n26598) );
  nand_x1_sg U55458 ( .A(n33923), .B(reg_iii_0[2]), .X(n26595) );
  nand_x1_sg U55459 ( .A(\filter_0/reg_i_0[2] ), .B(n31209), .X(n26596) );
  nand_x1_sg U55460 ( .A(n34025), .B(reg_iii_0[1]), .X(n26593) );
  nand_x1_sg U55461 ( .A(\filter_0/reg_i_0[1] ), .B(n32795), .X(n26594) );
  nand_x1_sg U55462 ( .A(n32224), .B(reg_iii_0[0]), .X(n26591) );
  nand_x1_sg U55463 ( .A(\filter_0/reg_i_0[0] ), .B(n32785), .X(n26592) );
  nand_x1_sg U55464 ( .A(n33911), .B(n28252), .X(n28250) );
  nand_x1_sg U55465 ( .A(\filter_0/reg_xor_w_mask[31] ), .B(n35073), .X(n28251) );
  nand_x1_sg U55466 ( .A(n28253), .B(n42478), .X(n28252) );
  nand_x1_sg U55467 ( .A(n34891), .B(o_mask[11]), .X(n27893) );
  nand_x1_sg U55468 ( .A(\filter_0/reg_o_mask[11] ), .B(n32475), .X(n27894) );
  nand_x1_sg U55469 ( .A(n33938), .B(o_mask[8]), .X(n27887) );
  nand_x1_sg U55470 ( .A(\filter_0/reg_o_mask[8] ), .B(n32478), .X(n27888) );
  nand_x1_sg U55471 ( .A(n32273), .B(o_mask[5]), .X(n27881) );
  nand_x1_sg U55472 ( .A(\filter_0/reg_o_mask[5] ), .B(n30739), .X(n27882) );
  nand_x1_sg U55473 ( .A(n34903), .B(o_mask[2]), .X(n27875) );
  nand_x1_sg U55474 ( .A(\filter_0/reg_o_mask[2] ), .B(n32471), .X(n27876) );
  nand_x1_sg U55475 ( .A(n31531), .B(n28247), .X(n28245) );
  nand_x1_sg U55476 ( .A(\filter_0/reg_xor_w_mask[30] ), .B(n32489), .X(n28246) );
  nand_x1_sg U55477 ( .A(n28248), .B(n42477), .X(n28247) );
  nand_x1_sg U55478 ( .A(n30386), .B(n28242), .X(n28240) );
  nand_x1_sg U55479 ( .A(\filter_0/reg_xor_w_mask[29] ), .B(n32438), .X(n28241) );
  nand_x1_sg U55480 ( .A(n28243), .B(n42476), .X(n28242) );
  nand_x1_sg U55481 ( .A(n30026), .B(o_mask[13]), .X(n27897) );
  nand_x1_sg U55482 ( .A(\filter_0/reg_o_mask[13] ), .B(n32882), .X(n27898) );
  nand_x1_sg U55483 ( .A(n34023), .B(o_mask[12]), .X(n27895) );
  nand_x1_sg U55484 ( .A(\filter_0/reg_o_mask[12] ), .B(n32860), .X(n27896) );
  nand_x1_sg U55485 ( .A(n30387), .B(o_mask[10]), .X(n27891) );
  nand_x1_sg U55486 ( .A(\filter_0/reg_o_mask[10] ), .B(n32474), .X(n27892) );
  nand_x1_sg U55487 ( .A(n34030), .B(o_mask[9]), .X(n27889) );
  nand_x1_sg U55488 ( .A(\filter_0/reg_o_mask[9] ), .B(n30247), .X(n27890) );
  nand_x1_sg U55489 ( .A(n34017), .B(o_mask[7]), .X(n27885) );
  nand_x1_sg U55490 ( .A(\filter_0/reg_o_mask[7] ), .B(n32869), .X(n27886) );
  nand_x1_sg U55491 ( .A(n32266), .B(o_mask[6]), .X(n27883) );
  nand_x1_sg U55492 ( .A(\filter_0/reg_o_mask[6] ), .B(n32806), .X(n27884) );
  nand_x1_sg U55493 ( .A(n30931), .B(o_mask[4]), .X(n27879) );
  nand_x1_sg U55494 ( .A(\filter_0/reg_o_mask[4] ), .B(n32870), .X(n27880) );
  nand_x1_sg U55495 ( .A(n33919), .B(o_mask[3]), .X(n27877) );
  nand_x1_sg U55496 ( .A(\filter_0/reg_o_mask[3] ), .B(n32468), .X(n27878) );
  nand_x1_sg U55497 ( .A(n33928), .B(o_mask[1]), .X(n27873) );
  nand_x1_sg U55498 ( .A(\filter_0/reg_o_mask[1] ), .B(n32488), .X(n27874) );
  nand_x1_sg U55499 ( .A(n32223), .B(o_mask[0]), .X(n27871) );
  nand_x1_sg U55500 ( .A(\filter_0/reg_o_mask[0] ), .B(n35069), .X(n27872) );
  nand_x1_sg U55501 ( .A(n31679), .B(n28237), .X(n28236) );
  nand_x1_sg U55502 ( .A(\filter_0/reg_xor_w_mask[28] ), .B(n31921), .X(n28235) );
  nand_x1_sg U55503 ( .A(n28238), .B(n42475), .X(n28237) );
  nand_x1_sg U55504 ( .A(n33913), .B(n28222), .X(n28221) );
  nand_x1_sg U55505 ( .A(\filter_0/reg_xor_w_mask[25] ), .B(n30768), .X(n28220) );
  nand_x1_sg U55506 ( .A(n28223), .B(n42472), .X(n28222) );
  nand_x1_sg U55507 ( .A(n33936), .B(n28207), .X(n28206) );
  nand_x1_sg U55508 ( .A(\filter_0/reg_xor_w_mask[22] ), .B(n30761), .X(n28205) );
  nand_x1_sg U55509 ( .A(n28208), .B(n42469), .X(n28207) );
  nand_x1_sg U55510 ( .A(n33939), .B(n28192), .X(n28191) );
  nand_x1_sg U55511 ( .A(\filter_0/reg_xor_w_mask[19] ), .B(n34688), .X(n28190) );
  nand_x1_sg U55512 ( .A(n28193), .B(n42466), .X(n28192) );
  nand_x1_sg U55513 ( .A(n33903), .B(n28177), .X(n28176) );
  nand_x1_sg U55514 ( .A(\filter_0/reg_xor_w_mask[16] ), .B(n34621), .X(n28175) );
  nand_x1_sg U55515 ( .A(n28178), .B(n42463), .X(n28177) );
  nand_x1_sg U55516 ( .A(n33940), .B(n28162), .X(n28161) );
  nand_x1_sg U55517 ( .A(\filter_0/reg_xor_w_mask[13] ), .B(n32787), .X(n28160) );
  nand_x1_sg U55518 ( .A(n28163), .B(n42460), .X(n28162) );
  nand_x1_sg U55519 ( .A(n33933), .B(n28042), .X(n28041) );
  nand_x1_sg U55520 ( .A(\filter_0/reg_xor_i_mask[21] ), .B(n32862), .X(n28040) );
  nand_x1_sg U55521 ( .A(n28043), .B(n42436), .X(n28042) );
  nand_x1_sg U55522 ( .A(n33899), .B(n28232), .X(n28231) );
  nand_x1_sg U55523 ( .A(\filter_0/reg_xor_w_mask[27] ), .B(n35075), .X(n28230) );
  nand_x1_sg U55524 ( .A(n28233), .B(n42474), .X(n28232) );
  nand_x1_sg U55525 ( .A(n33895), .B(n28227), .X(n28226) );
  nand_x1_sg U55526 ( .A(\filter_0/reg_xor_w_mask[26] ), .B(n32882), .X(n28225) );
  nand_x1_sg U55527 ( .A(n28228), .B(n42473), .X(n28227) );
  nand_x1_sg U55528 ( .A(n33931), .B(n28217), .X(n28216) );
  nand_x1_sg U55529 ( .A(\filter_0/reg_xor_w_mask[24] ), .B(n32817), .X(n28215) );
  nand_x1_sg U55530 ( .A(n28218), .B(n42471), .X(n28217) );
  nand_x1_sg U55531 ( .A(n33923), .B(n28212), .X(n28211) );
  nand_x1_sg U55532 ( .A(\filter_0/reg_xor_w_mask[23] ), .B(n32781), .X(n28210) );
  nand_x1_sg U55533 ( .A(n28213), .B(n42470), .X(n28212) );
  nand_x1_sg U55534 ( .A(n33889), .B(n28202), .X(n28201) );
  nand_x1_sg U55535 ( .A(\filter_0/reg_xor_w_mask[21] ), .B(n32827), .X(n28200) );
  nand_x1_sg U55536 ( .A(n28203), .B(n42468), .X(n28202) );
  nand_x1_sg U55537 ( .A(n33919), .B(n28197), .X(n28196) );
  nand_x1_sg U55538 ( .A(\filter_0/reg_xor_w_mask[20] ), .B(n32867), .X(n28195) );
  nand_x1_sg U55539 ( .A(n28198), .B(n42467), .X(n28197) );
  nand_x1_sg U55540 ( .A(n33914), .B(n28187), .X(n28186) );
  nand_x1_sg U55541 ( .A(\filter_0/reg_xor_w_mask[18] ), .B(n32812), .X(n28185) );
  nand_x1_sg U55542 ( .A(n28188), .B(n42465), .X(n28187) );
  nand_x1_sg U55543 ( .A(n33934), .B(n28182), .X(n28181) );
  nand_x1_sg U55544 ( .A(\filter_0/reg_xor_w_mask[17] ), .B(n32792), .X(n28180) );
  nand_x1_sg U55545 ( .A(n28183), .B(n42464), .X(n28182) );
  nand_x1_sg U55546 ( .A(n30204), .B(n28172), .X(n28171) );
  nand_x1_sg U55547 ( .A(\filter_0/reg_xor_w_mask[15] ), .B(n32822), .X(n28170) );
  nand_x1_sg U55548 ( .A(n28173), .B(n42462), .X(n28172) );
  nand_x1_sg U55549 ( .A(n33909), .B(n28167), .X(n28166) );
  nand_x1_sg U55550 ( .A(\filter_0/reg_xor_w_mask[14] ), .B(n32872), .X(n28165) );
  nand_x1_sg U55551 ( .A(n28168), .B(n42461), .X(n28167) );
  nand_x1_sg U55552 ( .A(n31684), .B(n28157), .X(n28156) );
  nand_x1_sg U55553 ( .A(\filter_0/reg_xor_w_mask[12] ), .B(n32791), .X(n28155) );
  nand_x1_sg U55554 ( .A(n28158), .B(n42459), .X(n28157) );
  nand_x1_sg U55555 ( .A(n33908), .B(n28152), .X(n28151) );
  nand_x1_sg U55556 ( .A(\filter_0/reg_xor_w_mask[11] ), .B(n32802), .X(n28150) );
  nand_x1_sg U55557 ( .A(n28153), .B(n42458), .X(n28152) );
  nand_x1_sg U55558 ( .A(n30035), .B(n28037), .X(n28036) );
  nand_x1_sg U55559 ( .A(\filter_0/reg_xor_i_mask[20] ), .B(n34620), .X(n28035) );
  nand_x1_sg U55560 ( .A(n28038), .B(n42435), .X(n28037) );
  nand_x1_sg U55561 ( .A(n30032), .B(n27942), .X(n27941) );
  nand_x1_sg U55562 ( .A(\filter_0/reg_xor_i_mask[1] ), .B(n35070), .X(n27940)
         );
  nand_x1_sg U55563 ( .A(n27943), .B(n42416), .X(n27942) );
  nand_x1_sg U55564 ( .A(n31682), .B(n27937), .X(n27936) );
  nand_x1_sg U55565 ( .A(\filter_0/reg_xor_i_mask[0] ), .B(n34621), .X(n27935)
         );
  nand_x1_sg U55566 ( .A(n27938), .B(n42415), .X(n27937) );
  nand_x1_sg U55567 ( .A(n34609), .B(reg_www_15[7]), .X(n27845) );
  nand_x1_sg U55568 ( .A(\filter_0/reg_w_15[7] ), .B(n32821), .X(n27846) );
  nand_x1_sg U55569 ( .A(n33912), .B(reg_www_15[6]), .X(n27843) );
  nand_x1_sg U55570 ( .A(\filter_0/reg_w_15[6] ), .B(n32812), .X(n27844) );
  nand_x1_sg U55571 ( .A(n31523), .B(reg_www_15[5]), .X(n27841) );
  nand_x1_sg U55572 ( .A(\filter_0/reg_w_15[5] ), .B(n32476), .X(n27842) );
  nand_x1_sg U55573 ( .A(n34603), .B(reg_www_15[4]), .X(n27839) );
  nand_x1_sg U55574 ( .A(\filter_0/reg_w_15[4] ), .B(n32870), .X(n27840) );
  nand_x1_sg U55575 ( .A(n31687), .B(reg_www_15[3]), .X(n27837) );
  nand_x1_sg U55576 ( .A(\filter_0/reg_w_15[3] ), .B(n34691), .X(n27838) );
  nand_x1_sg U55577 ( .A(n31242), .B(reg_www_15[2]), .X(n27835) );
  nand_x1_sg U55578 ( .A(\filter_0/reg_w_15[2] ), .B(n30772), .X(n27836) );
  nand_x1_sg U55579 ( .A(n30923), .B(reg_www_15[1]), .X(n27833) );
  nand_x1_sg U55580 ( .A(\filter_0/reg_w_15[1] ), .B(n32871), .X(n27834) );
  nand_x1_sg U55581 ( .A(n30925), .B(reg_www_15[0]), .X(n27831) );
  nand_x1_sg U55582 ( .A(\filter_0/reg_w_15[0] ), .B(n30732), .X(n27832) );
  nand_x1_sg U55583 ( .A(n33931), .B(reg_www_14[19]), .X(n27829) );
  nand_x1_sg U55584 ( .A(\filter_0/reg_w_14[19] ), .B(n32872), .X(n27830) );
  nand_x1_sg U55585 ( .A(n30159), .B(reg_www_14[18]), .X(n27827) );
  nand_x1_sg U55586 ( .A(\filter_0/reg_w_14[18] ), .B(n32461), .X(n27828) );
  nand_x1_sg U55587 ( .A(n34017), .B(reg_www_14[17]), .X(n27825) );
  nand_x1_sg U55588 ( .A(\filter_0/reg_w_14[17] ), .B(n32816), .X(n27826) );
  nand_x1_sg U55589 ( .A(n31525), .B(reg_www_14[16]), .X(n27823) );
  nand_x1_sg U55590 ( .A(\filter_0/reg_w_14[16] ), .B(n34626), .X(n27824) );
  nand_x1_sg U55591 ( .A(n34022), .B(reg_www_14[15]), .X(n27821) );
  nand_x1_sg U55592 ( .A(\filter_0/reg_w_14[15] ), .B(n30733), .X(n27822) );
  nand_x1_sg U55593 ( .A(n34030), .B(reg_www_14[14]), .X(n27819) );
  nand_x1_sg U55594 ( .A(\filter_0/reg_w_14[14] ), .B(n31296), .X(n27820) );
  nand_x1_sg U55595 ( .A(n29692), .B(reg_www_14[13]), .X(n27817) );
  nand_x1_sg U55596 ( .A(\filter_0/reg_w_14[13] ), .B(n34635), .X(n27818) );
  nand_x1_sg U55597 ( .A(n30933), .B(reg_www_14[12]), .X(n27815) );
  nand_x1_sg U55598 ( .A(\filter_0/reg_w_14[12] ), .B(n32461), .X(n27816) );
  nand_x1_sg U55599 ( .A(n33896), .B(reg_www_14[11]), .X(n27813) );
  nand_x1_sg U55600 ( .A(\filter_0/reg_w_14[11] ), .B(n34676), .X(n27814) );
  nand_x1_sg U55601 ( .A(n31517), .B(reg_www_14[10]), .X(n27811) );
  nand_x1_sg U55602 ( .A(\filter_0/reg_w_14[10] ), .B(n32871), .X(n27812) );
  nand_x1_sg U55603 ( .A(n31524), .B(reg_www_13[10]), .X(n27771) );
  nand_x1_sg U55604 ( .A(\filter_0/reg_w_13[10] ), .B(n32470), .X(n27772) );
  nand_x1_sg U55605 ( .A(n34026), .B(reg_www_13[9]), .X(n27769) );
  nand_x1_sg U55606 ( .A(\filter_0/reg_w_13[9] ), .B(n30744), .X(n27770) );
  nand_x1_sg U55607 ( .A(n32261), .B(reg_www_13[8]), .X(n27767) );
  nand_x1_sg U55608 ( .A(\filter_0/reg_w_13[8] ), .B(n31911), .X(n27768) );
  nand_x1_sg U55609 ( .A(n33912), .B(reg_www_13[7]), .X(n27765) );
  nand_x1_sg U55610 ( .A(\filter_0/reg_w_13[7] ), .B(n32807), .X(n27766) );
  nand_x1_sg U55611 ( .A(n33940), .B(reg_www_13[6]), .X(n27763) );
  nand_x1_sg U55612 ( .A(\filter_0/reg_w_13[6] ), .B(n32824), .X(n27764) );
  nand_x1_sg U55613 ( .A(n34907), .B(reg_www_13[5]), .X(n27761) );
  nand_x1_sg U55614 ( .A(\filter_0/reg_w_13[5] ), .B(n34692), .X(n27762) );
  nand_x1_sg U55615 ( .A(n32224), .B(reg_www_13[4]), .X(n27759) );
  nand_x1_sg U55616 ( .A(\filter_0/reg_w_13[4] ), .B(n31294), .X(n27760) );
  nand_x1_sg U55617 ( .A(n33921), .B(reg_www_13[3]), .X(n27757) );
  nand_x1_sg U55618 ( .A(\filter_0/reg_w_13[3] ), .B(n32792), .X(n27758) );
  nand_x1_sg U55619 ( .A(n33933), .B(reg_www_13[2]), .X(n27755) );
  nand_x1_sg U55620 ( .A(\filter_0/reg_w_13[2] ), .B(n32867), .X(n27756) );
  nand_x1_sg U55621 ( .A(n34022), .B(reg_www_13[1]), .X(n27753) );
  nand_x1_sg U55622 ( .A(\filter_0/reg_w_13[1] ), .B(n32882), .X(n27754) );
  nand_x1_sg U55623 ( .A(n30028), .B(reg_www_13[0]), .X(n27751) );
  nand_x1_sg U55624 ( .A(\filter_0/reg_w_13[0] ), .B(n30739), .X(n27752) );
  nand_x1_sg U55625 ( .A(n30159), .B(reg_www_12[19]), .X(n27749) );
  nand_x1_sg U55626 ( .A(\filter_0/reg_w_12[19] ), .B(n32482), .X(n27750) );
  nand_x1_sg U55627 ( .A(n34034), .B(reg_www_12[18]), .X(n27747) );
  nand_x1_sg U55628 ( .A(\filter_0/reg_w_12[18] ), .B(n32825), .X(n27748) );
  nand_x1_sg U55629 ( .A(n33925), .B(reg_www_12[17]), .X(n27745) );
  nand_x1_sg U55630 ( .A(\filter_0/reg_w_12[17] ), .B(n32861), .X(n27746) );
  nand_x1_sg U55631 ( .A(n35466), .B(reg_www_12[16]), .X(n27743) );
  nand_x1_sg U55632 ( .A(\filter_0/reg_w_12[16] ), .B(n34635), .X(n27744) );
  nand_x1_sg U55633 ( .A(n34008), .B(reg_www_12[15]), .X(n27741) );
  nand_x1_sg U55634 ( .A(\filter_0/reg_w_12[15] ), .B(n32810), .X(n27742) );
  nand_x1_sg U55635 ( .A(n31531), .B(reg_www_12[14]), .X(n27739) );
  nand_x1_sg U55636 ( .A(\filter_0/reg_w_12[14] ), .B(n34623), .X(n27740) );
  nand_x1_sg U55637 ( .A(n34035), .B(reg_www_12[13]), .X(n27737) );
  nand_x1_sg U55638 ( .A(\filter_0/reg_w_12[13] ), .B(n32479), .X(n27738) );
  nand_x1_sg U55639 ( .A(n31519), .B(reg_www_12[12]), .X(n27735) );
  nand_x1_sg U55640 ( .A(\filter_0/reg_w_12[12] ), .B(n34676), .X(n27736) );
  nand_x1_sg U55641 ( .A(n34013), .B(reg_www_12[5]), .X(n27721) );
  nand_x1_sg U55642 ( .A(\filter_0/reg_w_12[5] ), .B(n32483), .X(n27722) );
  nand_x1_sg U55643 ( .A(n31518), .B(reg_www_9[8]), .X(n27607) );
  nand_x1_sg U55644 ( .A(\filter_0/reg_w_9[8] ), .B(n32802), .X(n27608) );
  nand_x1_sg U55645 ( .A(n30629), .B(reg_www_9[7]), .X(n27605) );
  nand_x1_sg U55646 ( .A(\filter_0/reg_w_9[7] ), .B(n35073), .X(n27606) );
  nand_x1_sg U55647 ( .A(n33906), .B(reg_www_9[6]), .X(n27603) );
  nand_x1_sg U55648 ( .A(\filter_0/reg_w_9[6] ), .B(n32814), .X(n27604) );
  nand_x1_sg U55649 ( .A(n33892), .B(reg_www_9[5]), .X(n27601) );
  nand_x1_sg U55650 ( .A(\filter_0/reg_w_9[5] ), .B(n32825), .X(n27602) );
  nand_x1_sg U55651 ( .A(n32270), .B(reg_www_9[4]), .X(n27599) );
  nand_x1_sg U55652 ( .A(\filter_0/reg_w_9[4] ), .B(n34637), .X(n27600) );
  nand_x1_sg U55653 ( .A(n31527), .B(reg_www_9[3]), .X(n27597) );
  nand_x1_sg U55654 ( .A(\filter_0/reg_w_9[3] ), .B(n31292), .X(n27598) );
  nand_x1_sg U55655 ( .A(n34008), .B(reg_www_8[3]), .X(n27557) );
  nand_x1_sg U55656 ( .A(\filter_0/reg_w_8[3] ), .B(n34678), .X(n27558) );
  nand_x1_sg U55657 ( .A(n34009), .B(reg_www_8[2]), .X(n27555) );
  nand_x1_sg U55658 ( .A(\filter_0/reg_w_8[2] ), .B(n30249), .X(n27556) );
  nand_x1_sg U55659 ( .A(n34879), .B(reg_www_8[1]), .X(n27553) );
  nand_x1_sg U55660 ( .A(\filter_0/reg_w_8[1] ), .B(n31916), .X(n27554) );
  nand_x1_sg U55661 ( .A(n31685), .B(reg_www_8[0]), .X(n27551) );
  nand_x1_sg U55662 ( .A(\filter_0/reg_w_8[0] ), .B(n30252), .X(n27552) );
  nand_x1_sg U55663 ( .A(n34036), .B(reg_www_7[19]), .X(n27549) );
  nand_x1_sg U55664 ( .A(\filter_0/reg_w_7[19] ), .B(n32784), .X(n27550) );
  nand_x1_sg U55665 ( .A(n31519), .B(reg_www_7[18]), .X(n27547) );
  nand_x1_sg U55666 ( .A(\filter_0/reg_w_7[18] ), .B(n30741), .X(n27548) );
  nand_x1_sg U55667 ( .A(n31527), .B(reg_www_7[17]), .X(n27545) );
  nand_x1_sg U55668 ( .A(\filter_0/reg_w_7[17] ), .B(n35075), .X(n27546) );
  nand_x1_sg U55669 ( .A(n32258), .B(reg_www_7[16]), .X(n27543) );
  nand_x1_sg U55670 ( .A(\filter_0/reg_w_7[16] ), .B(n32795), .X(n27544) );
  nand_x1_sg U55671 ( .A(n31070), .B(reg_www_7[15]), .X(n27541) );
  nand_x1_sg U55672 ( .A(\filter_0/reg_w_7[15] ), .B(n32460), .X(n27542) );
  nand_x1_sg U55673 ( .A(n33936), .B(reg_www_7[14]), .X(n27539) );
  nand_x1_sg U55674 ( .A(\filter_0/reg_w_7[14] ), .B(n35074), .X(n27540) );
  nand_x1_sg U55675 ( .A(n30625), .B(reg_www_7[13]), .X(n27537) );
  nand_x1_sg U55676 ( .A(\filter_0/reg_w_7[13] ), .B(n32433), .X(n27538) );
  nand_x1_sg U55677 ( .A(n34881), .B(reg_www_7[12]), .X(n27535) );
  nand_x1_sg U55678 ( .A(\filter_0/reg_w_7[12] ), .B(n34648), .X(n27536) );
  nand_x1_sg U55679 ( .A(n33895), .B(reg_www_7[11]), .X(n27533) );
  nand_x1_sg U55680 ( .A(\filter_0/reg_w_7[11] ), .B(n34638), .X(n27534) );
  nand_x1_sg U55681 ( .A(n34016), .B(reg_www_5[12]), .X(n27455) );
  nand_x1_sg U55682 ( .A(\filter_0/reg_w_5[12] ), .B(n31293), .X(n27456) );
  nand_x1_sg U55683 ( .A(n31518), .B(reg_www_5[11]), .X(n27453) );
  nand_x1_sg U55684 ( .A(\filter_0/reg_w_5[11] ), .B(n32464), .X(n27454) );
  nand_x1_sg U55685 ( .A(n30925), .B(reg_www_5[10]), .X(n27451) );
  nand_x1_sg U55686 ( .A(\filter_0/reg_w_5[10] ), .B(n32484), .X(n27452) );
  nand_x1_sg U55687 ( .A(n33889), .B(reg_www_5[9]), .X(n27449) );
  nand_x1_sg U55688 ( .A(\filter_0/reg_w_5[9] ), .B(n32880), .X(n27450) );
  nand_x1_sg U55689 ( .A(n34880), .B(reg_www_5[8]), .X(n27447) );
  nand_x1_sg U55690 ( .A(\filter_0/reg_w_5[8] ), .B(n30733), .X(n27448) );
  nand_x1_sg U55691 ( .A(n33933), .B(reg_www_5[7]), .X(n27445) );
  nand_x1_sg U55692 ( .A(\filter_0/reg_w_5[7] ), .B(n32469), .X(n27446) );
  nand_x1_sg U55693 ( .A(n31065), .B(reg_www_5[6]), .X(n27443) );
  nand_x1_sg U55694 ( .A(\filter_0/reg_w_5[6] ), .B(n34678), .X(n27444) );
  nand_x1_sg U55695 ( .A(n29696), .B(reg_www_5[5]), .X(n27441) );
  nand_x1_sg U55696 ( .A(\filter_0/reg_w_5[5] ), .B(n32812), .X(n27442) );
  nand_x1_sg U55697 ( .A(n29689), .B(reg_www_5[4]), .X(n27439) );
  nand_x1_sg U55698 ( .A(\filter_0/reg_w_5[4] ), .B(n32435), .X(n27440) );
  nand_x1_sg U55699 ( .A(n34890), .B(reg_www_5[3]), .X(n27437) );
  nand_x1_sg U55700 ( .A(\filter_0/reg_w_5[3] ), .B(n30252), .X(n27438) );
  nand_x1_sg U55701 ( .A(n33912), .B(reg_www_5[2]), .X(n27435) );
  nand_x1_sg U55702 ( .A(\filter_0/reg_w_5[2] ), .B(n31296), .X(n27436) );
  nand_x1_sg U55703 ( .A(n31680), .B(reg_www_5[1]), .X(n27433) );
  nand_x1_sg U55704 ( .A(\filter_0/reg_w_5[1] ), .B(n32811), .X(n27434) );
  nand_x1_sg U55705 ( .A(n31243), .B(reg_www_4[7]), .X(n27405) );
  nand_x1_sg U55706 ( .A(\filter_0/reg_w_4[7] ), .B(n32437), .X(n27406) );
  nand_x1_sg U55707 ( .A(n35159), .B(reg_www_4[6]), .X(n27403) );
  nand_x1_sg U55708 ( .A(\filter_0/reg_w_4[6] ), .B(n34671), .X(n27404) );
  nand_x1_sg U55709 ( .A(n34041), .B(reg_www_4[5]), .X(n27401) );
  nand_x1_sg U55710 ( .A(\filter_0/reg_w_4[5] ), .B(n32859), .X(n27402) );
  nand_x1_sg U55711 ( .A(n31530), .B(reg_www_4[4]), .X(n27399) );
  nand_x1_sg U55712 ( .A(\filter_0/reg_w_4[4] ), .B(n32478), .X(n27400) );
  nand_x1_sg U55713 ( .A(n34033), .B(reg_www_4[3]), .X(n27397) );
  nand_x1_sg U55714 ( .A(\filter_0/reg_w_4[3] ), .B(n32822), .X(n27398) );
  nand_x1_sg U55715 ( .A(n31687), .B(reg_www_4[2]), .X(n27395) );
  nand_x1_sg U55716 ( .A(\filter_0/reg_w_4[2] ), .B(n34646), .X(n27396) );
  nand_x1_sg U55717 ( .A(n34034), .B(reg_www_4[1]), .X(n27393) );
  nand_x1_sg U55718 ( .A(\filter_0/reg_w_4[1] ), .B(n32861), .X(n27394) );
  nand_x1_sg U55719 ( .A(n34029), .B(reg_www_4[0]), .X(n27391) );
  nand_x1_sg U55720 ( .A(\filter_0/reg_w_4[0] ), .B(n32869), .X(n27392) );
  nand_x1_sg U55721 ( .A(n34889), .B(reg_www_3[19]), .X(n27389) );
  nand_x1_sg U55722 ( .A(\filter_0/reg_w_3[19] ), .B(n34648), .X(n27390) );
  nand_x1_sg U55723 ( .A(n33900), .B(reg_www_3[18]), .X(n27387) );
  nand_x1_sg U55724 ( .A(\filter_0/reg_w_3[18] ), .B(n32860), .X(n27388) );
  nand_x1_sg U55725 ( .A(n31527), .B(reg_www_3[17]), .X(n27385) );
  nand_x1_sg U55726 ( .A(\filter_0/reg_w_3[17] ), .B(n34625), .X(n27386) );
  nand_x1_sg U55727 ( .A(n32255), .B(reg_www_3[16]), .X(n27383) );
  nand_x1_sg U55728 ( .A(\filter_0/reg_w_3[16] ), .B(n34637), .X(n27384) );
  nand_x1_sg U55729 ( .A(n33890), .B(reg_www_3[15]), .X(n27381) );
  nand_x1_sg U55730 ( .A(\filter_0/reg_w_3[15] ), .B(n30773), .X(n27382) );
  nand_x1_sg U55731 ( .A(n30629), .B(reg_www_3[14]), .X(n27379) );
  nand_x1_sg U55732 ( .A(\filter_0/reg_w_3[14] ), .B(n32825), .X(n27380) );
  nand_x1_sg U55733 ( .A(n33913), .B(reg_www_3[13]), .X(n27377) );
  nand_x1_sg U55734 ( .A(\filter_0/reg_w_3[13] ), .B(n30735), .X(n27378) );
  nand_x1_sg U55735 ( .A(n33935), .B(reg_www_3[12]), .X(n27375) );
  nand_x1_sg U55736 ( .A(\filter_0/reg_w_3[12] ), .B(n32485), .X(n27376) );
  nand_x1_sg U55737 ( .A(n33906), .B(reg_www_3[11]), .X(n27373) );
  nand_x1_sg U55738 ( .A(\filter_0/reg_w_3[11] ), .B(n32478), .X(n27374) );
  nand_x1_sg U55739 ( .A(n31247), .B(reg_www_3[10]), .X(n27371) );
  nand_x1_sg U55740 ( .A(\filter_0/reg_w_3[10] ), .B(n32491), .X(n27372) );
  nand_x1_sg U55741 ( .A(n33899), .B(reg_www_3[9]), .X(n27369) );
  nand_x1_sg U55742 ( .A(\filter_0/reg_w_3[9] ), .B(n34686), .X(n27370) );
  nand_x1_sg U55743 ( .A(n31070), .B(reg_www_2[16]), .X(n27343) );
  nand_x1_sg U55744 ( .A(\filter_0/reg_w_2[16] ), .B(n34626), .X(n27344) );
  nand_x1_sg U55745 ( .A(n33897), .B(reg_www_2[15]), .X(n27341) );
  nand_x1_sg U55746 ( .A(\filter_0/reg_w_2[15] ), .B(n31918), .X(n27342) );
  nand_x1_sg U55747 ( .A(n31526), .B(reg_www_2[14]), .X(n27339) );
  nand_x1_sg U55748 ( .A(\filter_0/reg_w_2[14] ), .B(n31917), .X(n27340) );
  nand_x1_sg U55749 ( .A(n31064), .B(reg_www_2[13]), .X(n27337) );
  nand_x1_sg U55750 ( .A(\filter_0/reg_w_2[13] ), .B(n31293), .X(n27338) );
  nand_x1_sg U55751 ( .A(n31678), .B(reg_www_2[12]), .X(n27335) );
  nand_x1_sg U55752 ( .A(\filter_0/reg_w_2[12] ), .B(n32867), .X(n27336) );
  nand_x1_sg U55753 ( .A(n30925), .B(reg_www_2[11]), .X(n27333) );
  nand_x1_sg U55754 ( .A(\filter_0/reg_w_2[11] ), .B(n32801), .X(n27334) );
  nand_x1_sg U55755 ( .A(n34607), .B(reg_www_2[10]), .X(n27331) );
  nand_x1_sg U55756 ( .A(\filter_0/reg_w_2[10] ), .B(n32880), .X(n27332) );
  nand_x1_sg U55757 ( .A(n31520), .B(reg_www_0[5]), .X(n27241) );
  nand_x1_sg U55758 ( .A(\filter_0/reg_w_0[5] ), .B(n35075), .X(n27242) );
  nand_x1_sg U55759 ( .A(n31520), .B(reg_www_0[4]), .X(n27239) );
  nand_x1_sg U55760 ( .A(\filter_0/reg_w_0[4] ), .B(n32436), .X(n27240) );
  nand_x1_sg U55761 ( .A(n33923), .B(reg_www_0[3]), .X(n27237) );
  nand_x1_sg U55762 ( .A(\filter_0/reg_w_0[3] ), .B(n32481), .X(n27238) );
  nand_x1_sg U55763 ( .A(n34603), .B(reg_www_0[2]), .X(n27235) );
  nand_x1_sg U55764 ( .A(\filter_0/reg_w_0[2] ), .B(n32433), .X(n27236) );
  nand_x1_sg U55765 ( .A(n32270), .B(reg_www_0[1]), .X(n27233) );
  nand_x1_sg U55766 ( .A(\filter_0/reg_w_0[1] ), .B(n30744), .X(n27234) );
  nand_x1_sg U55767 ( .A(n31090), .B(reg_www_0[0]), .X(n27231) );
  nand_x1_sg U55768 ( .A(\filter_0/reg_w_0[0] ), .B(n31292), .X(n27232) );
  nand_x1_sg U55769 ( .A(n32276), .B(reg_iii_15[19]), .X(n27229) );
  nand_x1_sg U55770 ( .A(\filter_0/reg_i_15[19] ), .B(n34620), .X(n27230) );
  nand_x1_sg U55771 ( .A(n33894), .B(reg_iii_15[18]), .X(n27227) );
  nand_x1_sg U55772 ( .A(\filter_0/reg_i_15[18] ), .B(n30765), .X(n27228) );
  nand_x1_sg U55773 ( .A(n35264), .B(reg_iii_15[17]), .X(n27225) );
  nand_x1_sg U55774 ( .A(\filter_0/reg_i_15[17] ), .B(n32860), .X(n27226) );
  nand_x1_sg U55775 ( .A(n34029), .B(reg_iii_15[16]), .X(n27223) );
  nand_x1_sg U55776 ( .A(\filter_0/reg_i_15[16] ), .B(n32821), .X(n27224) );
  nand_x1_sg U55777 ( .A(n34885), .B(reg_iii_15[15]), .X(n27221) );
  nand_x1_sg U55778 ( .A(\filter_0/reg_i_15[15] ), .B(n32472), .X(n27222) );
  nand_x1_sg U55779 ( .A(n31079), .B(reg_iii_15[14]), .X(n27219) );
  nand_x1_sg U55780 ( .A(\filter_0/reg_i_15[14] ), .B(n32488), .X(n27220) );
  nand_x1_sg U55781 ( .A(n32267), .B(reg_iii_14[14]), .X(n27179) );
  nand_x1_sg U55782 ( .A(\filter_0/reg_i_14[14] ), .B(n32439), .X(n27180) );
  nand_x1_sg U55783 ( .A(n31532), .B(reg_iii_14[13]), .X(n27177) );
  nand_x1_sg U55784 ( .A(\filter_0/reg_i_14[13] ), .B(n30762), .X(n27178) );
  nand_x1_sg U55785 ( .A(n30210), .B(reg_iii_14[12]), .X(n27175) );
  nand_x1_sg U55786 ( .A(\filter_0/reg_i_14[12] ), .B(n32475), .X(n27176) );
  nand_x1_sg U55787 ( .A(n34038), .B(reg_iii_14[11]), .X(n27173) );
  nand_x1_sg U55788 ( .A(\filter_0/reg_i_14[11] ), .B(n32879), .X(n27174) );
  nand_x1_sg U55789 ( .A(n34023), .B(reg_iii_14[10]), .X(n27171) );
  nand_x1_sg U55790 ( .A(\filter_0/reg_i_14[10] ), .B(n35073), .X(n27172) );
  nand_x1_sg U55791 ( .A(n31522), .B(reg_iii_14[9]), .X(n27169) );
  nand_x1_sg U55792 ( .A(\filter_0/reg_i_14[9] ), .B(n32862), .X(n27170) );
  nand_x1_sg U55793 ( .A(n31683), .B(reg_iii_14[8]), .X(n27167) );
  nand_x1_sg U55794 ( .A(\filter_0/reg_i_14[8] ), .B(n31916), .X(n27168) );
  nand_x1_sg U55795 ( .A(n34913), .B(reg_iii_11[17]), .X(n27065) );
  nand_x1_sg U55796 ( .A(\filter_0/reg_i_11[17] ), .B(n32805), .X(n27066) );
  nand_x1_sg U55797 ( .A(n34029), .B(reg_iii_11[16]), .X(n27063) );
  nand_x1_sg U55798 ( .A(\filter_0/reg_i_11[16] ), .B(n32467), .X(n27064) );
  nand_x1_sg U55799 ( .A(n35466), .B(reg_iii_11[15]), .X(n27061) );
  nand_x1_sg U55800 ( .A(\filter_0/reg_i_11[15] ), .B(n31921), .X(n27062) );
  nand_x1_sg U55801 ( .A(n35264), .B(reg_iii_11[14]), .X(n27059) );
  nand_x1_sg U55802 ( .A(\filter_0/reg_i_11[14] ), .B(n32488), .X(n27060) );
  nand_x1_sg U55803 ( .A(n34034), .B(reg_iii_11[13]), .X(n27057) );
  nand_x1_sg U55804 ( .A(\filter_0/reg_i_11[13] ), .B(n32782), .X(n27058) );
  nand_x1_sg U55805 ( .A(n30209), .B(reg_iii_11[12]), .X(n27055) );
  nand_x1_sg U55806 ( .A(\filter_0/reg_i_11[12] ), .B(n35069), .X(n27056) );
  nand_x1_sg U55807 ( .A(n32264), .B(reg_iii_11[4]), .X(n27039) );
  nand_x1_sg U55808 ( .A(\filter_0/reg_i_11[4] ), .B(n34673), .X(n27040) );
  nand_x1_sg U55809 ( .A(n31069), .B(reg_iii_11[3]), .X(n27037) );
  nand_x1_sg U55810 ( .A(\filter_0/reg_i_11[3] ), .B(n34628), .X(n27038) );
  nand_x1_sg U55811 ( .A(n34606), .B(reg_iii_11[2]), .X(n27035) );
  nand_x1_sg U55812 ( .A(\filter_0/reg_i_11[2] ), .B(n34690), .X(n27036) );
  nand_x1_sg U55813 ( .A(n34040), .B(reg_iii_11[1]), .X(n27033) );
  nand_x1_sg U55814 ( .A(\filter_0/reg_i_11[1] ), .B(n31911), .X(n27034) );
  nand_x1_sg U55815 ( .A(n34017), .B(reg_iii_11[0]), .X(n27031) );
  nand_x1_sg U55816 ( .A(\filter_0/reg_i_11[0] ), .B(n34641), .X(n27032) );
  nand_x1_sg U55817 ( .A(n31680), .B(reg_iii_10[19]), .X(n27029) );
  nand_x1_sg U55818 ( .A(\filter_0/reg_i_10[19] ), .B(n32486), .X(n27030) );
  nand_x1_sg U55819 ( .A(n33903), .B(reg_iii_10[18]), .X(n27027) );
  nand_x1_sg U55820 ( .A(\filter_0/reg_i_10[18] ), .B(n32826), .X(n27028) );
  nand_x1_sg U55821 ( .A(n30931), .B(reg_iii_10[17]), .X(n27025) );
  nand_x1_sg U55822 ( .A(\filter_0/reg_i_10[17] ), .B(n32809), .X(n27026) );
  nand_x1_sg U55823 ( .A(n33902), .B(reg_iii_10[16]), .X(n27023) );
  nand_x1_sg U55824 ( .A(\filter_0/reg_i_10[16] ), .B(n34643), .X(n27024) );
  nand_x1_sg U55825 ( .A(n35264), .B(reg_iii_10[15]), .X(n27021) );
  nand_x1_sg U55826 ( .A(\filter_0/reg_i_10[15] ), .B(n32780), .X(n27022) );
  nand_x1_sg U55827 ( .A(n34014), .B(reg_iii_10[14]), .X(n27019) );
  nand_x1_sg U55828 ( .A(\filter_0/reg_i_10[14] ), .B(n32476), .X(n27020) );
  nand_x1_sg U55829 ( .A(n31084), .B(reg_iii_10[13]), .X(n27017) );
  nand_x1_sg U55830 ( .A(\filter_0/reg_i_10[13] ), .B(n35068), .X(n27018) );
  nand_x1_sg U55831 ( .A(n34014), .B(reg_iii_10[12]), .X(n27015) );
  nand_x1_sg U55832 ( .A(\filter_0/reg_i_10[12] ), .B(n34628), .X(n27016) );
  nand_x1_sg U55833 ( .A(n31075), .B(reg_iii_10[11]), .X(n27013) );
  nand_x1_sg U55834 ( .A(\filter_0/reg_i_10[11] ), .B(n34680), .X(n27014) );
  nand_x1_sg U55835 ( .A(n34909), .B(reg_iii_10[10]), .X(n27011) );
  nand_x1_sg U55836 ( .A(\filter_0/reg_i_10[10] ), .B(n32470), .X(n27012) );
  nand_x1_sg U55837 ( .A(n31523), .B(reg_iii_10[9]), .X(n27009) );
  nand_x1_sg U55838 ( .A(\filter_0/reg_i_10[9] ), .B(n30736), .X(n27010) );
  nand_x1_sg U55839 ( .A(n30210), .B(reg_iii_10[8]), .X(n27007) );
  nand_x1_sg U55840 ( .A(\filter_0/reg_i_10[8] ), .B(n30250), .X(n27008) );
  nand_x1_sg U55841 ( .A(n33920), .B(reg_iii_10[7]), .X(n27005) );
  nand_x1_sg U55842 ( .A(\filter_0/reg_i_10[7] ), .B(n31922), .X(n27006) );
  nand_x1_sg U55843 ( .A(n31080), .B(reg_iii_10[6]), .X(n27003) );
  nand_x1_sg U55844 ( .A(\filter_0/reg_i_10[6] ), .B(n32437), .X(n27004) );
  nand_x1_sg U55845 ( .A(n34891), .B(reg_iii_9[7]), .X(n26965) );
  nand_x1_sg U55846 ( .A(\filter_0/reg_i_9[7] ), .B(n32870), .X(n26966) );
  nand_x1_sg U55847 ( .A(n34038), .B(reg_iii_9[6]), .X(n26963) );
  nand_x1_sg U55848 ( .A(\filter_0/reg_i_9[6] ), .B(n32860), .X(n26964) );
  nand_x1_sg U55849 ( .A(n33897), .B(reg_iii_9[5]), .X(n26961) );
  nand_x1_sg U55850 ( .A(\filter_0/reg_i_9[5] ), .B(n35068), .X(n26962) );
  nand_x1_sg U55851 ( .A(n33921), .B(reg_iii_9[4]), .X(n26959) );
  nand_x1_sg U55852 ( .A(\filter_0/reg_i_9[4] ), .B(n32827), .X(n26960) );
  nand_x1_sg U55853 ( .A(n34033), .B(reg_iii_9[3]), .X(n26957) );
  nand_x1_sg U55854 ( .A(\filter_0/reg_i_9[3] ), .B(n30745), .X(n26958) );
  nand_x1_sg U55855 ( .A(n31517), .B(reg_iii_9[2]), .X(n26955) );
  nand_x1_sg U55856 ( .A(\filter_0/reg_i_9[2] ), .B(n30772), .X(n26956) );
  nand_x1_sg U55857 ( .A(n32266), .B(reg_iii_9[1]), .X(n26953) );
  nand_x1_sg U55858 ( .A(\filter_0/reg_i_9[1] ), .B(n34636), .X(n26954) );
  nand_x1_sg U55859 ( .A(n34886), .B(reg_iii_9[0]), .X(n26951) );
  nand_x1_sg U55860 ( .A(\filter_0/reg_i_9[0] ), .B(n32869), .X(n26952) );
  nand_x1_sg U55861 ( .A(n31681), .B(reg_iii_8[19]), .X(n26949) );
  nand_x1_sg U55862 ( .A(\filter_0/reg_i_8[19] ), .B(n32479), .X(n26950) );
  nand_x1_sg U55863 ( .A(n33920), .B(reg_iii_8[18]), .X(n26947) );
  nand_x1_sg U55864 ( .A(\filter_0/reg_i_8[18] ), .B(n32859), .X(n26948) );
  nand_x1_sg U55865 ( .A(n35412), .B(reg_iii_8[17]), .X(n26945) );
  nand_x1_sg U55866 ( .A(\filter_0/reg_i_8[17] ), .B(n31918), .X(n26946) );
  nand_x1_sg U55867 ( .A(n32272), .B(reg_iii_8[16]), .X(n26943) );
  nand_x1_sg U55868 ( .A(\filter_0/reg_i_8[16] ), .B(n32780), .X(n26944) );
  nand_x1_sg U55869 ( .A(n30629), .B(reg_iii_8[15]), .X(n26941) );
  nand_x1_sg U55870 ( .A(\filter_0/reg_i_8[15] ), .B(n34673), .X(n26942) );
  nand_x1_sg U55871 ( .A(n31074), .B(reg_iii_7[2]), .X(n26875) );
  nand_x1_sg U55872 ( .A(\filter_0/reg_i_7[2] ), .B(n32880), .X(n26876) );
  nand_x1_sg U55873 ( .A(n31090), .B(reg_iii_7[1]), .X(n26873) );
  nand_x1_sg U55874 ( .A(\filter_0/reg_i_7[1] ), .B(n34688), .X(n26874) );
  nand_x1_sg U55875 ( .A(n32223), .B(reg_iii_7[0]), .X(n26871) );
  nand_x1_sg U55876 ( .A(\filter_0/reg_i_7[0] ), .B(n30160), .X(n26872) );
  nand_x1_sg U55877 ( .A(n33907), .B(reg_iii_6[19]), .X(n26869) );
  nand_x1_sg U55878 ( .A(\filter_0/reg_i_6[19] ), .B(n32474), .X(n26870) );
  nand_x1_sg U55879 ( .A(n34608), .B(reg_iii_6[18]), .X(n26867) );
  nand_x1_sg U55880 ( .A(\filter_0/reg_i_6[18] ), .B(n32801), .X(n26868) );
  nand_x1_sg U55881 ( .A(n33935), .B(reg_iii_6[17]), .X(n26865) );
  nand_x1_sg U55882 ( .A(\filter_0/reg_i_6[17] ), .B(n30738), .X(n26866) );
  nand_x1_sg U55883 ( .A(n32267), .B(reg_iii_6[16]), .X(n26863) );
  nand_x1_sg U55884 ( .A(\filter_0/reg_i_6[16] ), .B(n32819), .X(n26864) );
  nand_x1_sg U55885 ( .A(n33925), .B(reg_iii_6[15]), .X(n26861) );
  nand_x1_sg U55886 ( .A(\filter_0/reg_i_6[15] ), .B(n30758), .X(n26862) );
  nand_x1_sg U55887 ( .A(n31687), .B(reg_iii_6[14]), .X(n26859) );
  nand_x1_sg U55888 ( .A(\filter_0/reg_i_6[14] ), .B(n32827), .X(n26860) );
  nand_x1_sg U55889 ( .A(n33929), .B(reg_iii_6[13]), .X(n26857) );
  nand_x1_sg U55890 ( .A(\filter_0/reg_i_6[13] ), .B(n34629), .X(n26858) );
  nand_x1_sg U55891 ( .A(n34904), .B(reg_iii_6[12]), .X(n26855) );
  nand_x1_sg U55892 ( .A(\filter_0/reg_i_6[12] ), .B(n34630), .X(n26856) );
  nand_x1_sg U55893 ( .A(n35265), .B(reg_iii_6[11]), .X(n26853) );
  nand_x1_sg U55894 ( .A(\filter_0/reg_i_6[11] ), .B(n34640), .X(n26854) );
  nand_x1_sg U55895 ( .A(n34018), .B(reg_iii_6[10]), .X(n26851) );
  nand_x1_sg U55896 ( .A(\filter_0/reg_i_6[10] ), .B(n30773), .X(n26852) );
  nand_x1_sg U55897 ( .A(n33939), .B(reg_iii_6[9]), .X(n26849) );
  nand_x1_sg U55898 ( .A(\filter_0/reg_i_6[9] ), .B(n30757), .X(n26850) );
  nand_x1_sg U55899 ( .A(n31069), .B(reg_iii_6[8]), .X(n26847) );
  nand_x1_sg U55900 ( .A(\filter_0/reg_i_6[8] ), .B(n34645), .X(n26848) );
  nand_x1_sg U55901 ( .A(n33939), .B(reg_iii_6[7]), .X(n26845) );
  nand_x1_sg U55902 ( .A(\filter_0/reg_i_6[7] ), .B(n34682), .X(n26846) );
  nand_x1_sg U55903 ( .A(n31516), .B(reg_iii_6[6]), .X(n26843) );
  nand_x1_sg U55904 ( .A(\filter_0/reg_i_6[6] ), .B(n32472), .X(n26844) );
  nand_x1_sg U55905 ( .A(n33924), .B(reg_iii_6[5]), .X(n26841) );
  nand_x1_sg U55906 ( .A(\filter_0/reg_i_6[5] ), .B(n30733), .X(n26842) );
  nand_x1_sg U55907 ( .A(n32271), .B(reg_iii_5[5]), .X(n26801) );
  nand_x1_sg U55908 ( .A(\filter_0/reg_i_5[5] ), .B(n32438), .X(n26802) );
  nand_x1_sg U55909 ( .A(n31531), .B(reg_iii_2[1]), .X(n26673) );
  nand_x1_sg U55910 ( .A(\filter_0/reg_i_2[1] ), .B(n31209), .X(n26674) );
  nand_x1_sg U55911 ( .A(n30386), .B(reg_iii_2[0]), .X(n26671) );
  nand_x1_sg U55912 ( .A(\filter_0/reg_i_2[0] ), .B(n34678), .X(n26672) );
  nand_x1_sg U55913 ( .A(n33929), .B(reg_iii_1[19]), .X(n26669) );
  nand_x1_sg U55914 ( .A(\filter_0/reg_i_1[19] ), .B(n35067), .X(n26670) );
  nand_x1_sg U55915 ( .A(n33907), .B(reg_iii_1[18]), .X(n26667) );
  nand_x1_sg U55916 ( .A(\filter_0/reg_i_1[18] ), .B(n32789), .X(n26668) );
  nand_x1_sg U55917 ( .A(n32259), .B(reg_iii_1[17]), .X(n26665) );
  nand_x1_sg U55918 ( .A(\filter_0/reg_i_1[17] ), .B(n30744), .X(n26666) );
  nand_x1_sg U55919 ( .A(n30256), .B(reg_iii_1[16]), .X(n26663) );
  nand_x1_sg U55920 ( .A(\filter_0/reg_i_1[16] ), .B(n30757), .X(n26664) );
  nand_x1_sg U55921 ( .A(n31530), .B(reg_iii_1[15]), .X(n26661) );
  nand_x1_sg U55922 ( .A(\filter_0/reg_i_1[15] ), .B(n32482), .X(n26662) );
  nand_x1_sg U55923 ( .A(n31684), .B(reg_iii_1[14]), .X(n26659) );
  nand_x1_sg U55924 ( .A(\filter_0/reg_i_1[14] ), .B(n32484), .X(n26660) );
  nand_x1_sg U55925 ( .A(n31682), .B(reg_iii_1[13]), .X(n26657) );
  nand_x1_sg U55926 ( .A(\filter_0/reg_i_1[13] ), .B(n31296), .X(n26658) );
  nand_x1_sg U55927 ( .A(n33930), .B(reg_iii_1[12]), .X(n26655) );
  nand_x1_sg U55928 ( .A(\filter_0/reg_i_1[12] ), .B(n32488), .X(n26656) );
  nand_x1_sg U55929 ( .A(n31080), .B(reg_iii_1[11]), .X(n26653) );
  nand_x1_sg U55930 ( .A(\filter_0/reg_i_1[11] ), .B(n34677), .X(n26654) );
  nand_x1_sg U55931 ( .A(n33893), .B(reg_iii_1[10]), .X(n26651) );
  nand_x1_sg U55932 ( .A(\filter_0/reg_i_1[10] ), .B(n31296), .X(n26652) );
  nand_x1_sg U55933 ( .A(n32273), .B(reg_iii_1[9]), .X(n26649) );
  nand_x1_sg U55934 ( .A(\filter_0/reg_i_1[9] ), .B(n32475), .X(n26650) );
  nand_x1_sg U55935 ( .A(n31688), .B(reg_iii_1[8]), .X(n26647) );
  nand_x1_sg U55936 ( .A(\filter_0/reg_i_1[8] ), .B(n34636), .X(n26648) );
  nand_x1_sg U55937 ( .A(n33909), .B(reg_iii_1[7]), .X(n26645) );
  nand_x1_sg U55938 ( .A(\filter_0/reg_i_1[7] ), .B(n30739), .X(n26646) );
  nand_x1_sg U55939 ( .A(n35159), .B(reg_iii_1[6]), .X(n26643) );
  nand_x1_sg U55940 ( .A(\filter_0/reg_i_1[6] ), .B(n32809), .X(n26644) );
  nand_x1_sg U55941 ( .A(n34033), .B(reg_iii_1[5]), .X(n26641) );
  nand_x1_sg U55942 ( .A(\filter_0/reg_i_1[5] ), .B(n32820), .X(n26642) );
  nand_x1_sg U55943 ( .A(n34018), .B(reg_iii_1[4]), .X(n26639) );
  nand_x1_sg U55944 ( .A(\filter_0/reg_i_1[4] ), .B(n35075), .X(n26640) );
  nand_x1_sg U55945 ( .A(n32260), .B(reg_iii_1[3]), .X(n26637) );
  nand_x1_sg U55946 ( .A(\filter_0/reg_i_1[3] ), .B(n34643), .X(n26638) );
  nand_x1_sg U55947 ( .A(n30209), .B(o_mask[29]), .X(n27929) );
  nand_x1_sg U55948 ( .A(\filter_0/reg_o_mask[29] ), .B(n32435), .X(n27930) );
  nand_x1_sg U55949 ( .A(n34890), .B(o_mask[26]), .X(n27923) );
  nand_x1_sg U55950 ( .A(\filter_0/reg_o_mask[26] ), .B(n31208), .X(n27924) );
  nand_x1_sg U55951 ( .A(n32255), .B(o_mask[23]), .X(n27917) );
  nand_x1_sg U55952 ( .A(\filter_0/reg_o_mask[23] ), .B(n32796), .X(n27918) );
  nand_x1_sg U55953 ( .A(n30025), .B(o_mask[20]), .X(n27911) );
  nand_x1_sg U55954 ( .A(\filter_0/reg_o_mask[20] ), .B(n32879), .X(n27912) );
  nand_x1_sg U55955 ( .A(n30027), .B(o_mask[17]), .X(n27905) );
  nand_x1_sg U55956 ( .A(\filter_0/reg_o_mask[17] ), .B(n31914), .X(n27906) );
  nand_x1_sg U55957 ( .A(n30028), .B(o_mask[14]), .X(n27899) );
  nand_x1_sg U55958 ( .A(\filter_0/reg_o_mask[14] ), .B(n32810), .X(n27900) );
  nand_x1_sg U55959 ( .A(n29702), .B(o_mask[31]), .X(n27933) );
  nand_x1_sg U55960 ( .A(\filter_0/reg_o_mask[31] ), .B(n32464), .X(n27934) );
  nand_x1_sg U55961 ( .A(n31525), .B(o_mask[30]), .X(n27931) );
  nand_x1_sg U55962 ( .A(\filter_0/reg_o_mask[30] ), .B(n32816), .X(n27932) );
  nand_x1_sg U55963 ( .A(n32278), .B(o_mask[28]), .X(n27927) );
  nand_x1_sg U55964 ( .A(\filter_0/reg_o_mask[28] ), .B(n32881), .X(n27928) );
  nand_x1_sg U55965 ( .A(n34024), .B(o_mask[27]), .X(n27925) );
  nand_x1_sg U55966 ( .A(\filter_0/reg_o_mask[27] ), .B(n32491), .X(n27926) );
  nand_x1_sg U55967 ( .A(n33919), .B(o_mask[25]), .X(n27921) );
  nand_x1_sg U55968 ( .A(\filter_0/reg_o_mask[25] ), .B(n32780), .X(n27922) );
  nand_x1_sg U55969 ( .A(n30210), .B(o_mask[24]), .X(n27919) );
  nand_x1_sg U55970 ( .A(\filter_0/reg_o_mask[24] ), .B(n32800), .X(n27920) );
  nand_x1_sg U55971 ( .A(n33899), .B(o_mask[22]), .X(n27915) );
  nand_x1_sg U55972 ( .A(\filter_0/reg_o_mask[22] ), .B(n30732), .X(n27916) );
  nand_x1_sg U55973 ( .A(n34885), .B(o_mask[21]), .X(n27913) );
  nand_x1_sg U55974 ( .A(\filter_0/reg_o_mask[21] ), .B(n32880), .X(n27914) );
  nand_x1_sg U55975 ( .A(n34040), .B(o_mask[19]), .X(n27909) );
  nand_x1_sg U55976 ( .A(\filter_0/reg_o_mask[19] ), .B(n32859), .X(n27910) );
  nand_x1_sg U55977 ( .A(n34016), .B(o_mask[18]), .X(n27907) );
  nand_x1_sg U55978 ( .A(\filter_0/reg_o_mask[18] ), .B(n32820), .X(n27908) );
  nand_x1_sg U55979 ( .A(n31527), .B(o_mask[16]), .X(n27903) );
  nand_x1_sg U55980 ( .A(\filter_0/reg_o_mask[16] ), .B(n32458), .X(n27904) );
  nand_x1_sg U55981 ( .A(n33918), .B(o_mask[15]), .X(n27901) );
  nand_x1_sg U55982 ( .A(\filter_0/reg_o_mask[15] ), .B(n32486), .X(n27902) );
  nor_x1_sg U55983 ( .A(n15312), .B(n15313), .X(n15310) );
  nor_x1_sg U55984 ( .A(\filter_0/reg_o_mask[10] ), .B(n32124), .X(n15313) );
  nor_x1_sg U55985 ( .A(\filter_0/reg_o_mask[8] ), .B(n32128), .X(n15312) );
  nand_x1_sg U55986 ( .A(n19602), .B(shifter_state[0]), .X(n19603) );
  nand_x1_sg U55987 ( .A(n19605), .B(n19606), .X(n19604) );
  nor_x1_sg U55988 ( .A(n19607), .B(n19602), .X(n19605) );
  nand_x1_sg U55989 ( .A(reg_ow_3[0]), .B(n33616), .X(n29062) );
  nand_x1_sg U55990 ( .A(reg_ow_3[1]), .B(n33616), .X(n29066) );
  nand_x1_sg U55991 ( .A(reg_ow_3[2]), .B(n33616), .X(n29068) );
  nand_x1_sg U55992 ( .A(reg_ow_3[3]), .B(n33615), .X(n29070) );
  nand_x1_sg U55993 ( .A(reg_ow_3[4]), .B(n33615), .X(n29072) );
  nand_x1_sg U55994 ( .A(reg_ow_3[5]), .B(n33616), .X(n29074) );
  nand_x1_sg U55995 ( .A(reg_ow_3[6]), .B(n33619), .X(n29076) );
  nand_x1_sg U55996 ( .A(n33465), .B(\filter_0/n8233 ), .X(n29077) );
  nand_x1_sg U55997 ( .A(reg_ow_3[7]), .B(n33620), .X(n29078) );
  nand_x1_sg U55998 ( .A(n33466), .B(\filter_0/n8232 ), .X(n29079) );
  nand_x1_sg U55999 ( .A(reg_ow_3[8]), .B(n33619), .X(n29080) );
  nand_x1_sg U56000 ( .A(n33465), .B(\filter_0/n8231 ), .X(n29081) );
  nand_x1_sg U56001 ( .A(reg_ow_3[9]), .B(n33615), .X(n29082) );
  nand_x1_sg U56002 ( .A(n33466), .B(\filter_0/n8230 ), .X(n29083) );
  nand_x1_sg U56003 ( .A(reg_ow_3[10]), .B(n33620), .X(n29084) );
  nand_x1_sg U56004 ( .A(n33467), .B(\filter_0/n8229 ), .X(n29085) );
  nand_x1_sg U56005 ( .A(reg_ow_3[11]), .B(n33621), .X(n29086) );
  nand_x1_sg U56006 ( .A(n33468), .B(\filter_0/n8228 ), .X(n29087) );
  nand_x1_sg U56007 ( .A(reg_ow_3[12]), .B(n33615), .X(n29088) );
  nand_x1_sg U56008 ( .A(n33468), .B(\filter_0/n8227 ), .X(n29089) );
  nand_x1_sg U56009 ( .A(reg_ow_3[13]), .B(n33621), .X(n29090) );
  nand_x1_sg U56010 ( .A(n33466), .B(\filter_0/n8226 ), .X(n29091) );
  nand_x1_sg U56011 ( .A(reg_ow_3[14]), .B(n33619), .X(n29092) );
  nand_x1_sg U56012 ( .A(n33467), .B(\filter_0/n8225 ), .X(n29093) );
  nand_x1_sg U56013 ( .A(reg_ow_3[15]), .B(n33621), .X(n29094) );
  nand_x1_sg U56014 ( .A(n29985), .B(\filter_0/n8224 ), .X(n29095) );
  nand_x1_sg U56015 ( .A(reg_ow_3[16]), .B(n33621), .X(n29096) );
  nand_x1_sg U56016 ( .A(n29985), .B(\filter_0/n8223 ), .X(n29097) );
  nand_x1_sg U56017 ( .A(reg_ow_3[17]), .B(n33620), .X(n29098) );
  nand_x1_sg U56018 ( .A(n33465), .B(\filter_0/n8222 ), .X(n29099) );
  nand_x1_sg U56019 ( .A(reg_ow_3[18]), .B(n33619), .X(n29100) );
  nand_x1_sg U56020 ( .A(n33465), .B(\filter_0/n8221 ), .X(n29101) );
  nand_x1_sg U56021 ( .A(reg_ow_3[19]), .B(n33620), .X(n29102) );
  nand_x1_sg U56022 ( .A(n33468), .B(\filter_0/n8220 ), .X(n29103) );
  nand_x1_sg U56023 ( .A(reg_ow_15[0]), .B(n33623), .X(n29275) );
  nand_x1_sg U56024 ( .A(reg_ow_15[1]), .B(n33627), .X(n29279) );
  nand_x1_sg U56025 ( .A(reg_ow_15[2]), .B(n33629), .X(n29281) );
  nand_x1_sg U56026 ( .A(reg_ow_15[3]), .B(n33627), .X(n29283) );
  nand_x1_sg U56027 ( .A(reg_ow_15[4]), .B(n33623), .X(n29285) );
  nand_x1_sg U56028 ( .A(reg_ow_15[5]), .B(n33624), .X(n29287) );
  nand_x1_sg U56029 ( .A(reg_ow_15[6]), .B(n33628), .X(n29289) );
  nand_x1_sg U56030 ( .A(n33407), .B(\filter_0/n8013 ), .X(n29290) );
  nand_x1_sg U56031 ( .A(reg_ow_15[7]), .B(n33624), .X(n29291) );
  nand_x1_sg U56032 ( .A(n33405), .B(\filter_0/n8012 ), .X(n29292) );
  nand_x1_sg U56033 ( .A(reg_ow_15[8]), .B(n33623), .X(n29293) );
  nand_x1_sg U56034 ( .A(n33405), .B(\filter_0/n8011 ), .X(n29294) );
  nand_x1_sg U56035 ( .A(reg_ow_15[9]), .B(n33624), .X(n29295) );
  nand_x1_sg U56036 ( .A(n29961), .B(\filter_0/n8010 ), .X(n29296) );
  nand_x1_sg U56037 ( .A(reg_ow_15[10]), .B(n33628), .X(n29297) );
  nand_x1_sg U56038 ( .A(n33406), .B(\filter_0/n8009 ), .X(n29298) );
  nand_x1_sg U56039 ( .A(reg_ow_15[11]), .B(n33627), .X(n29299) );
  nand_x1_sg U56040 ( .A(n29961), .B(\filter_0/n8008 ), .X(n29300) );
  nand_x1_sg U56041 ( .A(reg_ow_15[12]), .B(n33624), .X(n29301) );
  nand_x1_sg U56042 ( .A(n29961), .B(\filter_0/n8007 ), .X(n29302) );
  nand_x1_sg U56043 ( .A(reg_ow_15[13]), .B(n33627), .X(n29303) );
  nand_x1_sg U56044 ( .A(n33407), .B(\filter_0/n8006 ), .X(n29304) );
  nand_x1_sg U56045 ( .A(reg_ow_15[14]), .B(n33628), .X(n29305) );
  nand_x1_sg U56046 ( .A(n33406), .B(\filter_0/n8005 ), .X(n29306) );
  nand_x1_sg U56047 ( .A(reg_ow_15[15]), .B(n33628), .X(n29307) );
  nand_x1_sg U56048 ( .A(n33405), .B(\filter_0/n8004 ), .X(n29308) );
  nand_x1_sg U56049 ( .A(reg_ow_15[16]), .B(n33629), .X(n29309) );
  nand_x1_sg U56050 ( .A(n33407), .B(\filter_0/n8003 ), .X(n29310) );
  nand_x1_sg U56051 ( .A(reg_ow_15[17]), .B(n33629), .X(n29311) );
  nand_x1_sg U56052 ( .A(n33407), .B(\filter_0/n8002 ), .X(n29312) );
  nand_x1_sg U56053 ( .A(reg_ow_15[18]), .B(n33623), .X(n29313) );
  nand_x1_sg U56054 ( .A(n33408), .B(\filter_0/n8001 ), .X(n29314) );
  nand_x1_sg U56055 ( .A(reg_ow_15[19]), .B(n33629), .X(n29315) );
  nand_x1_sg U56056 ( .A(n33408), .B(\filter_0/n8000 ), .X(n29316) );
  nor_x1_sg U56057 ( .A(\filter_0/reg_o_mask[24] ), .B(n32126), .X(n15346) );
  nor_x1_sg U56058 ( .A(n15346), .B(n15347), .X(n15344) );
  nor_x1_sg U56059 ( .A(n32130), .B(\filter_0/reg_o_mask[28] ), .X(n15345) );
  nor_x1_sg U56060 ( .A(n32002), .B(n15297), .X(n15295) );
  nor_x1_sg U56061 ( .A(\filter_0/reg_o_mask[0] ), .B(n32126), .X(n15297) );
  nand_x1_sg U56062 ( .A(n29533), .B(n31878), .X(n29532) );
  nor_x1_sg U56063 ( .A(n31658), .B(n34063), .X(n29533) );
  nand_x1_sg U56064 ( .A(reg_ow_2[0]), .B(n33516), .X(n29019) );
  nand_x1_sg U56065 ( .A(reg_ow_2[1]), .B(n33515), .X(n29023) );
  nand_x1_sg U56066 ( .A(reg_ow_2[2]), .B(n33519), .X(n29025) );
  nand_x1_sg U56067 ( .A(reg_ow_2[3]), .B(n33520), .X(n29027) );
  nand_x1_sg U56068 ( .A(reg_ow_2[4]), .B(n33520), .X(n29029) );
  nand_x1_sg U56069 ( .A(reg_ow_2[5]), .B(n33516), .X(n29031) );
  nand_x1_sg U56070 ( .A(reg_ow_2[6]), .B(n33515), .X(n29033) );
  nand_x1_sg U56071 ( .A(n33317), .B(\filter_0/n8213 ), .X(n29034) );
  nand_x1_sg U56072 ( .A(reg_ow_2[7]), .B(n33516), .X(n29035) );
  nand_x1_sg U56073 ( .A(n33317), .B(\filter_0/n8212 ), .X(n29036) );
  nand_x1_sg U56074 ( .A(reg_ow_2[8]), .B(n33521), .X(n29037) );
  nand_x1_sg U56075 ( .A(n33318), .B(\filter_0/n8211 ), .X(n29038) );
  nand_x1_sg U56076 ( .A(reg_ow_2[9]), .B(n33516), .X(n29039) );
  nand_x1_sg U56077 ( .A(n33315), .B(\filter_0/n8210 ), .X(n29040) );
  nand_x1_sg U56078 ( .A(reg_ow_2[10]), .B(n33519), .X(n29041) );
  nand_x1_sg U56079 ( .A(n33317), .B(\filter_0/n8209 ), .X(n29042) );
  nand_x1_sg U56080 ( .A(reg_ow_2[11]), .B(n33521), .X(n29043) );
  nand_x1_sg U56081 ( .A(n33317), .B(\filter_0/n8208 ), .X(n29044) );
  nand_x1_sg U56082 ( .A(reg_ow_2[12]), .B(n33515), .X(n29045) );
  nand_x1_sg U56083 ( .A(n33316), .B(\filter_0/n8207 ), .X(n29046) );
  nand_x1_sg U56084 ( .A(reg_ow_2[13]), .B(n33520), .X(n29047) );
  nand_x1_sg U56085 ( .A(n29925), .B(\filter_0/n8206 ), .X(n29048) );
  nand_x1_sg U56086 ( .A(reg_ow_2[14]), .B(n33520), .X(n29049) );
  nand_x1_sg U56087 ( .A(n33318), .B(\filter_0/n8205 ), .X(n29050) );
  nand_x1_sg U56088 ( .A(reg_ow_2[15]), .B(n33521), .X(n29051) );
  nand_x1_sg U56089 ( .A(n29925), .B(\filter_0/n8204 ), .X(n29052) );
  nand_x1_sg U56090 ( .A(reg_ow_2[16]), .B(n33519), .X(n29053) );
  nand_x1_sg U56091 ( .A(n33316), .B(\filter_0/n8203 ), .X(n29054) );
  nand_x1_sg U56092 ( .A(reg_ow_2[17]), .B(n33519), .X(n29055) );
  nand_x1_sg U56093 ( .A(n33316), .B(\filter_0/n8202 ), .X(n29056) );
  nand_x1_sg U56094 ( .A(reg_ow_2[18]), .B(n33515), .X(n29057) );
  nand_x1_sg U56095 ( .A(n33315), .B(\filter_0/n8201 ), .X(n29058) );
  nand_x1_sg U56096 ( .A(reg_ow_2[19]), .B(n33521), .X(n29059) );
  nand_x1_sg U56097 ( .A(n33318), .B(\filter_0/n8200 ), .X(n29060) );
  nand_x1_sg U56098 ( .A(reg_ow_6[0]), .B(n33660), .X(n29191) );
  nand_x1_sg U56099 ( .A(reg_ow_6[1]), .B(n33656), .X(n29195) );
  nand_x1_sg U56100 ( .A(reg_ow_6[2]), .B(n33656), .X(n29197) );
  nand_x1_sg U56101 ( .A(reg_ow_6[3]), .B(n33660), .X(n29199) );
  nand_x1_sg U56102 ( .A(reg_ow_6[4]), .B(n33655), .X(n29201) );
  nand_x1_sg U56103 ( .A(reg_ow_6[5]), .B(n33659), .X(n29203) );
  nand_x1_sg U56104 ( .A(reg_ow_6[6]), .B(n33660), .X(n29205) );
  nand_x1_sg U56105 ( .A(n29973), .B(\filter_0/n8133 ), .X(n29206) );
  nand_x1_sg U56106 ( .A(reg_ow_6[7]), .B(n33659), .X(n29207) );
  nand_x1_sg U56107 ( .A(n33437), .B(\filter_0/n8132 ), .X(n29208) );
  nand_x1_sg U56108 ( .A(reg_ow_6[8]), .B(n33660), .X(n29209) );
  nand_x1_sg U56109 ( .A(n33436), .B(\filter_0/n8131 ), .X(n29210) );
  nand_x1_sg U56110 ( .A(reg_ow_6[9]), .B(n33661), .X(n29211) );
  nand_x1_sg U56111 ( .A(n33438), .B(\filter_0/n8130 ), .X(n29212) );
  nand_x1_sg U56112 ( .A(reg_ow_6[10]), .B(n33659), .X(n29213) );
  nand_x1_sg U56113 ( .A(n33435), .B(\filter_0/n8129 ), .X(n29214) );
  nand_x1_sg U56114 ( .A(reg_ow_6[11]), .B(n33655), .X(n29215) );
  nand_x1_sg U56115 ( .A(n33435), .B(\filter_0/n8128 ), .X(n29216) );
  nand_x1_sg U56116 ( .A(reg_ow_6[12]), .B(n33661), .X(n29217) );
  nand_x1_sg U56117 ( .A(n33438), .B(\filter_0/n8127 ), .X(n29218) );
  nand_x1_sg U56118 ( .A(reg_ow_6[13]), .B(n33655), .X(n29219) );
  nand_x1_sg U56119 ( .A(n33437), .B(\filter_0/n8126 ), .X(n29220) );
  nand_x1_sg U56120 ( .A(reg_ow_6[14]), .B(n33659), .X(n29221) );
  nand_x1_sg U56121 ( .A(n29973), .B(\filter_0/n8125 ), .X(n29222) );
  nand_x1_sg U56122 ( .A(reg_ow_6[15]), .B(n33661), .X(n29223) );
  nand_x1_sg U56123 ( .A(n33438), .B(\filter_0/n8124 ), .X(n29224) );
  nand_x1_sg U56124 ( .A(reg_ow_6[16]), .B(n33656), .X(n29225) );
  nand_x1_sg U56125 ( .A(n33436), .B(\filter_0/n8123 ), .X(n29226) );
  nand_x1_sg U56126 ( .A(reg_ow_6[17]), .B(n33656), .X(n29227) );
  nand_x1_sg U56127 ( .A(n33438), .B(\filter_0/n8122 ), .X(n29228) );
  nand_x1_sg U56128 ( .A(reg_ow_6[18]), .B(n33655), .X(n29229) );
  nand_x1_sg U56129 ( .A(n29973), .B(\filter_0/n8121 ), .X(n29230) );
  nand_x1_sg U56130 ( .A(reg_ow_6[19]), .B(n33661), .X(n29231) );
  nand_x1_sg U56131 ( .A(n33435), .B(\filter_0/n8120 ), .X(n29232) );
  nand_x1_sg U56132 ( .A(reg_ow_14[0]), .B(n33676), .X(n29318) );
  nand_x1_sg U56133 ( .A(reg_ow_14[1]), .B(n33677), .X(n29322) );
  nand_x1_sg U56134 ( .A(reg_ow_14[2]), .B(n33675), .X(n29324) );
  nand_x1_sg U56135 ( .A(reg_ow_14[3]), .B(n33672), .X(n29326) );
  nand_x1_sg U56136 ( .A(reg_ow_14[4]), .B(n33671), .X(n29328) );
  nand_x1_sg U56137 ( .A(reg_ow_14[5]), .B(n33672), .X(n29330) );
  nand_x1_sg U56138 ( .A(reg_ow_14[6]), .B(n33676), .X(n29332) );
  nand_x1_sg U56139 ( .A(n33312), .B(\filter_0/n8073 ), .X(n29333) );
  nand_x1_sg U56140 ( .A(reg_ow_14[7]), .B(n33677), .X(n29334) );
  nand_x1_sg U56141 ( .A(n29923), .B(\filter_0/n8072 ), .X(n29335) );
  nand_x1_sg U56142 ( .A(reg_ow_14[8]), .B(n33672), .X(n29336) );
  nand_x1_sg U56143 ( .A(n33312), .B(\filter_0/n8071 ), .X(n29337) );
  nand_x1_sg U56144 ( .A(reg_ow_14[9]), .B(n33672), .X(n29338) );
  nand_x1_sg U56145 ( .A(n33312), .B(\filter_0/n8070 ), .X(n29339) );
  nand_x1_sg U56146 ( .A(reg_ow_14[10]), .B(n33671), .X(n29340) );
  nand_x1_sg U56147 ( .A(n33311), .B(\filter_0/n8069 ), .X(n29341) );
  nand_x1_sg U56148 ( .A(reg_ow_14[11]), .B(n33675), .X(n29342) );
  nand_x1_sg U56149 ( .A(n33313), .B(\filter_0/n8068 ), .X(n29343) );
  nand_x1_sg U56150 ( .A(reg_ow_14[12]), .B(n33677), .X(n29344) );
  nand_x1_sg U56151 ( .A(n33311), .B(\filter_0/n8067 ), .X(n29345) );
  nand_x1_sg U56152 ( .A(reg_ow_14[13]), .B(n33675), .X(n29346) );
  nand_x1_sg U56153 ( .A(n33310), .B(\filter_0/n8066 ), .X(n29347) );
  nand_x1_sg U56154 ( .A(reg_ow_14[14]), .B(n33671), .X(n29348) );
  nand_x1_sg U56155 ( .A(n33312), .B(\filter_0/n8065 ), .X(n29349) );
  nand_x1_sg U56156 ( .A(reg_ow_14[15]), .B(n33676), .X(n29350) );
  nand_x1_sg U56157 ( .A(n33310), .B(\filter_0/n8064 ), .X(n29351) );
  nand_x1_sg U56158 ( .A(reg_ow_14[16]), .B(n33676), .X(n29352) );
  nand_x1_sg U56159 ( .A(n33313), .B(\filter_0/n8063 ), .X(n29353) );
  nand_x1_sg U56160 ( .A(reg_ow_14[17]), .B(n33671), .X(n29354) );
  nand_x1_sg U56161 ( .A(n29923), .B(\filter_0/n8062 ), .X(n29355) );
  nand_x1_sg U56162 ( .A(reg_ow_14[18]), .B(n33677), .X(n29356) );
  nand_x1_sg U56163 ( .A(n33310), .B(\filter_0/n8061 ), .X(n29357) );
  nand_x1_sg U56164 ( .A(reg_ow_14[19]), .B(n33675), .X(n29358) );
  nand_x1_sg U56165 ( .A(n33313), .B(\filter_0/n8060 ), .X(n29359) );
  nand_x1_sg U56166 ( .A(n31205), .B(n19601), .X(\shifter_0/n10884 ) );
  nand_x1_sg U56167 ( .A(n19602), .B(shifter_state[1]), .X(n19601) );
  nand_x1_sg U56168 ( .A(reg_ow_7[0]), .B(n33612), .X(n29233) );
  nand_x1_sg U56169 ( .A(reg_ow_7[2]), .B(n33611), .X(n29239) );
  nand_x1_sg U56170 ( .A(reg_ow_7[4]), .B(n33613), .X(n29243) );
  nand_x1_sg U56171 ( .A(reg_ow_7[6]), .B(n33607), .X(n29247) );
  nand_x1_sg U56172 ( .A(n33396), .B(\filter_0/n8153 ), .X(n29248) );
  nand_x1_sg U56173 ( .A(reg_ow_7[8]), .B(n33611), .X(n29251) );
  nand_x1_sg U56174 ( .A(n33398), .B(\filter_0/n8151 ), .X(n29252) );
  nand_x1_sg U56175 ( .A(reg_ow_7[10]), .B(n33613), .X(n29255) );
  nand_x1_sg U56176 ( .A(n33396), .B(\filter_0/n8149 ), .X(n29256) );
  nand_x1_sg U56177 ( .A(reg_ow_7[12]), .B(n33612), .X(n29259) );
  nand_x1_sg U56178 ( .A(n29957), .B(\filter_0/n8147 ), .X(n29260) );
  nand_x1_sg U56179 ( .A(reg_ow_7[14]), .B(n33613), .X(n29263) );
  nand_x1_sg U56180 ( .A(n33395), .B(\filter_0/n8145 ), .X(n29264) );
  nand_x1_sg U56181 ( .A(reg_ow_7[16]), .B(n33612), .X(n29267) );
  nand_x1_sg U56182 ( .A(n33397), .B(\filter_0/n8143 ), .X(n29268) );
  nand_x1_sg U56183 ( .A(reg_ow_7[18]), .B(n33611), .X(n29271) );
  nand_x1_sg U56184 ( .A(n33396), .B(\filter_0/n8141 ), .X(n29272) );
  nand_x1_sg U56185 ( .A(n29577), .B(n31658), .X(n29576) );
  nor_x1_sg U56186 ( .A(n31879), .B(n34062), .X(n29577) );
  nor_x1_sg U56187 ( .A(n35273), .B(n35154), .X(n15356) );
  nor_x1_sg U56188 ( .A(\filter_0/reg_o_mask[26] ), .B(n32122), .X(n15347) );
  nor_x1_sg U56189 ( .A(\filter_0/reg_o_mask[16] ), .B(n32127), .X(n15330) );
  nor_x1_sg U56190 ( .A(n35306), .B(n15352), .X(n15351) );
  nor_x1_sg U56191 ( .A(n32504), .B(\filter_0/reg_o_mask[31] ), .X(n15352) );
  nand_x1_sg U56192 ( .A(reg_ow_11[0]), .B(n33604), .X(n29445) );
  nand_x1_sg U56193 ( .A(reg_ow_11[2]), .B(n33605), .X(n29451) );
  nand_x1_sg U56194 ( .A(reg_ow_11[4]), .B(n33600), .X(n29455) );
  nand_x1_sg U56195 ( .A(reg_ow_11[6]), .B(n33599), .X(n29459) );
  nand_x1_sg U56196 ( .A(n33401), .B(\filter_0/n7993 ), .X(n29460) );
  nand_x1_sg U56197 ( .A(reg_ow_11[8]), .B(n33605), .X(n29463) );
  nand_x1_sg U56198 ( .A(n33402), .B(\filter_0/n7991 ), .X(n29464) );
  nand_x1_sg U56199 ( .A(reg_ow_11[10]), .B(n33600), .X(n29467) );
  nand_x1_sg U56200 ( .A(n33400), .B(\filter_0/n7989 ), .X(n29468) );
  nand_x1_sg U56201 ( .A(reg_ow_11[12]), .B(n33603), .X(n29471) );
  nand_x1_sg U56202 ( .A(n33401), .B(\filter_0/n7987 ), .X(n29472) );
  nand_x1_sg U56203 ( .A(reg_ow_11[14]), .B(n33605), .X(n29475) );
  nand_x1_sg U56204 ( .A(n33403), .B(\filter_0/n7985 ), .X(n29476) );
  nand_x1_sg U56205 ( .A(reg_ow_11[16]), .B(n33599), .X(n29479) );
  nand_x1_sg U56206 ( .A(n33401), .B(\filter_0/n7983 ), .X(n29480) );
  nand_x1_sg U56207 ( .A(reg_ow_11[18]), .B(n33605), .X(n29483) );
  nand_x1_sg U56208 ( .A(n33400), .B(\filter_0/n7981 ), .X(n29484) );
  nor_x1_sg U56209 ( .A(n32001), .B(n15330), .X(n15328) );
  nor_x1_sg U56210 ( .A(n32123), .B(\filter_0/reg_o_mask[18] ), .X(n15329) );
  nand_x1_sg U56211 ( .A(reg_ow_1[0]), .B(n33495), .X(n28976) );
  nand_x1_sg U56212 ( .A(reg_ow_1[1]), .B(n33497), .X(n28980) );
  nand_x1_sg U56213 ( .A(reg_ow_1[2]), .B(n33491), .X(n28982) );
  nand_x1_sg U56214 ( .A(reg_ow_1[3]), .B(n33497), .X(n28984) );
  nand_x1_sg U56215 ( .A(reg_ow_1[4]), .B(n33492), .X(n28986) );
  nand_x1_sg U56216 ( .A(reg_ow_1[5]), .B(n33491), .X(n28988) );
  nand_x1_sg U56217 ( .A(reg_ow_1[6]), .B(n33492), .X(n28990) );
  nand_x1_sg U56218 ( .A(n33305), .B(\filter_0/n8193 ), .X(n28991) );
  nand_x1_sg U56219 ( .A(reg_ow_1[7]), .B(n33495), .X(n28992) );
  nand_x1_sg U56220 ( .A(n33308), .B(\filter_0/n8192 ), .X(n28993) );
  nand_x1_sg U56221 ( .A(reg_ow_1[8]), .B(n33497), .X(n28994) );
  nand_x1_sg U56222 ( .A(n33306), .B(\filter_0/n8191 ), .X(n28995) );
  nand_x1_sg U56223 ( .A(reg_ow_1[9]), .B(n33496), .X(n28996) );
  nand_x1_sg U56224 ( .A(n29921), .B(\filter_0/n8190 ), .X(n28997) );
  nand_x1_sg U56225 ( .A(reg_ow_1[10]), .B(n33497), .X(n28998) );
  nand_x1_sg U56226 ( .A(n33306), .B(\filter_0/n8189 ), .X(n28999) );
  nand_x1_sg U56227 ( .A(reg_ow_1[11]), .B(n33491), .X(n29000) );
  nand_x1_sg U56228 ( .A(n33307), .B(\filter_0/n8188 ), .X(n29001) );
  nand_x1_sg U56229 ( .A(reg_ow_1[12]), .B(n33495), .X(n29002) );
  nand_x1_sg U56230 ( .A(n33308), .B(\filter_0/n8187 ), .X(n29003) );
  nand_x1_sg U56231 ( .A(reg_ow_1[13]), .B(n33496), .X(n29004) );
  nand_x1_sg U56232 ( .A(n33305), .B(\filter_0/n8186 ), .X(n29005) );
  nand_x1_sg U56233 ( .A(reg_ow_1[14]), .B(n33496), .X(n29006) );
  nand_x1_sg U56234 ( .A(n33308), .B(\filter_0/n8185 ), .X(n29007) );
  nand_x1_sg U56235 ( .A(reg_ow_1[15]), .B(n33496), .X(n29008) );
  nand_x1_sg U56236 ( .A(n29921), .B(\filter_0/n8184 ), .X(n29009) );
  nand_x1_sg U56237 ( .A(reg_ow_1[16]), .B(n33495), .X(n29010) );
  nand_x1_sg U56238 ( .A(n33308), .B(\filter_0/n8183 ), .X(n29011) );
  nand_x1_sg U56239 ( .A(reg_ow_1[17]), .B(n33491), .X(n29012) );
  nand_x1_sg U56240 ( .A(n33307), .B(\filter_0/n8182 ), .X(n29013) );
  nand_x1_sg U56241 ( .A(reg_ow_1[18]), .B(n33492), .X(n29014) );
  nand_x1_sg U56242 ( .A(n33307), .B(\filter_0/n8181 ), .X(n29015) );
  nand_x1_sg U56243 ( .A(reg_ow_1[19]), .B(n33492), .X(n29016) );
  nand_x1_sg U56244 ( .A(n33305), .B(\filter_0/n8180 ), .X(n29017) );
  nand_x1_sg U56245 ( .A(reg_ow_5[0]), .B(n33511), .X(n29149) );
  nand_x1_sg U56246 ( .A(reg_ow_5[1]), .B(n33507), .X(n29153) );
  nand_x1_sg U56247 ( .A(reg_ow_5[2]), .B(n33513), .X(n29155) );
  nand_x1_sg U56248 ( .A(reg_ow_5[3]), .B(n33508), .X(n29157) );
  nand_x1_sg U56249 ( .A(reg_ow_5[4]), .B(n33511), .X(n29159) );
  nand_x1_sg U56250 ( .A(reg_ow_5[5]), .B(n33513), .X(n29161) );
  nand_x1_sg U56251 ( .A(reg_ow_5[6]), .B(n33507), .X(n29163) );
  nand_x1_sg U56252 ( .A(n33460), .B(\filter_0/n8113 ), .X(n29164) );
  nand_x1_sg U56253 ( .A(reg_ow_5[7]), .B(n33508), .X(n29165) );
  nand_x1_sg U56254 ( .A(n33462), .B(\filter_0/n8112 ), .X(n29166) );
  nand_x1_sg U56255 ( .A(reg_ow_5[8]), .B(n33507), .X(n29167) );
  nand_x1_sg U56256 ( .A(n33461), .B(\filter_0/n8111 ), .X(n29168) );
  nand_x1_sg U56257 ( .A(reg_ow_5[9]), .B(n33512), .X(n29169) );
  nand_x1_sg U56258 ( .A(n33462), .B(\filter_0/n8110 ), .X(n29170) );
  nand_x1_sg U56259 ( .A(reg_ow_5[10]), .B(n33512), .X(n29171) );
  nand_x1_sg U56260 ( .A(n29983), .B(\filter_0/n8109 ), .X(n29172) );
  nand_x1_sg U56261 ( .A(reg_ow_5[11]), .B(n33508), .X(n29173) );
  nand_x1_sg U56262 ( .A(n33463), .B(\filter_0/n8108 ), .X(n29174) );
  nand_x1_sg U56263 ( .A(reg_ow_5[12]), .B(n33511), .X(n29175) );
  nand_x1_sg U56264 ( .A(n33461), .B(\filter_0/n8107 ), .X(n29176) );
  nand_x1_sg U56265 ( .A(reg_ow_5[13]), .B(n33511), .X(n29177) );
  nand_x1_sg U56266 ( .A(n33460), .B(\filter_0/n8106 ), .X(n29178) );
  nand_x1_sg U56267 ( .A(reg_ow_5[14]), .B(n33512), .X(n29179) );
  nand_x1_sg U56268 ( .A(n33463), .B(\filter_0/n8105 ), .X(n29180) );
  nand_x1_sg U56269 ( .A(reg_ow_5[15]), .B(n33513), .X(n29181) );
  nand_x1_sg U56270 ( .A(n33463), .B(\filter_0/n8104 ), .X(n29182) );
  nand_x1_sg U56271 ( .A(reg_ow_5[16]), .B(n33513), .X(n29183) );
  nand_x1_sg U56272 ( .A(n33460), .B(\filter_0/n8103 ), .X(n29184) );
  nand_x1_sg U56273 ( .A(reg_ow_5[17]), .B(n33507), .X(n29185) );
  nand_x1_sg U56274 ( .A(n33462), .B(\filter_0/n8102 ), .X(n29186) );
  nand_x1_sg U56275 ( .A(reg_ow_5[18]), .B(n33508), .X(n29187) );
  nand_x1_sg U56276 ( .A(n33461), .B(\filter_0/n8101 ), .X(n29188) );
  nand_x1_sg U56277 ( .A(reg_ow_5[19]), .B(n33512), .X(n29189) );
  nand_x1_sg U56278 ( .A(n29983), .B(\filter_0/n8100 ), .X(n29190) );
  nand_x1_sg U56279 ( .A(reg_ow_13[0]), .B(n33499), .X(n29360) );
  nand_x1_sg U56280 ( .A(reg_ow_13[1]), .B(n33505), .X(n29364) );
  nand_x1_sg U56281 ( .A(reg_ow_13[2]), .B(n33504), .X(n29366) );
  nand_x1_sg U56282 ( .A(reg_ow_13[3]), .B(n33499), .X(n29368) );
  nand_x1_sg U56283 ( .A(reg_ow_13[4]), .B(n33500), .X(n29370) );
  nand_x1_sg U56284 ( .A(reg_ow_13[5]), .B(n33500), .X(n29372) );
  nand_x1_sg U56285 ( .A(reg_ow_13[6]), .B(n33505), .X(n29374) );
  nand_x1_sg U56286 ( .A(n33441), .B(\filter_0/n8053 ), .X(n29375) );
  nand_x1_sg U56287 ( .A(reg_ow_13[7]), .B(n33504), .X(n29376) );
  nand_x1_sg U56288 ( .A(n33440), .B(\filter_0/n8052 ), .X(n29377) );
  nand_x1_sg U56289 ( .A(reg_ow_13[8]), .B(n33503), .X(n29378) );
  nand_x1_sg U56290 ( .A(n33440), .B(\filter_0/n8051 ), .X(n29379) );
  nand_x1_sg U56291 ( .A(reg_ow_13[9]), .B(n33500), .X(n29380) );
  nand_x1_sg U56292 ( .A(n29975), .B(\filter_0/n8050 ), .X(n29381) );
  nand_x1_sg U56293 ( .A(reg_ow_13[10]), .B(n33505), .X(n29382) );
  nand_x1_sg U56294 ( .A(n33443), .B(\filter_0/n8049 ), .X(n29383) );
  nand_x1_sg U56295 ( .A(reg_ow_13[11]), .B(n33499), .X(n29384) );
  nand_x1_sg U56296 ( .A(n33440), .B(\filter_0/n8048 ), .X(n29385) );
  nand_x1_sg U56297 ( .A(reg_ow_13[12]), .B(n33500), .X(n29386) );
  nand_x1_sg U56298 ( .A(n33440), .B(\filter_0/n8047 ), .X(n29387) );
  nand_x1_sg U56299 ( .A(reg_ow_13[13]), .B(n33499), .X(n29388) );
  nand_x1_sg U56300 ( .A(n33443), .B(\filter_0/n8046 ), .X(n29389) );
  nand_x1_sg U56301 ( .A(reg_ow_13[14]), .B(n33503), .X(n29390) );
  nand_x1_sg U56302 ( .A(n33441), .B(\filter_0/n8045 ), .X(n29391) );
  nand_x1_sg U56303 ( .A(reg_ow_13[15]), .B(n33503), .X(n29392) );
  nand_x1_sg U56304 ( .A(n33443), .B(\filter_0/n8044 ), .X(n29393) );
  nand_x1_sg U56305 ( .A(reg_ow_13[16]), .B(n33504), .X(n29394) );
  nand_x1_sg U56306 ( .A(n33443), .B(\filter_0/n8043 ), .X(n29395) );
  nand_x1_sg U56307 ( .A(reg_ow_13[17]), .B(n33505), .X(n29396) );
  nand_x1_sg U56308 ( .A(n33442), .B(\filter_0/n8042 ), .X(n29397) );
  nand_x1_sg U56309 ( .A(reg_ow_13[18]), .B(n33503), .X(n29398) );
  nand_x1_sg U56310 ( .A(n33441), .B(\filter_0/n8041 ), .X(n29399) );
  nand_x1_sg U56311 ( .A(reg_ow_13[19]), .B(n33504), .X(n29400) );
  nand_x1_sg U56312 ( .A(n33441), .B(\filter_0/n8040 ), .X(n29401) );
  nand_x1_sg U56313 ( .A(reg_ow_7[1]), .B(n33611), .X(n29237) );
  nand_x1_sg U56314 ( .A(reg_ow_7[3]), .B(n33612), .X(n29241) );
  nand_x1_sg U56315 ( .A(reg_ow_7[5]), .B(n33607), .X(n29245) );
  nand_x1_sg U56316 ( .A(reg_ow_7[7]), .B(n33608), .X(n29249) );
  nand_x1_sg U56317 ( .A(n33397), .B(\filter_0/n8152 ), .X(n29250) );
  nand_x1_sg U56318 ( .A(reg_ow_7[9]), .B(n33607), .X(n29253) );
  nand_x1_sg U56319 ( .A(n33395), .B(\filter_0/n8150 ), .X(n29254) );
  nand_x1_sg U56320 ( .A(reg_ow_7[11]), .B(n33608), .X(n29257) );
  nand_x1_sg U56321 ( .A(n33395), .B(\filter_0/n8148 ), .X(n29258) );
  nand_x1_sg U56322 ( .A(reg_ow_7[13]), .B(n33608), .X(n29261) );
  nand_x1_sg U56323 ( .A(n33398), .B(\filter_0/n8146 ), .X(n29262) );
  nand_x1_sg U56324 ( .A(reg_ow_7[15]), .B(n33613), .X(n29265) );
  nand_x1_sg U56325 ( .A(n33398), .B(\filter_0/n8144 ), .X(n29266) );
  nand_x1_sg U56326 ( .A(reg_ow_7[17]), .B(n33607), .X(n29269) );
  nand_x1_sg U56327 ( .A(n33397), .B(\filter_0/n8142 ), .X(n29270) );
  nand_x1_sg U56328 ( .A(reg_ow_7[19]), .B(n33608), .X(n29273) );
  nand_x1_sg U56329 ( .A(n33396), .B(\filter_0/n8140 ), .X(n29274) );
  nor_x1_sg U56330 ( .A(n32505), .B(\filter_0/reg_o_mask[15] ), .X(n15317) );
  nand_x1_sg U56331 ( .A(reg_ow_10[0]), .B(n33489), .X(n29490) );
  nand_x1_sg U56332 ( .A(reg_ow_10[2]), .B(n33487), .X(n29496) );
  nand_x1_sg U56333 ( .A(reg_ow_10[4]), .B(n33483), .X(n29500) );
  nand_x1_sg U56334 ( .A(reg_ow_10[6]), .B(n33483), .X(n29504) );
  nand_x1_sg U56335 ( .A(n33303), .B(\filter_0/n7973 ), .X(n29505) );
  nand_x1_sg U56336 ( .A(reg_ow_10[8]), .B(n33488), .X(n29508) );
  nand_x1_sg U56337 ( .A(n33303), .B(\filter_0/n7971 ), .X(n29509) );
  nand_x1_sg U56338 ( .A(reg_ow_10[10]), .B(n33484), .X(n29512) );
  nand_x1_sg U56339 ( .A(n33300), .B(\filter_0/n7969 ), .X(n29513) );
  nand_x1_sg U56340 ( .A(reg_ow_10[12]), .B(n33489), .X(n29516) );
  nand_x1_sg U56341 ( .A(n33302), .B(\filter_0/n7967 ), .X(n29517) );
  nand_x1_sg U56342 ( .A(reg_ow_10[14]), .B(n33484), .X(n29520) );
  nand_x1_sg U56343 ( .A(n33302), .B(\filter_0/n7965 ), .X(n29521) );
  nand_x1_sg U56344 ( .A(reg_ow_10[16]), .B(n33488), .X(n29524) );
  nand_x1_sg U56345 ( .A(n33302), .B(\filter_0/n7963 ), .X(n29525) );
  nand_x1_sg U56346 ( .A(reg_ow_10[18]), .B(n33487), .X(n29528) );
  nand_x1_sg U56347 ( .A(n29919), .B(\filter_0/n7961 ), .X(n29529) );
  nand_x1_sg U56348 ( .A(reg_ow_9[0]), .B(n33481), .X(n29534) );
  nand_x1_sg U56349 ( .A(reg_ow_9[2]), .B(n33476), .X(n29540) );
  nand_x1_sg U56350 ( .A(reg_ow_9[4]), .B(n33476), .X(n29544) );
  nand_x1_sg U56351 ( .A(reg_ow_9[6]), .B(n33480), .X(n29548) );
  nand_x1_sg U56352 ( .A(n33295), .B(\filter_0/n7953 ), .X(n29549) );
  nand_x1_sg U56353 ( .A(reg_ow_9[8]), .B(n33480), .X(n29552) );
  nand_x1_sg U56354 ( .A(n33295), .B(\filter_0/n7951 ), .X(n29553) );
  nand_x1_sg U56355 ( .A(reg_ow_9[10]), .B(n33476), .X(n29556) );
  nand_x1_sg U56356 ( .A(n33297), .B(\filter_0/n7949 ), .X(n29557) );
  nand_x1_sg U56357 ( .A(reg_ow_9[12]), .B(n33479), .X(n29560) );
  nand_x1_sg U56358 ( .A(n29917), .B(\filter_0/n7947 ), .X(n29561) );
  nand_x1_sg U56359 ( .A(reg_ow_9[14]), .B(n33475), .X(n29564) );
  nand_x1_sg U56360 ( .A(n33298), .B(\filter_0/n7945 ), .X(n29565) );
  nand_x1_sg U56361 ( .A(reg_ow_9[16]), .B(n33475), .X(n29568) );
  nand_x1_sg U56362 ( .A(n33295), .B(\filter_0/n7943 ), .X(n29569) );
  nand_x1_sg U56363 ( .A(reg_ow_9[18]), .B(n33475), .X(n29572) );
  nand_x1_sg U56364 ( .A(n33296), .B(\filter_0/n7941 ), .X(n29573) );
  nor_x1_sg U56365 ( .A(n32132), .B(\filter_0/reg_o_mask[4] ), .X(n15294) );
  nor_x1_sg U56366 ( .A(n15334), .B(n15335), .X(n15333) );
  nor_x1_sg U56367 ( .A(n32136), .B(\filter_0/reg_o_mask[22] ), .X(n15335) );
  nor_x1_sg U56368 ( .A(n32505), .B(\filter_0/reg_o_mask[23] ), .X(n15334) );
  nand_x1_sg U56369 ( .A(reg_ow_11[1]), .B(n33604), .X(n29449) );
  nand_x1_sg U56370 ( .A(reg_ow_11[3]), .B(n33603), .X(n29453) );
  nand_x1_sg U56371 ( .A(reg_ow_11[5]), .B(n33603), .X(n29457) );
  nand_x1_sg U56372 ( .A(reg_ow_11[7]), .B(n33600), .X(n29461) );
  nand_x1_sg U56373 ( .A(n33402), .B(\filter_0/n7992 ), .X(n29462) );
  nand_x1_sg U56374 ( .A(reg_ow_11[9]), .B(n33599), .X(n29465) );
  nand_x1_sg U56375 ( .A(n33401), .B(\filter_0/n7990 ), .X(n29466) );
  nand_x1_sg U56376 ( .A(reg_ow_11[11]), .B(n33599), .X(n29469) );
  nand_x1_sg U56377 ( .A(n33403), .B(\filter_0/n7988 ), .X(n29470) );
  nand_x1_sg U56378 ( .A(reg_ow_11[13]), .B(n33604), .X(n29473) );
  nand_x1_sg U56379 ( .A(n29959), .B(\filter_0/n7986 ), .X(n29474) );
  nand_x1_sg U56380 ( .A(reg_ow_11[15]), .B(n33603), .X(n29477) );
  nand_x1_sg U56381 ( .A(n33402), .B(\filter_0/n7984 ), .X(n29478) );
  nand_x1_sg U56382 ( .A(reg_ow_11[17]), .B(n33600), .X(n29481) );
  nand_x1_sg U56383 ( .A(n29959), .B(\filter_0/n7982 ), .X(n29482) );
  nand_x1_sg U56384 ( .A(reg_ow_11[19]), .B(n33604), .X(n29485) );
  nand_x1_sg U56385 ( .A(n33402), .B(\filter_0/n7980 ), .X(n29486) );
  nand_x1_sg U56386 ( .A(reg_ow_10[1]), .B(n33483), .X(n29494) );
  nand_x1_sg U56387 ( .A(reg_ow_10[3]), .B(n33487), .X(n29498) );
  nand_x1_sg U56388 ( .A(reg_ow_10[5]), .B(n33484), .X(n29502) );
  nand_x1_sg U56389 ( .A(reg_ow_10[7]), .B(n33488), .X(n29506) );
  nand_x1_sg U56390 ( .A(n33300), .B(\filter_0/n7972 ), .X(n29507) );
  nand_x1_sg U56391 ( .A(reg_ow_10[9]), .B(n33487), .X(n29510) );
  nand_x1_sg U56392 ( .A(n33301), .B(\filter_0/n7970 ), .X(n29511) );
  nand_x1_sg U56393 ( .A(reg_ow_10[11]), .B(n33489), .X(n29514) );
  nand_x1_sg U56394 ( .A(n33300), .B(\filter_0/n7968 ), .X(n29515) );
  nand_x1_sg U56395 ( .A(reg_ow_10[13]), .B(n33489), .X(n29518) );
  nand_x1_sg U56396 ( .A(n33301), .B(\filter_0/n7966 ), .X(n29519) );
  nand_x1_sg U56397 ( .A(reg_ow_10[15]), .B(n33488), .X(n29522) );
  nand_x1_sg U56398 ( .A(n33303), .B(\filter_0/n7964 ), .X(n29523) );
  nand_x1_sg U56399 ( .A(reg_ow_10[17]), .B(n33483), .X(n29526) );
  nand_x1_sg U56400 ( .A(n33302), .B(\filter_0/n7962 ), .X(n29527) );
  nand_x1_sg U56401 ( .A(reg_ow_10[19]), .B(n33484), .X(n29530) );
  nand_x1_sg U56402 ( .A(n29919), .B(\filter_0/n7960 ), .X(n29531) );
  nand_x1_sg U56403 ( .A(reg_ow_9[1]), .B(n33479), .X(n29538) );
  nand_x1_sg U56404 ( .A(reg_ow_9[3]), .B(n33480), .X(n29542) );
  nand_x1_sg U56405 ( .A(reg_ow_9[5]), .B(n33481), .X(n29546) );
  nand_x1_sg U56406 ( .A(reg_ow_9[7]), .B(n33479), .X(n29550) );
  nand_x1_sg U56407 ( .A(n29917), .B(\filter_0/n7952 ), .X(n29551) );
  nand_x1_sg U56408 ( .A(reg_ow_9[9]), .B(n33476), .X(n29554) );
  nand_x1_sg U56409 ( .A(n33296), .B(\filter_0/n7950 ), .X(n29555) );
  nand_x1_sg U56410 ( .A(reg_ow_9[11]), .B(n33481), .X(n29558) );
  nand_x1_sg U56411 ( .A(n33296), .B(\filter_0/n7948 ), .X(n29559) );
  nand_x1_sg U56412 ( .A(reg_ow_9[13]), .B(n33475), .X(n29562) );
  nand_x1_sg U56413 ( .A(n33298), .B(\filter_0/n7946 ), .X(n29563) );
  nand_x1_sg U56414 ( .A(reg_ow_9[15]), .B(n33479), .X(n29566) );
  nand_x1_sg U56415 ( .A(n33297), .B(\filter_0/n7944 ), .X(n29567) );
  nand_x1_sg U56416 ( .A(reg_ow_9[17]), .B(n33481), .X(n29570) );
  nand_x1_sg U56417 ( .A(n29917), .B(\filter_0/n7942 ), .X(n29571) );
  nand_x1_sg U56418 ( .A(reg_ow_9[19]), .B(n33480), .X(n29574) );
  nand_x1_sg U56419 ( .A(n33297), .B(\filter_0/n7940 ), .X(n29575) );
  nor_x1_sg U56420 ( .A(n32503), .B(\filter_0/reg_o_mask[7] ), .X(n15301) );
  nor_x1_sg U56421 ( .A(n15303), .B(n15304), .X(n15299) );
  nor_x1_sg U56422 ( .A(n15301), .B(n15302), .X(n15300) );
  nor_x1_sg U56423 ( .A(n32114), .B(\filter_0/reg_o_mask[5] ), .X(n15304) );
  nor_x1_sg U56424 ( .A(n15326), .B(n15327), .X(n15325) );
  nor_x1_sg U56425 ( .A(n32118), .B(\filter_0/reg_o_mask[17] ), .X(n15326) );
  nor_x1_sg U56426 ( .A(n32131), .B(\filter_0/reg_o_mask[20] ), .X(n15327) );
  nor_x1_sg U56427 ( .A(n32130), .B(\filter_0/reg_o_mask[12] ), .X(n15311) );
  nor_x1_sg U56428 ( .A(n32122), .B(\filter_0/reg_o_mask[2] ), .X(n15296) );
  nor_x1_sg U56429 ( .A(\filter_0/N13 ), .B(\filter_0/N14 ), .X(n15343) );
  nor_x1_sg U56430 ( .A(n35154), .B(\filter_0/N14 ), .X(n15348) );
  nand_x1_sg U56431 ( .A(n15343), .B(n31655), .X(n15090) );
  nand_x1_sg U56432 ( .A(n15348), .B(n31655), .X(n15105) );
  nor_x1_sg U56433 ( .A(n32119), .B(\filter_0/reg_o_mask[1] ), .X(n15293) );
  nor_x1_sg U56434 ( .A(n32206), .B(\filter_0/reg_o_mask[3] ), .X(n15303) );
  nor_x1_sg U56435 ( .A(n32135), .B(\filter_0/reg_o_mask[14] ), .X(n15318) );
  nor_x1_sg U56436 ( .A(n31656), .B(n35154), .X(n15355) );
  nor_x1_sg U56437 ( .A(n15353), .B(n15354), .X(n15350) );
  nor_x1_sg U56438 ( .A(n32207), .B(\filter_0/reg_o_mask[27] ), .X(n15354) );
  nor_x1_sg U56439 ( .A(n15101), .B(\filter_0/reg_o_mask[30] ), .X(n15353) );
  nor_x1_sg U56440 ( .A(n15336), .B(n15337), .X(n15332) );
  nor_x1_sg U56441 ( .A(n32116), .B(\filter_0/reg_o_mask[21] ), .X(n15337) );
  nor_x1_sg U56442 ( .A(n32205), .B(\filter_0/reg_o_mask[19] ), .X(n15336) );
  nor_x1_sg U56443 ( .A(n32118), .B(\filter_0/reg_o_mask[9] ), .X(n15309) );
  nor_x1_sg U56444 ( .A(n35268), .B(\filter_0/N13 ), .X(n15161) );
  nor_x1_sg U56445 ( .A(n32208), .B(\filter_0/reg_o_mask[11] ), .X(n15319) );
  nor_x1_sg U56446 ( .A(n15341), .B(n15342), .X(n15340) );
  nor_x1_sg U56447 ( .A(n32120), .B(\filter_0/reg_o_mask[25] ), .X(n15342) );
  nor_x1_sg U56448 ( .A(n32114), .B(\filter_0/reg_o_mask[29] ), .X(n15341) );
  nand_x1_sg U56449 ( .A(n15161), .B(n31656), .X(n15104) );
  nor_x1_sg U56450 ( .A(n32115), .B(\filter_0/reg_o_mask[13] ), .X(n15308) );
  nor_x1_sg U56451 ( .A(n32134), .B(\filter_0/reg_o_mask[6] ), .X(n15302) );
  nand_x1_sg U56452 ( .A(reg_ow_0[0]), .B(n33703), .X(n29621) );
  nand_x1_sg U56453 ( .A(reg_ow_0[1]), .B(n33704), .X(n29625) );
  nand_x1_sg U56454 ( .A(reg_ow_0[2]), .B(n33703), .X(n29627) );
  nand_x1_sg U56455 ( .A(reg_ow_0[3]), .B(n33703), .X(n29629) );
  nand_x1_sg U56456 ( .A(reg_ow_0[4]), .B(n33708), .X(n29631) );
  nand_x1_sg U56457 ( .A(reg_ow_0[5]), .B(n33709), .X(n29633) );
  nand_x1_sg U56458 ( .A(reg_ow_0[6]), .B(n33704), .X(n29635) );
  nand_x1_sg U56459 ( .A(n33391), .B(\filter_0/n8173 ), .X(n29636) );
  nand_x1_sg U56460 ( .A(reg_ow_0[7]), .B(n33704), .X(n29637) );
  nand_x1_sg U56461 ( .A(n33392), .B(\filter_0/n8172 ), .X(n29638) );
  nand_x1_sg U56462 ( .A(reg_ow_0[8]), .B(n33708), .X(n29639) );
  nand_x1_sg U56463 ( .A(n33392), .B(\filter_0/n8171 ), .X(n29640) );
  nand_x1_sg U56464 ( .A(reg_ow_0[9]), .B(n33704), .X(n29641) );
  nand_x1_sg U56465 ( .A(n33391), .B(\filter_0/n8170 ), .X(n29642) );
  nand_x1_sg U56466 ( .A(reg_ow_0[10]), .B(n33703), .X(n29643) );
  nand_x1_sg U56467 ( .A(n33390), .B(\filter_0/n8169 ), .X(n29644) );
  nand_x1_sg U56468 ( .A(reg_ow_0[11]), .B(n33707), .X(n29645) );
  nand_x1_sg U56469 ( .A(n33393), .B(\filter_0/n8168 ), .X(n29646) );
  nand_x1_sg U56470 ( .A(reg_ow_0[12]), .B(n33708), .X(n29647) );
  nand_x1_sg U56471 ( .A(n29955), .B(\filter_0/n8167 ), .X(n29648) );
  nand_x1_sg U56472 ( .A(reg_ow_0[13]), .B(n33709), .X(n29649) );
  nand_x1_sg U56473 ( .A(n33390), .B(\filter_0/n8166 ), .X(n29650) );
  nand_x1_sg U56474 ( .A(reg_ow_0[14]), .B(n33709), .X(n29651) );
  nand_x1_sg U56475 ( .A(n33391), .B(\filter_0/n8165 ), .X(n29652) );
  nand_x1_sg U56476 ( .A(reg_ow_0[15]), .B(n33707), .X(n29653) );
  nand_x1_sg U56477 ( .A(n33392), .B(\filter_0/n8164 ), .X(n29654) );
  nand_x1_sg U56478 ( .A(reg_ow_0[16]), .B(n33707), .X(n29655) );
  nand_x1_sg U56479 ( .A(n33392), .B(\filter_0/n8163 ), .X(n29656) );
  nand_x1_sg U56480 ( .A(reg_ow_0[17]), .B(n33708), .X(n29657) );
  nand_x1_sg U56481 ( .A(n33393), .B(\filter_0/n8162 ), .X(n29658) );
  nand_x1_sg U56482 ( .A(reg_ow_0[18]), .B(n33709), .X(n29659) );
  nand_x1_sg U56483 ( .A(n29955), .B(\filter_0/n8161 ), .X(n29660) );
  nand_x1_sg U56484 ( .A(reg_ow_0[19]), .B(n33707), .X(n29661) );
  nand_x1_sg U56485 ( .A(n29955), .B(\filter_0/n8160 ), .X(n29662) );
  nand_x1_sg U56486 ( .A(reg_ow_4[0]), .B(n33595), .X(n29105) );
  nand_x1_sg U56487 ( .A(reg_ow_4[1]), .B(n33591), .X(n29109) );
  nand_x1_sg U56488 ( .A(reg_ow_4[2]), .B(n33592), .X(n29111) );
  nand_x1_sg U56489 ( .A(reg_ow_4[3]), .B(n33595), .X(n29113) );
  nand_x1_sg U56490 ( .A(reg_ow_4[4]), .B(n33597), .X(n29115) );
  nand_x1_sg U56491 ( .A(reg_ow_4[5]), .B(n33591), .X(n29117) );
  nand_x1_sg U56492 ( .A(reg_ow_4[6]), .B(n33597), .X(n29119) );
  nand_x1_sg U56493 ( .A(n33456), .B(\filter_0/n8093 ), .X(n29120) );
  nand_x1_sg U56494 ( .A(reg_ow_4[7]), .B(n33596), .X(n29121) );
  nand_x1_sg U56495 ( .A(n33456), .B(\filter_0/n8092 ), .X(n29122) );
  nand_x1_sg U56496 ( .A(reg_ow_4[8]), .B(n33595), .X(n29123) );
  nand_x1_sg U56497 ( .A(n33455), .B(\filter_0/n8091 ), .X(n29124) );
  nand_x1_sg U56498 ( .A(reg_ow_4[9]), .B(n33592), .X(n29125) );
  nand_x1_sg U56499 ( .A(n33455), .B(\filter_0/n8090 ), .X(n29126) );
  nand_x1_sg U56500 ( .A(reg_ow_4[10]), .B(n33596), .X(n29127) );
  nand_x1_sg U56501 ( .A(n29981), .B(\filter_0/n8089 ), .X(n29128) );
  nand_x1_sg U56502 ( .A(reg_ow_4[11]), .B(n33596), .X(n29129) );
  nand_x1_sg U56503 ( .A(n33458), .B(\filter_0/n8088 ), .X(n29130) );
  nand_x1_sg U56504 ( .A(reg_ow_4[12]), .B(n33597), .X(n29131) );
  nand_x1_sg U56505 ( .A(n29981), .B(\filter_0/n8087 ), .X(n29132) );
  nand_x1_sg U56506 ( .A(reg_ow_4[13]), .B(n33596), .X(n29133) );
  nand_x1_sg U56507 ( .A(n33457), .B(\filter_0/n8086 ), .X(n29134) );
  nand_x1_sg U56508 ( .A(reg_ow_4[14]), .B(n33595), .X(n29135) );
  nand_x1_sg U56509 ( .A(n33455), .B(\filter_0/n8085 ), .X(n29136) );
  nand_x1_sg U56510 ( .A(reg_ow_4[15]), .B(n33592), .X(n29137) );
  nand_x1_sg U56511 ( .A(n33458), .B(\filter_0/n8084 ), .X(n29138) );
  nand_x1_sg U56512 ( .A(reg_ow_4[16]), .B(n33591), .X(n29139) );
  nand_x1_sg U56513 ( .A(n33457), .B(\filter_0/n8083 ), .X(n29140) );
  nand_x1_sg U56514 ( .A(reg_ow_4[17]), .B(n33597), .X(n29141) );
  nand_x1_sg U56515 ( .A(n29981), .B(\filter_0/n8082 ), .X(n29142) );
  nand_x1_sg U56516 ( .A(reg_ow_4[18]), .B(n33591), .X(n29143) );
  nand_x1_sg U56517 ( .A(n33457), .B(\filter_0/n8081 ), .X(n29144) );
  nand_x1_sg U56518 ( .A(reg_ow_4[19]), .B(n33592), .X(n29145) );
  nand_x1_sg U56519 ( .A(n33458), .B(\filter_0/n8080 ), .X(n29146) );
  nand_x1_sg U56520 ( .A(reg_oi_0[0]), .B(n33589), .X(n28922) );
  nand_x1_sg U56521 ( .A(reg_oi_0[1]), .B(n33584), .X(n28926) );
  nand_x1_sg U56522 ( .A(reg_oi_0[2]), .B(n33583), .X(n28928) );
  nand_x1_sg U56523 ( .A(reg_oi_0[3]), .B(n33583), .X(n28930) );
  nand_x1_sg U56524 ( .A(reg_oi_0[4]), .B(n33589), .X(n28932) );
  nand_x1_sg U56525 ( .A(reg_oi_0[5]), .B(n33583), .X(n28934) );
  nand_x1_sg U56526 ( .A(reg_oi_0[6]), .B(n33588), .X(n28936) );
  nand_x1_sg U56527 ( .A(n33452), .B(\filter_0/n7844 ), .X(n28937) );
  nand_x1_sg U56528 ( .A(reg_oi_0[7]), .B(n33587), .X(n28938) );
  nand_x1_sg U56529 ( .A(n33451), .B(\filter_0/n7843 ), .X(n28939) );
  nand_x1_sg U56530 ( .A(reg_oi_0[8]), .B(n33589), .X(n28940) );
  nand_x1_sg U56531 ( .A(n33452), .B(\filter_0/n7842 ), .X(n28941) );
  nand_x1_sg U56532 ( .A(reg_oi_0[9]), .B(n33584), .X(n28942) );
  nand_x1_sg U56533 ( .A(n33453), .B(\filter_0/n7841 ), .X(n28943) );
  nand_x1_sg U56534 ( .A(reg_oi_0[10]), .B(n33583), .X(n28944) );
  nand_x1_sg U56535 ( .A(n29979), .B(\filter_0/n7840 ), .X(n28945) );
  nand_x1_sg U56536 ( .A(reg_oi_0[11]), .B(n33587), .X(n28946) );
  nand_x1_sg U56537 ( .A(n33453), .B(\filter_0/n7839 ), .X(n28947) );
  nand_x1_sg U56538 ( .A(reg_oi_0[12]), .B(n33589), .X(n28948) );
  nand_x1_sg U56539 ( .A(n33450), .B(\filter_0/n7838 ), .X(n28949) );
  nand_x1_sg U56540 ( .A(reg_oi_0[13]), .B(n33584), .X(n28950) );
  nand_x1_sg U56541 ( .A(n33453), .B(\filter_0/n7837 ), .X(n28951) );
  nand_x1_sg U56542 ( .A(reg_oi_0[14]), .B(n33584), .X(n28952) );
  nand_x1_sg U56543 ( .A(n33451), .B(\filter_0/n7836 ), .X(n28953) );
  nand_x1_sg U56544 ( .A(reg_oi_0[15]), .B(n33587), .X(n28954) );
  nand_x1_sg U56545 ( .A(n29979), .B(\filter_0/n7835 ), .X(n28955) );
  nand_x1_sg U56546 ( .A(reg_oi_0[16]), .B(n33588), .X(n28956) );
  nand_x1_sg U56547 ( .A(n33450), .B(\filter_0/n7834 ), .X(n28957) );
  nand_x1_sg U56548 ( .A(reg_oi_0[17]), .B(n33587), .X(n28958) );
  nand_x1_sg U56549 ( .A(n33453), .B(\filter_0/n7833 ), .X(n28959) );
  nand_x1_sg U56550 ( .A(reg_oi_0[18]), .B(n33588), .X(n28960) );
  nand_x1_sg U56551 ( .A(n33451), .B(\filter_0/n7832 ), .X(n28961) );
  nand_x1_sg U56552 ( .A(reg_oi_0[19]), .B(n33588), .X(n28962) );
  nand_x1_sg U56553 ( .A(n29979), .B(\filter_0/n7831 ), .X(n28963) );
  nand_x1_sg U56554 ( .A(reg_oi_4[0]), .B(n33776), .X(n28406) );
  nand_x1_sg U56555 ( .A(reg_oi_4[1]), .B(n33773), .X(n28410) );
  nand_x1_sg U56556 ( .A(reg_oi_4[2]), .B(n33776), .X(n28412) );
  nand_x1_sg U56557 ( .A(reg_oi_4[3]), .B(n33776), .X(n28414) );
  nand_x1_sg U56558 ( .A(reg_oi_4[4]), .B(n33777), .X(n28416) );
  nand_x1_sg U56559 ( .A(reg_oi_4[5]), .B(n33772), .X(n28418) );
  nand_x1_sg U56560 ( .A(reg_oi_4[6]), .B(n33778), .X(n28420) );
  nand_x1_sg U56561 ( .A(n33386), .B(\filter_0/n7764 ), .X(n28421) );
  nand_x1_sg U56562 ( .A(reg_oi_4[7]), .B(n33777), .X(n28422) );
  nand_x1_sg U56563 ( .A(n33385), .B(\filter_0/n7763 ), .X(n28423) );
  nand_x1_sg U56564 ( .A(reg_oi_4[8]), .B(n33776), .X(n28424) );
  nand_x1_sg U56565 ( .A(n29953), .B(\filter_0/n7762 ), .X(n28425) );
  nand_x1_sg U56566 ( .A(reg_oi_4[9]), .B(n33773), .X(n28426) );
  nand_x1_sg U56567 ( .A(n29953), .B(\filter_0/n7761 ), .X(n28427) );
  nand_x1_sg U56568 ( .A(reg_oi_4[10]), .B(n33778), .X(n28428) );
  nand_x1_sg U56569 ( .A(n33385), .B(\filter_0/n7760 ), .X(n28429) );
  nand_x1_sg U56570 ( .A(reg_oi_4[11]), .B(n33772), .X(n28430) );
  nand_x1_sg U56571 ( .A(n33386), .B(\filter_0/n7759 ), .X(n28431) );
  nand_x1_sg U56572 ( .A(reg_oi_4[12]), .B(n33773), .X(n28432) );
  nand_x1_sg U56573 ( .A(n33387), .B(\filter_0/n7758 ), .X(n28433) );
  nand_x1_sg U56574 ( .A(reg_oi_4[13]), .B(n33772), .X(n28434) );
  nand_x1_sg U56575 ( .A(n33388), .B(\filter_0/n7757 ), .X(n28435) );
  nand_x1_sg U56576 ( .A(reg_oi_4[14]), .B(n33777), .X(n28436) );
  nand_x1_sg U56577 ( .A(n33388), .B(\filter_0/n7756 ), .X(n28437) );
  nand_x1_sg U56578 ( .A(reg_oi_4[15]), .B(n33778), .X(n28438) );
  nand_x1_sg U56579 ( .A(n29953), .B(\filter_0/n7755 ), .X(n28439) );
  nand_x1_sg U56580 ( .A(reg_oi_4[16]), .B(n33778), .X(n28440) );
  nand_x1_sg U56581 ( .A(n33388), .B(\filter_0/n7754 ), .X(n28441) );
  nand_x1_sg U56582 ( .A(reg_oi_4[17]), .B(n33773), .X(n28442) );
  nand_x1_sg U56583 ( .A(n33385), .B(\filter_0/n7753 ), .X(n28443) );
  nand_x1_sg U56584 ( .A(reg_oi_4[18]), .B(n33772), .X(n28444) );
  nand_x1_sg U56585 ( .A(n33386), .B(\filter_0/n7752 ), .X(n28445) );
  nand_x1_sg U56586 ( .A(reg_oi_4[19]), .B(n33777), .X(n28446) );
  nand_x1_sg U56587 ( .A(n33388), .B(\filter_0/n7751 ), .X(n28447) );
  nand_x1_sg U56588 ( .A(reg_oi_3[0]), .B(n33565), .X(n28363) );
  nand_x1_sg U56589 ( .A(reg_oi_3[1]), .B(n33560), .X(n28367) );
  nand_x1_sg U56590 ( .A(reg_oi_3[2]), .B(n33564), .X(n28369) );
  nand_x1_sg U56591 ( .A(reg_oi_3[3]), .B(n33563), .X(n28371) );
  nand_x1_sg U56592 ( .A(reg_oi_3[4]), .B(n33564), .X(n28373) );
  nand_x1_sg U56593 ( .A(reg_oi_3[5]), .B(n33559), .X(n28375) );
  nand_x1_sg U56594 ( .A(reg_oi_3[6]), .B(n33565), .X(n28377) );
  nand_x1_sg U56595 ( .A(n33445), .B(\filter_0/n7904 ), .X(n28378) );
  nand_x1_sg U56596 ( .A(reg_oi_3[7]), .B(n33563), .X(n28379) );
  nand_x1_sg U56597 ( .A(n33448), .B(\filter_0/n7903 ), .X(n28380) );
  nand_x1_sg U56598 ( .A(reg_oi_3[8]), .B(n33565), .X(n28381) );
  nand_x1_sg U56599 ( .A(n33448), .B(\filter_0/n7902 ), .X(n28382) );
  nand_x1_sg U56600 ( .A(reg_oi_3[9]), .B(n33564), .X(n28383) );
  nand_x1_sg U56601 ( .A(n33446), .B(\filter_0/n7901 ), .X(n28384) );
  nand_x1_sg U56602 ( .A(reg_oi_3[10]), .B(n33563), .X(n28385) );
  nand_x1_sg U56603 ( .A(n33447), .B(\filter_0/n7900 ), .X(n28386) );
  nand_x1_sg U56604 ( .A(reg_oi_3[11]), .B(n33564), .X(n28387) );
  nand_x1_sg U56605 ( .A(n29977), .B(\filter_0/n7899 ), .X(n28388) );
  nand_x1_sg U56606 ( .A(reg_oi_3[12]), .B(n33559), .X(n28389) );
  nand_x1_sg U56607 ( .A(n33446), .B(\filter_0/n7898 ), .X(n28390) );
  nand_x1_sg U56608 ( .A(reg_oi_3[13]), .B(n33560), .X(n28391) );
  nand_x1_sg U56609 ( .A(n33445), .B(\filter_0/n7897 ), .X(n28392) );
  nand_x1_sg U56610 ( .A(reg_oi_3[14]), .B(n33560), .X(n28393) );
  nand_x1_sg U56611 ( .A(n33446), .B(\filter_0/n7896 ), .X(n28394) );
  nand_x1_sg U56612 ( .A(reg_oi_3[15]), .B(n33560), .X(n28395) );
  nand_x1_sg U56613 ( .A(n33447), .B(\filter_0/n7895 ), .X(n28396) );
  nand_x1_sg U56614 ( .A(reg_oi_3[16]), .B(n33559), .X(n28397) );
  nand_x1_sg U56615 ( .A(n33445), .B(\filter_0/n7894 ), .X(n28398) );
  nand_x1_sg U56616 ( .A(reg_oi_3[17]), .B(n33565), .X(n28399) );
  nand_x1_sg U56617 ( .A(n33447), .B(\filter_0/n7893 ), .X(n28400) );
  nand_x1_sg U56618 ( .A(reg_oi_3[18]), .B(n33559), .X(n28401) );
  nand_x1_sg U56619 ( .A(n29977), .B(\filter_0/n7892 ), .X(n28402) );
  nand_x1_sg U56620 ( .A(reg_oi_3[19]), .B(n33563), .X(n28403) );
  nand_x1_sg U56621 ( .A(n33448), .B(\filter_0/n7891 ), .X(n28404) );
  nand_x1_sg U56622 ( .A(reg_oi_15[0]), .B(n33568), .X(n28576) );
  nand_x1_sg U56623 ( .A(reg_oi_15[1]), .B(n33572), .X(n28580) );
  nand_x1_sg U56624 ( .A(reg_oi_15[2]), .B(n33571), .X(n28582) );
  nand_x1_sg U56625 ( .A(reg_oi_15[3]), .B(n33571), .X(n28584) );
  nand_x1_sg U56626 ( .A(reg_oi_15[4]), .B(n33568), .X(n28586) );
  nand_x1_sg U56627 ( .A(reg_oi_15[5]), .B(n33568), .X(n28588) );
  nand_x1_sg U56628 ( .A(reg_oi_15[6]), .B(n33573), .X(n28590) );
  nand_x1_sg U56629 ( .A(n33383), .B(\filter_0/n7684 ), .X(n28591) );
  nand_x1_sg U56630 ( .A(reg_oi_15[7]), .B(n33567), .X(n28592) );
  nand_x1_sg U56631 ( .A(n33381), .B(\filter_0/n7683 ), .X(n28593) );
  nand_x1_sg U56632 ( .A(reg_oi_15[8]), .B(n33568), .X(n28594) );
  nand_x1_sg U56633 ( .A(n29951), .B(\filter_0/n7682 ), .X(n28595) );
  nand_x1_sg U56634 ( .A(reg_oi_15[9]), .B(n33573), .X(n28596) );
  nand_x1_sg U56635 ( .A(n29951), .B(\filter_0/n7681 ), .X(n28597) );
  nand_x1_sg U56636 ( .A(reg_oi_15[10]), .B(n33567), .X(n28598) );
  nand_x1_sg U56637 ( .A(n33382), .B(\filter_0/n7680 ), .X(n28599) );
  nand_x1_sg U56638 ( .A(reg_oi_15[11]), .B(n33572), .X(n28600) );
  nand_x1_sg U56639 ( .A(n33382), .B(\filter_0/n7679 ), .X(n28601) );
  nand_x1_sg U56640 ( .A(reg_oi_15[12]), .B(n33567), .X(n28602) );
  nand_x1_sg U56641 ( .A(n33383), .B(\filter_0/n7678 ), .X(n28603) );
  nand_x1_sg U56642 ( .A(reg_oi_15[13]), .B(n33572), .X(n28604) );
  nand_x1_sg U56643 ( .A(n33380), .B(\filter_0/n7677 ), .X(n28605) );
  nand_x1_sg U56644 ( .A(reg_oi_15[14]), .B(n33571), .X(n28606) );
  nand_x1_sg U56645 ( .A(n33383), .B(\filter_0/n7676 ), .X(n28607) );
  nand_x1_sg U56646 ( .A(reg_oi_15[15]), .B(n33573), .X(n28608) );
  nand_x1_sg U56647 ( .A(n33383), .B(\filter_0/n7675 ), .X(n28609) );
  nand_x1_sg U56648 ( .A(reg_oi_15[16]), .B(n33573), .X(n28610) );
  nand_x1_sg U56649 ( .A(n33381), .B(\filter_0/n7674 ), .X(n28611) );
  nand_x1_sg U56650 ( .A(reg_oi_15[17]), .B(n33572), .X(n28612) );
  nand_x1_sg U56651 ( .A(n33381), .B(\filter_0/n7673 ), .X(n28613) );
  nand_x1_sg U56652 ( .A(reg_oi_15[18]), .B(n33567), .X(n28614) );
  nand_x1_sg U56653 ( .A(n33382), .B(\filter_0/n7672 ), .X(n28615) );
  nand_x1_sg U56654 ( .A(reg_oi_15[19]), .B(n33571), .X(n28616) );
  nand_x1_sg U56655 ( .A(n29951), .B(\filter_0/n7671 ), .X(n28617) );
  nand_x1_sg U56656 ( .A(reg_oi_11[0]), .B(n33575), .X(n28746) );
  nand_x1_sg U56657 ( .A(reg_oi_11[1]), .B(n33576), .X(n28750) );
  nand_x1_sg U56658 ( .A(reg_oi_11[2]), .B(n33576), .X(n28752) );
  nand_x1_sg U56659 ( .A(reg_oi_11[3]), .B(n33580), .X(n28754) );
  nand_x1_sg U56660 ( .A(reg_oi_11[4]), .B(n33580), .X(n28756) );
  nand_x1_sg U56661 ( .A(reg_oi_11[5]), .B(n33579), .X(n28758) );
  nand_x1_sg U56662 ( .A(reg_oi_11[6]), .B(n33575), .X(n28760) );
  nand_x1_sg U56663 ( .A(n33378), .B(\filter_0/n7664 ), .X(n28761) );
  nand_x1_sg U56664 ( .A(reg_oi_11[7]), .B(n33580), .X(n28762) );
  nand_x1_sg U56665 ( .A(n29949), .B(\filter_0/n7663 ), .X(n28763) );
  nand_x1_sg U56666 ( .A(reg_oi_11[8]), .B(n33579), .X(n28764) );
  nand_x1_sg U56667 ( .A(n33377), .B(\filter_0/n7662 ), .X(n28765) );
  nand_x1_sg U56668 ( .A(reg_oi_11[9]), .B(n33579), .X(n28766) );
  nand_x1_sg U56669 ( .A(n33376), .B(\filter_0/n7661 ), .X(n28767) );
  nand_x1_sg U56670 ( .A(reg_oi_11[10]), .B(n33580), .X(n28768) );
  nand_x1_sg U56671 ( .A(n33377), .B(\filter_0/n7660 ), .X(n28769) );
  nand_x1_sg U56672 ( .A(reg_oi_11[11]), .B(n33575), .X(n28770) );
  nand_x1_sg U56673 ( .A(n33378), .B(\filter_0/n7659 ), .X(n28771) );
  nand_x1_sg U56674 ( .A(reg_oi_11[12]), .B(n33581), .X(n28772) );
  nand_x1_sg U56675 ( .A(n29949), .B(\filter_0/n7658 ), .X(n28773) );
  nand_x1_sg U56676 ( .A(reg_oi_11[13]), .B(n33576), .X(n28774) );
  nand_x1_sg U56677 ( .A(n33377), .B(\filter_0/n7657 ), .X(n28775) );
  nand_x1_sg U56678 ( .A(reg_oi_11[14]), .B(n33581), .X(n28776) );
  nand_x1_sg U56679 ( .A(n33375), .B(\filter_0/n7656 ), .X(n28777) );
  nand_x1_sg U56680 ( .A(reg_oi_11[15]), .B(n33579), .X(n28778) );
  nand_x1_sg U56681 ( .A(n33375), .B(\filter_0/n7655 ), .X(n28779) );
  nand_x1_sg U56682 ( .A(reg_oi_11[16]), .B(n33575), .X(n28780) );
  nand_x1_sg U56683 ( .A(n33376), .B(\filter_0/n7654 ), .X(n28781) );
  nand_x1_sg U56684 ( .A(reg_oi_11[17]), .B(n33581), .X(n28782) );
  nand_x1_sg U56685 ( .A(n33375), .B(\filter_0/n7653 ), .X(n28783) );
  nand_x1_sg U56686 ( .A(reg_oi_11[18]), .B(n33581), .X(n28784) );
  nand_x1_sg U56687 ( .A(n33375), .B(\filter_0/n7652 ), .X(n28785) );
  nand_x1_sg U56688 ( .A(reg_oi_11[19]), .B(n33576), .X(n28786) );
  nand_x1_sg U56689 ( .A(n33376), .B(\filter_0/n7651 ), .X(n28787) );
  nand_x1_sg U56690 ( .A(reg_ow_12[0]), .B(n33540), .X(n29402) );
  nand_x1_sg U56691 ( .A(reg_ow_12[2]), .B(n33539), .X(n29408) );
  nand_x1_sg U56692 ( .A(reg_ow_12[4]), .B(n33535), .X(n29412) );
  nand_x1_sg U56693 ( .A(reg_ow_12[6]), .B(n33535), .X(n29416) );
  nand_x1_sg U56694 ( .A(n33331), .B(\filter_0/n8033 ), .X(n29417) );
  nand_x1_sg U56695 ( .A(reg_ow_12[8]), .B(n33539), .X(n29420) );
  nand_x1_sg U56696 ( .A(n33330), .B(\filter_0/n8031 ), .X(n29421) );
  nand_x1_sg U56697 ( .A(reg_ow_12[10]), .B(n33536), .X(n29424) );
  nand_x1_sg U56698 ( .A(n33331), .B(\filter_0/n8029 ), .X(n29425) );
  nand_x1_sg U56699 ( .A(reg_ow_12[12]), .B(n33536), .X(n29428) );
  nand_x1_sg U56700 ( .A(n33332), .B(\filter_0/n8027 ), .X(n29429) );
  nand_x1_sg U56701 ( .A(reg_ow_12[14]), .B(n33536), .X(n29432) );
  nand_x1_sg U56702 ( .A(n33333), .B(\filter_0/n8025 ), .X(n29433) );
  nand_x1_sg U56703 ( .A(reg_ow_12[16]), .B(n33539), .X(n29436) );
  nand_x1_sg U56704 ( .A(n33333), .B(\filter_0/n8023 ), .X(n29437) );
  nand_x1_sg U56705 ( .A(reg_ow_12[18]), .B(n33540), .X(n29440) );
  nand_x1_sg U56706 ( .A(n33331), .B(\filter_0/n8021 ), .X(n29441) );
  nand_x1_sg U56707 ( .A(reg_ow_8[0]), .B(n33701), .X(n29578) );
  nand_x1_sg U56708 ( .A(reg_ow_8[2]), .B(n33699), .X(n29584) );
  nand_x1_sg U56709 ( .A(reg_ow_8[4]), .B(n33699), .X(n29588) );
  nand_x1_sg U56710 ( .A(reg_ow_8[6]), .B(n33695), .X(n29592) );
  nand_x1_sg U56711 ( .A(n29929), .B(\filter_0/n7933 ), .X(n29593) );
  nand_x1_sg U56712 ( .A(reg_ow_8[8]), .B(n33696), .X(n29596) );
  nand_x1_sg U56713 ( .A(n33327), .B(\filter_0/n7931 ), .X(n29597) );
  nand_x1_sg U56714 ( .A(reg_ow_8[10]), .B(n33696), .X(n29600) );
  nand_x1_sg U56715 ( .A(n33327), .B(\filter_0/n7929 ), .X(n29601) );
  nand_x1_sg U56716 ( .A(reg_ow_8[12]), .B(n33696), .X(n29604) );
  nand_x1_sg U56717 ( .A(n29929), .B(\filter_0/n7927 ), .X(n29605) );
  nand_x1_sg U56718 ( .A(reg_ow_8[14]), .B(n33701), .X(n29608) );
  nand_x1_sg U56719 ( .A(n33325), .B(\filter_0/n7925 ), .X(n29609) );
  nand_x1_sg U56720 ( .A(reg_ow_8[16]), .B(n33701), .X(n29612) );
  nand_x1_sg U56721 ( .A(n33326), .B(\filter_0/n7923 ), .X(n29613) );
  nand_x1_sg U56722 ( .A(reg_ow_8[18]), .B(n33699), .X(n29616) );
  nand_x1_sg U56723 ( .A(n33327), .B(\filter_0/n7921 ), .X(n29617) );
  nand_x1_sg U56724 ( .A(reg_oi_12[0]), .B(n33685), .X(n28703) );
  nand_x1_sg U56725 ( .A(reg_oi_12[2]), .B(n33679), .X(n28709) );
  nand_x1_sg U56726 ( .A(reg_oi_12[4]), .B(n33680), .X(n28713) );
  nand_x1_sg U56727 ( .A(reg_oi_12[6]), .B(n33680), .X(n28717) );
  nand_x1_sg U56728 ( .A(n29947), .B(\filter_0/n7704 ), .X(n28718) );
  nand_x1_sg U56729 ( .A(reg_oi_12[8]), .B(n33683), .X(n28721) );
  nand_x1_sg U56730 ( .A(n33373), .B(\filter_0/n7702 ), .X(n28722) );
  nand_x1_sg U56731 ( .A(reg_oi_12[10]), .B(n33680), .X(n28725) );
  nand_x1_sg U56732 ( .A(n33371), .B(\filter_0/n7700 ), .X(n28726) );
  nand_x1_sg U56733 ( .A(reg_oi_12[12]), .B(n33684), .X(n28729) );
  nand_x1_sg U56734 ( .A(n33373), .B(\filter_0/n7698 ), .X(n28730) );
  nand_x1_sg U56735 ( .A(reg_oi_12[14]), .B(n33685), .X(n28733) );
  nand_x1_sg U56736 ( .A(n33373), .B(\filter_0/n7696 ), .X(n28734) );
  nand_x1_sg U56737 ( .A(reg_oi_12[16]), .B(n33684), .X(n28737) );
  nand_x1_sg U56738 ( .A(n33370), .B(\filter_0/n7694 ), .X(n28738) );
  nand_x1_sg U56739 ( .A(reg_oi_12[18]), .B(n33685), .X(n28741) );
  nand_x1_sg U56740 ( .A(n33372), .B(\filter_0/n7692 ), .X(n28742) );
  nand_x1_sg U56741 ( .A(reg_oi_8[0]), .B(n33531), .X(n28879) );
  nand_x1_sg U56742 ( .A(reg_oi_8[2]), .B(n33527), .X(n28885) );
  nand_x1_sg U56743 ( .A(reg_oi_8[4]), .B(n33528), .X(n28889) );
  nand_x1_sg U56744 ( .A(reg_oi_8[6]), .B(n33531), .X(n28893) );
  nand_x1_sg U56745 ( .A(n33320), .B(\filter_0/n7604 ), .X(n28894) );
  nand_x1_sg U56746 ( .A(reg_oi_8[8]), .B(n33531), .X(n28897) );
  nand_x1_sg U56747 ( .A(n33322), .B(\filter_0/n7602 ), .X(n28898) );
  nand_x1_sg U56748 ( .A(reg_oi_8[10]), .B(n33528), .X(n28901) );
  nand_x1_sg U56749 ( .A(n33323), .B(\filter_0/n7600 ), .X(n28902) );
  nand_x1_sg U56750 ( .A(reg_oi_8[12]), .B(n33532), .X(n28905) );
  nand_x1_sg U56751 ( .A(n33323), .B(\filter_0/n7598 ), .X(n28906) );
  nand_x1_sg U56752 ( .A(reg_oi_8[14]), .B(n33528), .X(n28909) );
  nand_x1_sg U56753 ( .A(n33321), .B(\filter_0/n7596 ), .X(n28910) );
  nand_x1_sg U56754 ( .A(reg_oi_8[16]), .B(n33533), .X(n28913) );
  nand_x1_sg U56755 ( .A(n33320), .B(\filter_0/n7594 ), .X(n28914) );
  nand_x1_sg U56756 ( .A(reg_oi_8[18]), .B(n33527), .X(n28917) );
  nand_x1_sg U56757 ( .A(n33322), .B(\filter_0/n7592 ), .X(n28918) );
  nand_x1_sg U56758 ( .A(reg_oi_2[0]), .B(n33643), .X(n28320) );
  nand_x1_sg U56759 ( .A(reg_oi_2[1]), .B(n33640), .X(n28324) );
  nand_x1_sg U56760 ( .A(reg_oi_2[2]), .B(n33644), .X(n28326) );
  nand_x1_sg U56761 ( .A(reg_oi_2[3]), .B(n33643), .X(n28328) );
  nand_x1_sg U56762 ( .A(reg_oi_2[4]), .B(n33640), .X(n28330) );
  nand_x1_sg U56763 ( .A(reg_oi_2[5]), .B(n33639), .X(n28332) );
  nand_x1_sg U56764 ( .A(reg_oi_2[6]), .B(n33640), .X(n28334) );
  nand_x1_sg U56765 ( .A(n29945), .B(\filter_0/n7884 ), .X(n28335) );
  nand_x1_sg U56766 ( .A(reg_oi_2[7]), .B(n33639), .X(n28336) );
  nand_x1_sg U56767 ( .A(n33366), .B(\filter_0/n7883 ), .X(n28337) );
  nand_x1_sg U56768 ( .A(reg_oi_2[8]), .B(n33645), .X(n28338) );
  nand_x1_sg U56769 ( .A(n33365), .B(\filter_0/n7882 ), .X(n28339) );
  nand_x1_sg U56770 ( .A(reg_oi_2[9]), .B(n33643), .X(n28340) );
  nand_x1_sg U56771 ( .A(n33368), .B(\filter_0/n7881 ), .X(n28341) );
  nand_x1_sg U56772 ( .A(reg_oi_2[10]), .B(n33640), .X(n28342) );
  nand_x1_sg U56773 ( .A(n33366), .B(\filter_0/n7880 ), .X(n28343) );
  nand_x1_sg U56774 ( .A(reg_oi_2[11]), .B(n33645), .X(n28344) );
  nand_x1_sg U56775 ( .A(n33367), .B(\filter_0/n7879 ), .X(n28345) );
  nand_x1_sg U56776 ( .A(reg_oi_2[12]), .B(n33644), .X(n28346) );
  nand_x1_sg U56777 ( .A(n33366), .B(\filter_0/n7878 ), .X(n28347) );
  nand_x1_sg U56778 ( .A(reg_oi_2[13]), .B(n33644), .X(n28348) );
  nand_x1_sg U56779 ( .A(n33367), .B(\filter_0/n7877 ), .X(n28349) );
  nand_x1_sg U56780 ( .A(reg_oi_2[14]), .B(n33639), .X(n28350) );
  nand_x1_sg U56781 ( .A(n33365), .B(\filter_0/n7876 ), .X(n28351) );
  nand_x1_sg U56782 ( .A(reg_oi_2[15]), .B(n33643), .X(n28352) );
  nand_x1_sg U56783 ( .A(n29945), .B(\filter_0/n7875 ), .X(n28353) );
  nand_x1_sg U56784 ( .A(reg_oi_2[16]), .B(n33639), .X(n28354) );
  nand_x1_sg U56785 ( .A(n33368), .B(\filter_0/n7874 ), .X(n28355) );
  nand_x1_sg U56786 ( .A(reg_oi_2[17]), .B(n33645), .X(n28356) );
  nand_x1_sg U56787 ( .A(n33367), .B(\filter_0/n7873 ), .X(n28357) );
  nand_x1_sg U56788 ( .A(reg_oi_2[18]), .B(n33645), .X(n28358) );
  nand_x1_sg U56789 ( .A(n33365), .B(\filter_0/n7872 ), .X(n28359) );
  nand_x1_sg U56790 ( .A(reg_oi_2[19]), .B(n33644), .X(n28360) );
  nand_x1_sg U56791 ( .A(n33366), .B(\filter_0/n7871 ), .X(n28361) );
  nand_x1_sg U56792 ( .A(reg_oi_1[0]), .B(n33687), .X(n28276) );
  nand_x1_sg U56793 ( .A(reg_oi_1[1]), .B(n33691), .X(n28280) );
  nand_x1_sg U56794 ( .A(reg_oi_1[2]), .B(n33687), .X(n28282) );
  nand_x1_sg U56795 ( .A(reg_oi_1[3]), .B(n33692), .X(n28284) );
  nand_x1_sg U56796 ( .A(reg_oi_1[4]), .B(n33693), .X(n28286) );
  nand_x1_sg U56797 ( .A(reg_oi_1[5]), .B(n33691), .X(n28288) );
  nand_x1_sg U56798 ( .A(reg_oi_1[6]), .B(n33688), .X(n28290) );
  nand_x1_sg U56799 ( .A(n33353), .B(\filter_0/n7864 ), .X(n28291) );
  nand_x1_sg U56800 ( .A(reg_oi_1[7]), .B(n33688), .X(n28292) );
  nand_x1_sg U56801 ( .A(n33351), .B(\filter_0/n7863 ), .X(n28293) );
  nand_x1_sg U56802 ( .A(reg_oi_1[8]), .B(n33692), .X(n28294) );
  nand_x1_sg U56803 ( .A(n33351), .B(\filter_0/n7862 ), .X(n28295) );
  nand_x1_sg U56804 ( .A(reg_oi_1[9]), .B(n33687), .X(n28296) );
  nand_x1_sg U56805 ( .A(n29939), .B(\filter_0/n7861 ), .X(n28297) );
  nand_x1_sg U56806 ( .A(reg_oi_1[10]), .B(n33688), .X(n28298) );
  nand_x1_sg U56807 ( .A(n33350), .B(\filter_0/n7860 ), .X(n28299) );
  nand_x1_sg U56808 ( .A(reg_oi_1[11]), .B(n33687), .X(n28300) );
  nand_x1_sg U56809 ( .A(n33350), .B(\filter_0/n7859 ), .X(n28301) );
  nand_x1_sg U56810 ( .A(reg_oi_1[12]), .B(n33693), .X(n28302) );
  nand_x1_sg U56811 ( .A(n33352), .B(\filter_0/n7858 ), .X(n28303) );
  nand_x1_sg U56812 ( .A(reg_oi_1[13]), .B(n33688), .X(n28304) );
  nand_x1_sg U56813 ( .A(n33353), .B(\filter_0/n7857 ), .X(n28305) );
  nand_x1_sg U56814 ( .A(reg_oi_1[14]), .B(n33692), .X(n28306) );
  nand_x1_sg U56815 ( .A(n33352), .B(\filter_0/n7856 ), .X(n28307) );
  nand_x1_sg U56816 ( .A(reg_oi_1[15]), .B(n33693), .X(n28308) );
  nand_x1_sg U56817 ( .A(n33353), .B(\filter_0/n7855 ), .X(n28309) );
  nand_x1_sg U56818 ( .A(reg_oi_1[16]), .B(n33692), .X(n28310) );
  nand_x1_sg U56819 ( .A(n29939), .B(\filter_0/n7854 ), .X(n28311) );
  nand_x1_sg U56820 ( .A(reg_oi_1[17]), .B(n33691), .X(n28312) );
  nand_x1_sg U56821 ( .A(n33352), .B(\filter_0/n7853 ), .X(n28313) );
  nand_x1_sg U56822 ( .A(reg_oi_1[18]), .B(n33693), .X(n28314) );
  nand_x1_sg U56823 ( .A(n33351), .B(\filter_0/n7852 ), .X(n28315) );
  nand_x1_sg U56824 ( .A(reg_oi_1[19]), .B(n33691), .X(n28316) );
  nand_x1_sg U56825 ( .A(n33353), .B(\filter_0/n7851 ), .X(n28317) );
  nand_x1_sg U56826 ( .A(reg_oi_6[0]), .B(n33786), .X(n28492) );
  nand_x1_sg U56827 ( .A(reg_oi_6[1]), .B(n33781), .X(n28496) );
  nand_x1_sg U56828 ( .A(reg_oi_6[2]), .B(n33781), .X(n28498) );
  nand_x1_sg U56829 ( .A(reg_oi_6[3]), .B(n33780), .X(n28500) );
  nand_x1_sg U56830 ( .A(reg_oi_6[4]), .B(n33784), .X(n28502) );
  nand_x1_sg U56831 ( .A(reg_oi_6[5]), .B(n33780), .X(n28504) );
  nand_x1_sg U56832 ( .A(reg_oi_6[6]), .B(n33784), .X(n28506) );
  nand_x1_sg U56833 ( .A(n33470), .B(\filter_0/n7804 ), .X(n28507) );
  nand_x1_sg U56834 ( .A(reg_oi_6[7]), .B(n33785), .X(n28508) );
  nand_x1_sg U56835 ( .A(n33470), .B(\filter_0/n7803 ), .X(n28509) );
  nand_x1_sg U56836 ( .A(reg_oi_6[8]), .B(n33784), .X(n28510) );
  nand_x1_sg U56837 ( .A(n33472), .B(\filter_0/n7802 ), .X(n28511) );
  nand_x1_sg U56838 ( .A(reg_oi_6[9]), .B(n33781), .X(n28512) );
  nand_x1_sg U56839 ( .A(n33471), .B(\filter_0/n7801 ), .X(n28513) );
  nand_x1_sg U56840 ( .A(reg_oi_6[10]), .B(n33785), .X(n28514) );
  nand_x1_sg U56841 ( .A(n33472), .B(\filter_0/n7800 ), .X(n28515) );
  nand_x1_sg U56842 ( .A(reg_oi_6[11]), .B(n33786), .X(n28516) );
  nand_x1_sg U56843 ( .A(n33473), .B(\filter_0/n7799 ), .X(n28517) );
  nand_x1_sg U56844 ( .A(reg_oi_6[12]), .B(n33784), .X(n28518) );
  nand_x1_sg U56845 ( .A(n33473), .B(\filter_0/n7798 ), .X(n28519) );
  nand_x1_sg U56846 ( .A(reg_oi_6[13]), .B(n33785), .X(n28520) );
  nand_x1_sg U56847 ( .A(n33471), .B(\filter_0/n7797 ), .X(n28521) );
  nand_x1_sg U56848 ( .A(reg_oi_6[14]), .B(n33780), .X(n28522) );
  nand_x1_sg U56849 ( .A(n33471), .B(\filter_0/n7796 ), .X(n28523) );
  nand_x1_sg U56850 ( .A(reg_oi_6[15]), .B(n33786), .X(n28524) );
  nand_x1_sg U56851 ( .A(n29987), .B(\filter_0/n7795 ), .X(n28525) );
  nand_x1_sg U56852 ( .A(reg_oi_6[16]), .B(n33785), .X(n28526) );
  nand_x1_sg U56853 ( .A(n29987), .B(\filter_0/n7794 ), .X(n28527) );
  nand_x1_sg U56854 ( .A(reg_oi_6[17]), .B(n33781), .X(n28528) );
  nand_x1_sg U56855 ( .A(n33470), .B(\filter_0/n7793 ), .X(n28529) );
  nand_x1_sg U56856 ( .A(reg_oi_6[18]), .B(n33786), .X(n28530) );
  nand_x1_sg U56857 ( .A(n33472), .B(\filter_0/n7792 ), .X(n28531) );
  nand_x1_sg U56858 ( .A(reg_oi_6[19]), .B(n33780), .X(n28532) );
  nand_x1_sg U56859 ( .A(n33473), .B(\filter_0/n7791 ), .X(n28533) );
  nand_x1_sg U56860 ( .A(reg_oi_5[0]), .B(n33794), .X(n28450) );
  nand_x1_sg U56861 ( .A(reg_oi_5[1]), .B(n33793), .X(n28454) );
  nand_x1_sg U56862 ( .A(reg_oi_5[2]), .B(n33793), .X(n28456) );
  nand_x1_sg U56863 ( .A(reg_oi_5[3]), .B(n33792), .X(n28458) );
  nand_x1_sg U56864 ( .A(reg_oi_5[4]), .B(n33794), .X(n28460) );
  nand_x1_sg U56865 ( .A(reg_oi_5[5]), .B(n33788), .X(n28462) );
  nand_x1_sg U56866 ( .A(reg_oi_5[6]), .B(n33794), .X(n28464) );
  nand_x1_sg U56867 ( .A(n29937), .B(\filter_0/n7784 ), .X(n28465) );
  nand_x1_sg U56868 ( .A(reg_oi_5[7]), .B(n33788), .X(n28466) );
  nand_x1_sg U56869 ( .A(n29937), .B(\filter_0/n7783 ), .X(n28467) );
  nand_x1_sg U56870 ( .A(reg_oi_5[8]), .B(n33792), .X(n28468) );
  nand_x1_sg U56871 ( .A(n33347), .B(\filter_0/n7782 ), .X(n28469) );
  nand_x1_sg U56872 ( .A(reg_oi_5[9]), .B(n33794), .X(n28470) );
  nand_x1_sg U56873 ( .A(n33345), .B(\filter_0/n7781 ), .X(n28471) );
  nand_x1_sg U56874 ( .A(reg_oi_5[10]), .B(n33793), .X(n28472) );
  nand_x1_sg U56875 ( .A(n33345), .B(\filter_0/n7780 ), .X(n28473) );
  nand_x1_sg U56876 ( .A(reg_oi_5[11]), .B(n33788), .X(n28474) );
  nand_x1_sg U56877 ( .A(n33345), .B(\filter_0/n7779 ), .X(n28475) );
  nand_x1_sg U56878 ( .A(reg_oi_5[12]), .B(n33793), .X(n28476) );
  nand_x1_sg U56879 ( .A(n33347), .B(\filter_0/n7778 ), .X(n28477) );
  nand_x1_sg U56880 ( .A(reg_oi_5[13]), .B(n33789), .X(n28478) );
  nand_x1_sg U56881 ( .A(n33346), .B(\filter_0/n7777 ), .X(n28479) );
  nand_x1_sg U56882 ( .A(reg_oi_5[14]), .B(n33788), .X(n28480) );
  nand_x1_sg U56883 ( .A(n33348), .B(\filter_0/n7776 ), .X(n28481) );
  nand_x1_sg U56884 ( .A(reg_oi_5[15]), .B(n33789), .X(n28482) );
  nand_x1_sg U56885 ( .A(n33345), .B(\filter_0/n7775 ), .X(n28483) );
  nand_x1_sg U56886 ( .A(reg_oi_5[16]), .B(n33789), .X(n28484) );
  nand_x1_sg U56887 ( .A(n29937), .B(\filter_0/n7774 ), .X(n28485) );
  nand_x1_sg U56888 ( .A(reg_oi_5[17]), .B(n33792), .X(n28486) );
  nand_x1_sg U56889 ( .A(n33348), .B(\filter_0/n7773 ), .X(n28487) );
  nand_x1_sg U56890 ( .A(reg_oi_5[18]), .B(n33789), .X(n28488) );
  nand_x1_sg U56891 ( .A(n33347), .B(\filter_0/n7772 ), .X(n28489) );
  nand_x1_sg U56892 ( .A(reg_oi_5[19]), .B(n33792), .X(n28490) );
  nand_x1_sg U56893 ( .A(n33346), .B(\filter_0/n7771 ), .X(n28491) );
  nand_x1_sg U56894 ( .A(reg_oi_14[0]), .B(n33651), .X(n28619) );
  nand_x1_sg U56895 ( .A(reg_oi_14[1]), .B(n33648), .X(n28623) );
  nand_x1_sg U56896 ( .A(reg_oi_14[2]), .B(n33653), .X(n28625) );
  nand_x1_sg U56897 ( .A(reg_oi_14[3]), .B(n33652), .X(n28627) );
  nand_x1_sg U56898 ( .A(reg_oi_14[4]), .B(n33648), .X(n28629) );
  nand_x1_sg U56899 ( .A(reg_oi_14[5]), .B(n33651), .X(n28631) );
  nand_x1_sg U56900 ( .A(reg_oi_14[6]), .B(n33653), .X(n28633) );
  nand_x1_sg U56901 ( .A(n33362), .B(\filter_0/n7744 ), .X(n28634) );
  nand_x1_sg U56902 ( .A(reg_oi_14[7]), .B(n33647), .X(n28635) );
  nand_x1_sg U56903 ( .A(n33363), .B(\filter_0/n7743 ), .X(n28636) );
  nand_x1_sg U56904 ( .A(reg_oi_14[8]), .B(n33653), .X(n28637) );
  nand_x1_sg U56905 ( .A(n29943), .B(\filter_0/n7742 ), .X(n28638) );
  nand_x1_sg U56906 ( .A(reg_oi_14[9]), .B(n33651), .X(n28639) );
  nand_x1_sg U56907 ( .A(n33361), .B(\filter_0/n7741 ), .X(n28640) );
  nand_x1_sg U56908 ( .A(reg_oi_14[10]), .B(n33653), .X(n28641) );
  nand_x1_sg U56909 ( .A(n33360), .B(\filter_0/n7740 ), .X(n28642) );
  nand_x1_sg U56910 ( .A(reg_oi_14[11]), .B(n33648), .X(n28643) );
  nand_x1_sg U56911 ( .A(n33360), .B(\filter_0/n7739 ), .X(n28644) );
  nand_x1_sg U56912 ( .A(reg_oi_14[12]), .B(n33647), .X(n28645) );
  nand_x1_sg U56913 ( .A(n33363), .B(\filter_0/n7738 ), .X(n28646) );
  nand_x1_sg U56914 ( .A(reg_oi_14[13]), .B(n33652), .X(n28647) );
  nand_x1_sg U56915 ( .A(n29943), .B(\filter_0/n7737 ), .X(n28648) );
  nand_x1_sg U56916 ( .A(reg_oi_14[14]), .B(n33652), .X(n28649) );
  nand_x1_sg U56917 ( .A(n33363), .B(\filter_0/n7736 ), .X(n28650) );
  nand_x1_sg U56918 ( .A(reg_oi_14[15]), .B(n33648), .X(n28651) );
  nand_x1_sg U56919 ( .A(n33360), .B(\filter_0/n7735 ), .X(n28652) );
  nand_x1_sg U56920 ( .A(reg_oi_14[16]), .B(n33652), .X(n28653) );
  nand_x1_sg U56921 ( .A(n33362), .B(\filter_0/n7734 ), .X(n28654) );
  nand_x1_sg U56922 ( .A(reg_oi_14[17]), .B(n33647), .X(n28655) );
  nand_x1_sg U56923 ( .A(n33363), .B(\filter_0/n7733 ), .X(n28656) );
  nand_x1_sg U56924 ( .A(reg_oi_14[18]), .B(n33651), .X(n28657) );
  nand_x1_sg U56925 ( .A(n33361), .B(\filter_0/n7732 ), .X(n28658) );
  nand_x1_sg U56926 ( .A(reg_oi_14[19]), .B(n33647), .X(n28659) );
  nand_x1_sg U56927 ( .A(n33360), .B(\filter_0/n7731 ), .X(n28660) );
  nand_x1_sg U56928 ( .A(reg_oi_13[0]), .B(n33547), .X(n28661) );
  nand_x1_sg U56929 ( .A(reg_oi_13[1]), .B(n33548), .X(n28665) );
  nand_x1_sg U56930 ( .A(reg_oi_13[2]), .B(n33544), .X(n28667) );
  nand_x1_sg U56931 ( .A(reg_oi_13[3]), .B(n33544), .X(n28669) );
  nand_x1_sg U56932 ( .A(reg_oi_13[4]), .B(n33548), .X(n28671) );
  nand_x1_sg U56933 ( .A(reg_oi_13[5]), .B(n33543), .X(n28673) );
  nand_x1_sg U56934 ( .A(reg_oi_13[6]), .B(n33549), .X(n28675) );
  nand_x1_sg U56935 ( .A(n33343), .B(\filter_0/n7724 ), .X(n28676) );
  nand_x1_sg U56936 ( .A(reg_oi_13[7]), .B(n33543), .X(n28677) );
  nand_x1_sg U56937 ( .A(n29935), .B(\filter_0/n7723 ), .X(n28678) );
  nand_x1_sg U56938 ( .A(reg_oi_13[8]), .B(n33547), .X(n28679) );
  nand_x1_sg U56939 ( .A(n29935), .B(\filter_0/n7722 ), .X(n28680) );
  nand_x1_sg U56940 ( .A(reg_oi_13[9]), .B(n33544), .X(n28681) );
  nand_x1_sg U56941 ( .A(n33342), .B(\filter_0/n7721 ), .X(n28682) );
  nand_x1_sg U56942 ( .A(reg_oi_13[10]), .B(n33543), .X(n28683) );
  nand_x1_sg U56943 ( .A(n29935), .B(\filter_0/n7720 ), .X(n28684) );
  nand_x1_sg U56944 ( .A(reg_oi_13[11]), .B(n33549), .X(n28685) );
  nand_x1_sg U56945 ( .A(n33342), .B(\filter_0/n7719 ), .X(n28686) );
  nand_x1_sg U56946 ( .A(reg_oi_13[12]), .B(n33547), .X(n28687) );
  nand_x1_sg U56947 ( .A(n33340), .B(\filter_0/n7718 ), .X(n28688) );
  nand_x1_sg U56948 ( .A(reg_oi_13[13]), .B(n33548), .X(n28689) );
  nand_x1_sg U56949 ( .A(n33343), .B(\filter_0/n7717 ), .X(n28690) );
  nand_x1_sg U56950 ( .A(reg_oi_13[14]), .B(n33544), .X(n28691) );
  nand_x1_sg U56951 ( .A(n33340), .B(\filter_0/n7716 ), .X(n28692) );
  nand_x1_sg U56952 ( .A(reg_oi_13[15]), .B(n33549), .X(n28693) );
  nand_x1_sg U56953 ( .A(n33341), .B(\filter_0/n7715 ), .X(n28694) );
  nand_x1_sg U56954 ( .A(reg_oi_13[16]), .B(n33543), .X(n28695) );
  nand_x1_sg U56955 ( .A(n33340), .B(\filter_0/n7714 ), .X(n28696) );
  nand_x1_sg U56956 ( .A(reg_oi_13[17]), .B(n33547), .X(n28697) );
  nand_x1_sg U56957 ( .A(n33343), .B(\filter_0/n7713 ), .X(n28698) );
  nand_x1_sg U56958 ( .A(reg_oi_13[18]), .B(n33549), .X(n28699) );
  nand_x1_sg U56959 ( .A(n33342), .B(\filter_0/n7712 ), .X(n28700) );
  nand_x1_sg U56960 ( .A(reg_oi_13[19]), .B(n33548), .X(n28701) );
  nand_x1_sg U56961 ( .A(n33341), .B(\filter_0/n7711 ), .X(n28702) );
  nand_x1_sg U56962 ( .A(reg_oi_10[0]), .B(n33668), .X(n28791) );
  nand_x1_sg U56963 ( .A(reg_oi_10[1]), .B(n33663), .X(n28795) );
  nand_x1_sg U56964 ( .A(reg_oi_10[2]), .B(n33669), .X(n28797) );
  nand_x1_sg U56965 ( .A(reg_oi_10[3]), .B(n33668), .X(n28799) );
  nand_x1_sg U56966 ( .A(reg_oi_10[4]), .B(n33667), .X(n28801) );
  nand_x1_sg U56967 ( .A(reg_oi_10[5]), .B(n33663), .X(n28803) );
  nand_x1_sg U56968 ( .A(reg_oi_10[6]), .B(n33664), .X(n28805) );
  nand_x1_sg U56969 ( .A(n33356), .B(\filter_0/n7644 ), .X(n28806) );
  nand_x1_sg U56970 ( .A(reg_oi_10[7]), .B(n33664), .X(n28807) );
  nand_x1_sg U56971 ( .A(n33356), .B(\filter_0/n7643 ), .X(n28808) );
  nand_x1_sg U56972 ( .A(reg_oi_10[8]), .B(n33669), .X(n28809) );
  nand_x1_sg U56973 ( .A(n33358), .B(\filter_0/n7642 ), .X(n28810) );
  nand_x1_sg U56974 ( .A(reg_oi_10[9]), .B(n33663), .X(n28811) );
  nand_x1_sg U56975 ( .A(n33356), .B(\filter_0/n7641 ), .X(n28812) );
  nand_x1_sg U56976 ( .A(reg_oi_10[10]), .B(n33667), .X(n28813) );
  nand_x1_sg U56977 ( .A(n29941), .B(\filter_0/n7640 ), .X(n28814) );
  nand_x1_sg U56978 ( .A(reg_oi_10[11]), .B(n33664), .X(n28815) );
  nand_x1_sg U56979 ( .A(n33357), .B(\filter_0/n7639 ), .X(n28816) );
  nand_x1_sg U56980 ( .A(reg_oi_10[12]), .B(n33668), .X(n28817) );
  nand_x1_sg U56981 ( .A(n29941), .B(\filter_0/n7638 ), .X(n28818) );
  nand_x1_sg U56982 ( .A(reg_oi_10[13]), .B(n33668), .X(n28819) );
  nand_x1_sg U56983 ( .A(n29941), .B(\filter_0/n7637 ), .X(n28820) );
  nand_x1_sg U56984 ( .A(reg_oi_10[14]), .B(n33667), .X(n28821) );
  nand_x1_sg U56985 ( .A(n33358), .B(\filter_0/n7636 ), .X(n28822) );
  nand_x1_sg U56986 ( .A(reg_oi_10[15]), .B(n33664), .X(n28823) );
  nand_x1_sg U56987 ( .A(n33355), .B(\filter_0/n7635 ), .X(n28824) );
  nand_x1_sg U56988 ( .A(reg_oi_10[16]), .B(n33669), .X(n28825) );
  nand_x1_sg U56989 ( .A(n33358), .B(\filter_0/n7634 ), .X(n28826) );
  nand_x1_sg U56990 ( .A(reg_oi_10[17]), .B(n33663), .X(n28827) );
  nand_x1_sg U56991 ( .A(n33355), .B(\filter_0/n7633 ), .X(n28828) );
  nand_x1_sg U56992 ( .A(reg_oi_10[18]), .B(n33667), .X(n28829) );
  nand_x1_sg U56993 ( .A(n33357), .B(\filter_0/n7632 ), .X(n28830) );
  nand_x1_sg U56994 ( .A(reg_oi_10[19]), .B(n33669), .X(n28831) );
  nand_x1_sg U56995 ( .A(n33355), .B(\filter_0/n7631 ), .X(n28832) );
  nand_x1_sg U56996 ( .A(reg_oi_9[0]), .B(n33552), .X(n28835) );
  nand_x1_sg U56997 ( .A(reg_oi_9[1]), .B(n33556), .X(n28839) );
  nand_x1_sg U56998 ( .A(reg_oi_9[2]), .B(n33557), .X(n28841) );
  nand_x1_sg U56999 ( .A(reg_oi_9[3]), .B(n33551), .X(n28843) );
  nand_x1_sg U57000 ( .A(reg_oi_9[4]), .B(n33551), .X(n28845) );
  nand_x1_sg U57001 ( .A(reg_oi_9[5]), .B(n33555), .X(n28847) );
  nand_x1_sg U57002 ( .A(reg_oi_9[6]), .B(n33552), .X(n28849) );
  nand_x1_sg U57003 ( .A(n33338), .B(\filter_0/n7624 ), .X(n28850) );
  nand_x1_sg U57004 ( .A(reg_oi_9[7]), .B(n33552), .X(n28851) );
  nand_x1_sg U57005 ( .A(n29933), .B(\filter_0/n7623 ), .X(n28852) );
  nand_x1_sg U57006 ( .A(reg_oi_9[8]), .B(n33555), .X(n28853) );
  nand_x1_sg U57007 ( .A(n33337), .B(\filter_0/n7622 ), .X(n28854) );
  nand_x1_sg U57008 ( .A(reg_oi_9[9]), .B(n33555), .X(n28855) );
  nand_x1_sg U57009 ( .A(n33335), .B(\filter_0/n7621 ), .X(n28856) );
  nand_x1_sg U57010 ( .A(reg_oi_9[10]), .B(n33551), .X(n28857) );
  nand_x1_sg U57011 ( .A(n33337), .B(\filter_0/n7620 ), .X(n28858) );
  nand_x1_sg U57012 ( .A(reg_oi_9[11]), .B(n33557), .X(n28859) );
  nand_x1_sg U57013 ( .A(n33337), .B(\filter_0/n7619 ), .X(n28860) );
  nand_x1_sg U57014 ( .A(reg_oi_9[12]), .B(n33556), .X(n28861) );
  nand_x1_sg U57015 ( .A(n33336), .B(\filter_0/n7618 ), .X(n28862) );
  nand_x1_sg U57016 ( .A(reg_oi_9[13]), .B(n33556), .X(n28863) );
  nand_x1_sg U57017 ( .A(n33335), .B(\filter_0/n7617 ), .X(n28864) );
  nand_x1_sg U57018 ( .A(reg_oi_9[14]), .B(n33556), .X(n28865) );
  nand_x1_sg U57019 ( .A(n29933), .B(\filter_0/n7616 ), .X(n28866) );
  nand_x1_sg U57020 ( .A(reg_oi_9[15]), .B(n33552), .X(n28867) );
  nand_x1_sg U57021 ( .A(n33335), .B(\filter_0/n7615 ), .X(n28868) );
  nand_x1_sg U57022 ( .A(reg_oi_9[16]), .B(n33557), .X(n28869) );
  nand_x1_sg U57023 ( .A(n33336), .B(\filter_0/n7614 ), .X(n28870) );
  nand_x1_sg U57024 ( .A(reg_oi_9[17]), .B(n33551), .X(n28871) );
  nand_x1_sg U57025 ( .A(n33335), .B(\filter_0/n7613 ), .X(n28872) );
  nand_x1_sg U57026 ( .A(reg_oi_9[18]), .B(n33555), .X(n28873) );
  nand_x1_sg U57027 ( .A(n33338), .B(\filter_0/n7612 ), .X(n28874) );
  nand_x1_sg U57028 ( .A(reg_oi_9[19]), .B(n33557), .X(n28875) );
  nand_x1_sg U57029 ( .A(n33338), .B(\filter_0/n7611 ), .X(n28876) );
  nand_x1_sg U57030 ( .A(reg_ow_12[1]), .B(n33540), .X(n29406) );
  nand_x1_sg U57031 ( .A(reg_ow_12[3]), .B(n33541), .X(n29410) );
  nand_x1_sg U57032 ( .A(reg_ow_12[5]), .B(n33535), .X(n29414) );
  nand_x1_sg U57033 ( .A(reg_ow_12[7]), .B(n33539), .X(n29418) );
  nand_x1_sg U57034 ( .A(n33332), .B(\filter_0/n8032 ), .X(n29419) );
  nand_x1_sg U57035 ( .A(reg_ow_12[9]), .B(n33541), .X(n29422) );
  nand_x1_sg U57036 ( .A(n33331), .B(\filter_0/n8030 ), .X(n29423) );
  nand_x1_sg U57037 ( .A(reg_ow_12[11]), .B(n33541), .X(n29426) );
  nand_x1_sg U57038 ( .A(n29931), .B(\filter_0/n8028 ), .X(n29427) );
  nand_x1_sg U57039 ( .A(reg_ow_12[13]), .B(n33535), .X(n29430) );
  nand_x1_sg U57040 ( .A(n29931), .B(\filter_0/n8026 ), .X(n29431) );
  nand_x1_sg U57041 ( .A(reg_ow_12[15]), .B(n33541), .X(n29434) );
  nand_x1_sg U57042 ( .A(n33332), .B(\filter_0/n8024 ), .X(n29435) );
  nand_x1_sg U57043 ( .A(reg_ow_12[17]), .B(n33536), .X(n29438) );
  nand_x1_sg U57044 ( .A(n33333), .B(\filter_0/n8022 ), .X(n29439) );
  nand_x1_sg U57045 ( .A(reg_ow_12[19]), .B(n33540), .X(n29442) );
  nand_x1_sg U57046 ( .A(n33330), .B(\filter_0/n8020 ), .X(n29443) );
  nand_x1_sg U57047 ( .A(reg_ow_8[1]), .B(n33700), .X(n29582) );
  nand_x1_sg U57048 ( .A(reg_ow_8[3]), .B(n33700), .X(n29586) );
  nand_x1_sg U57049 ( .A(reg_ow_8[5]), .B(n33701), .X(n29590) );
  nand_x1_sg U57050 ( .A(reg_ow_8[7]), .B(n33695), .X(n29594) );
  nand_x1_sg U57051 ( .A(n33328), .B(\filter_0/n7932 ), .X(n29595) );
  nand_x1_sg U57052 ( .A(reg_ow_8[9]), .B(n33696), .X(n29598) );
  nand_x1_sg U57053 ( .A(n33326), .B(\filter_0/n7930 ), .X(n29599) );
  nand_x1_sg U57054 ( .A(reg_ow_8[11]), .B(n33700), .X(n29602) );
  nand_x1_sg U57055 ( .A(n33325), .B(\filter_0/n7928 ), .X(n29603) );
  nand_x1_sg U57056 ( .A(reg_ow_8[13]), .B(n33700), .X(n29606) );
  nand_x1_sg U57057 ( .A(n33326), .B(\filter_0/n7926 ), .X(n29607) );
  nand_x1_sg U57058 ( .A(reg_ow_8[15]), .B(n33695), .X(n29610) );
  nand_x1_sg U57059 ( .A(n33325), .B(\filter_0/n7924 ), .X(n29611) );
  nand_x1_sg U57060 ( .A(reg_ow_8[17]), .B(n33695), .X(n29614) );
  nand_x1_sg U57061 ( .A(n33328), .B(\filter_0/n7922 ), .X(n29615) );
  nand_x1_sg U57062 ( .A(reg_ow_8[19]), .B(n33699), .X(n29618) );
  nand_x1_sg U57063 ( .A(n33327), .B(\filter_0/n7920 ), .X(n29619) );
  nand_x1_sg U57064 ( .A(reg_oi_12[1]), .B(n33683), .X(n28707) );
  nand_x1_sg U57065 ( .A(reg_oi_12[3]), .B(n33679), .X(n28711) );
  nand_x1_sg U57066 ( .A(reg_oi_12[5]), .B(n33685), .X(n28715) );
  nand_x1_sg U57067 ( .A(reg_oi_12[7]), .B(n33679), .X(n28719) );
  nand_x1_sg U57068 ( .A(n33372), .B(\filter_0/n7703 ), .X(n28720) );
  nand_x1_sg U57069 ( .A(reg_oi_12[9]), .B(n33684), .X(n28723) );
  nand_x1_sg U57070 ( .A(n33373), .B(\filter_0/n7701 ), .X(n28724) );
  nand_x1_sg U57071 ( .A(reg_oi_12[11]), .B(n33679), .X(n28727) );
  nand_x1_sg U57072 ( .A(n29947), .B(\filter_0/n7699 ), .X(n28728) );
  nand_x1_sg U57073 ( .A(reg_oi_12[13]), .B(n33680), .X(n28731) );
  nand_x1_sg U57074 ( .A(n33370), .B(\filter_0/n7697 ), .X(n28732) );
  nand_x1_sg U57075 ( .A(reg_oi_12[15]), .B(n33683), .X(n28735) );
  nand_x1_sg U57076 ( .A(n33371), .B(\filter_0/n7695 ), .X(n28736) );
  nand_x1_sg U57077 ( .A(reg_oi_12[17]), .B(n33683), .X(n28739) );
  nand_x1_sg U57078 ( .A(n33371), .B(\filter_0/n7693 ), .X(n28740) );
  nand_x1_sg U57079 ( .A(reg_oi_12[19]), .B(n33684), .X(n28743) );
  nand_x1_sg U57080 ( .A(n33370), .B(\filter_0/n7691 ), .X(n28744) );
  nand_x1_sg U57081 ( .A(reg_oi_8[1]), .B(n33532), .X(n28883) );
  nand_x1_sg U57082 ( .A(reg_oi_8[3]), .B(n33533), .X(n28887) );
  nand_x1_sg U57083 ( .A(reg_oi_8[5]), .B(n33531), .X(n28891) );
  nand_x1_sg U57084 ( .A(reg_oi_8[7]), .B(n33533), .X(n28895) );
  nand_x1_sg U57085 ( .A(n33321), .B(\filter_0/n7603 ), .X(n28896) );
  nand_x1_sg U57086 ( .A(reg_oi_8[9]), .B(n33527), .X(n28899) );
  nand_x1_sg U57087 ( .A(n33320), .B(\filter_0/n7601 ), .X(n28900) );
  nand_x1_sg U57088 ( .A(reg_oi_8[11]), .B(n33528), .X(n28903) );
  nand_x1_sg U57089 ( .A(n29927), .B(\filter_0/n7599 ), .X(n28904) );
  nand_x1_sg U57090 ( .A(reg_oi_8[13]), .B(n33533), .X(n28907) );
  nand_x1_sg U57091 ( .A(n33320), .B(\filter_0/n7597 ), .X(n28908) );
  nand_x1_sg U57092 ( .A(reg_oi_8[15]), .B(n33527), .X(n28911) );
  nand_x1_sg U57093 ( .A(n33323), .B(\filter_0/n7595 ), .X(n28912) );
  nand_x1_sg U57094 ( .A(reg_oi_8[17]), .B(n33532), .X(n28915) );
  nand_x1_sg U57095 ( .A(n33321), .B(\filter_0/n7593 ), .X(n28916) );
  nand_x1_sg U57096 ( .A(reg_oi_8[19]), .B(n33532), .X(n28919) );
  nand_x1_sg U57097 ( .A(n33322), .B(\filter_0/n7591 ), .X(n28920) );
  nand_x1_sg U57098 ( .A(reg_oi_7[0]), .B(n33765), .X(n28534) );
  nand_x1_sg U57099 ( .A(reg_oi_7[2]), .B(n33764), .X(n28540) );
  nand_x1_sg U57100 ( .A(reg_oi_7[4]), .B(n33768), .X(n28544) );
  nand_x1_sg U57101 ( .A(reg_oi_7[6]), .B(n33764), .X(n28548) );
  nand_x1_sg U57102 ( .A(n33430), .B(\filter_0/n7824 ), .X(n28549) );
  nand_x1_sg U57103 ( .A(reg_oi_7[8]), .B(n33765), .X(n28552) );
  nand_x1_sg U57104 ( .A(n29971), .B(\filter_0/n7822 ), .X(n28553) );
  nand_x1_sg U57105 ( .A(reg_oi_7[10]), .B(n33769), .X(n28556) );
  nand_x1_sg U57106 ( .A(n33433), .B(\filter_0/n7820 ), .X(n28557) );
  nand_x1_sg U57107 ( .A(reg_oi_7[12]), .B(n33769), .X(n28560) );
  nand_x1_sg U57108 ( .A(n33431), .B(\filter_0/n7818 ), .X(n28561) );
  nand_x1_sg U57109 ( .A(reg_oi_7[14]), .B(n33770), .X(n28564) );
  nand_x1_sg U57110 ( .A(n33433), .B(\filter_0/n7816 ), .X(n28565) );
  nand_x1_sg U57111 ( .A(reg_oi_7[16]), .B(n33765), .X(n28568) );
  nand_x1_sg U57112 ( .A(n33432), .B(\filter_0/n7814 ), .X(n28569) );
  nand_x1_sg U57113 ( .A(reg_oi_7[18]), .B(n33769), .X(n28572) );
  nand_x1_sg U57114 ( .A(n29971), .B(\filter_0/n7812 ), .X(n28573) );
  nand_x1_sg U57115 ( .A(reg_oi_7[1]), .B(n33764), .X(n28538) );
  nand_x1_sg U57116 ( .A(reg_oi_7[3]), .B(n33770), .X(n28542) );
  nand_x1_sg U57117 ( .A(reg_oi_7[5]), .B(n33770), .X(n28546) );
  nand_x1_sg U57118 ( .A(reg_oi_7[7]), .B(n33770), .X(n28550) );
  nand_x1_sg U57119 ( .A(n33432), .B(\filter_0/n7823 ), .X(n28551) );
  nand_x1_sg U57120 ( .A(reg_oi_7[9]), .B(n33765), .X(n28554) );
  nand_x1_sg U57121 ( .A(n29971), .B(\filter_0/n7821 ), .X(n28555) );
  nand_x1_sg U57122 ( .A(reg_oi_7[11]), .B(n33764), .X(n28558) );
  nand_x1_sg U57123 ( .A(n33430), .B(\filter_0/n7819 ), .X(n28559) );
  nand_x1_sg U57124 ( .A(reg_oi_7[13]), .B(n33768), .X(n28562) );
  nand_x1_sg U57125 ( .A(n33433), .B(\filter_0/n7817 ), .X(n28563) );
  nand_x1_sg U57126 ( .A(reg_oi_7[15]), .B(n33768), .X(n28566) );
  nand_x1_sg U57127 ( .A(n33433), .B(\filter_0/n7815 ), .X(n28567) );
  nand_x1_sg U57128 ( .A(reg_oi_7[17]), .B(n33769), .X(n28570) );
  nand_x1_sg U57129 ( .A(n33432), .B(\filter_0/n7813 ), .X(n28571) );
  nand_x1_sg U57130 ( .A(reg_oi_7[19]), .B(n33768), .X(n28574) );
  nand_x1_sg U57131 ( .A(n33431), .B(\filter_0/n7811 ), .X(n28575) );
  nand_x1_sg U57132 ( .A(n20925), .B(n32938), .X(n20924) );
  nor_x1_sg U57133 ( .A(n20926), .B(n20927), .X(n20925) );
  nor_x1_sg U57134 ( .A(n20928), .B(n31709), .X(n20926) );
  nor_x1_sg U57135 ( .A(\shifter_0/w_pointer[0] ), .B(n42543), .X(n20927) );
  nand_x1_sg U57136 ( .A(\shifter_0/w_pointer[1] ), .B(n20940), .X(n20936) );
  nand_x1_sg U57137 ( .A(n31597), .B(n21336), .X(n21348) );
  nor_x1_sg U57138 ( .A(n32940), .B(n21576), .X(n21564) );
  nor_x1_sg U57139 ( .A(\shifter_0/i_pointer[0] ), .B(n42539), .X(n21576) );
  nor_x1_sg U57140 ( .A(\shifter_0/w_pointer[0] ), .B(n42544), .X(n20929) );
  nor_x1_sg U57141 ( .A(n21470), .B(n21471), .X(n21469) );
  nor_x1_sg U57142 ( .A(n21356), .B(n31668), .X(n21471) );
  nor_x1_sg U57143 ( .A(\shifter_0/i_pointer[0] ), .B(n42540), .X(n21470) );
  nor_x1_sg U57144 ( .A(n32935), .B(n21389), .X(n21377) );
  nor_x1_sg U57145 ( .A(n31595), .B(n42541), .X(n21389) );
  nand_x1_sg U57146 ( .A(n32509), .B(n20987), .X(n20986) );
  nand_x1_sg U57147 ( .A(n20992), .B(n31599), .X(n20989) );
  nor_x1_sg U57148 ( .A(n20913), .B(n20914), .X(n20912) );
  nor_x1_sg U57149 ( .A(\shifter_0/w_pointer[0] ), .B(n20916), .X(n20913) );
  nor_x1_sg U57150 ( .A(n20915), .B(n31709), .X(n20914) );
  nand_x1_sg U57151 ( .A(n32510), .B(n21661), .X(n21660) );
  nand_x1_sg U57152 ( .A(n21666), .B(n31599), .X(n21663) );
  nor_x1_sg U57153 ( .A(n21657), .B(n21658), .X(n21656) );
  nor_x1_sg U57154 ( .A(\shifter_0/i_pointer[0] ), .B(n21367), .X(n21657) );
  nor_x1_sg U57155 ( .A(n21359), .B(n31669), .X(n21658) );
  nor_x1_sg U57156 ( .A(n22211), .B(n35551), .X(n22210) );
  nand_x1_sg U57157 ( .A(n30255), .B(output_taken), .X(n22211) );
  nand_x1_sg U57158 ( .A(n22214), .B(n22215), .X(n22212) );
  nand_x1_sg U57159 ( .A(n34105), .B(state[1]), .X(n22213) );
  nor_x1_sg U57160 ( .A(state[1]), .B(state[0]), .X(n23632) );
  nand_x1_sg U57161 ( .A(i_0[2]), .B(n31946), .X(n22226) );
  nand_x1_sg U57162 ( .A(reg_i_0[2]), .B(n34463), .X(n22225) );
  nand_x1_sg U57163 ( .A(i_0[5]), .B(n31972), .X(n22232) );
  nand_x1_sg U57164 ( .A(reg_i_0[5]), .B(n34926), .X(n22231) );
  nand_x1_sg U57165 ( .A(i_0[8]), .B(n34483), .X(n22238) );
  nand_x1_sg U57166 ( .A(reg_i_0[8]), .B(n31277), .X(n22237) );
  nand_x1_sg U57167 ( .A(i_0[11]), .B(n30830), .X(n22244) );
  nand_x1_sg U57168 ( .A(reg_i_0[11]), .B(n34819), .X(n22243) );
  nand_x1_sg U57169 ( .A(i_0[14]), .B(n31262), .X(n22250) );
  nand_x1_sg U57170 ( .A(reg_i_0[14]), .B(n32981), .X(n22249) );
  nand_x1_sg U57171 ( .A(i_0[17]), .B(n33255), .X(n22256) );
  nand_x1_sg U57172 ( .A(reg_i_0[17]), .B(n30815), .X(n22255) );
  nand_x1_sg U57173 ( .A(i_1[0]), .B(n32944), .X(n22262) );
  nand_x1_sg U57174 ( .A(reg_i_1[0]), .B(n31927), .X(n22261) );
  nand_x1_sg U57175 ( .A(i_1[3]), .B(n34833), .X(n22268) );
  nand_x1_sg U57176 ( .A(reg_i_1[3]), .B(n34926), .X(n22267) );
  nand_x1_sg U57177 ( .A(i_1[6]), .B(n33247), .X(n22274) );
  nand_x1_sg U57178 ( .A(reg_i_1[6]), .B(n34928), .X(n22273) );
  nand_x1_sg U57179 ( .A(i_1[9]), .B(n31934), .X(n22280) );
  nand_x1_sg U57180 ( .A(reg_i_1[9]), .B(n30191), .X(n22279) );
  nand_x1_sg U57181 ( .A(i_1[12]), .B(n30383), .X(n22286) );
  nand_x1_sg U57182 ( .A(reg_i_1[12]), .B(n34809), .X(n22285) );
  nand_x1_sg U57183 ( .A(i_1[15]), .B(n31263), .X(n22292) );
  nand_x1_sg U57184 ( .A(reg_i_1[15]), .B(n31006), .X(n22291) );
  nand_x1_sg U57185 ( .A(i_1[18]), .B(n34505), .X(n22298) );
  nand_x1_sg U57186 ( .A(reg_i_1[18]), .B(n31017), .X(n22297) );
  nand_x1_sg U57187 ( .A(i_2[1]), .B(n31970), .X(n22304) );
  nand_x1_sg U57188 ( .A(reg_i_2[1]), .B(n31960), .X(n22303) );
  nand_x1_sg U57189 ( .A(i_2[4]), .B(n30810), .X(n22310) );
  nand_x1_sg U57190 ( .A(reg_i_2[4]), .B(n31282), .X(n22309) );
  nand_x1_sg U57191 ( .A(i_2[7]), .B(n34839), .X(n22316) );
  nand_x1_sg U57192 ( .A(reg_i_2[7]), .B(n34931), .X(n22315) );
  nand_x1_sg U57193 ( .A(i_2[10]), .B(n30813), .X(n22322) );
  nand_x1_sg U57194 ( .A(reg_i_2[10]), .B(n31961), .X(n22321) );
  nand_x1_sg U57195 ( .A(i_2[13]), .B(n29881), .X(n22328) );
  nand_x1_sg U57196 ( .A(reg_i_2[13]), .B(n32981), .X(n22327) );
  nand_x1_sg U57197 ( .A(i_2[16]), .B(n34845), .X(n22334) );
  nand_x1_sg U57198 ( .A(reg_i_2[16]), .B(n32077), .X(n22333) );
  nand_x1_sg U57199 ( .A(i_2[19]), .B(n34476), .X(n22340) );
  nand_x1_sg U57200 ( .A(reg_i_2[19]), .B(n32971), .X(n22339) );
  nand_x1_sg U57201 ( .A(i_3[2]), .B(n31973), .X(n22346) );
  nand_x1_sg U57202 ( .A(reg_i_3[2]), .B(n33840), .X(n22345) );
  nand_x1_sg U57203 ( .A(i_3[5]), .B(n34451), .X(n22352) );
  nand_x1_sg U57204 ( .A(reg_i_3[5]), .B(n32075), .X(n22351) );
  nand_x1_sg U57205 ( .A(i_3[8]), .B(n34842), .X(n22358) );
  nand_x1_sg U57206 ( .A(reg_i_3[8]), .B(n32978), .X(n22357) );
  nand_x1_sg U57207 ( .A(i_3[11]), .B(n34455), .X(n22364) );
  nand_x1_sg U57208 ( .A(reg_i_3[11]), .B(n32949), .X(n22363) );
  nand_x1_sg U57209 ( .A(i_3[14]), .B(n34462), .X(n22370) );
  nand_x1_sg U57210 ( .A(reg_i_3[14]), .B(n32092), .X(n22369) );
  nand_x1_sg U57211 ( .A(i_3[17]), .B(n34490), .X(n22376) );
  nand_x1_sg U57212 ( .A(reg_i_3[17]), .B(n31286), .X(n22375) );
  nand_x1_sg U57213 ( .A(i_4[0]), .B(n34455), .X(n22382) );
  nand_x1_sg U57214 ( .A(reg_i_4[0]), .B(n31286), .X(n22381) );
  nand_x1_sg U57215 ( .A(i_4[3]), .B(n34452), .X(n22388) );
  nand_x1_sg U57216 ( .A(reg_i_4[3]), .B(n32087), .X(n22387) );
  nand_x1_sg U57217 ( .A(i_4[6]), .B(n33257), .X(n22394) );
  nand_x1_sg U57218 ( .A(reg_i_4[6]), .B(n34529), .X(n22393) );
  nand_x1_sg U57219 ( .A(i_4[9]), .B(n30384), .X(n22400) );
  nand_x1_sg U57220 ( .A(reg_i_4[9]), .B(n35058), .X(n22399) );
  nand_x1_sg U57221 ( .A(i_4[12]), .B(n34481), .X(n22406) );
  nand_x1_sg U57222 ( .A(reg_i_4[12]), .B(n32969), .X(n22405) );
  nand_x1_sg U57223 ( .A(i_4[15]), .B(n30385), .X(n22412) );
  nand_x1_sg U57224 ( .A(reg_i_4[15]), .B(n31291), .X(n22411) );
  nand_x1_sg U57225 ( .A(i_4[18]), .B(n31933), .X(n22418) );
  nand_x1_sg U57226 ( .A(reg_i_4[18]), .B(n31961), .X(n22417) );
  nand_x1_sg U57227 ( .A(i_5[1]), .B(n34917), .X(n22424) );
  nand_x1_sg U57228 ( .A(reg_i_5[1]), .B(n32076), .X(n22423) );
  nand_x1_sg U57229 ( .A(i_5[4]), .B(n31964), .X(n22430) );
  nand_x1_sg U57230 ( .A(reg_i_5[4]), .B(n34508), .X(n22429) );
  nand_x1_sg U57231 ( .A(i_5[7]), .B(n31257), .X(n22436) );
  nand_x1_sg U57232 ( .A(reg_i_5[7]), .B(n34818), .X(n22435) );
  nand_x1_sg U57233 ( .A(i_5[10]), .B(n33238), .X(n22442) );
  nand_x1_sg U57234 ( .A(reg_i_5[10]), .B(n31102), .X(n22441) );
  nand_x1_sg U57235 ( .A(i_5[13]), .B(n31266), .X(n22448) );
  nand_x1_sg U57236 ( .A(reg_i_5[13]), .B(n32963), .X(n22447) );
  nand_x1_sg U57237 ( .A(i_5[16]), .B(n32945), .X(n22454) );
  nand_x1_sg U57238 ( .A(reg_i_5[16]), .B(n34820), .X(n22453) );
  nand_x1_sg U57239 ( .A(i_5[19]), .B(n30826), .X(n22460) );
  nand_x1_sg U57240 ( .A(reg_i_5[19]), .B(n32973), .X(n22459) );
  nand_x1_sg U57241 ( .A(i_6[2]), .B(n31937), .X(n22466) );
  nand_x1_sg U57242 ( .A(reg_i_6[2]), .B(n34926), .X(n22465) );
  nand_x1_sg U57243 ( .A(i_6[5]), .B(n30615), .X(n22472) );
  nand_x1_sg U57244 ( .A(reg_i_6[5]), .B(n35060), .X(n22471) );
  nand_x1_sg U57245 ( .A(i_6[8]), .B(n34844), .X(n22478) );
  nand_x1_sg U57246 ( .A(reg_i_6[8]), .B(n32953), .X(n22477) );
  nand_x1_sg U57247 ( .A(i_6[11]), .B(n31100), .X(n22484) );
  nand_x1_sg U57248 ( .A(reg_i_6[11]), .B(n34469), .X(n22483) );
  nand_x1_sg U57249 ( .A(i_6[14]), .B(n34476), .X(n22490) );
  nand_x1_sg U57250 ( .A(reg_i_6[14]), .B(n34529), .X(n22489) );
  nand_x1_sg U57251 ( .A(i_6[17]), .B(n34503), .X(n22496) );
  nand_x1_sg U57252 ( .A(reg_i_6[17]), .B(n32981), .X(n22495) );
  nand_x1_sg U57253 ( .A(i_7[0]), .B(n33250), .X(n22502) );
  nand_x1_sg U57254 ( .A(reg_i_7[0]), .B(n31928), .X(n22501) );
  nand_x1_sg U57255 ( .A(i_7[3]), .B(n33246), .X(n22508) );
  nand_x1_sg U57256 ( .A(reg_i_7[3]), .B(n34811), .X(n22507) );
  nand_x1_sg U57257 ( .A(i_7[6]), .B(n31944), .X(n22514) );
  nand_x1_sg U57258 ( .A(reg_i_7[6]), .B(n31210), .X(n22513) );
  nand_x1_sg U57259 ( .A(i_7[9]), .B(n31966), .X(n22520) );
  nand_x1_sg U57260 ( .A(reg_i_7[9]), .B(n30368), .X(n22519) );
  nand_x1_sg U57261 ( .A(i_7[12]), .B(n31946), .X(n22526) );
  nand_x1_sg U57262 ( .A(reg_i_7[12]), .B(n32974), .X(n22525) );
  nand_x1_sg U57263 ( .A(i_7[15]), .B(n31267), .X(n22532) );
  nand_x1_sg U57264 ( .A(reg_i_7[15]), .B(n32970), .X(n22531) );
  nand_x1_sg U57265 ( .A(i_7[18]), .B(n30383), .X(n22538) );
  nand_x1_sg U57266 ( .A(reg_i_7[18]), .B(n29905), .X(n22537) );
  nand_x1_sg U57267 ( .A(i_8[1]), .B(n34922), .X(n22544) );
  nand_x1_sg U57268 ( .A(reg_i_8[1]), .B(n30378), .X(n22543) );
  nand_x1_sg U57269 ( .A(i_8[4]), .B(n31262), .X(n22550) );
  nand_x1_sg U57270 ( .A(reg_i_8[4]), .B(n32084), .X(n22549) );
  nand_x1_sg U57271 ( .A(i_8[7]), .B(n33253), .X(n22556) );
  nand_x1_sg U57272 ( .A(reg_i_8[7]), .B(n34524), .X(n22555) );
  nand_x1_sg U57273 ( .A(i_8[10]), .B(n34454), .X(n22562) );
  nand_x1_sg U57274 ( .A(reg_i_8[10]), .B(n32961), .X(n22561) );
  nand_x1_sg U57275 ( .A(i_8[13]), .B(n34935), .X(n22568) );
  nand_x1_sg U57276 ( .A(reg_i_8[13]), .B(n32968), .X(n22567) );
  nand_x1_sg U57277 ( .A(i_8[16]), .B(n34503), .X(n22574) );
  nand_x1_sg U57278 ( .A(reg_i_8[16]), .B(n32960), .X(n22573) );
  nand_x1_sg U57279 ( .A(i_8[19]), .B(n29687), .X(n22580) );
  nand_x1_sg U57280 ( .A(reg_i_8[19]), .B(n34915), .X(n22579) );
  nand_x1_sg U57281 ( .A(i_9[2]), .B(n34918), .X(n22586) );
  nand_x1_sg U57282 ( .A(reg_i_9[2]), .B(n32086), .X(n22585) );
  nand_x1_sg U57283 ( .A(i_9[5]), .B(n31967), .X(n22592) );
  nand_x1_sg U57284 ( .A(reg_i_9[5]), .B(n34527), .X(n22591) );
  nand_x1_sg U57285 ( .A(i_9[8]), .B(n31628), .X(n22598) );
  nand_x1_sg U57286 ( .A(reg_i_9[8]), .B(n34929), .X(n22597) );
  nand_x1_sg U57287 ( .A(i_9[11]), .B(n33245), .X(n22604) );
  nand_x1_sg U57288 ( .A(reg_i_9[11]), .B(n34924), .X(n22603) );
  nand_x1_sg U57289 ( .A(i_9[14]), .B(n33229), .X(n22610) );
  nand_x1_sg U57290 ( .A(reg_i_9[14]), .B(n29906), .X(n22609) );
  nand_x1_sg U57291 ( .A(i_9[17]), .B(n34476), .X(n22616) );
  nand_x1_sg U57292 ( .A(reg_i_9[17]), .B(n34930), .X(n22615) );
  nand_x1_sg U57293 ( .A(i_10[0]), .B(n32184), .X(n22622) );
  nand_x1_sg U57294 ( .A(reg_i_10[0]), .B(n30819), .X(n22621) );
  nand_x1_sg U57295 ( .A(i_10[3]), .B(n34919), .X(n22628) );
  nand_x1_sg U57296 ( .A(reg_i_10[3]), .B(n34511), .X(n22627) );
  nand_x1_sg U57297 ( .A(i_10[6]), .B(n30616), .X(n22634) );
  nand_x1_sg U57298 ( .A(reg_i_10[6]), .B(n34464), .X(n22633) );
  nand_x1_sg U57299 ( .A(i_10[9]), .B(n30193), .X(n22640) );
  nand_x1_sg U57300 ( .A(reg_i_10[9]), .B(n33261), .X(n22639) );
  nand_x1_sg U57301 ( .A(i_10[12]), .B(n34456), .X(n22646) );
  nand_x1_sg U57302 ( .A(reg_i_10[12]), .B(n34529), .X(n22645) );
  nand_x1_sg U57303 ( .A(i_10[15]), .B(n31258), .X(n22652) );
  nand_x1_sg U57304 ( .A(reg_i_10[15]), .B(n31626), .X(n22651) );
  nand_x1_sg U57305 ( .A(i_10[18]), .B(n30824), .X(n22658) );
  nand_x1_sg U57306 ( .A(reg_i_10[18]), .B(n33840), .X(n22657) );
  nand_x1_sg U57307 ( .A(i_11[1]), .B(n34506), .X(n22664) );
  nand_x1_sg U57308 ( .A(reg_i_11[1]), .B(n32074), .X(n22663) );
  nand_x1_sg U57309 ( .A(i_11[4]), .B(n32179), .X(n22670) );
  nand_x1_sg U57310 ( .A(reg_i_11[4]), .B(n32975), .X(n22669) );
  nand_x1_sg U57311 ( .A(i_11[7]), .B(n34830), .X(n22676) );
  nand_x1_sg U57312 ( .A(reg_i_11[7]), .B(n31237), .X(n22675) );
  nand_x1_sg U57313 ( .A(i_11[10]), .B(n33258), .X(n22682) );
  nand_x1_sg U57314 ( .A(reg_i_11[10]), .B(n30191), .X(n22681) );
  nand_x1_sg U57315 ( .A(i_11[13]), .B(n34491), .X(n22688) );
  nand_x1_sg U57316 ( .A(reg_i_11[13]), .B(n34511), .X(n22687) );
  nand_x1_sg U57317 ( .A(i_11[16]), .B(n31972), .X(n22694) );
  nand_x1_sg U57318 ( .A(reg_i_11[16]), .B(n32962), .X(n22693) );
  nand_x1_sg U57319 ( .A(i_11[19]), .B(n34843), .X(n22700) );
  nand_x1_sg U57320 ( .A(reg_i_11[19]), .B(n32956), .X(n22699) );
  nand_x1_sg U57321 ( .A(i_12[2]), .B(n30828), .X(n22706) );
  nand_x1_sg U57322 ( .A(reg_i_12[2]), .B(n34522), .X(n22705) );
  nand_x1_sg U57323 ( .A(i_12[5]), .B(n34462), .X(n22712) );
  nand_x1_sg U57324 ( .A(reg_i_12[5]), .B(n32949), .X(n22711) );
  nand_x1_sg U57325 ( .A(i_12[8]), .B(n30382), .X(n22718) );
  nand_x1_sg U57326 ( .A(reg_i_12[8]), .B(n29798), .X(n22717) );
  nand_x1_sg U57327 ( .A(i_12[11]), .B(n33244), .X(n22724) );
  nand_x1_sg U57328 ( .A(reg_i_12[11]), .B(n34464), .X(n22723) );
  nand_x1_sg U57329 ( .A(i_12[14]), .B(n33227), .X(n22730) );
  nand_x1_sg U57330 ( .A(reg_i_12[14]), .B(n32072), .X(n22729) );
  nand_x1_sg U57331 ( .A(i_12[17]), .B(n31262), .X(n22736) );
  nand_x1_sg U57332 ( .A(reg_i_12[17]), .B(n34528), .X(n22735) );
  nand_x1_sg U57333 ( .A(i_13[0]), .B(n33223), .X(n22742) );
  nand_x1_sg U57334 ( .A(reg_i_13[0]), .B(n34923), .X(n22741) );
  nand_x1_sg U57335 ( .A(i_13[3]), .B(n31966), .X(n22748) );
  nand_x1_sg U57336 ( .A(reg_i_13[3]), .B(n30373), .X(n22747) );
  nand_x1_sg U57337 ( .A(i_13[6]), .B(n31972), .X(n22754) );
  nand_x1_sg U57338 ( .A(reg_i_13[6]), .B(n33273), .X(n22753) );
  nand_x1_sg U57339 ( .A(i_13[9]), .B(n30811), .X(n22760) );
  nand_x1_sg U57340 ( .A(reg_i_13[9]), .B(n32980), .X(n22759) );
  nand_x1_sg U57341 ( .A(i_13[12]), .B(n34479), .X(n22766) );
  nand_x1_sg U57342 ( .A(reg_i_13[12]), .B(n31285), .X(n22765) );
  nand_x1_sg U57343 ( .A(i_13[15]), .B(n34484), .X(n22772) );
  nand_x1_sg U57344 ( .A(reg_i_13[15]), .B(n34525), .X(n22771) );
  nand_x1_sg U57345 ( .A(i_13[18]), .B(n31970), .X(n22778) );
  nand_x1_sg U57346 ( .A(reg_i_13[18]), .B(n32956), .X(n22777) );
  nand_x1_sg U57347 ( .A(i_14[1]), .B(n34462), .X(n22784) );
  nand_x1_sg U57348 ( .A(reg_i_14[1]), .B(n32076), .X(n22783) );
  nand_x1_sg U57349 ( .A(i_14[4]), .B(n33223), .X(n22790) );
  nand_x1_sg U57350 ( .A(reg_i_14[4]), .B(n30823), .X(n22789) );
  nand_x1_sg U57351 ( .A(i_14[7]), .B(n33227), .X(n22796) );
  nand_x1_sg U57352 ( .A(reg_i_14[7]), .B(n32087), .X(n22795) );
  nand_x1_sg U57353 ( .A(i_14[10]), .B(n33916), .X(n22802) );
  nand_x1_sg U57354 ( .A(reg_i_14[10]), .B(n32082), .X(n22801) );
  nand_x1_sg U57355 ( .A(i_14[13]), .B(n33915), .X(n22808) );
  nand_x1_sg U57356 ( .A(reg_i_14[13]), .B(n34524), .X(n22807) );
  nand_x1_sg U57357 ( .A(i_14[16]), .B(n34451), .X(n22814) );
  nand_x1_sg U57358 ( .A(reg_i_14[16]), .B(n33260), .X(n22813) );
  nand_x1_sg U57359 ( .A(i_14[19]), .B(n30385), .X(n22820) );
  nand_x1_sg U57360 ( .A(reg_i_14[19]), .B(n34811), .X(n22819) );
  nand_x1_sg U57361 ( .A(i_15[2]), .B(n31967), .X(n22826) );
  nand_x1_sg U57362 ( .A(reg_i_15[2]), .B(n32950), .X(n22825) );
  nand_x1_sg U57363 ( .A(i_15[5]), .B(n32182), .X(n22832) );
  nand_x1_sg U57364 ( .A(reg_i_15[5]), .B(n31625), .X(n22831) );
  nand_x1_sg U57365 ( .A(i_15[8]), .B(n34491), .X(n22838) );
  nand_x1_sg U57366 ( .A(reg_i_15[8]), .B(n34809), .X(n22837) );
  nand_x1_sg U57367 ( .A(i_15[11]), .B(n30828), .X(n22844) );
  nand_x1_sg U57368 ( .A(reg_i_15[11]), .B(n32088), .X(n22843) );
  nand_x1_sg U57369 ( .A(i_15[14]), .B(n29901), .X(n22850) );
  nand_x1_sg U57370 ( .A(reg_i_15[14]), .B(n33263), .X(n22849) );
  nand_x1_sg U57371 ( .A(i_15[17]), .B(n31100), .X(n22856) );
  nand_x1_sg U57372 ( .A(reg_i_15[17]), .B(n32968), .X(n22855) );
  nand_x1_sg U57373 ( .A(w_0[0]), .B(n33244), .X(n22862) );
  nand_x1_sg U57374 ( .A(reg_w_0[0]), .B(n30371), .X(n22861) );
  nand_x1_sg U57375 ( .A(w_0[3]), .B(n31973), .X(n22868) );
  nand_x1_sg U57376 ( .A(reg_w_0[3]), .B(n31927), .X(n22867) );
  nand_x1_sg U57377 ( .A(w_0[6]), .B(n34506), .X(n22874) );
  nand_x1_sg U57378 ( .A(reg_w_0[6]), .B(n34471), .X(n22873) );
  nand_x1_sg U57379 ( .A(w_0[9]), .B(n31946), .X(n22880) );
  nand_x1_sg U57380 ( .A(reg_w_0[9]), .B(n32969), .X(n22879) );
  nand_x1_sg U57381 ( .A(w_0[12]), .B(n34457), .X(n22886) );
  nand_x1_sg U57382 ( .A(reg_w_0[12]), .B(n31954), .X(n22885) );
  nand_x1_sg U57383 ( .A(w_0[15]), .B(n34835), .X(n22892) );
  nand_x1_sg U57384 ( .A(reg_w_0[15]), .B(n33840), .X(n22891) );
  nand_x1_sg U57385 ( .A(w_0[18]), .B(n31106), .X(n22898) );
  nand_x1_sg U57386 ( .A(reg_w_0[18]), .B(n31003), .X(n22897) );
  nand_x1_sg U57387 ( .A(w_1[1]), .B(n32185), .X(n22904) );
  nand_x1_sg U57388 ( .A(reg_w_1[1]), .B(n30370), .X(n22903) );
  nand_x1_sg U57389 ( .A(w_1[4]), .B(n34480), .X(n22910) );
  nand_x1_sg U57390 ( .A(reg_w_1[4]), .B(n33273), .X(n22909) );
  nand_x1_sg U57391 ( .A(w_1[7]), .B(n33248), .X(n22916) );
  nand_x1_sg U57392 ( .A(reg_w_1[7]), .B(n32080), .X(n22915) );
  nand_x1_sg U57393 ( .A(w_1[10]), .B(n30801), .X(n22922) );
  nand_x1_sg U57394 ( .A(reg_w_1[10]), .B(n30371), .X(n22921) );
  nand_x1_sg U57395 ( .A(w_1[13]), .B(n33225), .X(n22928) );
  nand_x1_sg U57396 ( .A(reg_w_1[13]), .B(n31961), .X(n22927) );
  nand_x1_sg U57397 ( .A(w_1[16]), .B(n33230), .X(n22934) );
  nand_x1_sg U57398 ( .A(reg_w_1[16]), .B(n30373), .X(n22933) );
  nand_x1_sg U57399 ( .A(w_1[19]), .B(n34476), .X(n22940) );
  nand_x1_sg U57400 ( .A(reg_w_1[19]), .B(n32952), .X(n22939) );
  nand_x1_sg U57401 ( .A(w_2[2]), .B(n34827), .X(n22946) );
  nand_x1_sg U57402 ( .A(reg_w_2[2]), .B(n34825), .X(n22945) );
  nand_x1_sg U57403 ( .A(w_2[5]), .B(n33245), .X(n22952) );
  nand_x1_sg U57404 ( .A(reg_w_2[5]), .B(n30788), .X(n22951) );
  nand_x1_sg U57405 ( .A(w_2[8]), .B(n30802), .X(n22958) );
  nand_x1_sg U57406 ( .A(reg_w_2[8]), .B(n29751), .X(n22957) );
  nand_x1_sg U57407 ( .A(w_2[11]), .B(n34933), .X(n22964) );
  nand_x1_sg U57408 ( .A(reg_w_2[11]), .B(n34524), .X(n22963) );
  nand_x1_sg U57409 ( .A(w_2[14]), .B(n30825), .X(n22970) );
  nand_x1_sg U57410 ( .A(reg_w_2[14]), .B(n34466), .X(n22969) );
  nand_x1_sg U57411 ( .A(w_2[17]), .B(n33245), .X(n22976) );
  nand_x1_sg U57412 ( .A(reg_w_2[17]), .B(n32092), .X(n22975) );
  nand_x1_sg U57413 ( .A(w_3[0]), .B(n32180), .X(n22982) );
  nand_x1_sg U57414 ( .A(reg_w_3[0]), .B(n34826), .X(n22981) );
  nand_x1_sg U57415 ( .A(w_3[3]), .B(n30381), .X(n22988) );
  nand_x1_sg U57416 ( .A(reg_w_3[3]), .B(n32969), .X(n22987) );
  nand_x1_sg U57417 ( .A(w_3[6]), .B(n31936), .X(n22994) );
  nand_x1_sg U57418 ( .A(reg_w_3[6]), .B(n34473), .X(n22993) );
  nand_x1_sg U57419 ( .A(w_3[9]), .B(n34475), .X(n23000) );
  nand_x1_sg U57420 ( .A(reg_w_3[9]), .B(n33265), .X(n22999) );
  nand_x1_sg U57421 ( .A(w_3[12]), .B(n34934), .X(n23006) );
  nand_x1_sg U57422 ( .A(reg_w_3[12]), .B(n32075), .X(n23005) );
  nand_x1_sg U57423 ( .A(w_3[15]), .B(n33250), .X(n23012) );
  nand_x1_sg U57424 ( .A(reg_w_3[15]), .B(n29782), .X(n23011) );
  nand_x1_sg U57425 ( .A(w_3[18]), .B(n34479), .X(n23018) );
  nand_x1_sg U57426 ( .A(reg_w_3[18]), .B(n31958), .X(n23017) );
  nand_x1_sg U57427 ( .A(w_4[1]), .B(n31940), .X(n23024) );
  nand_x1_sg U57428 ( .A(reg_w_4[1]), .B(n34925), .X(n23023) );
  nand_x1_sg U57429 ( .A(w_4[4]), .B(n30383), .X(n23030) );
  nand_x1_sg U57430 ( .A(reg_w_4[4]), .B(n29907), .X(n23029) );
  nand_x1_sg U57431 ( .A(w_4[7]), .B(n33240), .X(n23036) );
  nand_x1_sg U57432 ( .A(reg_w_4[7]), .B(n34531), .X(n23035) );
  nand_x1_sg U57433 ( .A(w_4[10]), .B(n32946), .X(n23042) );
  nand_x1_sg U57434 ( .A(reg_w_4[10]), .B(n32979), .X(n23041) );
  nand_x1_sg U57435 ( .A(w_4[13]), .B(n33916), .X(n23048) );
  nand_x1_sg U57436 ( .A(reg_w_4[13]), .B(n34923), .X(n23047) );
  nand_x1_sg U57437 ( .A(w_4[16]), .B(n34922), .X(n23054) );
  nand_x1_sg U57438 ( .A(reg_w_4[16]), .B(n32080), .X(n23053) );
  nand_x1_sg U57439 ( .A(w_4[19]), .B(n31624), .X(n23060) );
  nand_x1_sg U57440 ( .A(reg_w_4[19]), .B(n34469), .X(n23059) );
  nand_x1_sg U57441 ( .A(w_5[2]), .B(n34490), .X(n23066) );
  nand_x1_sg U57442 ( .A(reg_w_5[2]), .B(n33267), .X(n23065) );
  nand_x1_sg U57443 ( .A(w_5[5]), .B(n30813), .X(n23072) );
  nand_x1_sg U57444 ( .A(reg_w_5[5]), .B(n34510), .X(n23071) );
  nand_x1_sg U57445 ( .A(w_5[8]), .B(n30825), .X(n23078) );
  nand_x1_sg U57446 ( .A(reg_w_5[8]), .B(n30614), .X(n23077) );
  nand_x1_sg U57447 ( .A(w_5[11]), .B(n29883), .X(n23084) );
  nand_x1_sg U57448 ( .A(reg_w_5[11]), .B(n30371), .X(n23083) );
  nand_x1_sg U57449 ( .A(w_5[14]), .B(n29879), .X(n23090) );
  nand_x1_sg U57450 ( .A(reg_w_5[14]), .B(n29784), .X(n23089) );
  nand_x1_sg U57451 ( .A(w_5[17]), .B(n33251), .X(n23096) );
  nand_x1_sg U57452 ( .A(reg_w_5[17]), .B(n34821), .X(n23095) );
  nand_x1_sg U57453 ( .A(w_6[0]), .B(n30806), .X(n23102) );
  nand_x1_sg U57454 ( .A(reg_w_6[0]), .B(n31017), .X(n23101) );
  nand_x1_sg U57455 ( .A(w_6[3]), .B(n30382), .X(n23108) );
  nand_x1_sg U57456 ( .A(reg_w_6[3]), .B(n30375), .X(n23107) );
  nand_x1_sg U57457 ( .A(w_6[6]), .B(n34503), .X(n23114) );
  nand_x1_sg U57458 ( .A(reg_w_6[6]), .B(n32963), .X(n23113) );
  nand_x1_sg U57459 ( .A(w_6[9]), .B(n33224), .X(n23120) );
  nand_x1_sg U57460 ( .A(reg_w_6[9]), .B(n34825), .X(n23119) );
  nand_x1_sg U57461 ( .A(w_6[12]), .B(n30612), .X(n23126) );
  nand_x1_sg U57462 ( .A(reg_w_6[12]), .B(n29754), .X(n23125) );
  nand_x1_sg U57463 ( .A(w_6[15]), .B(n30811), .X(n23132) );
  nand_x1_sg U57464 ( .A(reg_w_6[15]), .B(n31625), .X(n23131) );
  nand_x1_sg U57465 ( .A(w_6[18]), .B(n33252), .X(n23138) );
  nand_x1_sg U57466 ( .A(reg_w_6[18]), .B(n34524), .X(n23137) );
  nand_x1_sg U57467 ( .A(w_7[1]), .B(n30384), .X(n23144) );
  nand_x1_sg U57468 ( .A(reg_w_7[1]), .B(n32979), .X(n23143) );
  nand_x1_sg U57469 ( .A(w_7[4]), .B(n30832), .X(n23150) );
  nand_x1_sg U57470 ( .A(reg_w_7[4]), .B(n31286), .X(n23149) );
  nand_x1_sg U57471 ( .A(w_7[7]), .B(n30383), .X(n23156) );
  nand_x1_sg U57472 ( .A(reg_w_7[7]), .B(n34916), .X(n23155) );
  nand_x1_sg U57473 ( .A(w_7[10]), .B(n31968), .X(n23162) );
  nand_x1_sg U57474 ( .A(reg_w_7[10]), .B(n31011), .X(n23161) );
  nand_x1_sg U57475 ( .A(w_7[13]), .B(n33234), .X(n23168) );
  nand_x1_sg U57476 ( .A(reg_w_7[13]), .B(n31960), .X(n23167) );
  nand_x1_sg U57477 ( .A(w_7[16]), .B(n29895), .X(n23174) );
  nand_x1_sg U57478 ( .A(reg_w_7[16]), .B(n32974), .X(n23173) );
  nand_x1_sg U57479 ( .A(w_7[19]), .B(n30792), .X(n23180) );
  nand_x1_sg U57480 ( .A(reg_w_7[19]), .B(n32092), .X(n23179) );
  nand_x1_sg U57481 ( .A(w_8[2]), .B(n30612), .X(n23186) );
  nand_x1_sg U57482 ( .A(reg_w_8[2]), .B(n30790), .X(n23185) );
  nand_x1_sg U57483 ( .A(w_8[5]), .B(n34834), .X(n23192) );
  nand_x1_sg U57484 ( .A(reg_w_8[5]), .B(n30370), .X(n23191) );
  nand_x1_sg U57485 ( .A(w_8[8]), .B(n34478), .X(n23198) );
  nand_x1_sg U57486 ( .A(reg_w_8[8]), .B(n30614), .X(n23197) );
  nand_x1_sg U57487 ( .A(w_8[11]), .B(n32944), .X(n23204) );
  nand_x1_sg U57488 ( .A(reg_w_8[11]), .B(n32950), .X(n23203) );
  nand_x1_sg U57489 ( .A(w_8[14]), .B(n33240), .X(n23210) );
  nand_x1_sg U57490 ( .A(reg_w_8[14]), .B(n30818), .X(n23209) );
  nand_x1_sg U57491 ( .A(w_8[17]), .B(n34461), .X(n23216) );
  nand_x1_sg U57492 ( .A(reg_w_8[17]), .B(n32949), .X(n23215) );
  nand_x1_sg U57493 ( .A(w_9[0]), .B(n31949), .X(n23222) );
  nand_x1_sg U57494 ( .A(reg_w_9[0]), .B(n31282), .X(n23221) );
  nand_x1_sg U57495 ( .A(w_9[3]), .B(n31964), .X(n23228) );
  nand_x1_sg U57496 ( .A(reg_w_9[3]), .B(n32963), .X(n23227) );
  nand_x1_sg U57497 ( .A(w_9[6]), .B(n32941), .X(n23234) );
  nand_x1_sg U57498 ( .A(reg_w_9[6]), .B(n34509), .X(n23233) );
  nand_x1_sg U57499 ( .A(w_9[9]), .B(n30824), .X(n23240) );
  nand_x1_sg U57500 ( .A(reg_w_9[9]), .B(n32959), .X(n23239) );
  nand_x1_sg U57501 ( .A(w_9[12]), .B(n30619), .X(n23246) );
  nand_x1_sg U57502 ( .A(reg_w_9[12]), .B(n30790), .X(n23245) );
  nand_x1_sg U57503 ( .A(w_9[15]), .B(n31933), .X(n23252) );
  nand_x1_sg U57504 ( .A(reg_w_9[15]), .B(n34509), .X(n23251) );
  nand_x1_sg U57505 ( .A(w_9[18]), .B(n34454), .X(n23258) );
  nand_x1_sg U57506 ( .A(reg_w_9[18]), .B(n31290), .X(n23257) );
  nand_x1_sg U57507 ( .A(w_10[1]), .B(n32945), .X(n23264) );
  nand_x1_sg U57508 ( .A(reg_w_10[1]), .B(n31626), .X(n23263) );
  nand_x1_sg U57509 ( .A(w_10[4]), .B(n34485), .X(n23270) );
  nand_x1_sg U57510 ( .A(reg_w_10[4]), .B(n30375), .X(n23269) );
  nand_x1_sg U57511 ( .A(w_10[7]), .B(n34491), .X(n23276) );
  nand_x1_sg U57512 ( .A(reg_w_10[7]), .B(n31016), .X(n23275) );
  nand_x1_sg U57513 ( .A(w_10[10]), .B(n31970), .X(n23282) );
  nand_x1_sg U57514 ( .A(reg_w_10[10]), .B(n30130), .X(n23281) );
  nand_x1_sg U57515 ( .A(w_10[13]), .B(n31946), .X(n23288) );
  nand_x1_sg U57516 ( .A(reg_w_10[13]), .B(n30819), .X(n23287) );
  nand_x1_sg U57517 ( .A(w_10[16]), .B(n30379), .X(n23294) );
  nand_x1_sg U57518 ( .A(reg_w_10[16]), .B(n31957), .X(n23293) );
  nand_x1_sg U57519 ( .A(w_10[19]), .B(n32944), .X(n23300) );
  nand_x1_sg U57520 ( .A(reg_w_10[19]), .B(n32950), .X(n23299) );
  nand_x1_sg U57521 ( .A(w_11[2]), .B(n31099), .X(n23306) );
  nand_x1_sg U57522 ( .A(reg_w_11[2]), .B(n32964), .X(n23305) );
  nand_x1_sg U57523 ( .A(w_11[5]), .B(n33243), .X(n23312) );
  nand_x1_sg U57524 ( .A(reg_w_11[5]), .B(n35057), .X(n23311) );
  nand_x1_sg U57525 ( .A(w_11[8]), .B(n34829), .X(n23318) );
  nand_x1_sg U57526 ( .A(reg_w_11[8]), .B(n33270), .X(n23317) );
  nand_x1_sg U57527 ( .A(w_11[11]), .B(n34485), .X(n23324) );
  nand_x1_sg U57528 ( .A(reg_w_11[11]), .B(n32955), .X(n23323) );
  nand_x1_sg U57529 ( .A(w_11[14]), .B(n34481), .X(n23330) );
  nand_x1_sg U57530 ( .A(reg_w_11[14]), .B(n34528), .X(n23329) );
  nand_x1_sg U57531 ( .A(w_11[17]), .B(n32182), .X(n23336) );
  nand_x1_sg U57532 ( .A(reg_w_11[17]), .B(n33267), .X(n23335) );
  nand_x1_sg U57533 ( .A(w_12[0]), .B(n33253), .X(n23342) );
  nand_x1_sg U57534 ( .A(reg_w_12[0]), .B(n34531), .X(n23341) );
  nand_x1_sg U57535 ( .A(w_12[3]), .B(n34490), .X(n23348) );
  nand_x1_sg U57536 ( .A(reg_w_12[3]), .B(n31481), .X(n23347) );
  nand_x1_sg U57537 ( .A(w_12[6]), .B(n31271), .X(n23354) );
  nand_x1_sg U57538 ( .A(reg_w_12[6]), .B(n29780), .X(n23353) );
  nand_x1_sg U57539 ( .A(w_12[9]), .B(n31105), .X(n23360) );
  nand_x1_sg U57540 ( .A(reg_w_12[9]), .B(n30788), .X(n23359) );
  nand_x1_sg U57541 ( .A(w_12[12]), .B(n35053), .X(n23366) );
  nand_x1_sg U57542 ( .A(reg_w_12[12]), .B(n34931), .X(n23365) );
  nand_x1_sg U57543 ( .A(w_12[15]), .B(n33237), .X(n23372) );
  nand_x1_sg U57544 ( .A(reg_w_12[15]), .B(n31238), .X(n23371) );
  nand_x1_sg U57545 ( .A(w_12[18]), .B(n32948), .X(n23378) );
  nand_x1_sg U57546 ( .A(reg_w_12[18]), .B(n34509), .X(n23377) );
  nand_x1_sg U57547 ( .A(w_13[1]), .B(n33247), .X(n23384) );
  nand_x1_sg U57548 ( .A(reg_w_13[1]), .B(n31954), .X(n23383) );
  nand_x1_sg U57549 ( .A(w_13[4]), .B(n31969), .X(n23390) );
  nand_x1_sg U57550 ( .A(reg_w_13[4]), .B(n32090), .X(n23389) );
  nand_x1_sg U57551 ( .A(w_13[7]), .B(n35054), .X(n23396) );
  nand_x1_sg U57552 ( .A(reg_w_13[7]), .B(n32090), .X(n23395) );
  nand_x1_sg U57553 ( .A(w_13[10]), .B(n30807), .X(n23402) );
  nand_x1_sg U57554 ( .A(reg_w_13[10]), .B(n32970), .X(n23401) );
  nand_x1_sg U57555 ( .A(w_13[13]), .B(n31105), .X(n23408) );
  nand_x1_sg U57556 ( .A(reg_w_13[13]), .B(n34525), .X(n23407) );
  nand_x1_sg U57557 ( .A(w_13[16]), .B(n30619), .X(n23414) );
  nand_x1_sg U57558 ( .A(reg_w_13[16]), .B(n34471), .X(n23413) );
  nand_x1_sg U57559 ( .A(w_13[19]), .B(n34478), .X(n23420) );
  nand_x1_sg U57560 ( .A(reg_w_13[19]), .B(n31281), .X(n23419) );
  nand_x1_sg U57561 ( .A(w_14[2]), .B(n31968), .X(n23426) );
  nand_x1_sg U57562 ( .A(reg_w_14[2]), .B(n31291), .X(n23425) );
  nand_x1_sg U57563 ( .A(w_14[5]), .B(n31258), .X(n23432) );
  nand_x1_sg U57564 ( .A(reg_w_14[5]), .B(n34818), .X(n23431) );
  nand_x1_sg U57565 ( .A(w_14[8]), .B(n30830), .X(n23438) );
  nand_x1_sg U57566 ( .A(reg_w_14[8]), .B(n32955), .X(n23437) );
  nand_x1_sg U57567 ( .A(w_14[11]), .B(n30620), .X(n23444) );
  nand_x1_sg U57568 ( .A(reg_w_14[11]), .B(n34528), .X(n23443) );
  nand_x1_sg U57569 ( .A(w_14[14]), .B(n29873), .X(n23450) );
  nand_x1_sg U57570 ( .A(reg_w_14[14]), .B(n29792), .X(n23449) );
  nand_x1_sg U57571 ( .A(w_14[17]), .B(n34483), .X(n23456) );
  nand_x1_sg U57572 ( .A(reg_w_14[17]), .B(n30371), .X(n23455) );
  nand_x1_sg U57573 ( .A(w_15[0]), .B(n30807), .X(n23462) );
  nand_x1_sg U57574 ( .A(reg_w_15[0]), .B(n33263), .X(n23461) );
  nand_x1_sg U57575 ( .A(w_15[3]), .B(n33232), .X(n23468) );
  nand_x1_sg U57576 ( .A(reg_w_15[3]), .B(n31956), .X(n23467) );
  nand_x1_sg U57577 ( .A(w_15[6]), .B(n32948), .X(n23474) );
  nand_x1_sg U57578 ( .A(reg_w_15[6]), .B(n34814), .X(n23473) );
  nand_x1_sg U57579 ( .A(w_15[9]), .B(n34844), .X(n23480) );
  nand_x1_sg U57580 ( .A(reg_w_15[9]), .B(n32949), .X(n23479) );
  nand_x1_sg U57581 ( .A(w_15[12]), .B(n30381), .X(n23486) );
  nand_x1_sg U57582 ( .A(reg_w_15[12]), .B(n32973), .X(n23485) );
  nand_x1_sg U57583 ( .A(w_15[15]), .B(n34828), .X(n23492) );
  nand_x1_sg U57584 ( .A(reg_w_15[15]), .B(n32964), .X(n23491) );
  nand_x1_sg U57585 ( .A(w_15[18]), .B(n29885), .X(n23498) );
  nand_x1_sg U57586 ( .A(reg_w_15[18]), .B(n32974), .X(n23497) );
  nand_x1_sg U57587 ( .A(i_mask[1]), .B(n31936), .X(n23504) );
  nand_x1_sg U57588 ( .A(reg_i_mask[1]), .B(n32957), .X(n23503) );
  nand_x1_sg U57589 ( .A(i_mask[4]), .B(n34932), .X(n23510) );
  nand_x1_sg U57590 ( .A(reg_i_mask[4]), .B(n31012), .X(n23509) );
  nand_x1_sg U57591 ( .A(i_mask[7]), .B(n33916), .X(n23516) );
  nand_x1_sg U57592 ( .A(reg_i_mask[7]), .B(n30818), .X(n23515) );
  nand_x1_sg U57593 ( .A(i_mask[10]), .B(n34457), .X(n23522) );
  nand_x1_sg U57594 ( .A(reg_i_mask[10]), .B(n34526), .X(n23521) );
  nand_x1_sg U57595 ( .A(i_mask[13]), .B(n31945), .X(n23528) );
  nand_x1_sg U57596 ( .A(reg_i_mask[13]), .B(n30131), .X(n23527) );
  nand_x1_sg U57597 ( .A(i_mask[16]), .B(n30805), .X(n23534) );
  nand_x1_sg U57598 ( .A(reg_i_mask[16]), .B(n31960), .X(n23533) );
  nand_x1_sg U57599 ( .A(i_mask[19]), .B(n30127), .X(n23540) );
  nand_x1_sg U57600 ( .A(reg_i_mask[19]), .B(n34812), .X(n23539) );
  nand_x1_sg U57601 ( .A(i_mask[22]), .B(n29898), .X(n23546) );
  nand_x1_sg U57602 ( .A(reg_i_mask[22]), .B(n31480), .X(n23545) );
  nand_x1_sg U57603 ( .A(i_mask[25]), .B(n34505), .X(n23552) );
  nand_x1_sg U57604 ( .A(reg_i_mask[25]), .B(n33272), .X(n23551) );
  nand_x1_sg U57605 ( .A(i_mask[28]), .B(n34835), .X(n23558) );
  nand_x1_sg U57606 ( .A(reg_i_mask[28]), .B(n32955), .X(n23557) );
  nand_x1_sg U57607 ( .A(i_mask[31]), .B(n31100), .X(n23564) );
  nand_x1_sg U57608 ( .A(reg_i_mask[31]), .B(n30613), .X(n23563) );
  nand_x1_sg U57609 ( .A(w_mask[2]), .B(n30615), .X(n23570) );
  nand_x1_sg U57610 ( .A(reg_w_mask[2]), .B(n31291), .X(n23569) );
  nand_x1_sg U57611 ( .A(w_mask[5]), .B(n33251), .X(n23576) );
  nand_x1_sg U57612 ( .A(reg_w_mask[5]), .B(n34930), .X(n23575) );
  nand_x1_sg U57613 ( .A(w_mask[8]), .B(n34920), .X(n23582) );
  nand_x1_sg U57614 ( .A(reg_w_mask[8]), .B(n34810), .X(n23581) );
  nand_x1_sg U57615 ( .A(w_mask[11]), .B(n32185), .X(n23588) );
  nand_x1_sg U57616 ( .A(reg_w_mask[11]), .B(n32088), .X(n23587) );
  nand_x1_sg U57617 ( .A(w_mask[14]), .B(n33252), .X(n23594) );
  nand_x1_sg U57618 ( .A(reg_w_mask[14]), .B(n34816), .X(n23593) );
  nand_x1_sg U57619 ( .A(w_mask[17]), .B(n30809), .X(n23600) );
  nand_x1_sg U57620 ( .A(reg_w_mask[17]), .B(n33841), .X(n23599) );
  nand_x1_sg U57621 ( .A(w_mask[20]), .B(n32945), .X(n23606) );
  nand_x1_sg U57622 ( .A(reg_w_mask[20]), .B(n31290), .X(n23605) );
  nand_x1_sg U57623 ( .A(w_mask[23]), .B(n32182), .X(n23612) );
  nand_x1_sg U57624 ( .A(reg_w_mask[23]), .B(n34105), .X(n23611) );
  nand_x1_sg U57625 ( .A(w_mask[26]), .B(n30194), .X(n23618) );
  nand_x1_sg U57626 ( .A(reg_w_mask[26]), .B(n33272), .X(n23617) );
  nand_x1_sg U57627 ( .A(w_mask[29]), .B(n29897), .X(n23624) );
  nand_x1_sg U57628 ( .A(reg_w_mask[29]), .B(n31291), .X(n23623) );
  nand_x1_sg U57629 ( .A(input_taken), .B(n31954), .X(n23630) );
  nand_x1_sg U57630 ( .A(i_0[0]), .B(n31934), .X(n22222) );
  nand_x1_sg U57631 ( .A(reg_i_0[0]), .B(n33268), .X(n22221) );
  nand_x1_sg U57632 ( .A(i_0[1]), .B(n31963), .X(n22224) );
  nand_x1_sg U57633 ( .A(reg_i_0[1]), .B(n29798), .X(n22223) );
  nand_x1_sg U57634 ( .A(i_0[3]), .B(n31624), .X(n22228) );
  nand_x1_sg U57635 ( .A(reg_i_0[3]), .B(n32962), .X(n22227) );
  nand_x1_sg U57636 ( .A(i_0[4]), .B(n33239), .X(n22230) );
  nand_x1_sg U57637 ( .A(reg_i_0[4]), .B(n32976), .X(n22229) );
  nand_x1_sg U57638 ( .A(i_0[6]), .B(n35055), .X(n22234) );
  nand_x1_sg U57639 ( .A(reg_i_0[6]), .B(n34530), .X(n22233) );
  nand_x1_sg U57640 ( .A(i_0[7]), .B(n33234), .X(n22236) );
  nand_x1_sg U57641 ( .A(reg_i_0[7]), .B(n29907), .X(n22235) );
  nand_x1_sg U57642 ( .A(i_0[9]), .B(n31942), .X(n22240) );
  nand_x1_sg U57643 ( .A(reg_i_0[9]), .B(n31952), .X(n22239) );
  nand_x1_sg U57644 ( .A(i_0[10]), .B(n31943), .X(n22242) );
  nand_x1_sg U57645 ( .A(reg_i_0[10]), .B(n30212), .X(n22241) );
  nand_x1_sg U57646 ( .A(i_0[12]), .B(n33252), .X(n22246) );
  nand_x1_sg U57647 ( .A(reg_i_0[12]), .B(n33265), .X(n22245) );
  nand_x1_sg U57648 ( .A(i_0[13]), .B(n31940), .X(n22248) );
  nand_x1_sg U57649 ( .A(reg_i_0[13]), .B(n31958), .X(n22247) );
  nand_x1_sg U57650 ( .A(i_0[15]), .B(n33225), .X(n22252) );
  nand_x1_sg U57651 ( .A(reg_i_0[15]), .B(n34812), .X(n22251) );
  nand_x1_sg U57652 ( .A(i_0[16]), .B(n29885), .X(n22254) );
  nand_x1_sg U57653 ( .A(reg_i_0[16]), .B(n34825), .X(n22253) );
  nand_x1_sg U57654 ( .A(i_0[18]), .B(n34828), .X(n22258) );
  nand_x1_sg U57655 ( .A(reg_i_0[18]), .B(n31211), .X(n22257) );
  nand_x1_sg U57656 ( .A(i_0[19]), .B(n30826), .X(n22260) );
  nand_x1_sg U57657 ( .A(reg_i_0[19]), .B(n30190), .X(n22259) );
  nand_x1_sg U57658 ( .A(i_1[1]), .B(n31099), .X(n22264) );
  nand_x1_sg U57659 ( .A(reg_i_1[1]), .B(n31952), .X(n22263) );
  nand_x1_sg U57660 ( .A(i_1[2]), .B(n32180), .X(n22266) );
  nand_x1_sg U57661 ( .A(reg_i_1[2]), .B(n31007), .X(n22265) );
  nand_x1_sg U57662 ( .A(i_1[4]), .B(n35052), .X(n22270) );
  nand_x1_sg U57663 ( .A(reg_i_1[4]), .B(n30822), .X(n22269) );
  nand_x1_sg U57664 ( .A(i_1[5]), .B(n34479), .X(n22272) );
  nand_x1_sg U57665 ( .A(reg_i_1[5]), .B(n29906), .X(n22271) );
  nand_x1_sg U57666 ( .A(i_1[7]), .B(n30384), .X(n22276) );
  nand_x1_sg U57667 ( .A(reg_i_1[7]), .B(n33271), .X(n22275) );
  nand_x1_sg U57668 ( .A(i_1[8]), .B(n34452), .X(n22278) );
  nand_x1_sg U57669 ( .A(reg_i_1[8]), .B(n34463), .X(n22277) );
  nand_x1_sg U57670 ( .A(i_1[10]), .B(n31966), .X(n22282) );
  nand_x1_sg U57671 ( .A(reg_i_1[10]), .B(n31016), .X(n22281) );
  nand_x1_sg U57672 ( .A(i_1[11]), .B(n34506), .X(n22284) );
  nand_x1_sg U57673 ( .A(reg_i_1[11]), .B(n34813), .X(n22283) );
  nand_x1_sg U57674 ( .A(i_1[13]), .B(n31949), .X(n22288) );
  nand_x1_sg U57675 ( .A(reg_i_1[13]), .B(n32083), .X(n22287) );
  nand_x1_sg U57676 ( .A(i_1[14]), .B(n33915), .X(n22290) );
  nand_x1_sg U57677 ( .A(reg_i_1[14]), .B(n32086), .X(n22289) );
  nand_x1_sg U57678 ( .A(i_1[16]), .B(n34456), .X(n22294) );
  nand_x1_sg U57679 ( .A(reg_i_1[16]), .B(n34531), .X(n22293) );
  nand_x1_sg U57680 ( .A(i_1[17]), .B(n31938), .X(n22296) );
  nand_x1_sg U57681 ( .A(reg_i_1[17]), .B(n34472), .X(n22295) );
  nand_x1_sg U57682 ( .A(i_1[19]), .B(n29887), .X(n22300) );
  nand_x1_sg U57683 ( .A(reg_i_1[19]), .B(n34824), .X(n22299) );
  nand_x1_sg U57684 ( .A(i_2[0]), .B(n31942), .X(n22302) );
  nand_x1_sg U57685 ( .A(reg_i_2[0]), .B(n33266), .X(n22301) );
  nand_x1_sg U57686 ( .A(i_2[2]), .B(n31105), .X(n22306) );
  nand_x1_sg U57687 ( .A(reg_i_2[2]), .B(n32077), .X(n22305) );
  nand_x1_sg U57688 ( .A(i_2[3]), .B(n33256), .X(n22308) );
  nand_x1_sg U57689 ( .A(reg_i_2[3]), .B(n34106), .X(n22307) );
  nand_x1_sg U57690 ( .A(i_2[5]), .B(n34934), .X(n22312) );
  nand_x1_sg U57691 ( .A(reg_i_2[5]), .B(n34106), .X(n22311) );
  nand_x1_sg U57692 ( .A(i_2[6]), .B(n31627), .X(n22314) );
  nand_x1_sg U57693 ( .A(reg_i_2[6]), .B(n32091), .X(n22313) );
  nand_x1_sg U57694 ( .A(i_2[8]), .B(n31949), .X(n22318) );
  nand_x1_sg U57695 ( .A(reg_i_2[8]), .B(n34824), .X(n22317) );
  nand_x1_sg U57696 ( .A(i_2[9]), .B(n31933), .X(n22320) );
  nand_x1_sg U57697 ( .A(reg_i_2[9]), .B(n34467), .X(n22319) );
  nand_x1_sg U57698 ( .A(i_2[11]), .B(n34832), .X(n22324) );
  nand_x1_sg U57699 ( .A(reg_i_2[11]), .B(n30133), .X(n22323) );
  nand_x1_sg U57700 ( .A(i_2[12]), .B(n34456), .X(n22326) );
  nand_x1_sg U57701 ( .A(reg_i_2[12]), .B(n32980), .X(n22325) );
  nand_x1_sg U57702 ( .A(i_2[14]), .B(n33250), .X(n22330) );
  nand_x1_sg U57703 ( .A(reg_i_2[14]), .B(n34474), .X(n22329) );
  nand_x1_sg U57704 ( .A(i_2[15]), .B(n34489), .X(n22332) );
  nand_x1_sg U57705 ( .A(reg_i_2[15]), .B(n32964), .X(n22331) );
  nand_x1_sg U57706 ( .A(i_2[17]), .B(n33239), .X(n22336) );
  nand_x1_sg U57707 ( .A(reg_i_2[17]), .B(n32076), .X(n22335) );
  nand_x1_sg U57708 ( .A(i_2[18]), .B(n33250), .X(n22338) );
  nand_x1_sg U57709 ( .A(reg_i_2[18]), .B(n29788), .X(n22337) );
  nand_x1_sg U57710 ( .A(i_3[0]), .B(n34830), .X(n22342) );
  nand_x1_sg U57711 ( .A(reg_i_3[0]), .B(n32078), .X(n22341) );
  nand_x1_sg U57712 ( .A(i_3[1]), .B(n29875), .X(n22344) );
  nand_x1_sg U57713 ( .A(reg_i_3[1]), .B(n32970), .X(n22343) );
  nand_x1_sg U57714 ( .A(i_3[3]), .B(n31627), .X(n22348) );
  nand_x1_sg U57715 ( .A(reg_i_3[3]), .B(n31954), .X(n22347) );
  nand_x1_sg U57716 ( .A(i_3[4]), .B(n30830), .X(n22350) );
  nand_x1_sg U57717 ( .A(reg_i_3[4]), .B(n31017), .X(n22349) );
  nand_x1_sg U57718 ( .A(i_3[6]), .B(n32943), .X(n22354) );
  nand_x1_sg U57719 ( .A(reg_i_3[6]), .B(n34532), .X(n22353) );
  nand_x1_sg U57720 ( .A(i_3[7]), .B(n34827), .X(n22356) );
  nand_x1_sg U57721 ( .A(reg_i_3[7]), .B(n32966), .X(n22355) );
  nand_x1_sg U57722 ( .A(i_3[9]), .B(n33229), .X(n22360) );
  nand_x1_sg U57723 ( .A(reg_i_3[9]), .B(n34510), .X(n22359) );
  nand_x1_sg U57724 ( .A(i_3[10]), .B(n29898), .X(n22362) );
  nand_x1_sg U57725 ( .A(reg_i_3[10]), .B(n32976), .X(n22361) );
  nand_x1_sg U57726 ( .A(i_3[12]), .B(n31943), .X(n22366) );
  nand_x1_sg U57727 ( .A(reg_i_3[12]), .B(n34474), .X(n22365) );
  nand_x1_sg U57728 ( .A(i_3[13]), .B(n30793), .X(n22368) );
  nand_x1_sg U57729 ( .A(reg_i_3[13]), .B(n31286), .X(n22367) );
  nand_x1_sg U57730 ( .A(i_3[15]), .B(n34459), .X(n22372) );
  nand_x1_sg U57731 ( .A(reg_i_3[15]), .B(n32953), .X(n22371) );
  nand_x1_sg U57732 ( .A(i_3[16]), .B(n30801), .X(n22374) );
  nand_x1_sg U57733 ( .A(reg_i_3[16]), .B(n32975), .X(n22373) );
  nand_x1_sg U57734 ( .A(i_3[18]), .B(n33242), .X(n22378) );
  nand_x1_sg U57735 ( .A(reg_i_3[18]), .B(n31277), .X(n22377) );
  nand_x1_sg U57736 ( .A(i_3[19]), .B(n34932), .X(n22380) );
  nand_x1_sg U57737 ( .A(reg_i_3[19]), .B(n33841), .X(n22379) );
  nand_x1_sg U57738 ( .A(i_4[1]), .B(n33234), .X(n22384) );
  nand_x1_sg U57739 ( .A(reg_i_4[1]), .B(n34929), .X(n22383) );
  nand_x1_sg U57740 ( .A(i_4[2]), .B(n34840), .X(n22386) );
  nand_x1_sg U57741 ( .A(reg_i_4[2]), .B(n34923), .X(n22385) );
  nand_x1_sg U57742 ( .A(i_4[4]), .B(n33915), .X(n22390) );
  nand_x1_sg U57743 ( .A(reg_i_4[4]), .B(n34466), .X(n22389) );
  nand_x1_sg U57744 ( .A(i_4[5]), .B(n32947), .X(n22392) );
  nand_x1_sg U57745 ( .A(reg_i_4[5]), .B(n31017), .X(n22391) );
  nand_x1_sg U57746 ( .A(i_4[7]), .B(n31948), .X(n22396) );
  nand_x1_sg U57747 ( .A(reg_i_4[7]), .B(n32961), .X(n22395) );
  nand_x1_sg U57748 ( .A(i_4[8]), .B(n31974), .X(n22398) );
  nand_x1_sg U57749 ( .A(reg_i_4[8]), .B(n32071), .X(n22397) );
  nand_x1_sg U57750 ( .A(i_4[10]), .B(n29903), .X(n22402) );
  nand_x1_sg U57751 ( .A(reg_i_4[10]), .B(n30373), .X(n22401) );
  nand_x1_sg U57752 ( .A(i_4[11]), .B(n32947), .X(n22404) );
  nand_x1_sg U57753 ( .A(reg_i_4[11]), .B(n33261), .X(n22403) );
  nand_x1_sg U57754 ( .A(i_4[13]), .B(n34921), .X(n22408) );
  nand_x1_sg U57755 ( .A(reg_i_4[13]), .B(n35059), .X(n22407) );
  nand_x1_sg U57756 ( .A(i_4[14]), .B(n33239), .X(n22410) );
  nand_x1_sg U57757 ( .A(reg_i_4[14]), .B(n32087), .X(n22409) );
  nand_x1_sg U57758 ( .A(i_4[16]), .B(n33232), .X(n22414) );
  nand_x1_sg U57759 ( .A(reg_i_4[16]), .B(n30613), .X(n22413) );
  nand_x1_sg U57760 ( .A(i_4[17]), .B(n29898), .X(n22416) );
  nand_x1_sg U57761 ( .A(reg_i_4[17]), .B(n34815), .X(n22415) );
  nand_x1_sg U57762 ( .A(i_4[19]), .B(n31969), .X(n22420) );
  nand_x1_sg U57763 ( .A(reg_i_4[19]), .B(n32971), .X(n22419) );
  nand_x1_sg U57764 ( .A(i_5[0]), .B(n29901), .X(n22422) );
  nand_x1_sg U57765 ( .A(reg_i_5[0]), .B(n33270), .X(n22421) );
  nand_x1_sg U57766 ( .A(i_5[2]), .B(n33222), .X(n22426) );
  nand_x1_sg U57767 ( .A(reg_i_5[2]), .B(n34523), .X(n22425) );
  nand_x1_sg U57768 ( .A(i_5[3]), .B(n34504), .X(n22428) );
  nand_x1_sg U57769 ( .A(reg_i_5[3]), .B(n31003), .X(n22427) );
  nand_x1_sg U57770 ( .A(i_5[5]), .B(n31257), .X(n22432) );
  nand_x1_sg U57771 ( .A(reg_i_5[5]), .B(n31011), .X(n22431) );
  nand_x1_sg U57772 ( .A(i_5[6]), .B(n34456), .X(n22434) );
  nand_x1_sg U57773 ( .A(reg_i_5[6]), .B(n31480), .X(n22433) );
  nand_x1_sg U57774 ( .A(i_5[8]), .B(n33230), .X(n22438) );
  nand_x1_sg U57775 ( .A(reg_i_5[8]), .B(n31951), .X(n22437) );
  nand_x1_sg U57776 ( .A(i_5[9]), .B(n32941), .X(n22440) );
  nand_x1_sg U57777 ( .A(reg_i_5[9]), .B(n29796), .X(n22439) );
  nand_x1_sg U57778 ( .A(i_5[11]), .B(n33246), .X(n22444) );
  nand_x1_sg U57779 ( .A(reg_i_5[11]), .B(n35060), .X(n22443) );
  nand_x1_sg U57780 ( .A(i_5[12]), .B(n33237), .X(n22446) );
  nand_x1_sg U57781 ( .A(reg_i_5[12]), .B(n31011), .X(n22445) );
  nand_x1_sg U57782 ( .A(i_5[14]), .B(n30193), .X(n22450) );
  nand_x1_sg U57783 ( .A(reg_i_5[14]), .B(n30370), .X(n22449) );
  nand_x1_sg U57784 ( .A(i_5[15]), .B(n32941), .X(n22452) );
  nand_x1_sg U57785 ( .A(reg_i_5[15]), .B(n34826), .X(n22451) );
  nand_x1_sg U57786 ( .A(i_5[17]), .B(n30381), .X(n22456) );
  nand_x1_sg U57787 ( .A(reg_i_5[17]), .B(n34925), .X(n22455) );
  nand_x1_sg U57788 ( .A(i_5[18]), .B(n33915), .X(n22458) );
  nand_x1_sg U57789 ( .A(reg_i_5[18]), .B(n34463), .X(n22457) );
  nand_x1_sg U57790 ( .A(i_6[0]), .B(n34504), .X(n22462) );
  nand_x1_sg U57791 ( .A(reg_i_6[0]), .B(n30818), .X(n22461) );
  nand_x1_sg U57792 ( .A(i_6[1]), .B(n31271), .X(n22464) );
  nand_x1_sg U57793 ( .A(reg_i_6[1]), .B(n30790), .X(n22463) );
  nand_x1_sg U57794 ( .A(i_6[3]), .B(n30385), .X(n22468) );
  nand_x1_sg U57795 ( .A(reg_i_6[3]), .B(n31276), .X(n22467) );
  nand_x1_sg U57796 ( .A(i_6[4]), .B(n33235), .X(n22470) );
  nand_x1_sg U57797 ( .A(reg_i_6[4]), .B(n31625), .X(n22469) );
  nand_x1_sg U57798 ( .A(i_6[6]), .B(n32180), .X(n22474) );
  nand_x1_sg U57799 ( .A(reg_i_6[6]), .B(n32966), .X(n22473) );
  nand_x1_sg U57800 ( .A(i_6[7]), .B(n29893), .X(n22476) );
  nand_x1_sg U57801 ( .A(reg_i_6[7]), .B(n29907), .X(n22475) );
  nand_x1_sg U57802 ( .A(i_6[9]), .B(n30810), .X(n22480) );
  nand_x1_sg U57803 ( .A(reg_i_6[9]), .B(n34468), .X(n22479) );
  nand_x1_sg U57804 ( .A(i_6[10]), .B(n31967), .X(n22482) );
  nand_x1_sg U57805 ( .A(reg_i_6[10]), .B(n32967), .X(n22481) );
  nand_x1_sg U57806 ( .A(i_6[12]), .B(n31258), .X(n22486) );
  nand_x1_sg U57807 ( .A(reg_i_6[12]), .B(n34473), .X(n22485) );
  nand_x1_sg U57808 ( .A(i_6[13]), .B(n30803), .X(n22488) );
  nand_x1_sg U57809 ( .A(reg_i_6[13]), .B(n33268), .X(n22487) );
  nand_x1_sg U57810 ( .A(i_6[15]), .B(n29687), .X(n22492) );
  nand_x1_sg U57811 ( .A(reg_i_6[15]), .B(n35058), .X(n22491) );
  nand_x1_sg U57812 ( .A(i_6[16]), .B(n31257), .X(n22494) );
  nand_x1_sg U57813 ( .A(reg_i_6[16]), .B(n34467), .X(n22493) );
  nand_x1_sg U57814 ( .A(i_6[18]), .B(n30828), .X(n22498) );
  nand_x1_sg U57815 ( .A(reg_i_6[18]), .B(n29796), .X(n22497) );
  nand_x1_sg U57816 ( .A(i_6[19]), .B(n31271), .X(n22500) );
  nand_x1_sg U57817 ( .A(reg_i_6[19]), .B(n29752), .X(n22499) );
  nand_x1_sg U57818 ( .A(i_7[1]), .B(n30127), .X(n22504) );
  nand_x1_sg U57819 ( .A(reg_i_7[1]), .B(n32953), .X(n22503) );
  nand_x1_sg U57820 ( .A(i_7[2]), .B(n31099), .X(n22506) );
  nand_x1_sg U57821 ( .A(reg_i_7[2]), .B(n30378), .X(n22505) );
  nand_x1_sg U57822 ( .A(i_7[4]), .B(n30127), .X(n22510) );
  nand_x1_sg U57823 ( .A(reg_i_7[4]), .B(n34521), .X(n22509) );
  nand_x1_sg U57824 ( .A(i_7[5]), .B(n34480), .X(n22512) );
  nand_x1_sg U57825 ( .A(reg_i_7[5]), .B(n30613), .X(n22511) );
  nand_x1_sg U57826 ( .A(i_7[7]), .B(n33258), .X(n22516) );
  nand_x1_sg U57827 ( .A(reg_i_7[7]), .B(n30367), .X(n22515) );
  nand_x1_sg U57828 ( .A(i_7[8]), .B(n30381), .X(n22518) );
  nand_x1_sg U57829 ( .A(reg_i_7[8]), .B(n30823), .X(n22517) );
  nand_x1_sg U57830 ( .A(i_7[10]), .B(n29875), .X(n22522) );
  nand_x1_sg U57831 ( .A(reg_i_7[10]), .B(n29778), .X(n22521) );
  nand_x1_sg U57832 ( .A(i_7[11]), .B(n34829), .X(n22524) );
  nand_x1_sg U57833 ( .A(reg_i_7[11]), .B(n33266), .X(n22523) );
  nand_x1_sg U57834 ( .A(i_7[13]), .B(n29869), .X(n22528) );
  nand_x1_sg U57835 ( .A(reg_i_7[13]), .B(n29790), .X(n22527) );
  nand_x1_sg U57836 ( .A(i_7[14]), .B(n33242), .X(n22530) );
  nand_x1_sg U57837 ( .A(reg_i_7[14]), .B(n30190), .X(n22529) );
  nand_x1_sg U57838 ( .A(i_7[16]), .B(n30792), .X(n22534) );
  nand_x1_sg U57839 ( .A(reg_i_7[16]), .B(n34508), .X(n22533) );
  nand_x1_sg U57840 ( .A(i_7[17]), .B(n33257), .X(n22536) );
  nand_x1_sg U57841 ( .A(reg_i_7[17]), .B(n32979), .X(n22535) );
  nand_x1_sg U57842 ( .A(i_7[19]), .B(n33225), .X(n22540) );
  nand_x1_sg U57843 ( .A(reg_i_7[19]), .B(n34924), .X(n22539) );
  nand_x1_sg U57844 ( .A(i_8[0]), .B(n34917), .X(n22542) );
  nand_x1_sg U57845 ( .A(reg_i_8[0]), .B(n30820), .X(n22541) );
  nand_x1_sg U57846 ( .A(i_8[2]), .B(n32942), .X(n22546) );
  nand_x1_sg U57847 ( .A(reg_i_8[2]), .B(n31016), .X(n22545) );
  nand_x1_sg U57848 ( .A(i_8[3]), .B(n34920), .X(n22548) );
  nand_x1_sg U57849 ( .A(reg_i_8[3]), .B(n34813), .X(n22547) );
  nand_x1_sg U57850 ( .A(i_8[5]), .B(n29873), .X(n22552) );
  nand_x1_sg U57851 ( .A(reg_i_8[5]), .B(n29794), .X(n22551) );
  nand_x1_sg U57852 ( .A(i_8[6]), .B(n33255), .X(n22554) );
  nand_x1_sg U57853 ( .A(reg_i_8[6]), .B(n34915), .X(n22553) );
  nand_x1_sg U57854 ( .A(i_8[8]), .B(n34485), .X(n22558) );
  nand_x1_sg U57855 ( .A(reg_i_8[8]), .B(n35058), .X(n22557) );
  nand_x1_sg U57856 ( .A(i_8[9]), .B(n30806), .X(n22560) );
  nand_x1_sg U57857 ( .A(reg_i_8[9]), .B(n30823), .X(n22559) );
  nand_x1_sg U57858 ( .A(i_8[11]), .B(n30194), .X(n22564) );
  nand_x1_sg U57859 ( .A(reg_i_8[11]), .B(n34106), .X(n22563) );
  nand_x1_sg U57860 ( .A(i_8[12]), .B(n31973), .X(n22566) );
  nand_x1_sg U57861 ( .A(reg_i_8[12]), .B(n29907), .X(n22565) );
  nand_x1_sg U57862 ( .A(i_8[14]), .B(n31945), .X(n22570) );
  nand_x1_sg U57863 ( .A(reg_i_8[14]), .B(n32960), .X(n22569) );
  nand_x1_sg U57864 ( .A(i_8[15]), .B(n32941), .X(n22572) );
  nand_x1_sg U57865 ( .A(reg_i_8[15]), .B(n34526), .X(n22571) );
  nand_x1_sg U57866 ( .A(i_8[17]), .B(n31936), .X(n22576) );
  nand_x1_sg U57867 ( .A(reg_i_8[17]), .B(n30130), .X(n22575) );
  nand_x1_sg U57868 ( .A(i_8[18]), .B(n33255), .X(n22578) );
  nand_x1_sg U57869 ( .A(reg_i_8[18]), .B(n30819), .X(n22577) );
  nand_x1_sg U57870 ( .A(i_9[0]), .B(n29883), .X(n22582) );
  nand_x1_sg U57871 ( .A(reg_i_9[0]), .B(n29905), .X(n22581) );
  nand_x1_sg U57872 ( .A(i_9[1]), .B(n34488), .X(n22584) );
  nand_x1_sg U57873 ( .A(reg_i_9[1]), .B(n32978), .X(n22583) );
  nand_x1_sg U57874 ( .A(i_9[3]), .B(n31950), .X(n22588) );
  nand_x1_sg U57875 ( .A(reg_i_9[3]), .B(n34511), .X(n22587) );
  nand_x1_sg U57876 ( .A(i_9[4]), .B(n34922), .X(n22590) );
  nand_x1_sg U57877 ( .A(reg_i_9[4]), .B(n32071), .X(n22589) );
  nand_x1_sg U57878 ( .A(i_9[6]), .B(n31938), .X(n22594) );
  nand_x1_sg U57879 ( .A(reg_i_9[6]), .B(n31952), .X(n22593) );
  nand_x1_sg U57880 ( .A(i_9[7]), .B(n34475), .X(n22596) );
  nand_x1_sg U57881 ( .A(reg_i_9[7]), .B(n31102), .X(n22595) );
  nand_x1_sg U57882 ( .A(i_9[9]), .B(n31940), .X(n22600) );
  nand_x1_sg U57883 ( .A(reg_i_9[9]), .B(n33270), .X(n22599) );
  nand_x1_sg U57884 ( .A(i_9[10]), .B(n33256), .X(n22602) );
  nand_x1_sg U57885 ( .A(reg_i_9[10]), .B(n33270), .X(n22601) );
  nand_x1_sg U57886 ( .A(i_9[12]), .B(n31966), .X(n22606) );
  nand_x1_sg U57887 ( .A(reg_i_9[12]), .B(n31957), .X(n22605) );
  nand_x1_sg U57888 ( .A(i_9[13]), .B(n30192), .X(n22608) );
  nand_x1_sg U57889 ( .A(reg_i_9[13]), .B(n32954), .X(n22607) );
  nand_x1_sg U57890 ( .A(i_9[15]), .B(n33257), .X(n22612) );
  nand_x1_sg U57891 ( .A(reg_i_9[15]), .B(n30822), .X(n22611) );
  nand_x1_sg U57892 ( .A(i_9[16]), .B(n34505), .X(n22614) );
  nand_x1_sg U57893 ( .A(reg_i_9[16]), .B(n34105), .X(n22613) );
  nand_x1_sg U57894 ( .A(i_9[18]), .B(n35052), .X(n22618) );
  nand_x1_sg U57895 ( .A(reg_i_9[18]), .B(n32075), .X(n22617) );
  nand_x1_sg U57896 ( .A(i_9[19]), .B(n34837), .X(n22620) );
  nand_x1_sg U57897 ( .A(reg_i_9[19]), .B(n35059), .X(n22619) );
  nand_x1_sg U57898 ( .A(i_10[1]), .B(n33249), .X(n22624) );
  nand_x1_sg U57899 ( .A(reg_i_10[1]), .B(n33260), .X(n22623) );
  nand_x1_sg U57900 ( .A(i_10[2]), .B(n34935), .X(n22626) );
  nand_x1_sg U57901 ( .A(reg_i_10[2]), .B(n31238), .X(n22625) );
  nand_x1_sg U57902 ( .A(i_10[4]), .B(n34845), .X(n22630) );
  nand_x1_sg U57903 ( .A(reg_i_10[4]), .B(n30375), .X(n22629) );
  nand_x1_sg U57904 ( .A(i_10[5]), .B(n34457), .X(n22632) );
  nand_x1_sg U57905 ( .A(reg_i_10[5]), .B(n35060), .X(n22631) );
  nand_x1_sg U57906 ( .A(i_10[7]), .B(n29879), .X(n22636) );
  nand_x1_sg U57907 ( .A(reg_i_10[7]), .B(n32973), .X(n22635) );
  nand_x1_sg U57908 ( .A(i_10[8]), .B(n33228), .X(n22638) );
  nand_x1_sg U57909 ( .A(reg_i_10[8]), .B(n32078), .X(n22637) );
  nand_x1_sg U57910 ( .A(i_10[10]), .B(n34460), .X(n22642) );
  nand_x1_sg U57911 ( .A(reg_i_10[10]), .B(n31237), .X(n22641) );
  nand_x1_sg U57912 ( .A(i_10[11]), .B(n34933), .X(n22644) );
  nand_x1_sg U57913 ( .A(reg_i_10[11]), .B(n31962), .X(n22643) );
  nand_x1_sg U57914 ( .A(i_10[13]), .B(n30803), .X(n22648) );
  nand_x1_sg U57915 ( .A(reg_i_10[13]), .B(n30367), .X(n22647) );
  nand_x1_sg U57916 ( .A(i_10[14]), .B(n34481), .X(n22650) );
  nand_x1_sg U57917 ( .A(reg_i_10[14]), .B(n32091), .X(n22649) );
  nand_x1_sg U57918 ( .A(i_10[16]), .B(n29897), .X(n22654) );
  nand_x1_sg U57919 ( .A(reg_i_10[16]), .B(n29790), .X(n22653) );
  nand_x1_sg U57920 ( .A(i_10[17]), .B(n29897), .X(n22656) );
  nand_x1_sg U57921 ( .A(reg_i_10[17]), .B(n33261), .X(n22655) );
  nand_x1_sg U57922 ( .A(i_10[19]), .B(n30793), .X(n22660) );
  nand_x1_sg U57923 ( .A(reg_i_10[19]), .B(n35059), .X(n22659) );
  nand_x1_sg U57924 ( .A(i_11[0]), .B(n34917), .X(n22662) );
  nand_x1_sg U57925 ( .A(reg_i_11[0]), .B(n31012), .X(n22661) );
  nand_x1_sg U57926 ( .A(i_11[2]), .B(n30806), .X(n22666) );
  nand_x1_sg U57927 ( .A(reg_i_11[2]), .B(n34826), .X(n22665) );
  nand_x1_sg U57928 ( .A(i_11[3]), .B(n33238), .X(n22668) );
  nand_x1_sg U57929 ( .A(reg_i_11[3]), .B(n30789), .X(n22667) );
  nand_x1_sg U57930 ( .A(i_11[5]), .B(n34479), .X(n22672) );
  nand_x1_sg U57931 ( .A(reg_i_11[5]), .B(n30816), .X(n22671) );
  nand_x1_sg U57932 ( .A(i_11[6]), .B(n33248), .X(n22674) );
  nand_x1_sg U57933 ( .A(reg_i_11[6]), .B(n34916), .X(n22673) );
  nand_x1_sg U57934 ( .A(i_11[8]), .B(n34840), .X(n22678) );
  nand_x1_sg U57935 ( .A(reg_i_11[8]), .B(n32956), .X(n22677) );
  nand_x1_sg U57936 ( .A(i_11[9]), .B(n31272), .X(n22680) );
  nand_x1_sg U57937 ( .A(reg_i_11[9]), .B(n31276), .X(n22679) );
  nand_x1_sg U57938 ( .A(i_11[11]), .B(n30193), .X(n22684) );
  nand_x1_sg U57939 ( .A(reg_i_11[11]), .B(n30368), .X(n22683) );
  nand_x1_sg U57940 ( .A(i_11[12]), .B(n34486), .X(n22686) );
  nand_x1_sg U57941 ( .A(reg_i_11[12]), .B(n32088), .X(n22685) );
  nand_x1_sg U57942 ( .A(i_11[14]), .B(n34504), .X(n22690) );
  nand_x1_sg U57943 ( .A(reg_i_11[14]), .B(n30816), .X(n22689) );
  nand_x1_sg U57944 ( .A(i_11[15]), .B(n30612), .X(n22692) );
  nand_x1_sg U57945 ( .A(reg_i_11[15]), .B(n33268), .X(n22691) );
  nand_x1_sg U57946 ( .A(i_11[17]), .B(n31963), .X(n22696) );
  nand_x1_sg U57947 ( .A(reg_i_11[17]), .B(n34523), .X(n22695) );
  nand_x1_sg U57948 ( .A(i_11[18]), .B(n30619), .X(n22698) );
  nand_x1_sg U57949 ( .A(reg_i_11[18]), .B(n34931), .X(n22697) );
  nand_x1_sg U57950 ( .A(i_12[0]), .B(n34828), .X(n22702) );
  nand_x1_sg U57951 ( .A(reg_i_12[0]), .B(n32074), .X(n22701) );
  nand_x1_sg U57952 ( .A(i_12[1]), .B(n34460), .X(n22704) );
  nand_x1_sg U57953 ( .A(reg_i_12[1]), .B(n34810), .X(n22703) );
  nand_x1_sg U57954 ( .A(i_12[3]), .B(n34484), .X(n22708) );
  nand_x1_sg U57955 ( .A(reg_i_12[3]), .B(n32961), .X(n22707) );
  nand_x1_sg U57956 ( .A(i_12[4]), .B(n33237), .X(n22710) );
  nand_x1_sg U57957 ( .A(reg_i_12[4]), .B(n34510), .X(n22709) );
  nand_x1_sg U57958 ( .A(i_12[6]), .B(n34829), .X(n22714) );
  nand_x1_sg U57959 ( .A(reg_i_12[6]), .B(n33262), .X(n22713) );
  nand_x1_sg U57960 ( .A(i_12[7]), .B(n29897), .X(n22716) );
  nand_x1_sg U57961 ( .A(reg_i_12[7]), .B(n32980), .X(n22715) );
  nand_x1_sg U57962 ( .A(i_12[9]), .B(n31944), .X(n22720) );
  nand_x1_sg U57963 ( .A(reg_i_12[9]), .B(n31281), .X(n22719) );
  nand_x1_sg U57964 ( .A(i_12[10]), .B(n31628), .X(n22722) );
  nand_x1_sg U57965 ( .A(reg_i_12[10]), .B(n31958), .X(n22721) );
  nand_x1_sg U57966 ( .A(i_12[12]), .B(n34485), .X(n22726) );
  nand_x1_sg U57967 ( .A(reg_i_12[12]), .B(n34929), .X(n22725) );
  nand_x1_sg U57968 ( .A(i_12[13]), .B(n30384), .X(n22728) );
  nand_x1_sg U57969 ( .A(reg_i_12[13]), .B(n34813), .X(n22727) );
  nand_x1_sg U57970 ( .A(i_12[15]), .B(n34459), .X(n22732) );
  nand_x1_sg U57971 ( .A(reg_i_12[15]), .B(n31281), .X(n22731) );
  nand_x1_sg U57972 ( .A(i_12[16]), .B(n31934), .X(n22734) );
  nand_x1_sg U57973 ( .A(reg_i_12[16]), .B(n34510), .X(n22733) );
  nand_x1_sg U57974 ( .A(i_12[18]), .B(n34844), .X(n22738) );
  nand_x1_sg U57975 ( .A(reg_i_12[18]), .B(n31006), .X(n22737) );
  nand_x1_sg U57976 ( .A(i_12[19]), .B(n32943), .X(n22740) );
  nand_x1_sg U57977 ( .A(reg_i_12[19]), .B(n29786), .X(n22739) );
  nand_x1_sg U57978 ( .A(i_13[1]), .B(n31272), .X(n22744) );
  nand_x1_sg U57979 ( .A(reg_i_13[1]), .B(n32967), .X(n22743) );
  nand_x1_sg U57980 ( .A(i_13[2]), .B(n32946), .X(n22746) );
  nand_x1_sg U57981 ( .A(reg_i_13[2]), .B(n34816), .X(n22745) );
  nand_x1_sg U57982 ( .A(i_13[4]), .B(n31942), .X(n22750) );
  nand_x1_sg U57983 ( .A(reg_i_13[4]), .B(n34526), .X(n22749) );
  nand_x1_sg U57984 ( .A(i_13[5]), .B(n31948), .X(n22752) );
  nand_x1_sg U57985 ( .A(reg_i_13[5]), .B(n31928), .X(n22751) );
  nand_x1_sg U57986 ( .A(i_13[7]), .B(n31943), .X(n22756) );
  nand_x1_sg U57987 ( .A(reg_i_13[7]), .B(n31281), .X(n22755) );
  nand_x1_sg U57988 ( .A(i_13[8]), .B(n31939), .X(n22758) );
  nand_x1_sg U57989 ( .A(reg_i_13[8]), .B(n32077), .X(n22757) );
  nand_x1_sg U57990 ( .A(i_13[10]), .B(n32180), .X(n22762) );
  nand_x1_sg U57991 ( .A(reg_i_13[10]), .B(n31955), .X(n22761) );
  nand_x1_sg U57992 ( .A(i_13[11]), .B(n34460), .X(n22764) );
  nand_x1_sg U57993 ( .A(reg_i_13[11]), .B(n30367), .X(n22763) );
  nand_x1_sg U57994 ( .A(i_13[13]), .B(n31272), .X(n22768) );
  nand_x1_sg U57995 ( .A(reg_i_13[13]), .B(n34820), .X(n22767) );
  nand_x1_sg U57996 ( .A(i_13[14]), .B(n33247), .X(n22770) );
  nand_x1_sg U57997 ( .A(reg_i_13[14]), .B(n34811), .X(n22769) );
  nand_x1_sg U57998 ( .A(i_13[16]), .B(n30810), .X(n22774) );
  nand_x1_sg U57999 ( .A(reg_i_13[16]), .B(n34468), .X(n22773) );
  nand_x1_sg U58000 ( .A(i_13[17]), .B(n31963), .X(n22776) );
  nand_x1_sg U58001 ( .A(reg_i_13[17]), .B(n33265), .X(n22775) );
  nand_x1_sg U58002 ( .A(i_13[19]), .B(n29903), .X(n22780) );
  nand_x1_sg U58003 ( .A(reg_i_13[19]), .B(n29780), .X(n22779) );
  nand_x1_sg U58004 ( .A(i_14[0]), .B(n33235), .X(n22782) );
  nand_x1_sg U58005 ( .A(reg_i_14[0]), .B(n34821), .X(n22781) );
  nand_x1_sg U58006 ( .A(i_14[2]), .B(n30826), .X(n22786) );
  nand_x1_sg U58007 ( .A(reg_i_14[2]), .B(n30614), .X(n22785) );
  nand_x1_sg U58008 ( .A(i_14[3]), .B(n34461), .X(n22788) );
  nand_x1_sg U58009 ( .A(reg_i_14[3]), .B(n31927), .X(n22787) );
  nand_x1_sg U58010 ( .A(i_14[5]), .B(n33253), .X(n22792) );
  nand_x1_sg U58011 ( .A(reg_i_14[5]), .B(n30375), .X(n22791) );
  nand_x1_sg U58012 ( .A(i_14[6]), .B(n30829), .X(n22794) );
  nand_x1_sg U58013 ( .A(reg_i_14[6]), .B(n31956), .X(n22793) );
  nand_x1_sg U58014 ( .A(i_14[8]), .B(n32946), .X(n22798) );
  nand_x1_sg U58015 ( .A(reg_i_14[8]), .B(n34468), .X(n22797) );
  nand_x1_sg U58016 ( .A(i_14[9]), .B(n32945), .X(n22800) );
  nand_x1_sg U58017 ( .A(reg_i_14[9]), .B(n31237), .X(n22799) );
  nand_x1_sg U58018 ( .A(i_14[11]), .B(n31623), .X(n22804) );
  nand_x1_sg U58019 ( .A(reg_i_14[11]), .B(n30129), .X(n22803) );
  nand_x1_sg U58020 ( .A(i_14[12]), .B(n30194), .X(n22806) );
  nand_x1_sg U58021 ( .A(reg_i_14[12]), .B(n34819), .X(n22805) );
  nand_x1_sg U58022 ( .A(i_14[14]), .B(n32947), .X(n22810) );
  nand_x1_sg U58023 ( .A(reg_i_14[14]), .B(n34815), .X(n22809) );
  nand_x1_sg U58024 ( .A(i_14[15]), .B(n34506), .X(n22812) );
  nand_x1_sg U58025 ( .A(reg_i_14[15]), .B(n33262), .X(n22811) );
  nand_x1_sg U58026 ( .A(i_14[17]), .B(n30811), .X(n22816) );
  nand_x1_sg U58027 ( .A(reg_i_14[17]), .B(n32959), .X(n22815) );
  nand_x1_sg U58028 ( .A(i_14[18]), .B(n34935), .X(n22818) );
  nand_x1_sg U58029 ( .A(reg_i_14[18]), .B(n32082), .X(n22817) );
  nand_x1_sg U58030 ( .A(i_15[0]), .B(n31628), .X(n22822) );
  nand_x1_sg U58031 ( .A(reg_i_15[0]), .B(n34824), .X(n22821) );
  nand_x1_sg U58032 ( .A(i_15[1]), .B(n31949), .X(n22824) );
  nand_x1_sg U58033 ( .A(reg_i_15[1]), .B(n32076), .X(n22823) );
  nand_x1_sg U58034 ( .A(i_15[3]), .B(n31939), .X(n22828) );
  nand_x1_sg U58035 ( .A(reg_i_15[3]), .B(n31238), .X(n22827) );
  nand_x1_sg U58036 ( .A(i_15[4]), .B(n29871), .X(n22830) );
  nand_x1_sg U58037 ( .A(reg_i_15[4]), .B(n29794), .X(n22829) );
  nand_x1_sg U58038 ( .A(i_15[6]), .B(n34483), .X(n22834) );
  nand_x1_sg U58039 ( .A(reg_i_15[6]), .B(n31481), .X(n22833) );
  nand_x1_sg U58040 ( .A(i_15[7]), .B(n33223), .X(n22836) );
  nand_x1_sg U58041 ( .A(reg_i_15[7]), .B(n32978), .X(n22835) );
  nand_x1_sg U58042 ( .A(i_15[9]), .B(n31266), .X(n22840) );
  nand_x1_sg U58043 ( .A(reg_i_15[9]), .B(n31960), .X(n22839) );
  nand_x1_sg U58044 ( .A(i_15[10]), .B(n30379), .X(n22842) );
  nand_x1_sg U58045 ( .A(reg_i_15[10]), .B(n34521), .X(n22841) );
  nand_x1_sg U58046 ( .A(i_15[12]), .B(n31934), .X(n22846) );
  nand_x1_sg U58047 ( .A(reg_i_15[12]), .B(n31006), .X(n22845) );
  nand_x1_sg U58048 ( .A(i_15[13]), .B(n35055), .X(n22848) );
  nand_x1_sg U58049 ( .A(reg_i_15[13]), .B(n30814), .X(n22847) );
  nand_x1_sg U58050 ( .A(i_15[15]), .B(n31267), .X(n22852) );
  nand_x1_sg U58051 ( .A(reg_i_15[15]), .B(n34529), .X(n22851) );
  nand_x1_sg U58052 ( .A(i_15[16]), .B(n29871), .X(n22854) );
  nand_x1_sg U58053 ( .A(reg_i_15[16]), .B(n33268), .X(n22853) );
  nand_x1_sg U58054 ( .A(i_15[18]), .B(n34486), .X(n22858) );
  nand_x1_sg U58055 ( .A(reg_i_15[18]), .B(n33273), .X(n22857) );
  nand_x1_sg U58056 ( .A(i_15[19]), .B(n34833), .X(n22860) );
  nand_x1_sg U58057 ( .A(reg_i_15[19]), .B(n30191), .X(n22859) );
  nand_x1_sg U58058 ( .A(w_0[1]), .B(n34919), .X(n22864) );
  nand_x1_sg U58059 ( .A(reg_w_0[1]), .B(n34474), .X(n22863) );
  nand_x1_sg U58060 ( .A(w_0[2]), .B(n34838), .X(n22866) );
  nand_x1_sg U58061 ( .A(reg_w_0[2]), .B(n32083), .X(n22865) );
  nand_x1_sg U58062 ( .A(w_0[4]), .B(n30617), .X(n22870) );
  nand_x1_sg U58063 ( .A(reg_w_0[4]), .B(n34464), .X(n22869) );
  nand_x1_sg U58064 ( .A(w_0[5]), .B(n34842), .X(n22872) );
  nand_x1_sg U58065 ( .A(reg_w_0[5]), .B(n34527), .X(n22871) );
  nand_x1_sg U58066 ( .A(w_0[7]), .B(n34484), .X(n22876) );
  nand_x1_sg U58067 ( .A(reg_w_0[7]), .B(n32090), .X(n22875) );
  nand_x1_sg U58068 ( .A(w_0[8]), .B(n34830), .X(n22878) );
  nand_x1_sg U58069 ( .A(reg_w_0[8]), .B(n34820), .X(n22877) );
  nand_x1_sg U58070 ( .A(w_0[10]), .B(n29874), .X(n22882) );
  nand_x1_sg U58071 ( .A(reg_w_0[10]), .B(n31290), .X(n22881) );
  nand_x1_sg U58072 ( .A(w_0[11]), .B(n34486), .X(n22884) );
  nand_x1_sg U58073 ( .A(reg_w_0[11]), .B(n34463), .X(n22883) );
  nand_x1_sg U58074 ( .A(w_0[13]), .B(n33249), .X(n22888) );
  nand_x1_sg U58075 ( .A(reg_w_0[13]), .B(n34532), .X(n22887) );
  nand_x1_sg U58076 ( .A(w_0[14]), .B(n30805), .X(n22890) );
  nand_x1_sg U58077 ( .A(reg_w_0[14]), .B(n32975), .X(n22889) );
  nand_x1_sg U58078 ( .A(w_0[16]), .B(n32183), .X(n22894) );
  nand_x1_sg U58079 ( .A(reg_w_0[16]), .B(n31951), .X(n22893) );
  nand_x1_sg U58080 ( .A(w_0[17]), .B(n29889), .X(n22896) );
  nand_x1_sg U58081 ( .A(reg_w_0[17]), .B(n34812), .X(n22895) );
  nand_x1_sg U58082 ( .A(w_0[19]), .B(n32183), .X(n22900) );
  nand_x1_sg U58083 ( .A(reg_w_0[19]), .B(n32963), .X(n22899) );
  nand_x1_sg U58084 ( .A(w_1[0]), .B(n34452), .X(n22902) );
  nand_x1_sg U58085 ( .A(reg_w_1[0]), .B(n31625), .X(n22901) );
  nand_x1_sg U58086 ( .A(w_1[2]), .B(n34480), .X(n22906) );
  nand_x1_sg U58087 ( .A(reg_w_1[2]), .B(n32084), .X(n22905) );
  nand_x1_sg U58088 ( .A(w_1[3]), .B(n30809), .X(n22908) );
  nand_x1_sg U58089 ( .A(reg_w_1[3]), .B(n34826), .X(n22907) );
  nand_x1_sg U58090 ( .A(w_1[5]), .B(n33229), .X(n22912) );
  nand_x1_sg U58091 ( .A(reg_w_1[5]), .B(n32086), .X(n22911) );
  nand_x1_sg U58092 ( .A(w_1[6]), .B(n31948), .X(n22914) );
  nand_x1_sg U58093 ( .A(reg_w_1[6]), .B(n30614), .X(n22913) );
  nand_x1_sg U58094 ( .A(w_1[8]), .B(n31623), .X(n22918) );
  nand_x1_sg U58095 ( .A(reg_w_1[8]), .B(n32083), .X(n22917) );
  nand_x1_sg U58096 ( .A(w_1[9]), .B(n34457), .X(n22920) );
  nand_x1_sg U58097 ( .A(reg_w_1[9]), .B(n32952), .X(n22919) );
  nand_x1_sg U58098 ( .A(w_1[11]), .B(n32948), .X(n22924) );
  nand_x1_sg U58099 ( .A(reg_w_1[11]), .B(n30129), .X(n22923) );
  nand_x1_sg U58100 ( .A(w_1[12]), .B(n29901), .X(n22926) );
  nand_x1_sg U58101 ( .A(reg_w_1[12]), .B(n30367), .X(n22925) );
  nand_x1_sg U58102 ( .A(w_1[14]), .B(n29889), .X(n22930) );
  nand_x1_sg U58103 ( .A(reg_w_1[14]), .B(n29792), .X(n22929) );
  nand_x1_sg U58104 ( .A(w_1[15]), .B(n33242), .X(n22932) );
  nand_x1_sg U58105 ( .A(reg_w_1[15]), .B(n30212), .X(n22931) );
  nand_x1_sg U58106 ( .A(w_1[17]), .B(n31945), .X(n22936) );
  nand_x1_sg U58107 ( .A(reg_w_1[17]), .B(n32071), .X(n22935) );
  nand_x1_sg U58108 ( .A(w_1[18]), .B(n33232), .X(n22938) );
  nand_x1_sg U58109 ( .A(reg_w_1[18]), .B(n31211), .X(n22937) );
  nand_x1_sg U58110 ( .A(w_2[0]), .B(n31972), .X(n22942) );
  nand_x1_sg U58111 ( .A(reg_w_2[0]), .B(n31012), .X(n22941) );
  nand_x1_sg U58112 ( .A(w_2[1]), .B(n29891), .X(n22944) );
  nand_x1_sg U58113 ( .A(reg_w_2[1]), .B(n33841), .X(n22943) );
  nand_x1_sg U58114 ( .A(w_2[3]), .B(n34918), .X(n22948) );
  nand_x1_sg U58115 ( .A(reg_w_2[3]), .B(n30788), .X(n22947) );
  nand_x1_sg U58116 ( .A(w_2[4]), .B(n30192), .X(n22950) );
  nand_x1_sg U58117 ( .A(reg_w_2[4]), .B(n32072), .X(n22949) );
  nand_x1_sg U58118 ( .A(w_2[6]), .B(n33244), .X(n22954) );
  nand_x1_sg U58119 ( .A(reg_w_2[6]), .B(n32074), .X(n22953) );
  nand_x1_sg U58120 ( .A(w_2[7]), .B(n30828), .X(n22956) );
  nand_x1_sg U58121 ( .A(reg_w_2[7]), .B(n34815), .X(n22955) );
  nand_x1_sg U58122 ( .A(w_2[9]), .B(n31266), .X(n22960) );
  nand_x1_sg U58123 ( .A(reg_w_2[9]), .B(n34530), .X(n22959) );
  nand_x1_sg U58124 ( .A(w_2[10]), .B(n35053), .X(n22962) );
  nand_x1_sg U58125 ( .A(reg_w_2[10]), .B(n32081), .X(n22961) );
  nand_x1_sg U58126 ( .A(w_2[12]), .B(n31267), .X(n22966) );
  nand_x1_sg U58127 ( .A(reg_w_2[12]), .B(n34467), .X(n22965) );
  nand_x1_sg U58128 ( .A(w_2[13]), .B(n31933), .X(n22968) );
  nand_x1_sg U58129 ( .A(reg_w_2[13]), .B(n33267), .X(n22967) );
  nand_x1_sg U58130 ( .A(w_2[15]), .B(n30615), .X(n22972) );
  nand_x1_sg U58131 ( .A(reg_w_2[15]), .B(n31211), .X(n22971) );
  nand_x1_sg U58132 ( .A(w_2[16]), .B(n31968), .X(n22974) );
  nand_x1_sg U58133 ( .A(reg_w_2[16]), .B(n34521), .X(n22973) );
  nand_x1_sg U58134 ( .A(w_2[18]), .B(n32185), .X(n22978) );
  nand_x1_sg U58135 ( .A(reg_w_2[18]), .B(n31007), .X(n22977) );
  nand_x1_sg U58136 ( .A(w_2[19]), .B(n30194), .X(n22980) );
  nand_x1_sg U58137 ( .A(reg_w_2[19]), .B(n33266), .X(n22979) );
  nand_x1_sg U58138 ( .A(w_3[1]), .B(n32184), .X(n22984) );
  nand_x1_sg U58139 ( .A(reg_w_3[1]), .B(n32960), .X(n22983) );
  nand_x1_sg U58140 ( .A(w_3[2]), .B(n32942), .X(n22986) );
  nand_x1_sg U58141 ( .A(reg_w_3[2]), .B(n30190), .X(n22985) );
  nand_x1_sg U58142 ( .A(w_3[4]), .B(n34932), .X(n22990) );
  nand_x1_sg U58143 ( .A(reg_w_3[4]), .B(n30816), .X(n22989) );
  nand_x1_sg U58144 ( .A(w_3[5]), .B(n30617), .X(n22992) );
  nand_x1_sg U58145 ( .A(reg_w_3[5]), .B(n34928), .X(n22991) );
  nand_x1_sg U58146 ( .A(w_3[7]), .B(n32946), .X(n22996) );
  nand_x1_sg U58147 ( .A(reg_w_3[7]), .B(n30789), .X(n22995) );
  nand_x1_sg U58148 ( .A(w_3[8]), .B(n34837), .X(n22998) );
  nand_x1_sg U58149 ( .A(reg_w_3[8]), .B(n34464), .X(n22997) );
  nand_x1_sg U58150 ( .A(w_3[10]), .B(n33257), .X(n23002) );
  nand_x1_sg U58151 ( .A(reg_w_3[10]), .B(n32081), .X(n23001) );
  nand_x1_sg U58152 ( .A(w_3[11]), .B(n34460), .X(n23004) );
  nand_x1_sg U58153 ( .A(reg_w_3[11]), .B(n32082), .X(n23003) );
  nand_x1_sg U58154 ( .A(w_3[13]), .B(n31627), .X(n23008) );
  nand_x1_sg U58155 ( .A(reg_w_3[13]), .B(n34924), .X(n23007) );
  nand_x1_sg U58156 ( .A(w_3[14]), .B(n31100), .X(n23010) );
  nand_x1_sg U58157 ( .A(reg_w_3[14]), .B(n31282), .X(n23009) );
  nand_x1_sg U58158 ( .A(w_3[16]), .B(n29877), .X(n23014) );
  nand_x1_sg U58159 ( .A(reg_w_3[16]), .B(n32957), .X(n23013) );
  nand_x1_sg U58160 ( .A(w_3[17]), .B(n33245), .X(n23016) );
  nand_x1_sg U58161 ( .A(reg_w_3[17]), .B(n33260), .X(n23015) );
  nand_x1_sg U58162 ( .A(w_3[19]), .B(n30824), .X(n23020) );
  nand_x1_sg U58163 ( .A(reg_w_3[19]), .B(n34471), .X(n23019) );
  nand_x1_sg U58164 ( .A(w_4[0]), .B(n34918), .X(n23022) );
  nand_x1_sg U58165 ( .A(reg_w_4[0]), .B(n34930), .X(n23021) );
  nand_x1_sg U58166 ( .A(w_4[2]), .B(n33246), .X(n23026) );
  nand_x1_sg U58167 ( .A(reg_w_4[2]), .B(n31955), .X(n23025) );
  nand_x1_sg U58168 ( .A(w_4[3]), .B(n34920), .X(n23028) );
  nand_x1_sg U58169 ( .A(reg_w_4[3]), .B(n31003), .X(n23027) );
  nand_x1_sg U58170 ( .A(w_4[5]), .B(n31944), .X(n23032) );
  nand_x1_sg U58171 ( .A(reg_w_4[5]), .B(n31962), .X(n23031) );
  nand_x1_sg U58172 ( .A(w_4[6]), .B(n32179), .X(n23034) );
  nand_x1_sg U58173 ( .A(reg_w_4[6]), .B(n30814), .X(n23033) );
  nand_x1_sg U58174 ( .A(w_4[8]), .B(n34489), .X(n23038) );
  nand_x1_sg U58175 ( .A(reg_w_4[8]), .B(n31951), .X(n23037) );
  nand_x1_sg U58176 ( .A(w_4[9]), .B(n34921), .X(n23040) );
  nand_x1_sg U58177 ( .A(reg_w_4[9]), .B(n30822), .X(n23039) );
  nand_x1_sg U58178 ( .A(w_4[11]), .B(n32942), .X(n23044) );
  nand_x1_sg U58179 ( .A(reg_w_4[11]), .B(n30814), .X(n23043) );
  nand_x1_sg U58180 ( .A(w_4[12]), .B(n33233), .X(n23046) );
  nand_x1_sg U58181 ( .A(reg_w_4[12]), .B(n34472), .X(n23045) );
  nand_x1_sg U58182 ( .A(w_4[14]), .B(n30616), .X(n23050) );
  nand_x1_sg U58183 ( .A(reg_w_4[14]), .B(n34532), .X(n23049) );
  nand_x1_sg U58184 ( .A(w_4[15]), .B(n31258), .X(n23052) );
  nand_x1_sg U58185 ( .A(reg_w_4[15]), .B(n33272), .X(n23051) );
  nand_x1_sg U58186 ( .A(w_4[17]), .B(n34839), .X(n23056) );
  nand_x1_sg U58187 ( .A(reg_w_4[17]), .B(n35057), .X(n23055) );
  nand_x1_sg U58188 ( .A(w_4[18]), .B(n33240), .X(n23058) );
  nand_x1_sg U58189 ( .A(reg_w_4[18]), .B(n34821), .X(n23057) );
  nand_x1_sg U58190 ( .A(w_5[0]), .B(n31106), .X(n23062) );
  nand_x1_sg U58191 ( .A(reg_w_5[0]), .B(n31927), .X(n23061) );
  nand_x1_sg U58192 ( .A(w_5[1]), .B(n34459), .X(n23064) );
  nand_x1_sg U58193 ( .A(reg_w_5[1]), .B(n34925), .X(n23063) );
  nand_x1_sg U58194 ( .A(w_5[3]), .B(n34845), .X(n23068) );
  nand_x1_sg U58195 ( .A(reg_w_5[3]), .B(n32080), .X(n23067) );
  nand_x1_sg U58196 ( .A(w_5[4]), .B(n33238), .X(n23070) );
  nand_x1_sg U58197 ( .A(reg_w_5[4]), .B(n32969), .X(n23069) );
  nand_x1_sg U58198 ( .A(w_5[6]), .B(n31969), .X(n23074) );
  nand_x1_sg U58199 ( .A(reg_w_5[6]), .B(n34522), .X(n23073) );
  nand_x1_sg U58200 ( .A(w_5[7]), .B(n34935), .X(n23076) );
  nand_x1_sg U58201 ( .A(reg_w_5[7]), .B(n32966), .X(n23075) );
  nand_x1_sg U58202 ( .A(w_5[9]), .B(n31950), .X(n23080) );
  nand_x1_sg U58203 ( .A(reg_w_5[9]), .B(n34466), .X(n23079) );
  nand_x1_sg U58204 ( .A(w_5[10]), .B(n33222), .X(n23082) );
  nand_x1_sg U58205 ( .A(reg_w_5[10]), .B(n34472), .X(n23081) );
  nand_x1_sg U58206 ( .A(w_5[12]), .B(n32943), .X(n23086) );
  nand_x1_sg U58207 ( .A(reg_w_5[12]), .B(n30129), .X(n23085) );
  nand_x1_sg U58208 ( .A(w_5[13]), .B(n30801), .X(n23088) );
  nand_x1_sg U58209 ( .A(reg_w_5[13]), .B(n31285), .X(n23087) );
  nand_x1_sg U58210 ( .A(w_5[15]), .B(n35052), .X(n23092) );
  nand_x1_sg U58211 ( .A(reg_w_5[15]), .B(n34508), .X(n23091) );
  nand_x1_sg U58212 ( .A(w_5[16]), .B(n31106), .X(n23094) );
  nand_x1_sg U58213 ( .A(reg_w_5[16]), .B(n30814), .X(n23093) );
  nand_x1_sg U58214 ( .A(w_5[18]), .B(n30813), .X(n23098) );
  nand_x1_sg U58215 ( .A(reg_w_5[18]), .B(n31481), .X(n23097) );
  nand_x1_sg U58216 ( .A(w_5[19]), .B(n31105), .X(n23100) );
  nand_x1_sg U58217 ( .A(reg_w_5[19]), .B(n32968), .X(n23099) );
  nand_x1_sg U58218 ( .A(w_6[1]), .B(n29901), .X(n23104) );
  nand_x1_sg U58219 ( .A(reg_w_6[1]), .B(n31210), .X(n23103) );
  nand_x1_sg U58220 ( .A(w_6[2]), .B(n31973), .X(n23106) );
  nand_x1_sg U58221 ( .A(reg_w_6[2]), .B(n31951), .X(n23105) );
  nand_x1_sg U58222 ( .A(w_6[4]), .B(n32179), .X(n23110) );
  nand_x1_sg U58223 ( .A(reg_w_6[4]), .B(n29905), .X(n23109) );
  nand_x1_sg U58224 ( .A(w_6[5]), .B(n31937), .X(n23112) );
  nand_x1_sg U58225 ( .A(reg_w_6[5]), .B(n31285), .X(n23111) );
  nand_x1_sg U58226 ( .A(w_6[7]), .B(n31963), .X(n23116) );
  nand_x1_sg U58227 ( .A(reg_w_6[7]), .B(n34526), .X(n23115) );
  nand_x1_sg U58228 ( .A(w_6[8]), .B(n30801), .X(n23118) );
  nand_x1_sg U58229 ( .A(reg_w_6[8]), .B(n34928), .X(n23117) );
  nand_x1_sg U58230 ( .A(w_6[10]), .B(n31948), .X(n23122) );
  nand_x1_sg U58231 ( .A(reg_w_6[10]), .B(n33260), .X(n23121) );
  nand_x1_sg U58232 ( .A(w_6[11]), .B(n33246), .X(n23124) );
  nand_x1_sg U58233 ( .A(reg_w_6[11]), .B(n31277), .X(n23123) );
  nand_x1_sg U58234 ( .A(w_6[13]), .B(n34455), .X(n23128) );
  nand_x1_sg U58235 ( .A(reg_w_6[13]), .B(n30820), .X(n23127) );
  nand_x1_sg U58236 ( .A(w_6[14]), .B(n31936), .X(n23130) );
  nand_x1_sg U58237 ( .A(reg_w_6[14]), .B(n33263), .X(n23129) );
  nand_x1_sg U58238 ( .A(w_6[16]), .B(n31967), .X(n23134) );
  nand_x1_sg U58239 ( .A(reg_w_6[16]), .B(n34528), .X(n23133) );
  nand_x1_sg U58240 ( .A(w_6[17]), .B(n34834), .X(n23136) );
  nand_x1_sg U58241 ( .A(reg_w_6[17]), .B(n32075), .X(n23135) );
  nand_x1_sg U58242 ( .A(w_6[19]), .B(n34478), .X(n23140) );
  nand_x1_sg U58243 ( .A(reg_w_6[19]), .B(n32979), .X(n23139) );
  nand_x1_sg U58244 ( .A(w_7[0]), .B(n31969), .X(n23142) );
  nand_x1_sg U58245 ( .A(reg_w_7[0]), .B(n31956), .X(n23141) );
  nand_x1_sg U58246 ( .A(w_7[2]), .B(n29877), .X(n23146) );
  nand_x1_sg U58247 ( .A(reg_w_7[2]), .B(n33272), .X(n23145) );
  nand_x1_sg U58248 ( .A(w_7[3]), .B(n35053), .X(n23148) );
  nand_x1_sg U58249 ( .A(reg_w_7[3]), .B(n29754), .X(n23147) );
  nand_x1_sg U58250 ( .A(w_7[5]), .B(n34838), .X(n23152) );
  nand_x1_sg U58251 ( .A(reg_w_7[5]), .B(n34931), .X(n23151) );
  nand_x1_sg U58252 ( .A(w_7[6]), .B(n30193), .X(n23154) );
  nand_x1_sg U58253 ( .A(reg_w_7[6]), .B(n30191), .X(n23153) );
  nand_x1_sg U58254 ( .A(w_7[8]), .B(n31627), .X(n23158) );
  nand_x1_sg U58255 ( .A(reg_w_7[8]), .B(n32072), .X(n23157) );
  nand_x1_sg U58256 ( .A(w_7[9]), .B(n34934), .X(n23160) );
  nand_x1_sg U58257 ( .A(reg_w_7[9]), .B(n31285), .X(n23159) );
  nand_x1_sg U58258 ( .A(w_7[11]), .B(n33227), .X(n23164) );
  nand_x1_sg U58259 ( .A(reg_w_7[11]), .B(n35059), .X(n23163) );
  nand_x1_sg U58260 ( .A(w_7[12]), .B(n34837), .X(n23166) );
  nand_x1_sg U58261 ( .A(reg_w_7[12]), .B(n31007), .X(n23165) );
  nand_x1_sg U58262 ( .A(w_7[14]), .B(n34486), .X(n23170) );
  nand_x1_sg U58263 ( .A(reg_w_7[14]), .B(n34511), .X(n23169) );
  nand_x1_sg U58264 ( .A(w_7[15]), .B(n33258), .X(n23172) );
  nand_x1_sg U58265 ( .A(reg_w_7[15]), .B(n32091), .X(n23171) );
  nand_x1_sg U58266 ( .A(w_7[17]), .B(n34454), .X(n23176) );
  nand_x1_sg U58267 ( .A(reg_w_7[17]), .B(n31958), .X(n23175) );
  nand_x1_sg U58268 ( .A(w_7[18]), .B(n34844), .X(n23178) );
  nand_x1_sg U58269 ( .A(reg_w_7[18]), .B(n34814), .X(n23177) );
  nand_x1_sg U58270 ( .A(w_8[0]), .B(n29898), .X(n23182) );
  nand_x1_sg U58271 ( .A(reg_w_8[0]), .B(n33266), .X(n23181) );
  nand_x1_sg U58272 ( .A(w_8[1]), .B(n34838), .X(n23184) );
  nand_x1_sg U58273 ( .A(reg_w_8[1]), .B(n31277), .X(n23183) );
  nand_x1_sg U58274 ( .A(w_8[3]), .B(n34461), .X(n23188) );
  nand_x1_sg U58275 ( .A(reg_w_8[3]), .B(n34530), .X(n23187) );
  nand_x1_sg U58276 ( .A(w_8[4]), .B(n33256), .X(n23190) );
  nand_x1_sg U58277 ( .A(reg_w_8[4]), .B(n34816), .X(n23189) );
  nand_x1_sg U58278 ( .A(w_8[6]), .B(n34840), .X(n23194) );
  nand_x1_sg U58279 ( .A(reg_w_8[6]), .B(n30378), .X(n23193) );
  nand_x1_sg U58280 ( .A(w_8[7]), .B(n32943), .X(n23196) );
  nand_x1_sg U58281 ( .A(reg_w_8[7]), .B(n32980), .X(n23195) );
  nand_x1_sg U58282 ( .A(w_8[9]), .B(n31937), .X(n23200) );
  nand_x1_sg U58283 ( .A(reg_w_8[9]), .B(n33263), .X(n23199) );
  nand_x1_sg U58284 ( .A(w_8[10]), .B(n34839), .X(n23202) );
  nand_x1_sg U58285 ( .A(reg_w_8[10]), .B(n34530), .X(n23201) );
  nand_x1_sg U58286 ( .A(w_8[12]), .B(n33242), .X(n23206) );
  nand_x1_sg U58287 ( .A(reg_w_8[12]), .B(n32971), .X(n23205) );
  nand_x1_sg U58288 ( .A(w_8[13]), .B(n33230), .X(n23208) );
  nand_x1_sg U58289 ( .A(reg_w_8[13]), .B(n30815), .X(n23207) );
  nand_x1_sg U58290 ( .A(w_8[15]), .B(n34505), .X(n23212) );
  nand_x1_sg U58291 ( .A(reg_w_8[15]), .B(n31007), .X(n23211) );
  nand_x1_sg U58292 ( .A(w_8[16]), .B(n35054), .X(n23214) );
  nand_x1_sg U58293 ( .A(reg_w_8[16]), .B(n32091), .X(n23213) );
  nand_x1_sg U58294 ( .A(w_8[18]), .B(n32947), .X(n23218) );
  nand_x1_sg U58295 ( .A(reg_w_8[18]), .B(n34531), .X(n23217) );
  nand_x1_sg U58296 ( .A(w_8[19]), .B(n31106), .X(n23220) );
  nand_x1_sg U58297 ( .A(reg_w_8[19]), .B(n33261), .X(n23219) );
  nand_x1_sg U58298 ( .A(w_9[1]), .B(n30832), .X(n23224) );
  nand_x1_sg U58299 ( .A(reg_w_9[1]), .B(n33273), .X(n23223) );
  nand_x1_sg U58300 ( .A(w_9[2]), .B(n30792), .X(n23226) );
  nand_x1_sg U58301 ( .A(reg_w_9[2]), .B(n32087), .X(n23225) );
  nand_x1_sg U58302 ( .A(w_9[4]), .B(n34484), .X(n23230) );
  nand_x1_sg U58303 ( .A(reg_w_9[4]), .B(n32084), .X(n23229) );
  nand_x1_sg U58304 ( .A(w_9[5]), .B(n30809), .X(n23232) );
  nand_x1_sg U58305 ( .A(reg_w_9[5]), .B(n30373), .X(n23231) );
  nand_x1_sg U58306 ( .A(w_9[7]), .B(n30192), .X(n23236) );
  nand_x1_sg U58307 ( .A(reg_w_9[7]), .B(n35057), .X(n23235) );
  nand_x1_sg U58308 ( .A(w_9[8]), .B(n29891), .X(n23238) );
  nand_x1_sg U58309 ( .A(reg_w_9[8]), .B(n30368), .X(n23237) );
  nand_x1_sg U58310 ( .A(w_9[10]), .B(n33233), .X(n23242) );
  nand_x1_sg U58311 ( .A(reg_w_9[10]), .B(n31103), .X(n23241) );
  nand_x1_sg U58312 ( .A(w_9[11]), .B(n32944), .X(n23244) );
  nand_x1_sg U58313 ( .A(reg_w_9[11]), .B(n34472), .X(n23243) );
  nand_x1_sg U58314 ( .A(w_9[13]), .B(n34455), .X(n23248) );
  nand_x1_sg U58315 ( .A(reg_w_9[13]), .B(n31928), .X(n23247) );
  nand_x1_sg U58316 ( .A(w_9[14]), .B(n33256), .X(n23250) );
  nand_x1_sg U58317 ( .A(reg_w_9[14]), .B(n31016), .X(n23249) );
  nand_x1_sg U58318 ( .A(w_9[16]), .B(n34933), .X(n23254) );
  nand_x1_sg U58319 ( .A(reg_w_9[16]), .B(n32971), .X(n23253) );
  nand_x1_sg U58320 ( .A(w_9[17]), .B(n34833), .X(n23256) );
  nand_x1_sg U58321 ( .A(reg_w_9[17]), .B(n32090), .X(n23255) );
  nand_x1_sg U58322 ( .A(w_9[19]), .B(n29903), .X(n23260) );
  nand_x1_sg U58323 ( .A(reg_w_9[19]), .B(n30820), .X(n23259) );
  nand_x1_sg U58324 ( .A(w_10[0]), .B(n33228), .X(n23262) );
  nand_x1_sg U58325 ( .A(reg_w_10[0]), .B(n31238), .X(n23261) );
  nand_x1_sg U58326 ( .A(w_10[2]), .B(n31970), .X(n23266) );
  nand_x1_sg U58327 ( .A(reg_w_10[2]), .B(n29905), .X(n23265) );
  nand_x1_sg U58328 ( .A(w_10[3]), .B(n34490), .X(n23268) );
  nand_x1_sg U58329 ( .A(reg_w_10[3]), .B(n32080), .X(n23267) );
  nand_x1_sg U58330 ( .A(w_10[5]), .B(n30803), .X(n23272) );
  nand_x1_sg U58331 ( .A(reg_w_10[5]), .B(n34469), .X(n23271) );
  nand_x1_sg U58332 ( .A(w_10[6]), .B(n30615), .X(n23274) );
  nand_x1_sg U58333 ( .A(reg_w_10[6]), .B(n32974), .X(n23273) );
  nand_x1_sg U58334 ( .A(w_10[8]), .B(n30385), .X(n23278) );
  nand_x1_sg U58335 ( .A(reg_w_10[8]), .B(n33841), .X(n23277) );
  nand_x1_sg U58336 ( .A(w_10[9]), .B(n33252), .X(n23280) );
  nand_x1_sg U58337 ( .A(reg_w_10[9]), .B(n32981), .X(n23279) );
  nand_x1_sg U58338 ( .A(w_10[11]), .B(n31271), .X(n23284) );
  nand_x1_sg U58339 ( .A(reg_w_10[11]), .B(n32950), .X(n23283) );
  nand_x1_sg U58340 ( .A(w_10[12]), .B(n31950), .X(n23286) );
  nand_x1_sg U58341 ( .A(reg_w_10[12]), .B(n32957), .X(n23285) );
  nand_x1_sg U58342 ( .A(w_10[14]), .B(n31263), .X(n23290) );
  nand_x1_sg U58343 ( .A(reg_w_10[14]), .B(n33840), .X(n23289) );
  nand_x1_sg U58344 ( .A(w_10[15]), .B(n30619), .X(n23292) );
  nand_x1_sg U58345 ( .A(reg_w_10[15]), .B(n32078), .X(n23291) );
  nand_x1_sg U58346 ( .A(w_10[17]), .B(n29874), .X(n23296) );
  nand_x1_sg U58347 ( .A(reg_w_10[17]), .B(n30378), .X(n23295) );
  nand_x1_sg U58348 ( .A(w_10[18]), .B(n31964), .X(n23298) );
  nand_x1_sg U58349 ( .A(reg_w_10[18]), .B(n32074), .X(n23297) );
  nand_x1_sg U58350 ( .A(w_11[0]), .B(n31939), .X(n23302) );
  nand_x1_sg U58351 ( .A(reg_w_11[0]), .B(n31290), .X(n23301) );
  nand_x1_sg U58352 ( .A(w_11[1]), .B(n33255), .X(n23304) );
  nand_x1_sg U58353 ( .A(reg_w_11[1]), .B(n32955), .X(n23303) );
  nand_x1_sg U58354 ( .A(w_11[3]), .B(n33224), .X(n23308) );
  nand_x1_sg U58355 ( .A(reg_w_11[3]), .B(n34468), .X(n23307) );
  nand_x1_sg U58356 ( .A(w_11[4]), .B(n29869), .X(n23310) );
  nand_x1_sg U58357 ( .A(reg_w_11[4]), .B(n29798), .X(n23309) );
  nand_x1_sg U58358 ( .A(w_11[6]), .B(n33222), .X(n23314) );
  nand_x1_sg U58359 ( .A(reg_w_11[6]), .B(n29796), .X(n23313) );
  nand_x1_sg U58360 ( .A(w_11[7]), .B(n31938), .X(n23316) );
  nand_x1_sg U58361 ( .A(reg_w_11[7]), .B(n32970), .X(n23315) );
  nand_x1_sg U58362 ( .A(w_11[9]), .B(n34461), .X(n23320) );
  nand_x1_sg U58363 ( .A(reg_w_11[9]), .B(n32081), .X(n23319) );
  nand_x1_sg U58364 ( .A(w_11[10]), .B(n34921), .X(n23322) );
  nand_x1_sg U58365 ( .A(reg_w_11[10]), .B(n34523), .X(n23321) );
  nand_x1_sg U58366 ( .A(w_11[12]), .B(n30805), .X(n23326) );
  nand_x1_sg U58367 ( .A(reg_w_11[12]), .B(n34509), .X(n23325) );
  nand_x1_sg U58368 ( .A(w_11[13]), .B(n30825), .X(n23328) );
  nand_x1_sg U58369 ( .A(reg_w_11[13]), .B(n30788), .X(n23327) );
  nand_x1_sg U58370 ( .A(w_11[15]), .B(n35052), .X(n23332) );
  nand_x1_sg U58371 ( .A(reg_w_11[15]), .B(n29782), .X(n23331) );
  nand_x1_sg U58372 ( .A(w_11[16]), .B(n31263), .X(n23334) );
  nand_x1_sg U58373 ( .A(reg_w_11[16]), .B(n31276), .X(n23333) );
  nand_x1_sg U58374 ( .A(w_11[18]), .B(n32183), .X(n23338) );
  nand_x1_sg U58375 ( .A(reg_w_11[18]), .B(n31957), .X(n23337) );
  nand_x1_sg U58376 ( .A(w_11[19]), .B(n30805), .X(n23340) );
  nand_x1_sg U58377 ( .A(reg_w_11[19]), .B(n32078), .X(n23339) );
  nand_x1_sg U58378 ( .A(w_12[1]), .B(n30829), .X(n23344) );
  nand_x1_sg U58379 ( .A(reg_w_12[1]), .B(n31626), .X(n23343) );
  nand_x1_sg U58380 ( .A(w_12[2]), .B(n34462), .X(n23346) );
  nand_x1_sg U58381 ( .A(reg_w_12[2]), .B(n34527), .X(n23345) );
  nand_x1_sg U58382 ( .A(w_12[4]), .B(n31263), .X(n23350) );
  nand_x1_sg U58383 ( .A(reg_w_12[4]), .B(n34473), .X(n23349) );
  nand_x1_sg U58384 ( .A(w_12[5]), .B(n34842), .X(n23352) );
  nand_x1_sg U58385 ( .A(reg_w_12[5]), .B(n34810), .X(n23351) );
  nand_x1_sg U58386 ( .A(w_12[7]), .B(n31945), .X(n23356) );
  nand_x1_sg U58387 ( .A(reg_w_12[7]), .B(n31480), .X(n23355) );
  nand_x1_sg U58388 ( .A(w_12[8]), .B(n31267), .X(n23358) );
  nand_x1_sg U58389 ( .A(reg_w_12[8]), .B(n33271), .X(n23357) );
  nand_x1_sg U58390 ( .A(w_12[10]), .B(n34835), .X(n23362) );
  nand_x1_sg U58391 ( .A(reg_w_12[10]), .B(n29796), .X(n23361) );
  nand_x1_sg U58392 ( .A(w_12[11]), .B(n30807), .X(n23364) );
  nand_x1_sg U58393 ( .A(reg_w_12[11]), .B(n30815), .X(n23363) );
  nand_x1_sg U58394 ( .A(w_12[13]), .B(n30802), .X(n23368) );
  nand_x1_sg U58395 ( .A(reg_w_12[13]), .B(n32954), .X(n23367) );
  nand_x1_sg U58396 ( .A(w_12[14]), .B(n33251), .X(n23370) );
  nand_x1_sg U58397 ( .A(reg_w_12[14]), .B(n32973), .X(n23369) );
  nand_x1_sg U58398 ( .A(w_12[16]), .B(n30829), .X(n23374) );
  nand_x1_sg U58399 ( .A(reg_w_12[16]), .B(n31955), .X(n23373) );
  nand_x1_sg U58400 ( .A(w_12[17]), .B(n33224), .X(n23376) );
  nand_x1_sg U58401 ( .A(reg_w_12[17]), .B(n31928), .X(n23375) );
  nand_x1_sg U58402 ( .A(w_12[19]), .B(n30809), .X(n23380) );
  nand_x1_sg U58403 ( .A(reg_w_12[19]), .B(n34473), .X(n23379) );
  nand_x1_sg U58404 ( .A(w_13[0]), .B(n31940), .X(n23382) );
  nand_x1_sg U58405 ( .A(reg_w_13[0]), .B(n29906), .X(n23381) );
  nand_x1_sg U58406 ( .A(w_13[2]), .B(n34922), .X(n23386) );
  nand_x1_sg U58407 ( .A(reg_w_13[2]), .B(n32962), .X(n23385) );
  nand_x1_sg U58408 ( .A(w_13[3]), .B(n30382), .X(n23388) );
  nand_x1_sg U58409 ( .A(reg_w_13[3]), .B(n33262), .X(n23387) );
  nand_x1_sg U58410 ( .A(w_13[5]), .B(n34829), .X(n23392) );
  nand_x1_sg U58411 ( .A(reg_w_13[5]), .B(n32952), .X(n23391) );
  nand_x1_sg U58412 ( .A(w_13[6]), .B(n29895), .X(n23394) );
  nand_x1_sg U58413 ( .A(reg_w_13[6]), .B(n29906), .X(n23393) );
  nand_x1_sg U58414 ( .A(w_13[8]), .B(n29872), .X(n23398) );
  nand_x1_sg U58415 ( .A(reg_w_13[8]), .B(n34821), .X(n23397) );
  nand_x1_sg U58416 ( .A(w_13[9]), .B(n34475), .X(n23400) );
  nand_x1_sg U58417 ( .A(reg_w_13[9]), .B(n31011), .X(n23399) );
  nand_x1_sg U58418 ( .A(w_13[11]), .B(n31266), .X(n23404) );
  nand_x1_sg U58419 ( .A(reg_w_13[11]), .B(n34819), .X(n23403) );
  nand_x1_sg U58420 ( .A(w_13[12]), .B(n34843), .X(n23406) );
  nand_x1_sg U58421 ( .A(reg_w_13[12]), .B(n31282), .X(n23405) );
  nand_x1_sg U58422 ( .A(w_13[14]), .B(n30616), .X(n23410) );
  nand_x1_sg U58423 ( .A(reg_w_13[14]), .B(n34532), .X(n23409) );
  nand_x1_sg U58424 ( .A(w_13[15]), .B(n30802), .X(n23412) );
  nand_x1_sg U58425 ( .A(reg_w_13[15]), .B(n34106), .X(n23411) );
  nand_x1_sg U58426 ( .A(w_13[17]), .B(n33916), .X(n23416) );
  nand_x1_sg U58427 ( .A(reg_w_13[17]), .B(n31961), .X(n23415) );
  nand_x1_sg U58428 ( .A(w_13[18]), .B(n30617), .X(n23418) );
  nand_x1_sg U58429 ( .A(reg_w_13[18]), .B(n31012), .X(n23417) );
  nand_x1_sg U58430 ( .A(w_14[0]), .B(n33243), .X(n23422) );
  nand_x1_sg U58431 ( .A(reg_w_14[0]), .B(n31962), .X(n23421) );
  nand_x1_sg U58432 ( .A(w_14[1]), .B(n33247), .X(n23424) );
  nand_x1_sg U58433 ( .A(reg_w_14[1]), .B(n29778), .X(n23423) );
  nand_x1_sg U58434 ( .A(w_14[3]), .B(n34834), .X(n23428) );
  nand_x1_sg U58435 ( .A(reg_w_14[3]), .B(n34815), .X(n23427) );
  nand_x1_sg U58436 ( .A(w_14[4]), .B(n30824), .X(n23430) );
  nand_x1_sg U58437 ( .A(reg_w_14[4]), .B(n32954), .X(n23429) );
  nand_x1_sg U58438 ( .A(w_14[6]), .B(n34488), .X(n23434) );
  nand_x1_sg U58439 ( .A(reg_w_14[6]), .B(n31481), .X(n23433) );
  nand_x1_sg U58440 ( .A(w_14[7]), .B(n31943), .X(n23436) );
  nand_x1_sg U58441 ( .A(reg_w_14[7]), .B(n32071), .X(n23435) );
  nand_x1_sg U58442 ( .A(w_14[9]), .B(n34845), .X(n23440) );
  nand_x1_sg U58443 ( .A(reg_w_14[9]), .B(n34916), .X(n23439) );
  nand_x1_sg U58444 ( .A(w_14[10]), .B(n30793), .X(n23442) );
  nand_x1_sg U58445 ( .A(reg_w_14[10]), .B(n32957), .X(n23441) );
  nand_x1_sg U58446 ( .A(w_14[12]), .B(n34919), .X(n23446) );
  nand_x1_sg U58447 ( .A(reg_w_14[12]), .B(n34818), .X(n23445) );
  nand_x1_sg U58448 ( .A(w_14[13]), .B(n33228), .X(n23448) );
  nand_x1_sg U58449 ( .A(reg_w_14[13]), .B(n31955), .X(n23447) );
  nand_x1_sg U58450 ( .A(w_14[15]), .B(n30620), .X(n23452) );
  nand_x1_sg U58451 ( .A(reg_w_14[15]), .B(n31006), .X(n23451) );
  nand_x1_sg U58452 ( .A(w_14[16]), .B(n33248), .X(n23454) );
  nand_x1_sg U58453 ( .A(reg_w_14[16]), .B(n34105), .X(n23453) );
  nand_x1_sg U58454 ( .A(w_14[18]), .B(n34835), .X(n23458) );
  nand_x1_sg U58455 ( .A(reg_w_14[18]), .B(n30789), .X(n23457) );
  nand_x1_sg U58456 ( .A(w_14[19]), .B(n31257), .X(n23460) );
  nand_x1_sg U58457 ( .A(reg_w_14[19]), .B(n31210), .X(n23459) );
  nand_x1_sg U58458 ( .A(w_15[1]), .B(n30382), .X(n23464) );
  nand_x1_sg U58459 ( .A(reg_w_15[1]), .B(n31103), .X(n23463) );
  nand_x1_sg U58460 ( .A(w_15[2]), .B(n32184), .X(n23466) );
  nand_x1_sg U58461 ( .A(reg_w_15[2]), .B(n31103), .X(n23465) );
  nand_x1_sg U58462 ( .A(w_15[4]), .B(n34832), .X(n23470) );
  nand_x1_sg U58463 ( .A(reg_w_15[4]), .B(n32976), .X(n23469) );
  nand_x1_sg U58464 ( .A(w_15[5]), .B(n31942), .X(n23472) );
  nand_x1_sg U58465 ( .A(reg_w_15[5]), .B(n31237), .X(n23471) );
  nand_x1_sg U58466 ( .A(w_15[7]), .B(n34491), .X(n23476) );
  nand_x1_sg U58467 ( .A(reg_w_15[7]), .B(n32092), .X(n23475) );
  nand_x1_sg U58468 ( .A(w_15[8]), .B(n31099), .X(n23478) );
  nand_x1_sg U58469 ( .A(reg_w_15[8]), .B(n32081), .X(n23477) );
  nand_x1_sg U58470 ( .A(w_15[10]), .B(n33244), .X(n23482) );
  nand_x1_sg U58471 ( .A(reg_w_15[10]), .B(n30823), .X(n23481) );
  nand_x1_sg U58472 ( .A(w_15[11]), .B(n29903), .X(n23484) );
  nand_x1_sg U58473 ( .A(reg_w_15[11]), .B(n32962), .X(n23483) );
  nand_x1_sg U58474 ( .A(w_15[13]), .B(n33258), .X(n23488) );
  nand_x1_sg U58475 ( .A(reg_w_15[13]), .B(n31102), .X(n23487) );
  nand_x1_sg U58476 ( .A(w_15[14]), .B(n33249), .X(n23490) );
  nand_x1_sg U58477 ( .A(reg_w_15[14]), .B(n33271), .X(n23489) );
  nand_x1_sg U58478 ( .A(w_15[16]), .B(n30620), .X(n23494) );
  nand_x1_sg U58479 ( .A(reg_w_15[16]), .B(n34929), .X(n23493) );
  nand_x1_sg U58480 ( .A(w_15[17]), .B(n34489), .X(n23496) );
  nand_x1_sg U58481 ( .A(reg_w_15[17]), .B(n32086), .X(n23495) );
  nand_x1_sg U58482 ( .A(w_15[19]), .B(n34480), .X(n23500) );
  nand_x1_sg U58483 ( .A(reg_w_15[19]), .B(n31211), .X(n23499) );
  nand_x1_sg U58484 ( .A(i_mask[0]), .B(n31937), .X(n23502) );
  nand_x1_sg U58485 ( .A(reg_i_mask[0]), .B(n34522), .X(n23501) );
  nand_x1_sg U58486 ( .A(i_mask[2]), .B(n34489), .X(n23506) );
  nand_x1_sg U58487 ( .A(reg_i_mask[2]), .B(n30370), .X(n23505) );
  nand_x1_sg U58488 ( .A(i_mask[3]), .B(n31974), .X(n23508) );
  nand_x1_sg U58489 ( .A(reg_i_mask[3]), .B(n32082), .X(n23507) );
  nand_x1_sg U58490 ( .A(i_mask[5]), .B(n35054), .X(n23512) );
  nand_x1_sg U58491 ( .A(reg_i_mask[5]), .B(n34523), .X(n23511) );
  nand_x1_sg U58492 ( .A(i_mask[6]), .B(n35055), .X(n23514) );
  nand_x1_sg U58493 ( .A(reg_i_mask[6]), .B(n31480), .X(n23513) );
  nand_x1_sg U58494 ( .A(i_mask[8]), .B(n33249), .X(n23518) );
  nand_x1_sg U58495 ( .A(reg_i_mask[8]), .B(n34928), .X(n23517) );
  nand_x1_sg U58496 ( .A(i_mask[9]), .B(n29893), .X(n23520) );
  nand_x1_sg U58497 ( .A(reg_i_mask[9]), .B(n33262), .X(n23519) );
  nand_x1_sg U58498 ( .A(i_mask[11]), .B(n35054), .X(n23524) );
  nand_x1_sg U58499 ( .A(reg_i_mask[11]), .B(n30613), .X(n23523) );
  nand_x1_sg U58500 ( .A(i_mask[12]), .B(n33251), .X(n23526) );
  nand_x1_sg U58501 ( .A(reg_i_mask[12]), .B(n34474), .X(n23525) );
  nand_x1_sg U58502 ( .A(i_mask[14]), .B(n29887), .X(n23530) );
  nand_x1_sg U58503 ( .A(reg_i_mask[14]), .B(n33267), .X(n23529) );
  nand_x1_sg U58504 ( .A(i_mask[15]), .B(n34488), .X(n23532) );
  nand_x1_sg U58505 ( .A(reg_i_mask[15]), .B(n32975), .X(n23531) );
  nand_x1_sg U58506 ( .A(i_mask[17]), .B(n29872), .X(n23536) );
  nand_x1_sg U58507 ( .A(reg_i_mask[17]), .B(n32964), .X(n23535) );
  nand_x1_sg U58508 ( .A(i_mask[18]), .B(n34475), .X(n23538) );
  nand_x1_sg U58509 ( .A(reg_i_mask[18]), .B(n34809), .X(n23537) );
  nand_x1_sg U58510 ( .A(i_mask[20]), .B(n31623), .X(n23542) );
  nand_x1_sg U58511 ( .A(reg_i_mask[20]), .B(n29784), .X(n23541) );
  nand_x1_sg U58512 ( .A(i_mask[21]), .B(n31964), .X(n23544) );
  nand_x1_sg U58513 ( .A(reg_i_mask[21]), .B(n31957), .X(n23543) );
  nand_x1_sg U58514 ( .A(i_mask[23]), .B(n32942), .X(n23548) );
  nand_x1_sg U58515 ( .A(reg_i_mask[23]), .B(n33271), .X(n23547) );
  nand_x1_sg U58516 ( .A(i_mask[24]), .B(n34834), .X(n23550) );
  nand_x1_sg U58517 ( .A(reg_i_mask[24]), .B(n31952), .X(n23549) );
  nand_x1_sg U58518 ( .A(i_mask[26]), .B(n33253), .X(n23554) );
  nand_x1_sg U58519 ( .A(reg_i_mask[26]), .B(n29786), .X(n23553) );
  nand_x1_sg U58520 ( .A(i_mask[27]), .B(n34451), .X(n23556) );
  nand_x1_sg U58521 ( .A(reg_i_mask[27]), .B(n32077), .X(n23555) );
  nand_x1_sg U58522 ( .A(i_mask[29]), .B(n34830), .X(n23560) );
  nand_x1_sg U58523 ( .A(reg_i_mask[29]), .B(n31210), .X(n23559) );
  nand_x1_sg U58524 ( .A(i_mask[30]), .B(n34451), .X(n23562) );
  nand_x1_sg U58525 ( .A(reg_i_mask[30]), .B(n30368), .X(n23561) );
  nand_x1_sg U58526 ( .A(w_mask[0]), .B(n33233), .X(n23566) );
  nand_x1_sg U58527 ( .A(reg_w_mask[0]), .B(n30376), .X(n23565) );
  nand_x1_sg U58528 ( .A(w_mask[1]), .B(n33248), .X(n23568) );
  nand_x1_sg U58529 ( .A(reg_w_mask[1]), .B(n34812), .X(n23567) );
  nand_x1_sg U58530 ( .A(w_mask[3]), .B(n33235), .X(n23572) );
  nand_x1_sg U58531 ( .A(reg_w_mask[3]), .B(n32088), .X(n23571) );
  nand_x1_sg U58532 ( .A(w_mask[4]), .B(n34481), .X(n23574) );
  nand_x1_sg U58533 ( .A(reg_w_mask[4]), .B(n34467), .X(n23573) );
  nand_x1_sg U58534 ( .A(w_mask[6]), .B(n34839), .X(n23578) );
  nand_x1_sg U58535 ( .A(reg_w_mask[6]), .B(n32959), .X(n23577) );
  nand_x1_sg U58536 ( .A(w_mask[7]), .B(n32179), .X(n23580) );
  nand_x1_sg U58537 ( .A(reg_w_mask[7]), .B(n31102), .X(n23579) );
  nand_x1_sg U58538 ( .A(w_mask[9]), .B(n31939), .X(n23584) );
  nand_x1_sg U58539 ( .A(reg_w_mask[9]), .B(n34527), .X(n23583) );
  nand_x1_sg U58540 ( .A(w_mask[10]), .B(n31272), .X(n23586) );
  nand_x1_sg U58541 ( .A(reg_w_mask[10]), .B(n29788), .X(n23585) );
  nand_x1_sg U58542 ( .A(w_mask[12]), .B(n30616), .X(n23590) );
  nand_x1_sg U58543 ( .A(reg_w_mask[12]), .B(n32072), .X(n23589) );
  nand_x1_sg U58544 ( .A(w_mask[13]), .B(n30832), .X(n23592) );
  nand_x1_sg U58545 ( .A(reg_w_mask[13]), .B(n34820), .X(n23591) );
  nand_x1_sg U58546 ( .A(w_mask[15]), .B(n31262), .X(n23596) );
  nand_x1_sg U58547 ( .A(reg_w_mask[15]), .B(n34825), .X(n23595) );
  nand_x1_sg U58548 ( .A(w_mask[16]), .B(n32182), .X(n23598) );
  nand_x1_sg U58549 ( .A(reg_w_mask[16]), .B(n34469), .X(n23597) );
  nand_x1_sg U58550 ( .A(w_mask[18]), .B(n34843), .X(n23602) );
  nand_x1_sg U58551 ( .A(reg_w_mask[18]), .B(n34522), .X(n23601) );
  nand_x1_sg U58552 ( .A(w_mask[19]), .B(n34840), .X(n23604) );
  nand_x1_sg U58553 ( .A(reg_w_mask[19]), .B(n32978), .X(n23603) );
  nand_x1_sg U58554 ( .A(w_mask[21]), .B(n34827), .X(n23608) );
  nand_x1_sg U58555 ( .A(reg_w_mask[21]), .B(n34811), .X(n23607) );
  nand_x1_sg U58556 ( .A(w_mask[22]), .B(n30612), .X(n23610) );
  nand_x1_sg U58557 ( .A(reg_w_mask[22]), .B(n32967), .X(n23609) );
  nand_x1_sg U58558 ( .A(w_mask[24]), .B(n31624), .X(n23614) );
  nand_x1_sg U58559 ( .A(reg_w_mask[24]), .B(n35057), .X(n23613) );
  nand_x1_sg U58560 ( .A(w_mask[25]), .B(n33243), .X(n23616) );
  nand_x1_sg U58561 ( .A(reg_w_mask[25]), .B(n30818), .X(n23615) );
  nand_x1_sg U58562 ( .A(w_mask[27]), .B(n31974), .X(n23620) );
  nand_x1_sg U58563 ( .A(reg_w_mask[27]), .B(n34814), .X(n23619) );
  nand_x1_sg U58564 ( .A(w_mask[28]), .B(n29881), .X(n23622) );
  nand_x1_sg U58565 ( .A(reg_w_mask[28]), .B(n32956), .X(n23621) );
  nand_x1_sg U58566 ( .A(w_mask[30]), .B(n33243), .X(n23626) );
  nand_x1_sg U58567 ( .A(reg_w_mask[30]), .B(n33265), .X(n23625) );
  nand_x1_sg U58568 ( .A(w_mask[31]), .B(n34832), .X(n23628) );
  nand_x1_sg U58569 ( .A(reg_w_mask[31]), .B(n34816), .X(n23627) );
  inv_x1_sg U58570 ( .A(filter_input_ready), .X(n42413) );
  nor_x1_sg U58571 ( .A(n30200), .B(\shifter_0/pointer[1] ), .X(n19590) );
  nor_x1_sg U58572 ( .A(n34860), .B(\shifter_0/pointer[1] ), .X(n19589) );
  nand_x1_sg U58573 ( .A(filter_state[0]), .B(n42531), .X(n26587) );
  nand_x1_sg U58574 ( .A(reg_ow_15[19]), .B(n33070), .X(n20891) );
  nand_x1_sg U58575 ( .A(n34744), .B(\shifter_0/reg_w_15[19] ), .X(n20892) );
  nand_x1_sg U58576 ( .A(reg_ow_15[18]), .B(n33131), .X(n20889) );
  nand_x1_sg U58577 ( .A(n32676), .B(\shifter_0/reg_w_15[18] ), .X(n20890) );
  nand_x1_sg U58578 ( .A(reg_ow_15[15]), .B(n35043), .X(n20883) );
  nand_x1_sg U58579 ( .A(n34803), .B(\shifter_0/reg_w_15[15] ), .X(n20884) );
  nand_x1_sg U58580 ( .A(reg_ow_15[14]), .B(n35041), .X(n20881) );
  nand_x1_sg U58581 ( .A(n34109), .B(\shifter_0/reg_w_15[14] ), .X(n20882) );
  nand_x1_sg U58582 ( .A(reg_ow_15[13]), .B(n33095), .X(n20879) );
  nand_x1_sg U58583 ( .A(n32640), .B(\shifter_0/reg_w_15[13] ), .X(n20880) );
  nand_x1_sg U58584 ( .A(reg_ow_15[10]), .B(n29831), .X(n20873) );
  nand_x1_sg U58585 ( .A(n30641), .B(\shifter_0/reg_w_15[10] ), .X(n20874) );
  nand_x1_sg U58586 ( .A(reg_ow_15[7]), .B(n33044), .X(n20867) );
  nand_x1_sg U58587 ( .A(n34804), .B(\shifter_0/reg_w_15[7] ), .X(n20868) );
  nand_x1_sg U58588 ( .A(reg_ow_15[4]), .B(n33098), .X(n20861) );
  nand_x1_sg U58589 ( .A(n32706), .B(\shifter_0/reg_w_15[4] ), .X(n20862) );
  nand_x1_sg U58590 ( .A(reg_ow_15[1]), .B(n29836), .X(n20855) );
  nand_x1_sg U58591 ( .A(n34111), .B(\shifter_0/reg_w_15[1] ), .X(n20856) );
  nand_x1_sg U58592 ( .A(reg_ow_15[0]), .B(n35047), .X(n20853) );
  nand_x1_sg U58593 ( .A(n31235), .B(\shifter_0/reg_w_15[0] ), .X(n20854) );
  nand_x1_sg U58594 ( .A(reg_ow_3[19]), .B(n33057), .X(n20411) );
  nand_x1_sg U58595 ( .A(n32671), .B(\shifter_0/reg_w_3[19] ), .X(n20412) );
  nand_x1_sg U58596 ( .A(reg_ow_3[16]), .B(n33059), .X(n20405) );
  nand_x1_sg U58597 ( .A(n32658), .B(\shifter_0/reg_w_3[16] ), .X(n20406) );
  nand_x1_sg U58598 ( .A(reg_ow_3[15]), .B(n31572), .X(n20403) );
  nand_x1_sg U58599 ( .A(n32527), .B(\shifter_0/reg_w_3[15] ), .X(n20404) );
  nand_x1_sg U58600 ( .A(reg_ow_3[14]), .B(n29799), .X(n20401) );
  nand_x1_sg U58601 ( .A(n34415), .B(\shifter_0/reg_w_3[14] ), .X(n20402) );
  nand_x1_sg U58602 ( .A(reg_ow_3[11]), .B(n31580), .X(n20395) );
  nand_x1_sg U58603 ( .A(n31485), .B(\shifter_0/reg_w_3[11] ), .X(n20396) );
  nand_x1_sg U58604 ( .A(reg_ow_3[10]), .B(n30602), .X(n20393) );
  nand_x1_sg U58605 ( .A(n30688), .B(\shifter_0/reg_w_3[10] ), .X(n20394) );
  nand_x1_sg U58606 ( .A(reg_ow_3[7]), .B(n33099), .X(n20387) );
  nand_x1_sg U58607 ( .A(n32676), .B(\shifter_0/reg_w_3[7] ), .X(n20388) );
  nand_x1_sg U58608 ( .A(reg_ow_3[6]), .B(n33065), .X(n20385) );
  nand_x1_sg U58609 ( .A(n34968), .B(\shifter_0/reg_w_3[6] ), .X(n20386) );
  nand_x1_sg U58610 ( .A(reg_ow_3[5]), .B(n33082), .X(n20383) );
  nand_x1_sg U58611 ( .A(n34729), .B(\shifter_0/reg_w_3[5] ), .X(n20384) );
  nand_x1_sg U58612 ( .A(reg_ow_3[2]), .B(n33100), .X(n20377) );
  nand_x1_sg U58613 ( .A(n30697), .B(\shifter_0/reg_w_3[2] ), .X(n20378) );
  nand_x1_sg U58614 ( .A(reg_ow_3[1]), .B(n33050), .X(n20375) );
  nand_x1_sg U58615 ( .A(n32526), .B(\shifter_0/reg_w_3[1] ), .X(n20376) );
  nand_x1_sg U58616 ( .A(reg_ow_3[0]), .B(n35030), .X(n20373) );
  nand_x1_sg U58617 ( .A(n32660), .B(\shifter_0/reg_w_3[0] ), .X(n20374) );
  nand_x1_sg U58618 ( .A(reg_oi_15[19]), .B(n33063), .X(n20251) );
  nand_x1_sg U58619 ( .A(n34730), .B(\shifter_0/reg_i_15[19] ), .X(n20252) );
  nand_x1_sg U58620 ( .A(reg_oi_15[15]), .B(n33092), .X(n20243) );
  nand_x1_sg U58621 ( .A(n32685), .B(\shifter_0/reg_i_15[15] ), .X(n20244) );
  nand_x1_sg U58622 ( .A(reg_oi_15[14]), .B(n33089), .X(n20241) );
  nand_x1_sg U58623 ( .A(n32903), .B(\shifter_0/reg_i_15[14] ), .X(n20242) );
  nand_x1_sg U58624 ( .A(reg_oi_15[13]), .B(n33110), .X(n20239) );
  nand_x1_sg U58625 ( .A(n34744), .B(\shifter_0/reg_i_15[13] ), .X(n20240) );
  nand_x1_sg U58626 ( .A(reg_oi_15[10]), .B(n33102), .X(n20233) );
  nand_x1_sg U58627 ( .A(n34966), .B(\shifter_0/reg_i_15[10] ), .X(n20234) );
  nand_x1_sg U58628 ( .A(reg_oi_15[7]), .B(n33083), .X(n20227) );
  nand_x1_sg U58629 ( .A(n34733), .B(\shifter_0/reg_i_15[7] ), .X(n20228) );
  nand_x1_sg U58630 ( .A(reg_oi_15[1]), .B(n31562), .X(n20215) );
  nand_x1_sg U58631 ( .A(n34731), .B(\shifter_0/reg_i_15[1] ), .X(n20216) );
  nand_x1_sg U58632 ( .A(reg_oi_15[0]), .B(n35017), .X(n20213) );
  nand_x1_sg U58633 ( .A(n32704), .B(\shifter_0/reg_i_15[0] ), .X(n20214) );
  nand_x1_sg U58634 ( .A(reg_oi_3[19]), .B(n35022), .X(n19771) );
  nand_x1_sg U58635 ( .A(n31482), .B(\shifter_0/reg_i_3[19] ), .X(n19772) );
  nand_x1_sg U58636 ( .A(reg_oi_3[16]), .B(n33061), .X(n19765) );
  nand_x1_sg U58637 ( .A(n32527), .B(\shifter_0/reg_i_3[16] ), .X(n19766) );
  nand_x1_sg U58638 ( .A(reg_oi_3[15]), .B(n31571), .X(n19763) );
  nand_x1_sg U58639 ( .A(n34099), .B(\shifter_0/reg_i_3[15] ), .X(n19764) );
  nand_x1_sg U58640 ( .A(reg_oi_3[14]), .B(n29804), .X(n19761) );
  nand_x1_sg U58641 ( .A(n32654), .B(\shifter_0/reg_i_3[14] ), .X(n19762) );
  nand_x1_sg U58642 ( .A(reg_oi_3[11]), .B(n33822), .X(n19755) );
  nand_x1_sg U58643 ( .A(n32639), .B(\shifter_0/reg_i_3[11] ), .X(n19756) );
  nand_x1_sg U58644 ( .A(reg_oi_3[10]), .B(n33057), .X(n19753) );
  nand_x1_sg U58645 ( .A(n31859), .B(\shifter_0/reg_i_3[10] ), .X(n19754) );
  nand_x1_sg U58646 ( .A(reg_oi_3[7]), .B(n33074), .X(n19747) );
  nand_x1_sg U58647 ( .A(n32666), .B(\shifter_0/reg_i_3[7] ), .X(n19748) );
  nand_x1_sg U58648 ( .A(reg_oi_3[6]), .B(n31587), .X(n19745) );
  nand_x1_sg U58649 ( .A(n34727), .B(\shifter_0/reg_i_3[6] ), .X(n19746) );
  nand_x1_sg U58650 ( .A(reg_oi_3[5]), .B(n31578), .X(n19743) );
  nand_x1_sg U58651 ( .A(n34749), .B(\shifter_0/reg_i_3[5] ), .X(n19744) );
  nand_x1_sg U58652 ( .A(reg_oi_3[2]), .B(n31215), .X(n19737) );
  nand_x1_sg U58653 ( .A(n32902), .B(\shifter_0/reg_i_3[2] ), .X(n19738) );
  nand_x1_sg U58654 ( .A(reg_oi_3[1]), .B(n33100), .X(n19735) );
  nand_x1_sg U58655 ( .A(n32680), .B(\shifter_0/reg_i_3[1] ), .X(n19736) );
  nand_x1_sg U58656 ( .A(reg_oi_3[0]), .B(n33066), .X(n19733) );
  nand_x1_sg U58657 ( .A(n30854), .B(\shifter_0/reg_i_3[0] ), .X(n19734) );
  nand_x1_sg U58658 ( .A(reg_ow_8[19]), .B(n35024), .X(n20611) );
  nand_x1_sg U58659 ( .A(n34743), .B(\shifter_0/reg_w_8[19] ), .X(n20612) );
  nand_x1_sg U58660 ( .A(reg_ow_8[18]), .B(n29810), .X(n20609) );
  nand_x1_sg U58661 ( .A(n31488), .B(\shifter_0/reg_w_8[18] ), .X(n20610) );
  nand_x1_sg U58662 ( .A(reg_ow_8[17]), .B(n31580), .X(n20607) );
  nand_x1_sg U58663 ( .A(n34098), .B(\shifter_0/reg_w_8[17] ), .X(n20608) );
  nand_x1_sg U58664 ( .A(reg_ow_8[16]), .B(n31569), .X(n20605) );
  nand_x1_sg U58665 ( .A(n31487), .B(\shifter_0/reg_w_8[16] ), .X(n20606) );
  nand_x1_sg U58666 ( .A(reg_ow_8[15]), .B(n35045), .X(n20603) );
  nand_x1_sg U58667 ( .A(n30216), .B(\shifter_0/reg_w_8[15] ), .X(n20604) );
  nand_x1_sg U58668 ( .A(reg_ow_8[14]), .B(n33119), .X(n20601) );
  nand_x1_sg U58669 ( .A(n34108), .B(\shifter_0/reg_w_8[14] ), .X(n20602) );
  nand_x1_sg U58670 ( .A(reg_ow_8[13]), .B(n33124), .X(n20599) );
  nand_x1_sg U58671 ( .A(n34101), .B(\shifter_0/reg_w_8[13] ), .X(n20600) );
  nand_x1_sg U58672 ( .A(reg_ow_8[12]), .B(n33044), .X(n20597) );
  nand_x1_sg U58673 ( .A(n30689), .B(\shifter_0/reg_w_8[12] ), .X(n20598) );
  nand_x1_sg U58674 ( .A(reg_ow_8[11]), .B(n33054), .X(n20595) );
  nand_x1_sg U58675 ( .A(n34104), .B(\shifter_0/reg_w_8[11] ), .X(n20596) );
  nand_x1_sg U58676 ( .A(reg_ow_8[10]), .B(n35041), .X(n20593) );
  nand_x1_sg U58677 ( .A(n31860), .B(\shifter_0/reg_w_8[10] ), .X(n20594) );
  nand_x1_sg U58678 ( .A(reg_ow_8[9]), .B(n35024), .X(n20591) );
  nand_x1_sg U58679 ( .A(n30640), .B(\shifter_0/reg_w_8[9] ), .X(n20592) );
  nand_x1_sg U58680 ( .A(reg_ow_8[8]), .B(n35039), .X(n20589) );
  nand_x1_sg U58681 ( .A(n32673), .B(\shifter_0/reg_w_8[8] ), .X(n20590) );
  nand_x1_sg U58682 ( .A(reg_ow_8[7]), .B(n33077), .X(n20587) );
  nand_x1_sg U58683 ( .A(n32521), .B(\shifter_0/reg_w_8[7] ), .X(n20588) );
  nand_x1_sg U58684 ( .A(reg_ow_8[6]), .B(n35019), .X(n20585) );
  nand_x1_sg U58685 ( .A(n32693), .B(\shifter_0/reg_w_8[6] ), .X(n20586) );
  nand_x1_sg U58686 ( .A(reg_ow_8[5]), .B(n31567), .X(n20583) );
  nand_x1_sg U58687 ( .A(n34965), .B(\shifter_0/reg_w_8[5] ), .X(n20584) );
  nand_x1_sg U58688 ( .A(reg_ow_8[4]), .B(n33090), .X(n20581) );
  nand_x1_sg U58689 ( .A(n32681), .B(\shifter_0/reg_w_8[4] ), .X(n20582) );
  nand_x1_sg U58690 ( .A(reg_ow_8[3]), .B(n33078), .X(n20579) );
  nand_x1_sg U58691 ( .A(n32700), .B(\shifter_0/reg_w_8[3] ), .X(n20580) );
  nand_x1_sg U58692 ( .A(reg_ow_8[2]), .B(n35025), .X(n20577) );
  nand_x1_sg U58693 ( .A(n34102), .B(\shifter_0/reg_w_8[2] ), .X(n20578) );
  nand_x1_sg U58694 ( .A(reg_ow_8[1]), .B(n29807), .X(n20575) );
  nand_x1_sg U58695 ( .A(n31485), .B(\shifter_0/reg_w_8[1] ), .X(n20576) );
  nand_x1_sg U58696 ( .A(reg_ow_8[0]), .B(n31571), .X(n20573) );
  nand_x1_sg U58697 ( .A(n32693), .B(\shifter_0/reg_w_8[0] ), .X(n20574) );
  nand_x1_sg U58698 ( .A(reg_oi_8[19]), .B(n33053), .X(n19971) );
  nand_x1_sg U58699 ( .A(n31988), .B(\shifter_0/reg_i_8[19] ), .X(n19972) );
  nand_x1_sg U58700 ( .A(reg_oi_8[16]), .B(n33095), .X(n19965) );
  nand_x1_sg U58701 ( .A(n32526), .B(\shifter_0/reg_i_8[16] ), .X(n19966) );
  nand_x1_sg U58702 ( .A(reg_oi_8[15]), .B(n31576), .X(n19963) );
  nand_x1_sg U58703 ( .A(n30681), .B(\shifter_0/reg_i_8[15] ), .X(n19964) );
  nand_x1_sg U58704 ( .A(reg_oi_8[14]), .B(n33131), .X(n19961) );
  nand_x1_sg U58705 ( .A(n34743), .B(\shifter_0/reg_i_8[14] ), .X(n19962) );
  nand_x1_sg U58706 ( .A(reg_oi_8[13]), .B(n29829), .X(n19959) );
  nand_x1_sg U58707 ( .A(n31985), .B(\shifter_0/reg_i_8[13] ), .X(n19960) );
  nand_x1_sg U58708 ( .A(reg_oi_8[12]), .B(n31213), .X(n19957) );
  nand_x1_sg U58709 ( .A(n32646), .B(\shifter_0/reg_i_8[12] ), .X(n19958) );
  nand_x1_sg U58710 ( .A(reg_oi_8[11]), .B(n33054), .X(n19955) );
  nand_x1_sg U58711 ( .A(n32661), .B(\shifter_0/reg_i_8[11] ), .X(n19956) );
  nand_x1_sg U58712 ( .A(reg_oi_8[10]), .B(n31578), .X(n19953) );
  nand_x1_sg U58713 ( .A(n32666), .B(\shifter_0/reg_i_8[10] ), .X(n19954) );
  nand_x1_sg U58714 ( .A(reg_oi_8[9]), .B(n33116), .X(n19951) );
  nand_x1_sg U58715 ( .A(n34754), .B(\shifter_0/reg_i_8[9] ), .X(n19952) );
  nand_x1_sg U58716 ( .A(reg_oi_8[8]), .B(n35050), .X(n19949) );
  nand_x1_sg U58717 ( .A(n32694), .B(\shifter_0/reg_i_8[8] ), .X(n19950) );
  nand_x1_sg U58718 ( .A(reg_ow_6[19]), .B(n33112), .X(n20531) );
  nand_x1_sg U58719 ( .A(n34412), .B(\shifter_0/reg_w_6[19] ), .X(n20532) );
  nand_x1_sg U58720 ( .A(reg_ow_6[16]), .B(n35016), .X(n20525) );
  nand_x1_sg U58721 ( .A(n32904), .B(\shifter_0/reg_w_6[16] ), .X(n20526) );
  nand_x1_sg U58722 ( .A(reg_ow_6[15]), .B(n31213), .X(n20523) );
  nand_x1_sg U58723 ( .A(n34747), .B(\shifter_0/reg_w_6[15] ), .X(n20524) );
  nand_x1_sg U58724 ( .A(reg_ow_6[14]), .B(n33047), .X(n20521) );
  nand_x1_sg U58725 ( .A(n34103), .B(\shifter_0/reg_w_6[14] ), .X(n20522) );
  nand_x1_sg U58726 ( .A(reg_ow_6[11]), .B(n29807), .X(n20515) );
  nand_x1_sg U58727 ( .A(n30853), .B(\shifter_0/reg_w_6[11] ), .X(n20516) );
  nand_x1_sg U58728 ( .A(reg_ow_6[10]), .B(n33131), .X(n20513) );
  nand_x1_sg U58729 ( .A(n34962), .B(\shifter_0/reg_w_6[10] ), .X(n20514) );
  nand_x1_sg U58730 ( .A(reg_ow_6[7]), .B(n33063), .X(n20507) );
  nand_x1_sg U58731 ( .A(n32690), .B(\shifter_0/reg_w_6[7] ), .X(n20508) );
  nand_x1_sg U58732 ( .A(reg_ow_6[6]), .B(n33112), .X(n20505) );
  nand_x1_sg U58733 ( .A(n34960), .B(\shifter_0/reg_w_6[6] ), .X(n20506) );
  nand_x1_sg U58734 ( .A(reg_ow_6[5]), .B(n33104), .X(n20503) );
  nand_x1_sg U58735 ( .A(n34108), .B(\shifter_0/reg_w_6[5] ), .X(n20504) );
  nand_x1_sg U58736 ( .A(reg_ow_6[2]), .B(n29821), .X(n20497) );
  nand_x1_sg U58737 ( .A(n32670), .B(\shifter_0/reg_w_6[2] ), .X(n20498) );
  nand_x1_sg U58738 ( .A(reg_ow_6[1]), .B(n33105), .X(n20495) );
  nand_x1_sg U58739 ( .A(n32663), .B(\shifter_0/reg_w_6[1] ), .X(n20496) );
  nand_x1_sg U58740 ( .A(reg_ow_6[0]), .B(n31570), .X(n20493) );
  nand_x1_sg U58741 ( .A(n32657), .B(\shifter_0/reg_w_6[0] ), .X(n20494) );
  nand_x1_sg U58742 ( .A(reg_ow_2[19]), .B(n33071), .X(n20371) );
  nand_x1_sg U58743 ( .A(n34727), .B(\shifter_0/reg_w_2[19] ), .X(n20372) );
  nand_x1_sg U58744 ( .A(reg_ow_2[16]), .B(n33097), .X(n20365) );
  nand_x1_sg U58745 ( .A(n32904), .B(\shifter_0/reg_w_2[16] ), .X(n20366) );
  nand_x1_sg U58746 ( .A(reg_ow_2[15]), .B(n33061), .X(n20363) );
  nand_x1_sg U58747 ( .A(n30694), .B(\shifter_0/reg_w_2[15] ), .X(n20364) );
  nand_x1_sg U58748 ( .A(reg_ow_2[14]), .B(n35024), .X(n20361) );
  nand_x1_sg U58749 ( .A(n34110), .B(\shifter_0/reg_w_2[14] ), .X(n20362) );
  nand_x1_sg U58750 ( .A(reg_ow_2[11]), .B(n31590), .X(n20355) );
  nand_x1_sg U58751 ( .A(n32525), .B(\shifter_0/reg_w_2[11] ), .X(n20356) );
  nand_x1_sg U58752 ( .A(reg_ow_2[10]), .B(n30973), .X(n20353) );
  nand_x1_sg U58753 ( .A(n32700), .B(\shifter_0/reg_w_2[10] ), .X(n20354) );
  nand_x1_sg U58754 ( .A(reg_ow_2[7]), .B(n33058), .X(n20347) );
  nand_x1_sg U58755 ( .A(n34098), .B(\shifter_0/reg_w_2[7] ), .X(n20348) );
  nand_x1_sg U58756 ( .A(reg_ow_2[6]), .B(n31579), .X(n20345) );
  nand_x1_sg U58757 ( .A(n32693), .B(\shifter_0/reg_w_2[6] ), .X(n20346) );
  nand_x1_sg U58758 ( .A(reg_ow_2[5]), .B(n33102), .X(n20343) );
  nand_x1_sg U58759 ( .A(n34104), .B(\shifter_0/reg_w_2[5] ), .X(n20344) );
  nand_x1_sg U58760 ( .A(reg_ow_2[2]), .B(n31583), .X(n20337) );
  nand_x1_sg U58761 ( .A(n34738), .B(\shifter_0/reg_w_2[2] ), .X(n20338) );
  nand_x1_sg U58762 ( .A(reg_ow_2[1]), .B(n33080), .X(n20335) );
  nand_x1_sg U58763 ( .A(n34415), .B(\shifter_0/reg_w_2[1] ), .X(n20336) );
  nand_x1_sg U58764 ( .A(reg_ow_2[0]), .B(n35026), .X(n20333) );
  nand_x1_sg U58765 ( .A(n34968), .B(\shifter_0/reg_w_2[0] ), .X(n20334) );
  nand_x1_sg U58766 ( .A(reg_oi_6[19]), .B(n33049), .X(n19891) );
  nand_x1_sg U58767 ( .A(n31985), .B(\shifter_0/reg_i_6[19] ), .X(n19892) );
  nand_x1_sg U58768 ( .A(reg_oi_6[16]), .B(n33046), .X(n19885) );
  nand_x1_sg U58769 ( .A(n30692), .B(\shifter_0/reg_i_6[16] ), .X(n19886) );
  nand_x1_sg U58770 ( .A(reg_oi_6[15]), .B(n33081), .X(n19883) );
  nand_x1_sg U58771 ( .A(n32654), .B(\shifter_0/reg_i_6[15] ), .X(n19884) );
  nand_x1_sg U58772 ( .A(reg_oi_6[14]), .B(n33097), .X(n19881) );
  nand_x1_sg U58773 ( .A(n30702), .B(\shifter_0/reg_i_6[14] ), .X(n19882) );
  nand_x1_sg U58774 ( .A(reg_oi_6[11]), .B(n31566), .X(n19875) );
  nand_x1_sg U58775 ( .A(n32636), .B(\shifter_0/reg_i_6[11] ), .X(n19876) );
  nand_x1_sg U58776 ( .A(reg_oi_6[10]), .B(n31563), .X(n19873) );
  nand_x1_sg U58777 ( .A(n32695), .B(\shifter_0/reg_i_6[10] ), .X(n19874) );
  nand_x1_sg U58778 ( .A(reg_oi_6[7]), .B(n33105), .X(n19867) );
  nand_x1_sg U58779 ( .A(n32699), .B(\shifter_0/reg_i_6[7] ), .X(n19868) );
  nand_x1_sg U58780 ( .A(reg_oi_6[6]), .B(n33104), .X(n19865) );
  nand_x1_sg U58781 ( .A(n34727), .B(\shifter_0/reg_i_6[6] ), .X(n19866) );
  nand_x1_sg U58782 ( .A(reg_oi_6[5]), .B(n31576), .X(n19863) );
  nand_x1_sg U58783 ( .A(n34728), .B(\shifter_0/reg_i_6[5] ), .X(n19864) );
  nand_x1_sg U58784 ( .A(reg_oi_6[2]), .B(n31587), .X(n19857) );
  nand_x1_sg U58785 ( .A(n34958), .B(\shifter_0/reg_i_6[2] ), .X(n19858) );
  nand_x1_sg U58786 ( .A(reg_oi_6[1]), .B(n31573), .X(n19855) );
  nand_x1_sg U58787 ( .A(n32699), .B(\shifter_0/reg_i_6[1] ), .X(n19856) );
  nand_x1_sg U58788 ( .A(reg_oi_6[0]), .B(n33104), .X(n19853) );
  nand_x1_sg U58789 ( .A(n30693), .B(\shifter_0/reg_i_6[0] ), .X(n19854) );
  nand_x1_sg U58790 ( .A(reg_oi_2[19]), .B(n35036), .X(n19731) );
  nand_x1_sg U58791 ( .A(n32697), .B(\shifter_0/reg_i_2[19] ), .X(n19732) );
  nand_x1_sg U58792 ( .A(reg_oi_2[16]), .B(n35039), .X(n19725) );
  nand_x1_sg U58793 ( .A(n32690), .B(\shifter_0/reg_i_2[16] ), .X(n19726) );
  nand_x1_sg U58794 ( .A(reg_oi_2[15]), .B(n33098), .X(n19723) );
  nand_x1_sg U58795 ( .A(n32644), .B(\shifter_0/reg_i_2[15] ), .X(n19724) );
  nand_x1_sg U58796 ( .A(reg_oi_2[14]), .B(n30974), .X(n19721) );
  nand_x1_sg U58797 ( .A(n31475), .B(\shifter_0/reg_i_2[14] ), .X(n19722) );
  nand_x1_sg U58798 ( .A(reg_oi_2[11]), .B(n33090), .X(n19715) );
  nand_x1_sg U58799 ( .A(n34109), .B(\shifter_0/reg_i_2[11] ), .X(n19716) );
  nand_x1_sg U58800 ( .A(reg_oi_2[10]), .B(n33116), .X(n19713) );
  nand_x1_sg U58801 ( .A(n34966), .B(\shifter_0/reg_i_2[10] ), .X(n19714) );
  nand_x1_sg U58802 ( .A(reg_oi_2[7]), .B(n35044), .X(n19707) );
  nand_x1_sg U58803 ( .A(n31986), .B(\shifter_0/reg_i_2[7] ), .X(n19708) );
  nand_x1_sg U58804 ( .A(reg_oi_2[6]), .B(n31215), .X(n19705) );
  nand_x1_sg U58805 ( .A(n30684), .B(\shifter_0/reg_i_2[6] ), .X(n19706) );
  nand_x1_sg U58806 ( .A(reg_oi_2[5]), .B(n33050), .X(n19703) );
  nand_x1_sg U58807 ( .A(n34414), .B(\shifter_0/reg_i_2[5] ), .X(n19704) );
  nand_x1_sg U58808 ( .A(reg_oi_2[2]), .B(n31563), .X(n19697) );
  nand_x1_sg U58809 ( .A(n31989), .B(\shifter_0/reg_i_2[2] ), .X(n19698) );
  nand_x1_sg U58810 ( .A(reg_oi_2[1]), .B(n31564), .X(n19695) );
  nand_x1_sg U58811 ( .A(n32647), .B(\shifter_0/reg_i_2[1] ), .X(n19696) );
  nand_x1_sg U58812 ( .A(reg_oi_2[0]), .B(n31215), .X(n19693) );
  nand_x1_sg U58813 ( .A(n32642), .B(\shifter_0/reg_i_2[0] ), .X(n19694) );
  nand_x1_sg U58814 ( .A(reg_ow_15[17]), .B(n31111), .X(n20887) );
  nand_x1_sg U58815 ( .A(n30697), .B(\shifter_0/reg_w_15[17] ), .X(n20888) );
  nand_x1_sg U58816 ( .A(reg_ow_15[16]), .B(n33124), .X(n20885) );
  nand_x1_sg U58817 ( .A(n32680), .B(\shifter_0/reg_w_15[16] ), .X(n20886) );
  nand_x1_sg U58818 ( .A(reg_ow_15[12]), .B(n29822), .X(n20877) );
  nand_x1_sg U58819 ( .A(n30688), .B(\shifter_0/reg_w_15[12] ), .X(n20878) );
  nand_x1_sg U58820 ( .A(reg_ow_15[11]), .B(n33070), .X(n20875) );
  nand_x1_sg U58821 ( .A(n34108), .B(\shifter_0/reg_w_15[11] ), .X(n20876) );
  nand_x1_sg U58822 ( .A(reg_ow_15[9]), .B(n35023), .X(n20871) );
  nand_x1_sg U58823 ( .A(n32699), .B(\shifter_0/reg_w_15[9] ), .X(n20872) );
  nand_x1_sg U58824 ( .A(reg_ow_15[8]), .B(n31562), .X(n20869) );
  nand_x1_sg U58825 ( .A(n32660), .B(\shifter_0/reg_w_15[8] ), .X(n20870) );
  nand_x1_sg U58826 ( .A(reg_ow_15[6]), .B(n29818), .X(n20865) );
  nand_x1_sg U58827 ( .A(n32688), .B(\shifter_0/reg_w_15[6] ), .X(n20866) );
  nand_x1_sg U58828 ( .A(reg_ow_15[5]), .B(n35015), .X(n20863) );
  nand_x1_sg U58829 ( .A(n34967), .B(\shifter_0/reg_w_15[5] ), .X(n20864) );
  nand_x1_sg U58830 ( .A(reg_ow_15[3]), .B(n35020), .X(n20859) );
  nand_x1_sg U58831 ( .A(n32641), .B(\shifter_0/reg_w_15[3] ), .X(n20860) );
  nand_x1_sg U58832 ( .A(reg_ow_15[2]), .B(n31568), .X(n20857) );
  nand_x1_sg U58833 ( .A(n34744), .B(\shifter_0/reg_w_15[2] ), .X(n20858) );
  nand_x1_sg U58834 ( .A(reg_ow_14[19]), .B(n33118), .X(n20851) );
  nand_x1_sg U58835 ( .A(n31476), .B(\shifter_0/reg_w_14[19] ), .X(n20852) );
  nand_x1_sg U58836 ( .A(reg_ow_14[16]), .B(n33082), .X(n20845) );
  nand_x1_sg U58837 ( .A(n32646), .B(\shifter_0/reg_w_14[16] ), .X(n20846) );
  nand_x1_sg U58838 ( .A(reg_ow_14[15]), .B(n35030), .X(n20843) );
  nand_x1_sg U58839 ( .A(n32652), .B(\shifter_0/reg_w_14[15] ), .X(n20844) );
  nand_x1_sg U58840 ( .A(reg_ow_14[14]), .B(n33104), .X(n20841) );
  nand_x1_sg U58841 ( .A(n32697), .B(\shifter_0/reg_w_14[14] ), .X(n20842) );
  nand_x1_sg U58842 ( .A(reg_ow_14[11]), .B(n33131), .X(n20835) );
  nand_x1_sg U58843 ( .A(n34412), .B(\shifter_0/reg_w_14[11] ), .X(n20836) );
  nand_x1_sg U58844 ( .A(reg_ow_14[10]), .B(n30974), .X(n20833) );
  nand_x1_sg U58845 ( .A(n29761), .B(\shifter_0/reg_w_14[10] ), .X(n20834) );
  nand_x1_sg U58846 ( .A(reg_ow_14[7]), .B(n29827), .X(n20827) );
  nand_x1_sg U58847 ( .A(n34413), .B(\shifter_0/reg_w_14[7] ), .X(n20828) );
  nand_x1_sg U58848 ( .A(reg_ow_14[6]), .B(n35036), .X(n20825) );
  nand_x1_sg U58849 ( .A(n30046), .B(\shifter_0/reg_w_14[6] ), .X(n20826) );
  nand_x1_sg U58850 ( .A(reg_ow_14[5]), .B(n29807), .X(n20823) );
  nand_x1_sg U58851 ( .A(n31989), .B(\shifter_0/reg_w_14[5] ), .X(n20824) );
  nand_x1_sg U58852 ( .A(reg_ow_14[2]), .B(n29836), .X(n20817) );
  nand_x1_sg U58853 ( .A(n32641), .B(\shifter_0/reg_w_14[2] ), .X(n20818) );
  nand_x1_sg U58854 ( .A(reg_ow_14[1]), .B(n33100), .X(n20815) );
  nand_x1_sg U58855 ( .A(n34752), .B(\shifter_0/reg_w_14[1] ), .X(n20816) );
  nand_x1_sg U58856 ( .A(reg_ow_14[0]), .B(n33066), .X(n20813) );
  nand_x1_sg U58857 ( .A(n32692), .B(\shifter_0/reg_w_14[0] ), .X(n20814) );
  nand_x1_sg U58858 ( .A(reg_ow_13[19]), .B(n31564), .X(n20811) );
  nand_x1_sg U58859 ( .A(n30690), .B(\shifter_0/reg_w_13[19] ), .X(n20812) );
  nand_x1_sg U58860 ( .A(reg_ow_13[16]), .B(n33117), .X(n20805) );
  nand_x1_sg U58861 ( .A(n32642), .B(\shifter_0/reg_w_13[16] ), .X(n20806) );
  nand_x1_sg U58862 ( .A(reg_ow_13[15]), .B(n33121), .X(n20803) );
  nand_x1_sg U58863 ( .A(n31475), .B(\shifter_0/reg_w_13[15] ), .X(n20804) );
  nand_x1_sg U58864 ( .A(reg_ow_13[14]), .B(n33105), .X(n20801) );
  nand_x1_sg U58865 ( .A(n30642), .B(\shifter_0/reg_w_13[14] ), .X(n20802) );
  nand_x1_sg U58866 ( .A(reg_ow_13[11]), .B(n31578), .X(n20795) );
  nand_x1_sg U58867 ( .A(n31475), .B(\shifter_0/reg_w_13[11] ), .X(n20796) );
  nand_x1_sg U58868 ( .A(reg_ow_13[0]), .B(n33073), .X(n20773) );
  nand_x1_sg U58869 ( .A(n30698), .B(\shifter_0/reg_w_13[0] ), .X(n20774) );
  nand_x1_sg U58870 ( .A(reg_ow_12[19]), .B(n29821), .X(n20771) );
  nand_x1_sg U58871 ( .A(n31472), .B(\shifter_0/reg_w_12[19] ), .X(n20772) );
  nand_x1_sg U58872 ( .A(reg_ow_12[16]), .B(n31579), .X(n20765) );
  nand_x1_sg U58873 ( .A(n34748), .B(\shifter_0/reg_w_12[16] ), .X(n20766) );
  nand_x1_sg U58874 ( .A(reg_ow_12[15]), .B(n31563), .X(n20763) );
  nand_x1_sg U58875 ( .A(n34754), .B(\shifter_0/reg_w_12[15] ), .X(n20764) );
  nand_x1_sg U58876 ( .A(reg_ow_12[14]), .B(n31576), .X(n20761) );
  nand_x1_sg U58877 ( .A(n31486), .B(\shifter_0/reg_w_12[14] ), .X(n20762) );
  nand_x1_sg U58878 ( .A(reg_ow_12[11]), .B(n31584), .X(n20755) );
  nand_x1_sg U58879 ( .A(n32706), .B(\shifter_0/reg_w_12[11] ), .X(n20756) );
  nand_x1_sg U58880 ( .A(reg_ow_12[10]), .B(n33106), .X(n20753) );
  nand_x1_sg U58881 ( .A(n30681), .B(\shifter_0/reg_w_12[10] ), .X(n20754) );
  nand_x1_sg U58882 ( .A(reg_ow_12[7]), .B(n33068), .X(n20747) );
  nand_x1_sg U58883 ( .A(n32660), .B(\shifter_0/reg_w_12[7] ), .X(n20748) );
  nand_x1_sg U58884 ( .A(reg_ow_12[6]), .B(n33058), .X(n20745) );
  nand_x1_sg U58885 ( .A(n32702), .B(\shifter_0/reg_w_12[6] ), .X(n20746) );
  nand_x1_sg U58886 ( .A(reg_ow_12[5]), .B(n33819), .X(n20743) );
  nand_x1_sg U58887 ( .A(n34739), .B(\shifter_0/reg_w_12[5] ), .X(n20744) );
  nand_x1_sg U58888 ( .A(reg_ow_12[2]), .B(n33077), .X(n20737) );
  nand_x1_sg U58889 ( .A(n34728), .B(\shifter_0/reg_w_12[2] ), .X(n20738) );
  nand_x1_sg U58890 ( .A(reg_ow_12[1]), .B(n31566), .X(n20735) );
  nand_x1_sg U58891 ( .A(n32685), .B(\shifter_0/reg_w_12[1] ), .X(n20736) );
  nand_x1_sg U58892 ( .A(reg_ow_12[0]), .B(n30605), .X(n20733) );
  nand_x1_sg U58893 ( .A(n32668), .B(\shifter_0/reg_w_12[0] ), .X(n20734) );
  nand_x1_sg U58894 ( .A(reg_ow_11[19]), .B(n31579), .X(n20731) );
  nand_x1_sg U58895 ( .A(n32689), .B(\shifter_0/reg_w_11[19] ), .X(n20732) );
  nand_x1_sg U58896 ( .A(reg_ow_11[16]), .B(n33049), .X(n20725) );
  nand_x1_sg U58897 ( .A(n32522), .B(\shifter_0/reg_w_11[16] ), .X(n20726) );
  nand_x1_sg U58898 ( .A(reg_ow_11[15]), .B(n33056), .X(n20723) );
  nand_x1_sg U58899 ( .A(n32683), .B(\shifter_0/reg_w_11[15] ), .X(n20724) );
  nand_x1_sg U58900 ( .A(reg_ow_11[14]), .B(n31214), .X(n20721) );
  nand_x1_sg U58901 ( .A(n32654), .B(\shifter_0/reg_w_11[14] ), .X(n20722) );
  nand_x1_sg U58902 ( .A(reg_ow_11[11]), .B(n31215), .X(n20715) );
  nand_x1_sg U58903 ( .A(n32695), .B(\shifter_0/reg_w_11[11] ), .X(n20716) );
  nand_x1_sg U58904 ( .A(reg_ow_11[10]), .B(n33114), .X(n20713) );
  nand_x1_sg U58905 ( .A(n32705), .B(\shifter_0/reg_w_11[10] ), .X(n20714) );
  nand_x1_sg U58906 ( .A(reg_ow_11[0]), .B(n35042), .X(n20693) );
  nand_x1_sg U58907 ( .A(n31233), .B(\shifter_0/reg_w_11[0] ), .X(n20694) );
  nand_x1_sg U58908 ( .A(reg_ow_9[19]), .B(n33088), .X(n20651) );
  nand_x1_sg U58909 ( .A(n32641), .B(\shifter_0/reg_w_9[19] ), .X(n20652) );
  nand_x1_sg U58910 ( .A(reg_ow_9[16]), .B(n33052), .X(n20645) );
  nand_x1_sg U58911 ( .A(n32646), .B(\shifter_0/reg_w_9[16] ), .X(n20646) );
  nand_x1_sg U58912 ( .A(reg_ow_9[15]), .B(n33050), .X(n20643) );
  nand_x1_sg U58913 ( .A(n31858), .B(\shifter_0/reg_w_9[15] ), .X(n20644) );
  nand_x1_sg U58914 ( .A(reg_ow_9[14]), .B(n35048), .X(n20641) );
  nand_x1_sg U58915 ( .A(n34099), .B(\shifter_0/reg_w_9[14] ), .X(n20642) );
  nand_x1_sg U58916 ( .A(reg_ow_9[11]), .B(n31578), .X(n20635) );
  nand_x1_sg U58917 ( .A(n30044), .B(\shifter_0/reg_w_9[11] ), .X(n20636) );
  nand_x1_sg U58918 ( .A(reg_ow_9[10]), .B(n33062), .X(n20633) );
  nand_x1_sg U58919 ( .A(n31861), .B(\shifter_0/reg_w_9[10] ), .X(n20634) );
  nand_x1_sg U58920 ( .A(reg_ow_9[7]), .B(n31569), .X(n20627) );
  nand_x1_sg U58921 ( .A(n32700), .B(\shifter_0/reg_w_9[7] ), .X(n20628) );
  nand_x1_sg U58922 ( .A(reg_ow_9[6]), .B(n33044), .X(n20625) );
  nand_x1_sg U58923 ( .A(n34734), .B(\shifter_0/reg_w_9[6] ), .X(n20626) );
  nand_x1_sg U58924 ( .A(reg_ow_9[5]), .B(n33094), .X(n20623) );
  nand_x1_sg U58925 ( .A(n34101), .B(\shifter_0/reg_w_9[5] ), .X(n20624) );
  nand_x1_sg U58926 ( .A(reg_ow_9[2]), .B(n29804), .X(n20617) );
  nand_x1_sg U58927 ( .A(n34962), .B(\shifter_0/reg_w_9[2] ), .X(n20618) );
  nand_x1_sg U58928 ( .A(reg_ow_9[1]), .B(n33069), .X(n20615) );
  nand_x1_sg U58929 ( .A(n32682), .B(\shifter_0/reg_w_9[1] ), .X(n20616) );
  nand_x1_sg U58930 ( .A(reg_ow_9[0]), .B(n29804), .X(n20613) );
  nand_x1_sg U58931 ( .A(n34415), .B(\shifter_0/reg_w_9[0] ), .X(n20614) );
  nand_x1_sg U58932 ( .A(reg_ow_5[19]), .B(n29826), .X(n20491) );
  nand_x1_sg U58933 ( .A(n34104), .B(\shifter_0/reg_w_5[19] ), .X(n20492) );
  nand_x1_sg U58934 ( .A(reg_ow_5[16]), .B(n35016), .X(n20485) );
  nand_x1_sg U58935 ( .A(n32644), .B(\shifter_0/reg_w_5[16] ), .X(n20486) );
  nand_x1_sg U58936 ( .A(reg_ow_5[15]), .B(n33099), .X(n20483) );
  nand_x1_sg U58937 ( .A(n32672), .B(\shifter_0/reg_w_5[15] ), .X(n20484) );
  nand_x1_sg U58938 ( .A(reg_ow_5[14]), .B(n33109), .X(n20481) );
  nand_x1_sg U58939 ( .A(n30854), .B(\shifter_0/reg_w_5[14] ), .X(n20482) );
  nand_x1_sg U58940 ( .A(reg_ow_5[11]), .B(n30973), .X(n20475) );
  nand_x1_sg U58941 ( .A(n32707), .B(\shifter_0/reg_w_5[11] ), .X(n20476) );
  nand_x1_sg U58942 ( .A(reg_ow_5[10]), .B(n31573), .X(n20473) );
  nand_x1_sg U58943 ( .A(n32524), .B(\shifter_0/reg_w_5[10] ), .X(n20474) );
  nand_x1_sg U58944 ( .A(reg_ow_5[7]), .B(n35038), .X(n20467) );
  nand_x1_sg U58945 ( .A(n34962), .B(\shifter_0/reg_w_5[7] ), .X(n20468) );
  nand_x1_sg U58946 ( .A(reg_ow_5[6]), .B(n31213), .X(n20465) );
  nand_x1_sg U58947 ( .A(n32669), .B(\shifter_0/reg_w_5[6] ), .X(n20466) );
  nand_x1_sg U58948 ( .A(reg_ow_5[5]), .B(n33093), .X(n20463) );
  nand_x1_sg U58949 ( .A(n34737), .B(\shifter_0/reg_w_5[5] ), .X(n20464) );
  nand_x1_sg U58950 ( .A(reg_ow_5[2]), .B(n30243), .X(n20457) );
  nand_x1_sg U58951 ( .A(n31858), .B(\shifter_0/reg_w_5[2] ), .X(n20458) );
  nand_x1_sg U58952 ( .A(reg_ow_5[1]), .B(n29825), .X(n20455) );
  nand_x1_sg U58953 ( .A(n32666), .B(\shifter_0/reg_w_5[1] ), .X(n20456) );
  nand_x1_sg U58954 ( .A(reg_ow_5[0]), .B(n31573), .X(n20453) );
  nand_x1_sg U58955 ( .A(n32680), .B(\shifter_0/reg_w_5[0] ), .X(n20454) );
  nand_x1_sg U58956 ( .A(reg_ow_3[18]), .B(n31570), .X(n20409) );
  nand_x1_sg U58957 ( .A(n34804), .B(\shifter_0/reg_w_3[18] ), .X(n20410) );
  nand_x1_sg U58958 ( .A(reg_ow_3[17]), .B(n33063), .X(n20407) );
  nand_x1_sg U58959 ( .A(n32688), .B(\shifter_0/reg_w_3[17] ), .X(n20408) );
  nand_x1_sg U58960 ( .A(reg_ow_3[13]), .B(n35017), .X(n20399) );
  nand_x1_sg U58961 ( .A(n30696), .B(\shifter_0/reg_w_3[13] ), .X(n20400) );
  nand_x1_sg U58962 ( .A(reg_ow_3[12]), .B(n35028), .X(n20397) );
  nand_x1_sg U58963 ( .A(n34098), .B(\shifter_0/reg_w_3[12] ), .X(n20398) );
  nand_x1_sg U58964 ( .A(reg_ow_3[9]), .B(n33095), .X(n20391) );
  nand_x1_sg U58965 ( .A(n30046), .B(\shifter_0/reg_w_3[9] ), .X(n20392) );
  nand_x1_sg U58966 ( .A(reg_ow_3[8]), .B(n33111), .X(n20389) );
  nand_x1_sg U58967 ( .A(n32525), .B(\shifter_0/reg_w_3[8] ), .X(n20390) );
  nand_x1_sg U58968 ( .A(reg_ow_3[4]), .B(n33109), .X(n20381) );
  nand_x1_sg U58969 ( .A(n34960), .B(\shifter_0/reg_w_3[4] ), .X(n20382) );
  nand_x1_sg U58970 ( .A(reg_ow_3[3]), .B(n35036), .X(n20379) );
  nand_x1_sg U58971 ( .A(n32669), .B(\shifter_0/reg_w_3[3] ), .X(n20380) );
  nand_x1_sg U58972 ( .A(reg_oi_15[16]), .B(n35049), .X(n20245) );
  nand_x1_sg U58973 ( .A(n30688), .B(\shifter_0/reg_i_15[16] ), .X(n20246) );
  nand_x1_sg U58974 ( .A(reg_oi_15[12]), .B(n31582), .X(n20237) );
  nand_x1_sg U58975 ( .A(n34753), .B(\shifter_0/reg_i_15[12] ), .X(n20238) );
  nand_x1_sg U58976 ( .A(reg_oi_15[11]), .B(n35029), .X(n20235) );
  nand_x1_sg U58977 ( .A(n32664), .B(\shifter_0/reg_i_15[11] ), .X(n20236) );
  nand_x1_sg U58978 ( .A(reg_oi_15[9]), .B(n29836), .X(n20231) );
  nand_x1_sg U58979 ( .A(n34414), .B(\shifter_0/reg_i_15[9] ), .X(n20232) );
  nand_x1_sg U58980 ( .A(reg_oi_15[8]), .B(n35020), .X(n20229) );
  nand_x1_sg U58981 ( .A(n34730), .B(\shifter_0/reg_i_15[8] ), .X(n20230) );
  nand_x1_sg U58982 ( .A(reg_oi_15[6]), .B(n29830), .X(n20225) );
  nand_x1_sg U58983 ( .A(n32701), .B(\shifter_0/reg_i_15[6] ), .X(n20226) );
  nand_x1_sg U58984 ( .A(reg_oi_15[5]), .B(n31565), .X(n20223) );
  nand_x1_sg U58985 ( .A(n32682), .B(\shifter_0/reg_i_15[5] ), .X(n20224) );
  nand_x1_sg U58986 ( .A(reg_oi_15[3]), .B(n31567), .X(n20219) );
  nand_x1_sg U58987 ( .A(n32663), .B(\shifter_0/reg_i_15[3] ), .X(n20220) );
  nand_x1_sg U58988 ( .A(reg_oi_14[19]), .B(n35038), .X(n20211) );
  nand_x1_sg U58989 ( .A(n30698), .B(\shifter_0/reg_i_14[19] ), .X(n20212) );
  nand_x1_sg U58990 ( .A(reg_oi_14[15]), .B(n33123), .X(n20203) );
  nand_x1_sg U58991 ( .A(n34104), .B(\shifter_0/reg_i_14[15] ), .X(n20204) );
  nand_x1_sg U58992 ( .A(reg_oi_14[7]), .B(n35028), .X(n20187) );
  nand_x1_sg U58993 ( .A(n32692), .B(\shifter_0/reg_i_14[7] ), .X(n20188) );
  nand_x1_sg U58994 ( .A(reg_oi_14[6]), .B(n31566), .X(n20185) );
  nand_x1_sg U58995 ( .A(n31472), .B(\shifter_0/reg_i_14[6] ), .X(n20186) );
  nand_x1_sg U58996 ( .A(reg_oi_13[15]), .B(n33107), .X(n20163) );
  nand_x1_sg U58997 ( .A(n32526), .B(\shifter_0/reg_i_13[15] ), .X(n20164) );
  nand_x1_sg U58998 ( .A(reg_oi_13[14]), .B(n35025), .X(n20161) );
  nand_x1_sg U58999 ( .A(n32661), .B(\shifter_0/reg_i_13[14] ), .X(n20162) );
  nand_x1_sg U59000 ( .A(reg_oi_13[11]), .B(n29799), .X(n20155) );
  nand_x1_sg U59001 ( .A(n32521), .B(\shifter_0/reg_i_13[11] ), .X(n20156) );
  nand_x1_sg U59002 ( .A(reg_oi_13[10]), .B(n33117), .X(n20153) );
  nand_x1_sg U59003 ( .A(n32657), .B(\shifter_0/reg_i_13[10] ), .X(n20154) );
  nand_x1_sg U59004 ( .A(reg_oi_13[7]), .B(n33073), .X(n20147) );
  nand_x1_sg U59005 ( .A(n34751), .B(\shifter_0/reg_i_13[7] ), .X(n20148) );
  nand_x1_sg U59006 ( .A(reg_oi_13[6]), .B(n35015), .X(n20145) );
  nand_x1_sg U59007 ( .A(n32678), .B(\shifter_0/reg_i_13[6] ), .X(n20146) );
  nand_x1_sg U59008 ( .A(reg_oi_13[5]), .B(n31591), .X(n20143) );
  nand_x1_sg U59009 ( .A(n32690), .B(\shifter_0/reg_i_13[5] ), .X(n20144) );
  nand_x1_sg U59010 ( .A(reg_oi_13[3]), .B(n31585), .X(n20139) );
  nand_x1_sg U59011 ( .A(n32669), .B(\shifter_0/reg_i_13[3] ), .X(n20140) );
  nand_x1_sg U59012 ( .A(reg_oi_13[1]), .B(n30240), .X(n20135) );
  nand_x1_sg U59013 ( .A(n34738), .B(\shifter_0/reg_i_13[1] ), .X(n20136) );
  nand_x1_sg U59014 ( .A(reg_oi_13[0]), .B(n33051), .X(n20133) );
  nand_x1_sg U59015 ( .A(n32661), .B(\shifter_0/reg_i_13[0] ), .X(n20134) );
  nand_x1_sg U59016 ( .A(reg_oi_12[19]), .B(n35023), .X(n20131) );
  nand_x1_sg U59017 ( .A(n30684), .B(\shifter_0/reg_i_12[19] ), .X(n20132) );
  nand_x1_sg U59018 ( .A(reg_oi_12[15]), .B(n29827), .X(n20123) );
  nand_x1_sg U59019 ( .A(n34109), .B(\shifter_0/reg_i_12[15] ), .X(n20124) );
  nand_x1_sg U59020 ( .A(reg_oi_12[14]), .B(n31590), .X(n20121) );
  nand_x1_sg U59021 ( .A(n30682), .B(\shifter_0/reg_i_12[14] ), .X(n20122) );
  nand_x1_sg U59022 ( .A(reg_oi_12[11]), .B(n29821), .X(n20115) );
  nand_x1_sg U59023 ( .A(n34959), .B(\shifter_0/reg_i_12[11] ), .X(n20116) );
  nand_x1_sg U59024 ( .A(reg_oi_12[10]), .B(n29827), .X(n20113) );
  nand_x1_sg U59025 ( .A(n34801), .B(\shifter_0/reg_i_12[10] ), .X(n20114) );
  nand_x1_sg U59026 ( .A(reg_oi_12[3]), .B(n33051), .X(n20099) );
  nand_x1_sg U59027 ( .A(n32659), .B(\shifter_0/reg_i_12[3] ), .X(n20100) );
  nand_x1_sg U59028 ( .A(reg_oi_12[1]), .B(n33110), .X(n20095) );
  nand_x1_sg U59029 ( .A(n31860), .B(\shifter_0/reg_i_12[1] ), .X(n20096) );
  nand_x1_sg U59030 ( .A(reg_oi_12[0]), .B(n33071), .X(n20093) );
  nand_x1_sg U59031 ( .A(n32677), .B(\shifter_0/reg_i_12[0] ), .X(n20094) );
  nand_x1_sg U59032 ( .A(reg_oi_11[19]), .B(n33059), .X(n20091) );
  nand_x1_sg U59033 ( .A(n32652), .B(\shifter_0/reg_i_11[19] ), .X(n20092) );
  nand_x1_sg U59034 ( .A(reg_oi_11[15]), .B(n29826), .X(n20083) );
  nand_x1_sg U59035 ( .A(n34964), .B(\shifter_0/reg_i_11[15] ), .X(n20084) );
  nand_x1_sg U59036 ( .A(reg_oi_11[14]), .B(n33086), .X(n20081) );
  nand_x1_sg U59037 ( .A(n34101), .B(\shifter_0/reg_i_11[14] ), .X(n20082) );
  nand_x1_sg U59038 ( .A(reg_oi_11[11]), .B(n35049), .X(n20075) );
  nand_x1_sg U59039 ( .A(n32525), .B(\shifter_0/reg_i_11[11] ), .X(n20076) );
  nand_x1_sg U59040 ( .A(reg_oi_11[10]), .B(n31569), .X(n20073) );
  nand_x1_sg U59041 ( .A(n34725), .B(\shifter_0/reg_i_11[10] ), .X(n20074) );
  nand_x1_sg U59042 ( .A(reg_oi_11[7]), .B(n33099), .X(n20067) );
  nand_x1_sg U59043 ( .A(n34961), .B(\shifter_0/reg_i_11[7] ), .X(n20068) );
  nand_x1_sg U59044 ( .A(reg_oi_9[19]), .B(n33100), .X(n20011) );
  nand_x1_sg U59045 ( .A(n32676), .B(\shifter_0/reg_i_9[19] ), .X(n20012) );
  nand_x1_sg U59046 ( .A(reg_oi_9[15]), .B(n29824), .X(n20003) );
  nand_x1_sg U59047 ( .A(n30701), .B(\shifter_0/reg_i_9[15] ), .X(n20004) );
  nand_x1_sg U59048 ( .A(reg_oi_9[14]), .B(n33124), .X(n20001) );
  nand_x1_sg U59049 ( .A(n31861), .B(\shifter_0/reg_i_9[14] ), .X(n20002) );
  nand_x1_sg U59050 ( .A(reg_oi_9[11]), .B(n33822), .X(n19995) );
  nand_x1_sg U59051 ( .A(n32678), .B(\shifter_0/reg_i_9[11] ), .X(n19996) );
  nand_x1_sg U59052 ( .A(reg_oi_9[10]), .B(n35043), .X(n19993) );
  nand_x1_sg U59053 ( .A(n32901), .B(\shifter_0/reg_i_9[10] ), .X(n19994) );
  nand_x1_sg U59054 ( .A(reg_oi_9[7]), .B(n31214), .X(n19987) );
  nand_x1_sg U59055 ( .A(n34967), .B(\shifter_0/reg_i_9[7] ), .X(n19988) );
  nand_x1_sg U59056 ( .A(reg_oi_9[6]), .B(n33085), .X(n19985) );
  nand_x1_sg U59057 ( .A(n32648), .B(\shifter_0/reg_i_9[6] ), .X(n19986) );
  nand_x1_sg U59058 ( .A(reg_oi_9[5]), .B(n33050), .X(n19983) );
  nand_x1_sg U59059 ( .A(n32639), .B(\shifter_0/reg_i_9[5] ), .X(n19984) );
  nand_x1_sg U59060 ( .A(reg_oi_9[3]), .B(n33097), .X(n19979) );
  nand_x1_sg U59061 ( .A(n30044), .B(\shifter_0/reg_i_9[3] ), .X(n19980) );
  nand_x1_sg U59062 ( .A(reg_oi_9[1]), .B(n35028), .X(n19975) );
  nand_x1_sg U59063 ( .A(n31861), .B(\shifter_0/reg_i_9[1] ), .X(n19976) );
  nand_x1_sg U59064 ( .A(reg_oi_9[0]), .B(n33075), .X(n19973) );
  nand_x1_sg U59065 ( .A(n34958), .B(\shifter_0/reg_i_9[0] ), .X(n19974) );
  nand_x1_sg U59066 ( .A(reg_oi_5[19]), .B(n33041), .X(n19851) );
  nand_x1_sg U59067 ( .A(n32640), .B(\shifter_0/reg_i_5[19] ), .X(n19852) );
  nand_x1_sg U59068 ( .A(reg_oi_5[16]), .B(n33107), .X(n19845) );
  nand_x1_sg U59069 ( .A(n31859), .B(\shifter_0/reg_i_5[16] ), .X(n19846) );
  nand_x1_sg U59070 ( .A(reg_oi_5[15]), .B(n30240), .X(n19843) );
  nand_x1_sg U59071 ( .A(n31858), .B(\shifter_0/reg_i_5[15] ), .X(n19844) );
  nand_x1_sg U59072 ( .A(reg_oi_5[14]), .B(n33064), .X(n19841) );
  nand_x1_sg U59073 ( .A(n32648), .B(\shifter_0/reg_i_5[14] ), .X(n19842) );
  nand_x1_sg U59074 ( .A(reg_oi_5[11]), .B(n33071), .X(n19835) );
  nand_x1_sg U59075 ( .A(n30680), .B(\shifter_0/reg_i_5[11] ), .X(n19836) );
  nand_x1_sg U59076 ( .A(reg_oi_5[10]), .B(n31570), .X(n19833) );
  nand_x1_sg U59077 ( .A(n34961), .B(\shifter_0/reg_i_5[10] ), .X(n19834) );
  nand_x1_sg U59078 ( .A(reg_oi_3[18]), .B(n35045), .X(n19769) );
  nand_x1_sg U59079 ( .A(n32668), .B(\shifter_0/reg_i_3[18] ), .X(n19770) );
  nand_x1_sg U59080 ( .A(reg_oi_3[17]), .B(n35022), .X(n19767) );
  nand_x1_sg U59081 ( .A(n32699), .B(\shifter_0/reg_i_3[17] ), .X(n19768) );
  nand_x1_sg U59082 ( .A(reg_oi_3[13]), .B(n35038), .X(n19759) );
  nand_x1_sg U59083 ( .A(n34110), .B(\shifter_0/reg_i_3[13] ), .X(n19760) );
  nand_x1_sg U59084 ( .A(reg_oi_3[12]), .B(n33076), .X(n19757) );
  nand_x1_sg U59085 ( .A(n32647), .B(\shifter_0/reg_i_3[12] ), .X(n19758) );
  nand_x1_sg U59086 ( .A(reg_oi_3[9]), .B(n29821), .X(n19751) );
  nand_x1_sg U59087 ( .A(n30681), .B(\shifter_0/reg_i_3[9] ), .X(n19752) );
  nand_x1_sg U59088 ( .A(reg_oi_3[8]), .B(n31563), .X(n19749) );
  nand_x1_sg U59089 ( .A(n32687), .B(\shifter_0/reg_i_3[8] ), .X(n19750) );
  nand_x1_sg U59090 ( .A(reg_oi_3[4]), .B(n35021), .X(n19741) );
  nand_x1_sg U59091 ( .A(n32521), .B(\shifter_0/reg_i_3[4] ), .X(n19742) );
  nand_x1_sg U59092 ( .A(reg_oi_3[3]), .B(n33092), .X(n19739) );
  nand_x1_sg U59093 ( .A(n32524), .B(\shifter_0/reg_i_3[3] ), .X(n19740) );
  nand_x1_sg U59094 ( .A(reg_ow_1[19]), .B(n33066), .X(n20331) );
  nand_x1_sg U59095 ( .A(n32668), .B(\shifter_0/reg_w_1[19] ), .X(n20332) );
  nand_x1_sg U59096 ( .A(reg_ow_1[16]), .B(n35050), .X(n20325) );
  nand_x1_sg U59097 ( .A(n32653), .B(\shifter_0/reg_w_1[16] ), .X(n20326) );
  nand_x1_sg U59098 ( .A(reg_ow_1[15]), .B(n33113), .X(n20323) );
  nand_x1_sg U59099 ( .A(n32660), .B(\shifter_0/reg_w_1[15] ), .X(n20324) );
  nand_x1_sg U59100 ( .A(reg_ow_1[14]), .B(n35048), .X(n20321) );
  nand_x1_sg U59101 ( .A(n30693), .B(\shifter_0/reg_w_1[14] ), .X(n20322) );
  nand_x1_sg U59102 ( .A(reg_ow_1[7]), .B(n31576), .X(n20307) );
  nand_x1_sg U59103 ( .A(n31235), .B(\shifter_0/reg_w_1[7] ), .X(n20308) );
  nand_x1_sg U59104 ( .A(reg_ow_1[6]), .B(n35019), .X(n20305) );
  nand_x1_sg U59105 ( .A(n34110), .B(\shifter_0/reg_w_1[6] ), .X(n20306) );
  nand_x1_sg U59106 ( .A(reg_ow_1[5]), .B(n35028), .X(n20303) );
  nand_x1_sg U59107 ( .A(n32706), .B(\shifter_0/reg_w_1[5] ), .X(n20304) );
  nand_x1_sg U59108 ( .A(reg_ow_1[2]), .B(n31212), .X(n20297) );
  nand_x1_sg U59109 ( .A(n31988), .B(\shifter_0/reg_w_1[2] ), .X(n20298) );
  nand_x1_sg U59110 ( .A(reg_ow_1[1]), .B(n31568), .X(n20295) );
  nand_x1_sg U59111 ( .A(n32664), .B(\shifter_0/reg_w_1[1] ), .X(n20296) );
  nand_x1_sg U59112 ( .A(reg_ow_1[0]), .B(n35023), .X(n20293) );
  nand_x1_sg U59113 ( .A(n32524), .B(\shifter_0/reg_w_1[0] ), .X(n20294) );
  nand_x1_sg U59114 ( .A(reg_oi_14[18]), .B(n31579), .X(n20209) );
  nand_x1_sg U59115 ( .A(n32522), .B(\shifter_0/reg_i_14[18] ), .X(n20210) );
  nand_x1_sg U59116 ( .A(reg_oi_14[17]), .B(n31581), .X(n20207) );
  nand_x1_sg U59117 ( .A(n34730), .B(\shifter_0/reg_i_14[17] ), .X(n20208) );
  nand_x1_sg U59118 ( .A(reg_oi_13[4]), .B(n33076), .X(n20141) );
  nand_x1_sg U59119 ( .A(n32682), .B(\shifter_0/reg_i_13[4] ), .X(n20142) );
  nand_x1_sg U59120 ( .A(reg_oi_13[2]), .B(n33049), .X(n20137) );
  nand_x1_sg U59121 ( .A(n32639), .B(\shifter_0/reg_i_13[2] ), .X(n20138) );
  nand_x1_sg U59122 ( .A(reg_oi_12[18]), .B(n31213), .X(n20129) );
  nand_x1_sg U59123 ( .A(n32675), .B(\shifter_0/reg_i_12[18] ), .X(n20130) );
  nand_x1_sg U59124 ( .A(reg_oi_12[17]), .B(n33075), .X(n20127) );
  nand_x1_sg U59125 ( .A(n34733), .B(\shifter_0/reg_i_12[17] ), .X(n20128) );
  nand_x1_sg U59126 ( .A(reg_oi_12[4]), .B(n33820), .X(n20101) );
  nand_x1_sg U59127 ( .A(n30853), .B(\shifter_0/reg_i_12[4] ), .X(n20102) );
  nand_x1_sg U59128 ( .A(reg_oi_12[2]), .B(n33820), .X(n20097) );
  nand_x1_sg U59129 ( .A(n30215), .B(\shifter_0/reg_i_12[2] ), .X(n20098) );
  nand_x1_sg U59130 ( .A(reg_oi_11[18]), .B(n33109), .X(n20089) );
  nand_x1_sg U59131 ( .A(n30692), .B(\shifter_0/reg_i_11[18] ), .X(n20090) );
  nand_x1_sg U59132 ( .A(reg_oi_11[17]), .B(n35047), .X(n20087) );
  nand_x1_sg U59133 ( .A(n32659), .B(\shifter_0/reg_i_11[17] ), .X(n20088) );
  nand_x1_sg U59134 ( .A(reg_oi_10[17]), .B(n33128), .X(n20047) );
  nand_x1_sg U59135 ( .A(n32525), .B(\shifter_0/reg_i_10[17] ), .X(n20048) );
  nand_x1_sg U59136 ( .A(reg_oi_10[4]), .B(n33111), .X(n20021) );
  nand_x1_sg U59137 ( .A(n31236), .B(\shifter_0/reg_i_10[4] ), .X(n20022) );
  nand_x1_sg U59138 ( .A(reg_oi_10[2]), .B(n33117), .X(n20017) );
  nand_x1_sg U59139 ( .A(n32653), .B(\shifter_0/reg_i_10[2] ), .X(n20018) );
  nand_x1_sg U59140 ( .A(reg_oi_9[18]), .B(n33062), .X(n20009) );
  nand_x1_sg U59141 ( .A(n32652), .B(\shifter_0/reg_i_9[18] ), .X(n20010) );
  nand_x1_sg U59142 ( .A(reg_oi_9[17]), .B(n33044), .X(n20007) );
  nand_x1_sg U59143 ( .A(n34101), .B(\shifter_0/reg_i_9[17] ), .X(n20008) );
  nand_x1_sg U59144 ( .A(reg_oi_9[4]), .B(n29822), .X(n19981) );
  nand_x1_sg U59145 ( .A(n34968), .B(\shifter_0/reg_i_9[4] ), .X(n19982) );
  nand_x1_sg U59146 ( .A(reg_oi_9[2]), .B(n35016), .X(n19977) );
  nand_x1_sg U59147 ( .A(n32694), .B(\shifter_0/reg_i_9[2] ), .X(n19978) );
  nand_x1_sg U59148 ( .A(reg_oi_1[11]), .B(n33102), .X(n19675) );
  nand_x1_sg U59149 ( .A(n32696), .B(\shifter_0/reg_i_1[11] ), .X(n19676) );
  nand_x1_sg U59150 ( .A(reg_oi_1[10]), .B(n33070), .X(n19673) );
  nand_x1_sg U59151 ( .A(n31859), .B(\shifter_0/reg_i_1[10] ), .X(n19674) );
  nand_x1_sg U59152 ( .A(reg_oi_1[7]), .B(n35035), .X(n19667) );
  nand_x1_sg U59153 ( .A(n32675), .B(\shifter_0/reg_i_1[7] ), .X(n19668) );
  nand_x1_sg U59154 ( .A(reg_oi_1[6]), .B(n31212), .X(n19665) );
  nand_x1_sg U59155 ( .A(n32665), .B(\shifter_0/reg_i_1[6] ), .X(n19666) );
  nand_x1_sg U59156 ( .A(reg_oi_1[5]), .B(n30246), .X(n19663) );
  nand_x1_sg U59157 ( .A(n34110), .B(\shifter_0/reg_i_1[5] ), .X(n19664) );
  nand_x1_sg U59158 ( .A(reg_oi_1[2]), .B(n33061), .X(n19657) );
  nand_x1_sg U59159 ( .A(n32664), .B(\shifter_0/reg_i_1[2] ), .X(n19658) );
  nand_x1_sg U59160 ( .A(reg_oi_1[1]), .B(n33130), .X(n19655) );
  nand_x1_sg U59161 ( .A(n32696), .B(\shifter_0/reg_i_1[1] ), .X(n19656) );
  nand_x1_sg U59162 ( .A(reg_oi_1[0]), .B(n29833), .X(n19653) );
  nand_x1_sg U59163 ( .A(n30043), .B(\shifter_0/reg_i_1[0] ), .X(n19654) );
  nand_x1_sg U59164 ( .A(reg_ow_10[19]), .B(n35035), .X(n20691) );
  nand_x1_sg U59165 ( .A(n30215), .B(\shifter_0/reg_w_10[19] ), .X(n20692) );
  nand_x1_sg U59166 ( .A(reg_ow_10[18]), .B(n35042), .X(n20689) );
  nand_x1_sg U59167 ( .A(n31986), .B(\shifter_0/reg_w_10[18] ), .X(n20690) );
  nand_x1_sg U59168 ( .A(reg_ow_10[17]), .B(n33130), .X(n20687) );
  nand_x1_sg U59169 ( .A(n32649), .B(\shifter_0/reg_w_10[17] ), .X(n20688) );
  nand_x1_sg U59170 ( .A(reg_ow_10[16]), .B(n33123), .X(n20685) );
  nand_x1_sg U59171 ( .A(n34738), .B(\shifter_0/reg_w_10[16] ), .X(n20686) );
  nand_x1_sg U59172 ( .A(reg_ow_10[15]), .B(n35043), .X(n20683) );
  nand_x1_sg U59173 ( .A(n34746), .B(\shifter_0/reg_w_10[15] ), .X(n20684) );
  nand_x1_sg U59174 ( .A(reg_ow_10[14]), .B(n35022), .X(n20681) );
  nand_x1_sg U59175 ( .A(n32676), .B(\shifter_0/reg_w_10[14] ), .X(n20682) );
  nand_x1_sg U59176 ( .A(reg_ow_10[13]), .B(n35046), .X(n20679) );
  nand_x1_sg U59177 ( .A(n34742), .B(\shifter_0/reg_w_10[13] ), .X(n20680) );
  nand_x1_sg U59178 ( .A(reg_ow_10[12]), .B(n33046), .X(n20677) );
  nand_x1_sg U59179 ( .A(n32678), .B(\shifter_0/reg_w_10[12] ), .X(n20678) );
  nand_x1_sg U59180 ( .A(reg_ow_10[11]), .B(n33085), .X(n20675) );
  nand_x1_sg U59181 ( .A(n32522), .B(\shifter_0/reg_w_10[11] ), .X(n20676) );
  nand_x1_sg U59182 ( .A(reg_ow_10[1]), .B(n33081), .X(n20655) );
  nand_x1_sg U59183 ( .A(n31860), .B(\shifter_0/reg_w_10[1] ), .X(n20656) );
  nand_x1_sg U59184 ( .A(reg_ow_10[0]), .B(n35018), .X(n20653) );
  nand_x1_sg U59185 ( .A(n32672), .B(\shifter_0/reg_w_10[0] ), .X(n20654) );
  nand_x1_sg U59186 ( .A(reg_oi_10[16]), .B(n30602), .X(n20045) );
  nand_x1_sg U59187 ( .A(n30046), .B(\shifter_0/reg_i_10[16] ), .X(n20046) );
  nand_x1_sg U59188 ( .A(reg_oi_10[15]), .B(n29827), .X(n20043) );
  nand_x1_sg U59189 ( .A(n34739), .B(\shifter_0/reg_i_10[15] ), .X(n20044) );
  nand_x1_sg U59190 ( .A(reg_oi_10[14]), .B(n30241), .X(n20041) );
  nand_x1_sg U59191 ( .A(n34102), .B(\shifter_0/reg_i_10[14] ), .X(n20042) );
  nand_x1_sg U59192 ( .A(reg_oi_10[13]), .B(n31584), .X(n20039) );
  nand_x1_sg U59193 ( .A(n32656), .B(\shifter_0/reg_i_10[13] ), .X(n20040) );
  nand_x1_sg U59194 ( .A(reg_oi_10[12]), .B(n33083), .X(n20037) );
  nand_x1_sg U59195 ( .A(n32640), .B(\shifter_0/reg_i_10[12] ), .X(n20038) );
  nand_x1_sg U59196 ( .A(reg_oi_10[11]), .B(n30243), .X(n20035) );
  nand_x1_sg U59197 ( .A(n34111), .B(\shifter_0/reg_i_10[11] ), .X(n20036) );
  nand_x1_sg U59198 ( .A(reg_oi_10[10]), .B(n33056), .X(n20033) );
  nand_x1_sg U59199 ( .A(n34959), .B(\shifter_0/reg_i_10[10] ), .X(n20034) );
  nand_x1_sg U59200 ( .A(reg_oi_10[9]), .B(n35018), .X(n20031) );
  nand_x1_sg U59201 ( .A(n30043), .B(\shifter_0/reg_i_10[9] ), .X(n20032) );
  nand_x1_sg U59202 ( .A(reg_oi_10[8]), .B(n33113), .X(n20029) );
  nand_x1_sg U59203 ( .A(n32661), .B(\shifter_0/reg_i_10[8] ), .X(n20030) );
  nand_x1_sg U59204 ( .A(reg_oi_10[7]), .B(n29801), .X(n20027) );
  nand_x1_sg U59205 ( .A(n32687), .B(\shifter_0/reg_i_10[7] ), .X(n20028) );
  nand_x1_sg U59206 ( .A(reg_oi_10[6]), .B(n33101), .X(n20025) );
  nand_x1_sg U59207 ( .A(n32677), .B(\shifter_0/reg_i_10[6] ), .X(n20026) );
  nand_x1_sg U59208 ( .A(reg_oi_10[5]), .B(n35029), .X(n20023) );
  nand_x1_sg U59209 ( .A(n34103), .B(\shifter_0/reg_i_10[5] ), .X(n20024) );
  nand_x1_sg U59210 ( .A(reg_oi_10[3]), .B(n29815), .X(n20019) );
  nand_x1_sg U59211 ( .A(n34412), .B(\shifter_0/reg_i_10[3] ), .X(n20020) );
  nand_x1_sg U59212 ( .A(reg_oi_10[1]), .B(n35039), .X(n20015) );
  nand_x1_sg U59213 ( .A(n32903), .B(\shifter_0/reg_i_10[1] ), .X(n20016) );
  nand_x1_sg U59214 ( .A(reg_oi_10[0]), .B(n29799), .X(n20013) );
  nand_x1_sg U59215 ( .A(n30688), .B(\shifter_0/reg_i_10[0] ), .X(n20014) );
  nand_x1_sg U59216 ( .A(reg_ow_14[18]), .B(n33129), .X(n20849) );
  nand_x1_sg U59217 ( .A(n32902), .B(\shifter_0/reg_w_14[18] ), .X(n20850) );
  nand_x1_sg U59218 ( .A(reg_ow_14[17]), .B(n33092), .X(n20847) );
  nand_x1_sg U59219 ( .A(n34737), .B(\shifter_0/reg_w_14[17] ), .X(n20848) );
  nand_x1_sg U59220 ( .A(reg_ow_14[13]), .B(n33129), .X(n20839) );
  nand_x1_sg U59221 ( .A(n32702), .B(\shifter_0/reg_w_14[13] ), .X(n20840) );
  nand_x1_sg U59222 ( .A(reg_ow_14[12]), .B(n33086), .X(n20837) );
  nand_x1_sg U59223 ( .A(n34960), .B(\shifter_0/reg_w_14[12] ), .X(n20838) );
  nand_x1_sg U59224 ( .A(reg_ow_14[9]), .B(n31585), .X(n20831) );
  nand_x1_sg U59225 ( .A(n31858), .B(\shifter_0/reg_w_14[9] ), .X(n20832) );
  nand_x1_sg U59226 ( .A(reg_ow_14[8]), .B(n33059), .X(n20829) );
  nand_x1_sg U59227 ( .A(n32651), .B(\shifter_0/reg_w_14[8] ), .X(n20830) );
  nand_x1_sg U59228 ( .A(reg_ow_14[4]), .B(n33058), .X(n20821) );
  nand_x1_sg U59229 ( .A(n31236), .B(\shifter_0/reg_w_14[4] ), .X(n20822) );
  nand_x1_sg U59230 ( .A(reg_ow_14[3]), .B(n33101), .X(n20819) );
  nand_x1_sg U59231 ( .A(n32705), .B(\shifter_0/reg_w_14[3] ), .X(n20820) );
  nand_x1_sg U59232 ( .A(reg_ow_13[18]), .B(n33125), .X(n20809) );
  nand_x1_sg U59233 ( .A(n32689), .B(\shifter_0/reg_w_13[18] ), .X(n20810) );
  nand_x1_sg U59234 ( .A(reg_ow_13[17]), .B(n33130), .X(n20807) );
  nand_x1_sg U59235 ( .A(n32651), .B(\shifter_0/reg_w_13[17] ), .X(n20808) );
  nand_x1_sg U59236 ( .A(reg_ow_13[13]), .B(n30241), .X(n20799) );
  nand_x1_sg U59237 ( .A(n34108), .B(\shifter_0/reg_w_13[13] ), .X(n20800) );
  nand_x1_sg U59238 ( .A(reg_ow_13[12]), .B(n33047), .X(n20797) );
  nand_x1_sg U59239 ( .A(n34749), .B(\shifter_0/reg_w_13[12] ), .X(n20798) );
  nand_x1_sg U59240 ( .A(reg_ow_12[18]), .B(n33089), .X(n20769) );
  nand_x1_sg U59241 ( .A(n34746), .B(\shifter_0/reg_w_12[18] ), .X(n20770) );
  nand_x1_sg U59242 ( .A(reg_ow_12[17]), .B(n31577), .X(n20767) );
  nand_x1_sg U59243 ( .A(n31476), .B(\shifter_0/reg_w_12[17] ), .X(n20768) );
  nand_x1_sg U59244 ( .A(reg_ow_12[13]), .B(n29822), .X(n20759) );
  nand_x1_sg U59245 ( .A(n32644), .B(\shifter_0/reg_w_12[13] ), .X(n20760) );
  nand_x1_sg U59246 ( .A(reg_ow_12[12]), .B(n33058), .X(n20757) );
  nand_x1_sg U59247 ( .A(n32681), .B(\shifter_0/reg_w_12[12] ), .X(n20758) );
  nand_x1_sg U59248 ( .A(reg_ow_12[9]), .B(n35018), .X(n20751) );
  nand_x1_sg U59249 ( .A(n34801), .B(\shifter_0/reg_w_12[9] ), .X(n20752) );
  nand_x1_sg U59250 ( .A(reg_ow_12[8]), .B(n29799), .X(n20749) );
  nand_x1_sg U59251 ( .A(n34736), .B(\shifter_0/reg_w_12[8] ), .X(n20750) );
  nand_x1_sg U59252 ( .A(reg_ow_12[4]), .B(n31568), .X(n20741) );
  nand_x1_sg U59253 ( .A(n32672), .B(\shifter_0/reg_w_12[4] ), .X(n20742) );
  nand_x1_sg U59254 ( .A(reg_ow_12[3]), .B(n33129), .X(n20739) );
  nand_x1_sg U59255 ( .A(n34965), .B(\shifter_0/reg_w_12[3] ), .X(n20740) );
  nand_x1_sg U59256 ( .A(reg_ow_11[18]), .B(n30605), .X(n20729) );
  nand_x1_sg U59257 ( .A(n32524), .B(\shifter_0/reg_w_11[18] ), .X(n20730) );
  nand_x1_sg U59258 ( .A(reg_ow_11[17]), .B(n35017), .X(n20727) );
  nand_x1_sg U59259 ( .A(n32651), .B(\shifter_0/reg_w_11[17] ), .X(n20728) );
  nand_x1_sg U59260 ( .A(reg_ow_11[13]), .B(n29804), .X(n20719) );
  nand_x1_sg U59261 ( .A(n34964), .B(\shifter_0/reg_w_11[13] ), .X(n20720) );
  nand_x1_sg U59262 ( .A(reg_ow_11[12]), .B(n31572), .X(n20717) );
  nand_x1_sg U59263 ( .A(n30046), .B(\shifter_0/reg_w_11[12] ), .X(n20718) );
  nand_x1_sg U59264 ( .A(reg_ow_11[9]), .B(n31591), .X(n20711) );
  nand_x1_sg U59265 ( .A(n32690), .B(\shifter_0/reg_w_11[9] ), .X(n20712) );
  nand_x1_sg U59266 ( .A(reg_ow_9[18]), .B(n33112), .X(n20649) );
  nand_x1_sg U59267 ( .A(n32657), .B(\shifter_0/reg_w_9[18] ), .X(n20650) );
  nand_x1_sg U59268 ( .A(reg_ow_9[17]), .B(n35050), .X(n20647) );
  nand_x1_sg U59269 ( .A(n34958), .B(\shifter_0/reg_w_9[17] ), .X(n20648) );
  nand_x1_sg U59270 ( .A(reg_ow_9[13]), .B(n35040), .X(n20639) );
  nand_x1_sg U59271 ( .A(n30694), .B(\shifter_0/reg_w_9[13] ), .X(n20640) );
  nand_x1_sg U59272 ( .A(reg_ow_9[12]), .B(n33107), .X(n20637) );
  nand_x1_sg U59273 ( .A(n34747), .B(\shifter_0/reg_w_9[12] ), .X(n20638) );
  nand_x1_sg U59274 ( .A(reg_ow_9[9]), .B(n33075), .X(n20631) );
  nand_x1_sg U59275 ( .A(n32901), .B(\shifter_0/reg_w_9[9] ), .X(n20632) );
  nand_x1_sg U59276 ( .A(reg_ow_9[8]), .B(n31567), .X(n20629) );
  nand_x1_sg U59277 ( .A(n34748), .B(\shifter_0/reg_w_9[8] ), .X(n20630) );
  nand_x1_sg U59278 ( .A(reg_ow_9[4]), .B(n30241), .X(n20621) );
  nand_x1_sg U59279 ( .A(n30044), .B(\shifter_0/reg_w_9[4] ), .X(n20622) );
  nand_x1_sg U59280 ( .A(reg_ow_9[3]), .B(n33089), .X(n20619) );
  nand_x1_sg U59281 ( .A(n32675), .B(\shifter_0/reg_w_9[3] ), .X(n20620) );
  nand_x1_sg U59282 ( .A(reg_ow_6[18]), .B(n35048), .X(n20529) );
  nand_x1_sg U59283 ( .A(n34734), .B(\shifter_0/reg_w_6[18] ), .X(n20530) );
  nand_x1_sg U59284 ( .A(reg_ow_6[17]), .B(n31581), .X(n20527) );
  nand_x1_sg U59285 ( .A(n32521), .B(\shifter_0/reg_w_6[17] ), .X(n20528) );
  nand_x1_sg U59286 ( .A(reg_ow_6[13]), .B(n33125), .X(n20519) );
  nand_x1_sg U59287 ( .A(n34733), .B(\shifter_0/reg_w_6[13] ), .X(n20520) );
  nand_x1_sg U59288 ( .A(reg_ow_6[12]), .B(n33123), .X(n20517) );
  nand_x1_sg U59289 ( .A(n30697), .B(\shifter_0/reg_w_6[12] ), .X(n20518) );
  nand_x1_sg U59290 ( .A(reg_ow_6[9]), .B(n33112), .X(n20511) );
  nand_x1_sg U59291 ( .A(n30694), .B(\shifter_0/reg_w_6[9] ), .X(n20512) );
  nand_x1_sg U59292 ( .A(reg_ow_6[8]), .B(n33107), .X(n20509) );
  nand_x1_sg U59293 ( .A(n34738), .B(\shifter_0/reg_w_6[8] ), .X(n20510) );
  nand_x1_sg U59294 ( .A(reg_ow_6[4]), .B(n31212), .X(n20501) );
  nand_x1_sg U59295 ( .A(n31482), .B(\shifter_0/reg_w_6[4] ), .X(n20502) );
  nand_x1_sg U59296 ( .A(reg_ow_6[3]), .B(n35030), .X(n20499) );
  nand_x1_sg U59297 ( .A(n32687), .B(\shifter_0/reg_w_6[3] ), .X(n20500) );
  nand_x1_sg U59298 ( .A(reg_ow_5[18]), .B(n31577), .X(n20489) );
  nand_x1_sg U59299 ( .A(n34754), .B(\shifter_0/reg_w_5[18] ), .X(n20490) );
  nand_x1_sg U59300 ( .A(reg_ow_5[17]), .B(n33821), .X(n20487) );
  nand_x1_sg U59301 ( .A(n34103), .B(\shifter_0/reg_w_5[17] ), .X(n20488) );
  nand_x1_sg U59302 ( .A(reg_ow_5[13]), .B(n33042), .X(n20479) );
  nand_x1_sg U59303 ( .A(n32696), .B(\shifter_0/reg_w_5[13] ), .X(n20480) );
  nand_x1_sg U59304 ( .A(reg_ow_5[12]), .B(n35021), .X(n20477) );
  nand_x1_sg U59305 ( .A(n34747), .B(\shifter_0/reg_w_5[12] ), .X(n20478) );
  nand_x1_sg U59306 ( .A(reg_ow_5[9]), .B(n33080), .X(n20471) );
  nand_x1_sg U59307 ( .A(n32689), .B(\shifter_0/reg_w_5[9] ), .X(n20472) );
  nand_x1_sg U59308 ( .A(reg_ow_5[8]), .B(n33051), .X(n20469) );
  nand_x1_sg U59309 ( .A(n30693), .B(\shifter_0/reg_w_5[8] ), .X(n20470) );
  nand_x1_sg U59310 ( .A(reg_ow_5[4]), .B(n33110), .X(n20461) );
  nand_x1_sg U59311 ( .A(n30216), .B(\shifter_0/reg_w_5[4] ), .X(n20462) );
  nand_x1_sg U59312 ( .A(reg_ow_5[3]), .B(n35018), .X(n20459) );
  nand_x1_sg U59313 ( .A(n32692), .B(\shifter_0/reg_w_5[3] ), .X(n20460) );
  nand_x1_sg U59314 ( .A(reg_ow_4[19]), .B(n33074), .X(n20451) );
  nand_x1_sg U59315 ( .A(n31990), .B(\shifter_0/reg_w_4[19] ), .X(n20452) );
  nand_x1_sg U59316 ( .A(reg_ow_4[18]), .B(n33122), .X(n20449) );
  nand_x1_sg U59317 ( .A(n32637), .B(\shifter_0/reg_w_4[18] ), .X(n20450) );
  nand_x1_sg U59318 ( .A(reg_ow_4[17]), .B(n35041), .X(n20447) );
  nand_x1_sg U59319 ( .A(n34743), .B(\shifter_0/reg_w_4[17] ), .X(n20448) );
  nand_x1_sg U59320 ( .A(reg_ow_4[16]), .B(n31565), .X(n20445) );
  nand_x1_sg U59321 ( .A(n32644), .B(\shifter_0/reg_w_4[16] ), .X(n20446) );
  nand_x1_sg U59322 ( .A(reg_ow_4[15]), .B(n31566), .X(n20443) );
  nand_x1_sg U59323 ( .A(n32668), .B(\shifter_0/reg_w_4[15] ), .X(n20444) );
  nand_x1_sg U59324 ( .A(reg_ow_4[14]), .B(n35040), .X(n20441) );
  nand_x1_sg U59325 ( .A(n30640), .B(\shifter_0/reg_w_4[14] ), .X(n20442) );
  nand_x1_sg U59326 ( .A(reg_ow_4[13]), .B(n35037), .X(n20439) );
  nand_x1_sg U59327 ( .A(n30640), .B(\shifter_0/reg_w_4[13] ), .X(n20440) );
  nand_x1_sg U59328 ( .A(reg_ow_4[3]), .B(n35029), .X(n20419) );
  nand_x1_sg U59329 ( .A(n30692), .B(\shifter_0/reg_w_4[3] ), .X(n20420) );
  nand_x1_sg U59330 ( .A(reg_ow_4[2]), .B(n35021), .X(n20417) );
  nand_x1_sg U59331 ( .A(n32641), .B(\shifter_0/reg_w_4[2] ), .X(n20418) );
  nand_x1_sg U59332 ( .A(reg_ow_4[1]), .B(n33065), .X(n20415) );
  nand_x1_sg U59333 ( .A(n32684), .B(\shifter_0/reg_w_4[1] ), .X(n20416) );
  nand_x1_sg U59334 ( .A(reg_ow_4[0]), .B(n33074), .X(n20413) );
  nand_x1_sg U59335 ( .A(n34736), .B(\shifter_0/reg_w_4[0] ), .X(n20414) );
  nand_x1_sg U59336 ( .A(reg_ow_2[18]), .B(n35023), .X(n20369) );
  nand_x1_sg U59337 ( .A(n32671), .B(\shifter_0/reg_w_2[18] ), .X(n20370) );
  nand_x1_sg U59338 ( .A(reg_ow_2[17]), .B(n33064), .X(n20367) );
  nand_x1_sg U59339 ( .A(n31990), .B(\shifter_0/reg_w_2[17] ), .X(n20368) );
  nand_x1_sg U59340 ( .A(reg_ow_2[13]), .B(n33059), .X(n20359) );
  nand_x1_sg U59341 ( .A(n34746), .B(\shifter_0/reg_w_2[13] ), .X(n20360) );
  nand_x1_sg U59342 ( .A(reg_ow_2[12]), .B(n33042), .X(n20357) );
  nand_x1_sg U59343 ( .A(n32684), .B(\shifter_0/reg_w_2[12] ), .X(n20358) );
  nand_x1_sg U59344 ( .A(reg_ow_2[9]), .B(n29824), .X(n20351) );
  nand_x1_sg U59345 ( .A(n31990), .B(\shifter_0/reg_w_2[9] ), .X(n20352) );
  nand_x1_sg U59346 ( .A(reg_ow_2[8]), .B(n33106), .X(n20349) );
  nand_x1_sg U59347 ( .A(n32706), .B(\shifter_0/reg_w_2[8] ), .X(n20350) );
  nand_x1_sg U59348 ( .A(reg_ow_2[4]), .B(n29813), .X(n20341) );
  nand_x1_sg U59349 ( .A(n32901), .B(\shifter_0/reg_w_2[4] ), .X(n20342) );
  nand_x1_sg U59350 ( .A(reg_ow_2[3]), .B(n31569), .X(n20339) );
  nand_x1_sg U59351 ( .A(n31985), .B(\shifter_0/reg_w_2[3] ), .X(n20340) );
  nand_x1_sg U59352 ( .A(reg_ow_1[18]), .B(n33125), .X(n20329) );
  nand_x1_sg U59353 ( .A(n32678), .B(\shifter_0/reg_w_1[18] ), .X(n20330) );
  nand_x1_sg U59354 ( .A(reg_ow_1[17]), .B(n33082), .X(n20327) );
  nand_x1_sg U59355 ( .A(n30215), .B(\shifter_0/reg_w_1[17] ), .X(n20328) );
  nand_x1_sg U59356 ( .A(reg_ow_1[8]), .B(n33069), .X(n20309) );
  nand_x1_sg U59357 ( .A(n31476), .B(\shifter_0/reg_w_1[8] ), .X(n20310) );
  nand_x1_sg U59358 ( .A(reg_ow_1[4]), .B(n29810), .X(n20301) );
  nand_x1_sg U59359 ( .A(n34729), .B(\shifter_0/reg_w_1[4] ), .X(n20302) );
  nand_x1_sg U59360 ( .A(reg_ow_1[3]), .B(n33122), .X(n20299) );
  nand_x1_sg U59361 ( .A(n32656), .B(\shifter_0/reg_w_1[3] ), .X(n20300) );
  nand_x1_sg U59362 ( .A(reg_ow_0[15]), .B(n31577), .X(n20283) );
  nand_x1_sg U59363 ( .A(n32687), .B(\shifter_0/reg_w_0[15] ), .X(n20284) );
  nand_x1_sg U59364 ( .A(reg_ow_0[14]), .B(n33081), .X(n20281) );
  nand_x1_sg U59365 ( .A(n32645), .B(\shifter_0/reg_w_0[14] ), .X(n20282) );
  nand_x1_sg U59366 ( .A(reg_ow_0[13]), .B(n31565), .X(n20279) );
  nand_x1_sg U59367 ( .A(n30684), .B(\shifter_0/reg_w_0[13] ), .X(n20280) );
  nand_x1_sg U59368 ( .A(reg_ow_0[12]), .B(n29830), .X(n20277) );
  nand_x1_sg U59369 ( .A(n30686), .B(\shifter_0/reg_w_0[12] ), .X(n20278) );
  nand_x1_sg U59370 ( .A(reg_ow_0[11]), .B(n33052), .X(n20275) );
  nand_x1_sg U59371 ( .A(n32522), .B(\shifter_0/reg_w_0[11] ), .X(n20276) );
  nand_x1_sg U59372 ( .A(reg_ow_0[10]), .B(n29830), .X(n20273) );
  nand_x1_sg U59373 ( .A(n32663), .B(\shifter_0/reg_w_0[10] ), .X(n20274) );
  nand_x1_sg U59374 ( .A(reg_ow_0[9]), .B(n30240), .X(n20271) );
  nand_x1_sg U59375 ( .A(n32636), .B(\shifter_0/reg_w_0[9] ), .X(n20272) );
  nand_x1_sg U59376 ( .A(reg_ow_0[8]), .B(n33094), .X(n20269) );
  nand_x1_sg U59377 ( .A(n30642), .B(\shifter_0/reg_w_0[8] ), .X(n20270) );
  nand_x1_sg U59378 ( .A(reg_ow_0[7]), .B(n29833), .X(n20267) );
  nand_x1_sg U59379 ( .A(n34732), .B(\shifter_0/reg_w_0[7] ), .X(n20268) );
  nand_x1_sg U59380 ( .A(reg_ow_0[6]), .B(n33094), .X(n20265) );
  nand_x1_sg U59381 ( .A(n32647), .B(\shifter_0/reg_w_0[6] ), .X(n20266) );
  nand_x1_sg U59382 ( .A(reg_ow_0[5]), .B(n35026), .X(n20263) );
  nand_x1_sg U59383 ( .A(n34744), .B(\shifter_0/reg_w_0[5] ), .X(n20264) );
  nand_x1_sg U59384 ( .A(reg_ow_0[4]), .B(n35050), .X(n20261) );
  nand_x1_sg U59385 ( .A(n34098), .B(\shifter_0/reg_w_0[4] ), .X(n20262) );
  nand_x1_sg U59386 ( .A(reg_ow_0[3]), .B(n33821), .X(n20259) );
  nand_x1_sg U59387 ( .A(n34964), .B(\shifter_0/reg_w_0[3] ), .X(n20260) );
  nand_x1_sg U59388 ( .A(reg_ow_0[2]), .B(n29813), .X(n20257) );
  nand_x1_sg U59389 ( .A(n32695), .B(\shifter_0/reg_w_0[2] ), .X(n20258) );
  nand_x1_sg U59390 ( .A(reg_ow_0[1]), .B(n33090), .X(n20255) );
  nand_x1_sg U59391 ( .A(n30680), .B(\shifter_0/reg_w_0[1] ), .X(n20256) );
  nand_x1_sg U59392 ( .A(reg_ow_0[0]), .B(n33097), .X(n20253) );
  nand_x1_sg U59393 ( .A(n32688), .B(\shifter_0/reg_w_0[0] ), .X(n20254) );
  nand_x1_sg U59394 ( .A(reg_oi_14[16]), .B(n35035), .X(n20205) );
  nand_x1_sg U59395 ( .A(n34803), .B(\shifter_0/reg_i_14[16] ), .X(n20206) );
  nand_x1_sg U59396 ( .A(reg_oi_14[9]), .B(n33066), .X(n20191) );
  nand_x1_sg U59397 ( .A(n31472), .B(\shifter_0/reg_i_14[9] ), .X(n20192) );
  nand_x1_sg U59398 ( .A(reg_oi_14[8]), .B(n33047), .X(n20189) );
  nand_x1_sg U59399 ( .A(n32701), .B(\shifter_0/reg_i_14[8] ), .X(n20190) );
  nand_x1_sg U59400 ( .A(reg_oi_13[16]), .B(n35026), .X(n20165) );
  nand_x1_sg U59401 ( .A(n32652), .B(\shifter_0/reg_i_13[16] ), .X(n20166) );
  nand_x1_sg U59402 ( .A(reg_oi_13[13]), .B(n33121), .X(n20159) );
  nand_x1_sg U59403 ( .A(n31476), .B(\shifter_0/reg_i_13[13] ), .X(n20160) );
  nand_x1_sg U59404 ( .A(reg_oi_13[12]), .B(n31564), .X(n20157) );
  nand_x1_sg U59405 ( .A(n34966), .B(\shifter_0/reg_i_13[12] ), .X(n20158) );
  nand_x1_sg U59406 ( .A(reg_oi_13[9]), .B(n33124), .X(n20151) );
  nand_x1_sg U59407 ( .A(n32903), .B(\shifter_0/reg_i_13[9] ), .X(n20152) );
  nand_x1_sg U59408 ( .A(reg_oi_13[8]), .B(n31590), .X(n20149) );
  nand_x1_sg U59409 ( .A(n34737), .B(\shifter_0/reg_i_13[8] ), .X(n20150) );
  nand_x1_sg U59410 ( .A(reg_oi_12[16]), .B(n29801), .X(n20125) );
  nand_x1_sg U59411 ( .A(n32683), .B(\shifter_0/reg_i_12[16] ), .X(n20126) );
  nand_x1_sg U59412 ( .A(reg_oi_12[13]), .B(n29818), .X(n20119) );
  nand_x1_sg U59413 ( .A(n34959), .B(\shifter_0/reg_i_12[13] ), .X(n20120) );
  nand_x1_sg U59414 ( .A(reg_oi_12[12]), .B(n33065), .X(n20117) );
  nand_x1_sg U59415 ( .A(n30686), .B(\shifter_0/reg_i_12[12] ), .X(n20118) );
  nand_x1_sg U59416 ( .A(reg_oi_12[9]), .B(n30602), .X(n20111) );
  nand_x1_sg U59417 ( .A(n34752), .B(\shifter_0/reg_i_12[9] ), .X(n20112) );
  nand_x1_sg U59418 ( .A(reg_oi_11[16]), .B(n33116), .X(n20085) );
  nand_x1_sg U59419 ( .A(n31475), .B(\shifter_0/reg_i_11[16] ), .X(n20086) );
  nand_x1_sg U59420 ( .A(reg_oi_11[13]), .B(n33075), .X(n20079) );
  nand_x1_sg U59421 ( .A(n31235), .B(\shifter_0/reg_i_11[13] ), .X(n20080) );
  nand_x1_sg U59422 ( .A(reg_oi_11[12]), .B(n30240), .X(n20077) );
  nand_x1_sg U59423 ( .A(n34964), .B(\shifter_0/reg_i_11[12] ), .X(n20078) );
  nand_x1_sg U59424 ( .A(reg_oi_11[9]), .B(n33078), .X(n20071) );
  nand_x1_sg U59425 ( .A(n32656), .B(\shifter_0/reg_i_11[9] ), .X(n20072) );
  nand_x1_sg U59426 ( .A(reg_oi_11[8]), .B(n31214), .X(n20069) );
  nand_x1_sg U59427 ( .A(n32673), .B(\shifter_0/reg_i_11[8] ), .X(n20070) );
  nand_x1_sg U59428 ( .A(reg_oi_9[16]), .B(n33094), .X(n20005) );
  nand_x1_sg U59429 ( .A(n34961), .B(\shifter_0/reg_i_9[16] ), .X(n20006) );
  nand_x1_sg U59430 ( .A(reg_oi_9[13]), .B(n33118), .X(n19999) );
  nand_x1_sg U59431 ( .A(n34749), .B(\shifter_0/reg_i_9[13] ), .X(n20000) );
  nand_x1_sg U59432 ( .A(reg_oi_9[12]), .B(n33085), .X(n19997) );
  nand_x1_sg U59433 ( .A(n34743), .B(\shifter_0/reg_i_9[12] ), .X(n19998) );
  nand_x1_sg U59434 ( .A(reg_oi_9[9]), .B(n35042), .X(n19991) );
  nand_x1_sg U59435 ( .A(n32653), .B(\shifter_0/reg_i_9[9] ), .X(n19992) );
  nand_x1_sg U59436 ( .A(reg_oi_9[8]), .B(n33045), .X(n19989) );
  nand_x1_sg U59437 ( .A(n31860), .B(\shifter_0/reg_i_9[8] ), .X(n19990) );
  nand_x1_sg U59438 ( .A(reg_oi_6[18]), .B(n31111), .X(n19889) );
  nand_x1_sg U59439 ( .A(n32649), .B(\shifter_0/reg_i_6[18] ), .X(n19890) );
  nand_x1_sg U59440 ( .A(reg_oi_6[17]), .B(n29831), .X(n19887) );
  nand_x1_sg U59441 ( .A(n32637), .B(\shifter_0/reg_i_6[17] ), .X(n19888) );
  nand_x1_sg U59442 ( .A(reg_oi_6[13]), .B(n33076), .X(n19879) );
  nand_x1_sg U59443 ( .A(n31988), .B(\shifter_0/reg_i_6[13] ), .X(n19880) );
  nand_x1_sg U59444 ( .A(reg_oi_6[12]), .B(n33090), .X(n19877) );
  nand_x1_sg U59445 ( .A(n34966), .B(\shifter_0/reg_i_6[12] ), .X(n19878) );
  nand_x1_sg U59446 ( .A(reg_oi_6[9]), .B(n33061), .X(n19871) );
  nand_x1_sg U59447 ( .A(n32665), .B(\shifter_0/reg_i_6[9] ), .X(n19872) );
  nand_x1_sg U59448 ( .A(reg_oi_6[8]), .B(n33074), .X(n19869) );
  nand_x1_sg U59449 ( .A(n34731), .B(\shifter_0/reg_i_6[8] ), .X(n19870) );
  nand_x1_sg U59450 ( .A(reg_oi_6[4]), .B(n30563), .X(n19861) );
  nand_x1_sg U59451 ( .A(n30045), .B(\shifter_0/reg_i_6[4] ), .X(n19862) );
  nand_x1_sg U59452 ( .A(reg_oi_6[3]), .B(n31586), .X(n19859) );
  nand_x1_sg U59453 ( .A(n31986), .B(\shifter_0/reg_i_6[3] ), .X(n19860) );
  nand_x1_sg U59454 ( .A(reg_oi_5[18]), .B(n33085), .X(n19849) );
  nand_x1_sg U59455 ( .A(n32701), .B(\shifter_0/reg_i_5[18] ), .X(n19850) );
  nand_x1_sg U59456 ( .A(reg_oi_5[17]), .B(n31583), .X(n19847) );
  nand_x1_sg U59457 ( .A(n34731), .B(\shifter_0/reg_i_5[17] ), .X(n19848) );
  nand_x1_sg U59458 ( .A(reg_oi_5[13]), .B(n33126), .X(n19839) );
  nand_x1_sg U59459 ( .A(n30686), .B(\shifter_0/reg_i_5[13] ), .X(n19840) );
  nand_x1_sg U59460 ( .A(reg_oi_5[12]), .B(n35038), .X(n19837) );
  nand_x1_sg U59461 ( .A(n32705), .B(\shifter_0/reg_i_5[12] ), .X(n19838) );
  nand_x1_sg U59462 ( .A(reg_oi_5[9]), .B(n33053), .X(n19831) );
  nand_x1_sg U59463 ( .A(n31232), .B(\shifter_0/reg_i_5[9] ), .X(n19832) );
  nand_x1_sg U59464 ( .A(reg_oi_4[19]), .B(n33076), .X(n19811) );
  nand_x1_sg U59465 ( .A(n34725), .B(\shifter_0/reg_i_4[19] ), .X(n19812) );
  nand_x1_sg U59466 ( .A(reg_oi_4[18]), .B(n30246), .X(n19809) );
  nand_x1_sg U59467 ( .A(n34730), .B(\shifter_0/reg_i_4[18] ), .X(n19810) );
  nand_x1_sg U59468 ( .A(reg_oi_4[17]), .B(n33054), .X(n19807) );
  nand_x1_sg U59469 ( .A(n34732), .B(\shifter_0/reg_i_4[17] ), .X(n19808) );
  nand_x1_sg U59470 ( .A(reg_oi_4[16]), .B(n31583), .X(n19805) );
  nand_x1_sg U59471 ( .A(n32688), .B(\shifter_0/reg_i_4[16] ), .X(n19806) );
  nand_x1_sg U59472 ( .A(reg_oi_4[15]), .B(n35029), .X(n19803) );
  nand_x1_sg U59473 ( .A(n30689), .B(\shifter_0/reg_i_4[15] ), .X(n19804) );
  nand_x1_sg U59474 ( .A(reg_oi_4[14]), .B(n33820), .X(n19801) );
  nand_x1_sg U59475 ( .A(n32670), .B(\shifter_0/reg_i_4[14] ), .X(n19802) );
  nand_x1_sg U59476 ( .A(reg_oi_4[13]), .B(n33129), .X(n19799) );
  nand_x1_sg U59477 ( .A(n32673), .B(\shifter_0/reg_i_4[13] ), .X(n19800) );
  nand_x1_sg U59478 ( .A(reg_oi_4[12]), .B(n33046), .X(n19797) );
  nand_x1_sg U59479 ( .A(n31236), .B(\shifter_0/reg_i_4[12] ), .X(n19798) );
  nand_x1_sg U59480 ( .A(reg_oi_4[11]), .B(n33068), .X(n19795) );
  nand_x1_sg U59481 ( .A(n32707), .B(\shifter_0/reg_i_4[11] ), .X(n19796) );
  nand_x1_sg U59482 ( .A(reg_oi_4[10]), .B(n33080), .X(n19793) );
  nand_x1_sg U59483 ( .A(n34751), .B(\shifter_0/reg_i_4[10] ), .X(n19794) );
  nand_x1_sg U59484 ( .A(reg_oi_4[9]), .B(n33098), .X(n19791) );
  nand_x1_sg U59485 ( .A(n34741), .B(\shifter_0/reg_i_4[9] ), .X(n19792) );
  nand_x1_sg U59486 ( .A(reg_oi_4[8]), .B(n31585), .X(n19789) );
  nand_x1_sg U59487 ( .A(n34753), .B(\shifter_0/reg_i_4[8] ), .X(n19790) );
  nand_x1_sg U59488 ( .A(reg_oi_4[7]), .B(n29833), .X(n19787) );
  nand_x1_sg U59489 ( .A(n31488), .B(\shifter_0/reg_i_4[7] ), .X(n19788) );
  nand_x1_sg U59490 ( .A(reg_oi_4[6]), .B(n33077), .X(n19785) );
  nand_x1_sg U59491 ( .A(n32677), .B(\shifter_0/reg_i_4[6] ), .X(n19786) );
  nand_x1_sg U59492 ( .A(reg_oi_4[5]), .B(n33086), .X(n19783) );
  nand_x1_sg U59493 ( .A(n30696), .B(\shifter_0/reg_i_4[5] ), .X(n19784) );
  nand_x1_sg U59494 ( .A(reg_oi_4[4]), .B(n33057), .X(n19781) );
  nand_x1_sg U59495 ( .A(n32649), .B(\shifter_0/reg_i_4[4] ), .X(n19782) );
  nand_x1_sg U59496 ( .A(reg_oi_4[3]), .B(n33092), .X(n19779) );
  nand_x1_sg U59497 ( .A(n30682), .B(\shifter_0/reg_i_4[3] ), .X(n19780) );
  nand_x1_sg U59498 ( .A(reg_oi_4[2]), .B(n31111), .X(n19777) );
  nand_x1_sg U59499 ( .A(n34741), .B(\shifter_0/reg_i_4[2] ), .X(n19778) );
  nand_x1_sg U59500 ( .A(reg_oi_4[1]), .B(n31586), .X(n19775) );
  nand_x1_sg U59501 ( .A(n32664), .B(\shifter_0/reg_i_4[1] ), .X(n19776) );
  nand_x1_sg U59502 ( .A(reg_oi_4[0]), .B(n29836), .X(n19773) );
  nand_x1_sg U59503 ( .A(n31488), .B(\shifter_0/reg_i_4[0] ), .X(n19774) );
  nand_x1_sg U59504 ( .A(reg_oi_2[18]), .B(n33821), .X(n19729) );
  nand_x1_sg U59505 ( .A(n32704), .B(\shifter_0/reg_i_2[18] ), .X(n19730) );
  nand_x1_sg U59506 ( .A(reg_oi_2[17]), .B(n31562), .X(n19727) );
  nand_x1_sg U59507 ( .A(n32704), .B(\shifter_0/reg_i_2[17] ), .X(n19728) );
  nand_x1_sg U59508 ( .A(reg_oi_2[13]), .B(n33052), .X(n19719) );
  nand_x1_sg U59509 ( .A(n30692), .B(\shifter_0/reg_i_2[13] ), .X(n19720) );
  nand_x1_sg U59510 ( .A(reg_oi_2[12]), .B(n33819), .X(n19717) );
  nand_x1_sg U59511 ( .A(n34111), .B(\shifter_0/reg_i_2[12] ), .X(n19718) );
  nand_x1_sg U59512 ( .A(reg_oi_2[8]), .B(n33064), .X(n19709) );
  nand_x1_sg U59513 ( .A(n31986), .B(\shifter_0/reg_i_2[8] ), .X(n19710) );
  nand_x1_sg U59514 ( .A(reg_oi_2[4]), .B(n33101), .X(n19701) );
  nand_x1_sg U59515 ( .A(n31485), .B(\shifter_0/reg_i_2[4] ), .X(n19702) );
  nand_x1_sg U59516 ( .A(reg_oi_2[3]), .B(n33083), .X(n19699) );
  nand_x1_sg U59517 ( .A(n31988), .B(\shifter_0/reg_i_2[3] ), .X(n19700) );
  nand_x1_sg U59518 ( .A(reg_oi_1[9]), .B(n30974), .X(n19671) );
  nand_x1_sg U59519 ( .A(n32649), .B(\shifter_0/reg_i_1[9] ), .X(n19672) );
  nand_x1_sg U59520 ( .A(reg_oi_1[8]), .B(n33081), .X(n19669) );
  nand_x1_sg U59521 ( .A(n32694), .B(\shifter_0/reg_i_1[8] ), .X(n19670) );
  nand_x1_sg U59522 ( .A(reg_oi_1[4]), .B(n31564), .X(n19661) );
  nand_x1_sg U59523 ( .A(n32654), .B(\shifter_0/reg_i_1[4] ), .X(n19662) );
  nand_x1_sg U59524 ( .A(reg_oi_1[3]), .B(n31587), .X(n19659) );
  nand_x1_sg U59525 ( .A(n32645), .B(\shifter_0/reg_i_1[3] ), .X(n19660) );
  nand_x1_sg U59526 ( .A(reg_oi_0[19]), .B(n33088), .X(n19651) );
  nand_x1_sg U59527 ( .A(n32707), .B(\shifter_0/reg_i_0[19] ), .X(n19652) );
  nand_x1_sg U59528 ( .A(reg_oi_0[18]), .B(n31591), .X(n19649) );
  nand_x1_sg U59529 ( .A(n34801), .B(\shifter_0/reg_i_0[18] ), .X(n19650) );
  nand_x1_sg U59530 ( .A(reg_oi_0[17]), .B(n35037), .X(n19647) );
  nand_x1_sg U59531 ( .A(n34102), .B(\shifter_0/reg_i_0[17] ), .X(n19648) );
  nand_x1_sg U59532 ( .A(reg_oi_0[16]), .B(n29810), .X(n19645) );
  nand_x1_sg U59533 ( .A(n31487), .B(\shifter_0/reg_i_0[16] ), .X(n19646) );
  nand_x1_sg U59534 ( .A(reg_oi_0[15]), .B(n35044), .X(n19643) );
  nand_x1_sg U59535 ( .A(n32648), .B(\shifter_0/reg_i_0[15] ), .X(n19644) );
  nand_x1_sg U59536 ( .A(reg_oi_0[14]), .B(n29829), .X(n19641) );
  nand_x1_sg U59537 ( .A(n31989), .B(\shifter_0/reg_i_0[14] ), .X(n19642) );
  nand_x1_sg U59538 ( .A(reg_oi_0[13]), .B(n35046), .X(n19639) );
  nand_x1_sg U59539 ( .A(n30045), .B(\shifter_0/reg_i_0[13] ), .X(n19640) );
  nand_x1_sg U59540 ( .A(reg_oi_0[12]), .B(n29831), .X(n19637) );
  nand_x1_sg U59541 ( .A(n30702), .B(\shifter_0/reg_i_0[12] ), .X(n19638) );
  nand_x1_sg U59542 ( .A(reg_oi_0[11]), .B(n33128), .X(n19635) );
  nand_x1_sg U59543 ( .A(n32684), .B(\shifter_0/reg_i_0[11] ), .X(n19636) );
  nand_x1_sg U59544 ( .A(reg_oi_0[10]), .B(n33093), .X(n19633) );
  nand_x1_sg U59545 ( .A(n30640), .B(\shifter_0/reg_i_0[10] ), .X(n19634) );
  nand_x1_sg U59546 ( .A(reg_oi_0[9]), .B(n33101), .X(n19631) );
  nand_x1_sg U59547 ( .A(n34732), .B(\shifter_0/reg_i_0[9] ), .X(n19632) );
  nand_x1_sg U59548 ( .A(reg_oi_0[8]), .B(n29810), .X(n19629) );
  nand_x1_sg U59549 ( .A(n34736), .B(\shifter_0/reg_i_0[8] ), .X(n19630) );
  nand_x1_sg U59550 ( .A(reg_oi_0[7]), .B(n35027), .X(n19627) );
  nand_x1_sg U59551 ( .A(n30680), .B(\shifter_0/reg_i_0[7] ), .X(n19628) );
  nand_x1_sg U59552 ( .A(reg_oi_0[6]), .B(n35037), .X(n19625) );
  nand_x1_sg U59553 ( .A(n34103), .B(\shifter_0/reg_i_0[6] ), .X(n19626) );
  nand_x1_sg U59554 ( .A(reg_oi_0[5]), .B(n33064), .X(n19623) );
  nand_x1_sg U59555 ( .A(n32700), .B(\shifter_0/reg_i_0[5] ), .X(n19624) );
  nand_x1_sg U59556 ( .A(reg_oi_0[4]), .B(n31585), .X(n19621) );
  nand_x1_sg U59557 ( .A(n31482), .B(\shifter_0/reg_i_0[4] ), .X(n19622) );
  nand_x1_sg U59558 ( .A(reg_oi_0[3]), .B(n33073), .X(n19619) );
  nand_x1_sg U59559 ( .A(n34802), .B(\shifter_0/reg_i_0[3] ), .X(n19620) );
  nand_x1_sg U59560 ( .A(reg_oi_0[2]), .B(n29818), .X(n19617) );
  nand_x1_sg U59561 ( .A(n30641), .B(\shifter_0/reg_i_0[2] ), .X(n19618) );
  nand_x1_sg U59562 ( .A(reg_oi_0[1]), .B(n33125), .X(n19615) );
  nand_x1_sg U59563 ( .A(n32904), .B(\shifter_0/reg_i_0[1] ), .X(n19616) );
  nand_x1_sg U59564 ( .A(reg_oi_0[0]), .B(n35045), .X(n19613) );
  nand_x1_sg U59565 ( .A(n31486), .B(\shifter_0/reg_i_0[0] ), .X(n19614) );
  nand_x1_sg U59566 ( .A(reg_oi_8[18]), .B(n33073), .X(n19969) );
  nand_x1_sg U59567 ( .A(n34413), .B(\shifter_0/reg_i_8[18] ), .X(n19970) );
  nand_x1_sg U59568 ( .A(reg_oi_8[17]), .B(n33062), .X(n19967) );
  nand_x1_sg U59569 ( .A(n34748), .B(\shifter_0/reg_i_8[17] ), .X(n19968) );
  nand_x1_sg U59570 ( .A(reg_oi_15[17]), .B(n33122), .X(n20247) );
  nand_x1_sg U59571 ( .A(n34802), .B(n30453), .X(n20248) );
  nand_x1_sg U59572 ( .A(reg_oi_15[2]), .B(n33106), .X(n20217) );
  nand_x1_sg U59573 ( .A(n31488), .B(n30447), .X(n20218) );
  nand_x1_sg U59574 ( .A(reg_oi_7[18]), .B(n33068), .X(n19929) );
  nand_x1_sg U59575 ( .A(n32647), .B(n30404), .X(n19930) );
  nand_x1_sg U59576 ( .A(reg_oi_7[17]), .B(n33078), .X(n19927) );
  nand_x1_sg U59577 ( .A(n34414), .B(n30403), .X(n19928) );
  nand_x1_sg U59578 ( .A(reg_oi_7[2]), .B(n31568), .X(n19897) );
  nand_x1_sg U59579 ( .A(n32526), .B(n30402), .X(n19898) );
  nand_x1_sg U59580 ( .A(reg_oi_15[18]), .B(n33042), .X(n20249) );
  nand_x1_sg U59581 ( .A(n31861), .B(\shifter_0/reg_i_15[18] ), .X(n20250) );
  nand_x1_sg U59582 ( .A(reg_oi_15[4]), .B(n33056), .X(n20221) );
  nand_x1_sg U59583 ( .A(n32665), .B(\shifter_0/reg_i_15[4] ), .X(n20222) );
  nand_x1_sg U59584 ( .A(reg_oi_7[4]), .B(n33049), .X(n19901) );
  nand_x1_sg U59585 ( .A(n32651), .B(\shifter_0/reg_i_7[4] ), .X(n19902) );
  nand_x1_sg U59586 ( .A(reg_ow_7[19]), .B(n31572), .X(n20571) );
  nand_x1_sg U59587 ( .A(n30685), .B(\shifter_0/reg_w_7[19] ), .X(n20572) );
  nand_x1_sg U59588 ( .A(reg_ow_7[18]), .B(n31214), .X(n20569) );
  nand_x1_sg U59589 ( .A(n30702), .B(\shifter_0/reg_w_7[18] ), .X(n20570) );
  nand_x1_sg U59590 ( .A(reg_ow_7[17]), .B(n31582), .X(n20567) );
  nand_x1_sg U59591 ( .A(n32663), .B(\shifter_0/reg_w_7[17] ), .X(n20568) );
  nand_x1_sg U59592 ( .A(reg_ow_7[16]), .B(n33106), .X(n20565) );
  nand_x1_sg U59593 ( .A(n32637), .B(\shifter_0/reg_w_7[16] ), .X(n20566) );
  nand_x1_sg U59594 ( .A(reg_ow_7[15]), .B(n33051), .X(n20563) );
  nand_x1_sg U59595 ( .A(n34739), .B(\shifter_0/reg_w_7[15] ), .X(n20564) );
  nand_x1_sg U59596 ( .A(reg_ow_7[14]), .B(n33057), .X(n20561) );
  nand_x1_sg U59597 ( .A(n32666), .B(\shifter_0/reg_w_7[14] ), .X(n20562) );
  nand_x1_sg U59598 ( .A(reg_ow_7[13]), .B(n35042), .X(n20559) );
  nand_x1_sg U59599 ( .A(n32636), .B(\shifter_0/reg_w_7[13] ), .X(n20560) );
  nand_x1_sg U59600 ( .A(reg_ow_7[12]), .B(n35025), .X(n20557) );
  nand_x1_sg U59601 ( .A(n34729), .B(\shifter_0/reg_w_7[12] ), .X(n20558) );
  nand_x1_sg U59602 ( .A(reg_ow_7[2]), .B(n35049), .X(n20537) );
  nand_x1_sg U59603 ( .A(n30685), .B(\shifter_0/reg_w_7[2] ), .X(n20538) );
  nand_x1_sg U59604 ( .A(reg_ow_7[1]), .B(n31581), .X(n20535) );
  nand_x1_sg U59605 ( .A(n30689), .B(\shifter_0/reg_w_7[1] ), .X(n20536) );
  nand_x1_sg U59606 ( .A(reg_ow_7[0]), .B(n33071), .X(n20533) );
  nand_x1_sg U59607 ( .A(n32902), .B(\shifter_0/reg_w_7[0] ), .X(n20534) );
  nand_x1_sg U59608 ( .A(reg_oi_7[16]), .B(n35026), .X(n19925) );
  nand_x1_sg U59609 ( .A(n34965), .B(\shifter_0/reg_i_7[16] ), .X(n19926) );
  nand_x1_sg U59610 ( .A(reg_oi_7[15]), .B(n33822), .X(n19923) );
  nand_x1_sg U59611 ( .A(n34753), .B(\shifter_0/reg_i_7[15] ), .X(n19924) );
  nand_x1_sg U59612 ( .A(reg_oi_7[14]), .B(n33128), .X(n19921) );
  nand_x1_sg U59613 ( .A(n34733), .B(\shifter_0/reg_i_7[14] ), .X(n19922) );
  nand_x1_sg U59614 ( .A(reg_oi_7[13]), .B(n33121), .X(n19919) );
  nand_x1_sg U59615 ( .A(n32683), .B(\shifter_0/reg_i_7[13] ), .X(n19920) );
  nand_x1_sg U59616 ( .A(reg_oi_7[12]), .B(n33088), .X(n19917) );
  nand_x1_sg U59617 ( .A(n31486), .B(\shifter_0/reg_i_7[12] ), .X(n19918) );
  nand_x1_sg U59618 ( .A(reg_oi_7[11]), .B(n29813), .X(n19915) );
  nand_x1_sg U59619 ( .A(n34099), .B(\shifter_0/reg_i_7[11] ), .X(n19916) );
  nand_x1_sg U59620 ( .A(reg_oi_7[10]), .B(n33119), .X(n19913) );
  nand_x1_sg U59621 ( .A(n32675), .B(\shifter_0/reg_i_7[10] ), .X(n19914) );
  nand_x1_sg U59622 ( .A(reg_oi_7[9]), .B(n33046), .X(n19911) );
  nand_x1_sg U59623 ( .A(n32671), .B(\shifter_0/reg_i_7[9] ), .X(n19912) );
  nand_x1_sg U59624 ( .A(reg_oi_7[8]), .B(n29818), .X(n19909) );
  nand_x1_sg U59625 ( .A(n34749), .B(\shifter_0/reg_i_7[8] ), .X(n19910) );
  nand_x1_sg U59626 ( .A(reg_oi_7[7]), .B(n35027), .X(n19907) );
  nand_x1_sg U59627 ( .A(n34739), .B(\shifter_0/reg_i_7[7] ), .X(n19908) );
  nand_x1_sg U59628 ( .A(reg_oi_7[6]), .B(n33110), .X(n19905) );
  nand_x1_sg U59629 ( .A(n30701), .B(\shifter_0/reg_i_7[6] ), .X(n19906) );
  nand_x1_sg U59630 ( .A(reg_oi_7[5]), .B(n33078), .X(n19903) );
  nand_x1_sg U59631 ( .A(n32648), .B(\shifter_0/reg_i_7[5] ), .X(n19904) );
  nand_x1_sg U59632 ( .A(reg_oi_7[3]), .B(n31562), .X(n19899) );
  nand_x1_sg U59633 ( .A(n32527), .B(\shifter_0/reg_i_7[3] ), .X(n19900) );
  nand_x1_sg U59634 ( .A(reg_oi_7[1]), .B(n30973), .X(n19895) );
  nand_x1_sg U59635 ( .A(n30641), .B(\shifter_0/reg_i_7[1] ), .X(n19896) );
  nand_x1_sg U59636 ( .A(reg_oi_7[0]), .B(n35020), .X(n19893) );
  nand_x1_sg U59637 ( .A(n34753), .B(\shifter_0/reg_i_7[0] ), .X(n19894) );
  nand_x1_sg U59638 ( .A(reg_ow_10[10]), .B(n29831), .X(n20673) );
  nand_x1_sg U59639 ( .A(n32659), .B(\shifter_0/reg_w_10[10] ), .X(n20674) );
  nand_x1_sg U59640 ( .A(reg_ow_10[9]), .B(n33087), .X(n20671) );
  nand_x1_sg U59641 ( .A(n32903), .B(\shifter_0/reg_w_10[9] ), .X(n20672) );
  nand_x1_sg U59642 ( .A(reg_ow_10[8]), .B(n35047), .X(n20669) );
  nand_x1_sg U59643 ( .A(n31485), .B(\shifter_0/reg_w_10[8] ), .X(n20670) );
  nand_x1_sg U59644 ( .A(reg_ow_10[7]), .B(n35030), .X(n20667) );
  nand_x1_sg U59645 ( .A(n32659), .B(\shifter_0/reg_w_10[7] ), .X(n20668) );
  nand_x1_sg U59646 ( .A(reg_ow_10[6]), .B(n33068), .X(n20665) );
  nand_x1_sg U59647 ( .A(n30696), .B(\shifter_0/reg_w_10[6] ), .X(n20666) );
  nand_x1_sg U59648 ( .A(reg_ow_10[5]), .B(n33093), .X(n20663) );
  nand_x1_sg U59649 ( .A(n29761), .B(\shifter_0/reg_w_10[5] ), .X(n20664) );
  nand_x1_sg U59650 ( .A(reg_ow_10[4]), .B(n33109), .X(n20661) );
  nand_x1_sg U59651 ( .A(n32672), .B(\shifter_0/reg_w_10[4] ), .X(n20662) );
  nand_x1_sg U59652 ( .A(reg_ow_10[3]), .B(n33119), .X(n20659) );
  nand_x1_sg U59653 ( .A(n34099), .B(\shifter_0/reg_w_10[3] ), .X(n20660) );
  nand_x1_sg U59654 ( .A(reg_ow_10[2]), .B(n31586), .X(n20657) );
  nand_x1_sg U59655 ( .A(n32681), .B(\shifter_0/reg_w_10[2] ), .X(n20658) );
  nand_x1_sg U59656 ( .A(reg_oi_10[19]), .B(n33093), .X(n20051) );
  nand_x1_sg U59657 ( .A(n34109), .B(\shifter_0/reg_i_10[19] ), .X(n20052) );
  nand_x1_sg U59658 ( .A(reg_ow_1[11]), .B(n31580), .X(n20315) );
  nand_x1_sg U59659 ( .A(n34734), .B(\shifter_0/reg_w_1[11] ), .X(n20316) );
  nand_x1_sg U59660 ( .A(reg_ow_1[10]), .B(n29815), .X(n20313) );
  nand_x1_sg U59661 ( .A(n30216), .B(\shifter_0/reg_w_1[10] ), .X(n20314) );
  nand_x1_sg U59662 ( .A(reg_oi_14[4]), .B(n31571), .X(n20181) );
  nand_x1_sg U59663 ( .A(n34734), .B(\shifter_0/reg_i_14[4] ), .X(n20182) );
  nand_x1_sg U59664 ( .A(reg_oi_14[2]), .B(n33070), .X(n20177) );
  nand_x1_sg U59665 ( .A(n34752), .B(\shifter_0/reg_i_14[2] ), .X(n20178) );
  nand_x1_sg U59666 ( .A(reg_oi_13[18]), .B(n33045), .X(n20169) );
  nand_x1_sg U59667 ( .A(n30701), .B(\shifter_0/reg_i_13[18] ), .X(n20170) );
  nand_x1_sg U59668 ( .A(reg_oi_13[17]), .B(n33111), .X(n20167) );
  nand_x1_sg U59669 ( .A(n30696), .B(\shifter_0/reg_i_13[17] ), .X(n20168) );
  nand_x1_sg U59670 ( .A(reg_oi_11[4]), .B(n35043), .X(n20061) );
  nand_x1_sg U59671 ( .A(n32640), .B(\shifter_0/reg_i_11[4] ), .X(n20062) );
  nand_x1_sg U59672 ( .A(reg_oi_11[2]), .B(n31573), .X(n20057) );
  nand_x1_sg U59673 ( .A(n32636), .B(\shifter_0/reg_i_11[2] ), .X(n20058) );
  nand_x1_sg U59674 ( .A(reg_oi_10[18]), .B(n33083), .X(n20049) );
  nand_x1_sg U59675 ( .A(n34802), .B(\shifter_0/reg_i_10[18] ), .X(n20050) );
  nand_x1_sg U59676 ( .A(reg_oi_1[19]), .B(n33130), .X(n19691) );
  nand_x1_sg U59677 ( .A(n29772), .B(\shifter_0/reg_i_1[19] ), .X(n19692) );
  nand_x1_sg U59678 ( .A(reg_oi_1[16]), .B(n33126), .X(n19685) );
  nand_x1_sg U59679 ( .A(n32671), .B(\shifter_0/reg_i_1[16] ), .X(n19686) );
  nand_x1_sg U59680 ( .A(reg_oi_1[15]), .B(n33099), .X(n19683) );
  nand_x1_sg U59681 ( .A(n32656), .B(\shifter_0/reg_i_1[15] ), .X(n19684) );
  nand_x1_sg U59682 ( .A(reg_oi_1[14]), .B(n29801), .X(n19681) );
  nand_x1_sg U59683 ( .A(n34803), .B(\shifter_0/reg_i_1[14] ), .X(n19682) );
  nand_x1_sg U59684 ( .A(reg_ow_13[10]), .B(n33069), .X(n20793) );
  nand_x1_sg U59685 ( .A(n32642), .B(\shifter_0/reg_w_13[10] ), .X(n20794) );
  nand_x1_sg U59686 ( .A(reg_ow_13[7]), .B(n29826), .X(n20787) );
  nand_x1_sg U59687 ( .A(n32689), .B(\shifter_0/reg_w_13[7] ), .X(n20788) );
  nand_x1_sg U59688 ( .A(reg_ow_13[6]), .B(n31587), .X(n20785) );
  nand_x1_sg U59689 ( .A(n32665), .B(\shifter_0/reg_w_13[6] ), .X(n20786) );
  nand_x1_sg U59690 ( .A(reg_ow_13[5]), .B(n35046), .X(n20783) );
  nand_x1_sg U59691 ( .A(n31486), .B(\shifter_0/reg_w_13[5] ), .X(n20784) );
  nand_x1_sg U59692 ( .A(reg_ow_13[2]), .B(n31590), .X(n20777) );
  nand_x1_sg U59693 ( .A(n32697), .B(\shifter_0/reg_w_13[2] ), .X(n20778) );
  nand_x1_sg U59694 ( .A(reg_ow_13[1]), .B(n33080), .X(n20775) );
  nand_x1_sg U59695 ( .A(n32701), .B(\shifter_0/reg_w_13[1] ), .X(n20776) );
  nand_x1_sg U59696 ( .A(reg_ow_11[7]), .B(n31570), .X(n20707) );
  nand_x1_sg U59697 ( .A(n34804), .B(\shifter_0/reg_w_11[7] ), .X(n20708) );
  nand_x1_sg U59698 ( .A(reg_ow_11[6]), .B(n33069), .X(n20705) );
  nand_x1_sg U59699 ( .A(n32902), .B(\shifter_0/reg_w_11[6] ), .X(n20706) );
  nand_x1_sg U59700 ( .A(reg_ow_11[5]), .B(n33121), .X(n20703) );
  nand_x1_sg U59701 ( .A(n32692), .B(\shifter_0/reg_w_11[5] ), .X(n20704) );
  nand_x1_sg U59702 ( .A(reg_ow_11[2]), .B(n33114), .X(n20697) );
  nand_x1_sg U59703 ( .A(n31859), .B(\shifter_0/reg_w_11[2] ), .X(n20698) );
  nand_x1_sg U59704 ( .A(reg_ow_11[1]), .B(n31586), .X(n20695) );
  nand_x1_sg U59705 ( .A(n32702), .B(\shifter_0/reg_w_11[1] ), .X(n20696) );
  nand_x1_sg U59706 ( .A(reg_oi_14[14]), .B(n31584), .X(n20201) );
  nand_x1_sg U59707 ( .A(n30682), .B(\shifter_0/reg_i_14[14] ), .X(n20202) );
  nand_x1_sg U59708 ( .A(reg_oi_14[11]), .B(n33095), .X(n20195) );
  nand_x1_sg U59709 ( .A(n30690), .B(\shifter_0/reg_i_14[11] ), .X(n20196) );
  nand_x1_sg U59710 ( .A(reg_oi_14[10]), .B(n33087), .X(n20193) );
  nand_x1_sg U59711 ( .A(n32673), .B(\shifter_0/reg_i_14[10] ), .X(n20194) );
  nand_x1_sg U59712 ( .A(reg_oi_14[5]), .B(n35037), .X(n20183) );
  nand_x1_sg U59713 ( .A(n32642), .B(\shifter_0/reg_i_14[5] ), .X(n20184) );
  nand_x1_sg U59714 ( .A(reg_oi_14[3]), .B(n33128), .X(n20179) );
  nand_x1_sg U59715 ( .A(n30690), .B(\shifter_0/reg_i_14[3] ), .X(n20180) );
  nand_x1_sg U59716 ( .A(reg_oi_14[1]), .B(n35016), .X(n20175) );
  nand_x1_sg U59717 ( .A(n30701), .B(\shifter_0/reg_i_14[1] ), .X(n20176) );
  nand_x1_sg U59718 ( .A(reg_oi_14[0]), .B(n35046), .X(n20173) );
  nand_x1_sg U59719 ( .A(n32684), .B(\shifter_0/reg_i_14[0] ), .X(n20174) );
  nand_x1_sg U59720 ( .A(reg_oi_13[19]), .B(n33126), .X(n20171) );
  nand_x1_sg U59721 ( .A(n30684), .B(\shifter_0/reg_i_13[19] ), .X(n20172) );
  nand_x1_sg U59722 ( .A(reg_oi_12[7]), .B(n30246), .X(n20107) );
  nand_x1_sg U59723 ( .A(n32693), .B(\shifter_0/reg_i_12[7] ), .X(n20108) );
  nand_x1_sg U59724 ( .A(reg_oi_12[6]), .B(n33119), .X(n20105) );
  nand_x1_sg U59725 ( .A(n32685), .B(\shifter_0/reg_i_12[6] ), .X(n20106) );
  nand_x1_sg U59726 ( .A(reg_oi_12[5]), .B(n35039), .X(n20103) );
  nand_x1_sg U59727 ( .A(n32639), .B(\shifter_0/reg_i_12[5] ), .X(n20104) );
  nand_x1_sg U59728 ( .A(reg_oi_11[6]), .B(n33053), .X(n20065) );
  nand_x1_sg U59729 ( .A(n31232), .B(\shifter_0/reg_i_11[6] ), .X(n20066) );
  nand_x1_sg U59730 ( .A(reg_oi_11[5]), .B(n35020), .X(n20063) );
  nand_x1_sg U59731 ( .A(n32682), .B(\shifter_0/reg_i_11[5] ), .X(n20064) );
  nand_x1_sg U59732 ( .A(reg_oi_11[3]), .B(n31565), .X(n20059) );
  nand_x1_sg U59733 ( .A(n34742), .B(\shifter_0/reg_i_11[3] ), .X(n20060) );
  nand_x1_sg U59734 ( .A(reg_oi_11[1]), .B(n35017), .X(n20055) );
  nand_x1_sg U59735 ( .A(n32904), .B(\shifter_0/reg_i_11[1] ), .X(n20056) );
  nand_x1_sg U59736 ( .A(reg_oi_11[0]), .B(n33118), .X(n20053) );
  nand_x1_sg U59737 ( .A(n32646), .B(\shifter_0/reg_i_11[0] ), .X(n20054) );
  nand_x1_sg U59738 ( .A(reg_oi_5[7]), .B(n30563), .X(n19827) );
  nand_x1_sg U59739 ( .A(n32658), .B(\shifter_0/reg_i_5[7] ), .X(n19828) );
  nand_x1_sg U59740 ( .A(reg_oi_5[6]), .B(n33122), .X(n19825) );
  nand_x1_sg U59741 ( .A(n30854), .B(\shifter_0/reg_i_5[6] ), .X(n19826) );
  nand_x1_sg U59742 ( .A(reg_oi_5[5]), .B(n33118), .X(n19823) );
  nand_x1_sg U59743 ( .A(n34748), .B(\shifter_0/reg_i_5[5] ), .X(n19824) );
  nand_x1_sg U59744 ( .A(reg_oi_5[2]), .B(n29807), .X(n19817) );
  nand_x1_sg U59745 ( .A(n31487), .B(\shifter_0/reg_i_5[2] ), .X(n19818) );
  nand_x1_sg U59746 ( .A(reg_oi_5[1]), .B(n33062), .X(n19815) );
  nand_x1_sg U59747 ( .A(n34751), .B(\shifter_0/reg_i_5[1] ), .X(n19816) );
  nand_x1_sg U59748 ( .A(reg_oi_5[0]), .B(n33123), .X(n19813) );
  nand_x1_sg U59749 ( .A(n32637), .B(\shifter_0/reg_i_5[0] ), .X(n19814) );
  nand_x1_sg U59750 ( .A(reg_oi_8[4]), .B(n33082), .X(n19941) );
  nand_x1_sg U59751 ( .A(n29761), .B(\shifter_0/reg_i_8[4] ), .X(n19942) );
  nand_x1_sg U59752 ( .A(reg_oi_8[2]), .B(n33045), .X(n19937) );
  nand_x1_sg U59753 ( .A(n32696), .B(\shifter_0/reg_i_8[2] ), .X(n19938) );
  nand_x1_sg U59754 ( .A(reg_oi_8[7]), .B(n33821), .X(n19947) );
  nand_x1_sg U59755 ( .A(n32707), .B(\shifter_0/reg_i_8[7] ), .X(n19948) );
  nand_x1_sg U59756 ( .A(reg_oi_8[6]), .B(n33047), .X(n19945) );
  nand_x1_sg U59757 ( .A(n34728), .B(\shifter_0/reg_i_8[6] ), .X(n19946) );
  nand_x1_sg U59758 ( .A(reg_oi_8[5]), .B(n30605), .X(n19943) );
  nand_x1_sg U59759 ( .A(n32695), .B(\shifter_0/reg_i_8[5] ), .X(n19944) );
  nand_x1_sg U59760 ( .A(reg_oi_8[3]), .B(n35025), .X(n19939) );
  nand_x1_sg U59761 ( .A(n32705), .B(\shifter_0/reg_i_8[3] ), .X(n19940) );
  nand_x1_sg U59762 ( .A(reg_oi_8[1]), .B(n33113), .X(n19935) );
  nand_x1_sg U59763 ( .A(n32681), .B(\shifter_0/reg_i_8[1] ), .X(n19936) );
  nand_x1_sg U59764 ( .A(reg_oi_8[0]), .B(n33042), .X(n19933) );
  nand_x1_sg U59765 ( .A(n32653), .B(\shifter_0/reg_i_8[0] ), .X(n19934) );
  nand_x1_sg U59766 ( .A(reg_ow_13[9]), .B(n33819), .X(n20791) );
  nand_x1_sg U59767 ( .A(n34968), .B(\shifter_0/reg_w_13[9] ), .X(n20792) );
  nand_x1_sg U59768 ( .A(reg_ow_13[8]), .B(n33086), .X(n20789) );
  nand_x1_sg U59769 ( .A(n34413), .B(\shifter_0/reg_w_13[8] ), .X(n20790) );
  nand_x1_sg U59770 ( .A(reg_ow_13[4]), .B(n35015), .X(n20781) );
  nand_x1_sg U59771 ( .A(n32669), .B(\shifter_0/reg_w_13[4] ), .X(n20782) );
  nand_x1_sg U59772 ( .A(reg_ow_13[3]), .B(n33102), .X(n20779) );
  nand_x1_sg U59773 ( .A(n32527), .B(\shifter_0/reg_w_13[3] ), .X(n20780) );
  nand_x1_sg U59774 ( .A(reg_ow_11[8]), .B(n33117), .X(n20709) );
  nand_x1_sg U59775 ( .A(n34742), .B(\shifter_0/reg_w_11[8] ), .X(n20710) );
  nand_x1_sg U59776 ( .A(reg_ow_11[4]), .B(n31582), .X(n20701) );
  nand_x1_sg U59777 ( .A(n31232), .B(\shifter_0/reg_w_11[4] ), .X(n20702) );
  nand_x1_sg U59778 ( .A(reg_ow_11[3]), .B(n35022), .X(n20699) );
  nand_x1_sg U59779 ( .A(n34754), .B(\shifter_0/reg_w_11[3] ), .X(n20700) );
  nand_x1_sg U59780 ( .A(reg_ow_4[12]), .B(n31582), .X(n20437) );
  nand_x1_sg U59781 ( .A(n30045), .B(\shifter_0/reg_w_4[12] ), .X(n20438) );
  nand_x1_sg U59782 ( .A(reg_ow_4[11]), .B(n33822), .X(n20435) );
  nand_x1_sg U59783 ( .A(n32670), .B(\shifter_0/reg_w_4[11] ), .X(n20436) );
  nand_x1_sg U59784 ( .A(reg_ow_4[10]), .B(n33041), .X(n20433) );
  nand_x1_sg U59785 ( .A(n32683), .B(\shifter_0/reg_w_4[10] ), .X(n20434) );
  nand_x1_sg U59786 ( .A(reg_ow_4[9]), .B(n31567), .X(n20431) );
  nand_x1_sg U59787 ( .A(n31487), .B(\shifter_0/reg_w_4[9] ), .X(n20432) );
  nand_x1_sg U59788 ( .A(reg_ow_4[8]), .B(n33114), .X(n20429) );
  nand_x1_sg U59789 ( .A(n30702), .B(\shifter_0/reg_w_4[8] ), .X(n20430) );
  nand_x1_sg U59790 ( .A(reg_ow_4[7]), .B(n33098), .X(n20427) );
  nand_x1_sg U59791 ( .A(n32645), .B(\shifter_0/reg_w_4[7] ), .X(n20428) );
  nand_x1_sg U59792 ( .A(reg_ow_4[6]), .B(n29824), .X(n20425) );
  nand_x1_sg U59793 ( .A(n31232), .B(\shifter_0/reg_w_4[6] ), .X(n20426) );
  nand_x1_sg U59794 ( .A(reg_ow_4[5]), .B(n33105), .X(n20423) );
  nand_x1_sg U59795 ( .A(n30685), .B(\shifter_0/reg_w_4[5] ), .X(n20424) );
  nand_x1_sg U59796 ( .A(reg_ow_4[4]), .B(n33045), .X(n20421) );
  nand_x1_sg U59797 ( .A(n32685), .B(\shifter_0/reg_w_4[4] ), .X(n20422) );
  nand_x1_sg U59798 ( .A(reg_ow_1[13]), .B(n33087), .X(n20319) );
  nand_x1_sg U59799 ( .A(n30642), .B(\shifter_0/reg_w_1[13] ), .X(n20320) );
  nand_x1_sg U59800 ( .A(reg_ow_1[12]), .B(n35019), .X(n20317) );
  nand_x1_sg U59801 ( .A(n32677), .B(\shifter_0/reg_w_1[12] ), .X(n20318) );
  nand_x1_sg U59802 ( .A(reg_ow_1[9]), .B(n33052), .X(n20311) );
  nand_x1_sg U59803 ( .A(n32658), .B(\shifter_0/reg_w_1[9] ), .X(n20312) );
  nand_x1_sg U59804 ( .A(reg_ow_0[19]), .B(n29826), .X(n20291) );
  nand_x1_sg U59805 ( .A(n32694), .B(\shifter_0/reg_w_0[19] ), .X(n20292) );
  nand_x1_sg U59806 ( .A(reg_ow_0[18]), .B(n31571), .X(n20289) );
  nand_x1_sg U59807 ( .A(n30853), .B(\shifter_0/reg_w_0[18] ), .X(n20290) );
  nand_x1_sg U59808 ( .A(reg_ow_0[17]), .B(n33056), .X(n20287) );
  nand_x1_sg U59809 ( .A(n34741), .B(\shifter_0/reg_w_0[17] ), .X(n20288) );
  nand_x1_sg U59810 ( .A(reg_ow_0[16]), .B(n35041), .X(n20285) );
  nand_x1_sg U59811 ( .A(n30698), .B(\shifter_0/reg_w_0[16] ), .X(n20286) );
  nand_x1_sg U59812 ( .A(reg_oi_14[13]), .B(n33063), .X(n20199) );
  nand_x1_sg U59813 ( .A(n32645), .B(\shifter_0/reg_i_14[13] ), .X(n20200) );
  nand_x1_sg U59814 ( .A(reg_oi_14[12]), .B(n33053), .X(n20197) );
  nand_x1_sg U59815 ( .A(n31989), .B(\shifter_0/reg_i_14[12] ), .X(n20198) );
  nand_x1_sg U59816 ( .A(reg_oi_12[8]), .B(n30563), .X(n20109) );
  nand_x1_sg U59817 ( .A(n34729), .B(\shifter_0/reg_i_12[8] ), .X(n20110) );
  nand_x1_sg U59818 ( .A(reg_oi_5[8]), .B(n33041), .X(n19829) );
  nand_x1_sg U59819 ( .A(n34967), .B(\shifter_0/reg_i_5[8] ), .X(n19830) );
  nand_x1_sg U59820 ( .A(reg_oi_5[4]), .B(n33114), .X(n19821) );
  nand_x1_sg U59821 ( .A(n34804), .B(\shifter_0/reg_i_5[4] ), .X(n19822) );
  nand_x1_sg U59822 ( .A(reg_oi_5[3]), .B(n29813), .X(n19819) );
  nand_x1_sg U59823 ( .A(n31233), .B(\shifter_0/reg_i_5[3] ), .X(n19820) );
  nand_x1_sg U59824 ( .A(reg_oi_2[9]), .B(n29830), .X(n19711) );
  nand_x1_sg U59825 ( .A(n32702), .B(\shifter_0/reg_i_2[9] ), .X(n19712) );
  nand_x1_sg U59826 ( .A(reg_oi_1[18]), .B(n29801), .X(n19689) );
  nand_x1_sg U59827 ( .A(n31233), .B(\shifter_0/reg_i_1[18] ), .X(n19690) );
  nand_x1_sg U59828 ( .A(reg_oi_1[17]), .B(n35040), .X(n19687) );
  nand_x1_sg U59829 ( .A(n32658), .B(\shifter_0/reg_i_1[17] ), .X(n19688) );
  nand_x1_sg U59830 ( .A(reg_oi_1[13]), .B(n29822), .X(n19679) );
  nand_x1_sg U59831 ( .A(n32670), .B(\shifter_0/reg_i_1[13] ), .X(n19680) );
  nand_x1_sg U59832 ( .A(reg_oi_1[12]), .B(n33089), .X(n19677) );
  nand_x1_sg U59833 ( .A(n30043), .B(\shifter_0/reg_i_1[12] ), .X(n19678) );
  nand_x1_sg U59834 ( .A(reg_ow_7[11]), .B(n29824), .X(n20555) );
  nand_x1_sg U59835 ( .A(n32657), .B(\shifter_0/reg_w_7[11] ), .X(n20556) );
  nand_x1_sg U59836 ( .A(reg_ow_7[10]), .B(n31584), .X(n20553) );
  nand_x1_sg U59837 ( .A(n30680), .B(\shifter_0/reg_w_7[10] ), .X(n20554) );
  nand_x1_sg U59838 ( .A(reg_ow_7[9]), .B(n35015), .X(n20551) );
  nand_x1_sg U59839 ( .A(n34102), .B(\shifter_0/reg_w_7[9] ), .X(n20552) );
  nand_x1_sg U59840 ( .A(reg_ow_7[8]), .B(n33088), .X(n20549) );
  nand_x1_sg U59841 ( .A(n34803), .B(\shifter_0/reg_w_7[8] ), .X(n20550) );
  nand_x1_sg U59842 ( .A(reg_ow_7[7]), .B(n33111), .X(n20547) );
  nand_x1_sg U59843 ( .A(n34725), .B(\shifter_0/reg_w_7[7] ), .X(n20548) );
  nand_x1_sg U59844 ( .A(reg_ow_7[6]), .B(n31583), .X(n20545) );
  nand_x1_sg U59845 ( .A(n31235), .B(\shifter_0/reg_w_7[6] ), .X(n20546) );
  nand_x1_sg U59846 ( .A(reg_ow_7[5]), .B(n35044), .X(n20543) );
  nand_x1_sg U59847 ( .A(n32704), .B(\shifter_0/reg_w_7[5] ), .X(n20544) );
  nand_x1_sg U59848 ( .A(reg_ow_7[4]), .B(n33087), .X(n20541) );
  nand_x1_sg U59849 ( .A(n30044), .B(\shifter_0/reg_w_7[4] ), .X(n20542) );
  nand_x1_sg U59850 ( .A(reg_ow_7[3]), .B(n33116), .X(n20539) );
  nand_x1_sg U59851 ( .A(n32680), .B(\shifter_0/reg_w_7[3] ), .X(n20540) );
  nand_x1_sg U59852 ( .A(reg_oi_7[19]), .B(n35045), .X(n19931) );
  nand_x1_sg U59853 ( .A(n34111), .B(\shifter_0/reg_i_7[19] ), .X(n19932) );
  nand_x1_sg U59854 ( .A(filter_output_shifter_input_taken), .B(n32901), .X(
        n19610) );
  nand_x1_sg U59855 ( .A(n19594), .B(n31599), .X(n20895) );
  nand_x1_sg U59856 ( .A(n35266), .B(n20897), .X(n20896) );
  nand_x1_sg U59857 ( .A(n32517), .B(n32219), .X(n20897) );
  nor_x1_sg U59858 ( .A(n35258), .B(\filter_0/i_pointer[3] ), .X(n15045) );
  nor_x1_sg U59859 ( .A(n35256), .B(\filter_0/w_pointer[3] ), .X(n15178) );
  nor_x1_sg U59860 ( .A(\filter_0/i_pointer[0] ), .B(n35269), .X(n28834) );
  nand_x1_sg U59861 ( .A(\filter_0/w_pointer[2] ), .B(n32210), .X(n28973) );
  nand_x1_sg U59862 ( .A(n31123), .B(n32212), .X(n28975) );
  nand_x1_sg U59863 ( .A(n31118), .B(n32211), .X(n28275) );
  nand_x1_sg U59864 ( .A(n32886), .B(\filter_0/n8243 ), .X(n28968) );
  nand_x1_sg U59865 ( .A(n31657), .B(n28259), .X(n28969) );
  nor_x1_sg U59866 ( .A(\mask_0/state[0] ), .B(n42529), .X(n26575) );
  nand_x1_sg U59867 ( .A(n42526), .B(n34869), .X(n26349) );
  nand_x1_sg U59868 ( .A(o_mask[31]), .B(n30961), .X(n26348) );
  inv_x1_sg U59869 ( .A(n26351), .X(n42526) );
  nand_x1_sg U59870 ( .A(n42525), .B(n31250), .X(n26354) );
  nand_x1_sg U59871 ( .A(o_mask[30]), .B(n33856), .X(n26353) );
  inv_x1_sg U59872 ( .A(n26355), .X(n42525) );
  nand_x1_sg U59873 ( .A(n42524), .B(n34871), .X(n26357) );
  nand_x1_sg U59874 ( .A(o_mask[29]), .B(n30953), .X(n26356) );
  inv_x1_sg U59875 ( .A(n26358), .X(n42524) );
  nand_x1_sg U59876 ( .A(n42523), .B(n31044), .X(n26360) );
  nand_x1_sg U59877 ( .A(o_mask[28]), .B(n30956), .X(n26359) );
  inv_x1_sg U59878 ( .A(n26361), .X(n42523) );
  nand_x1_sg U59879 ( .A(n42522), .B(n31747), .X(n26363) );
  nand_x1_sg U59880 ( .A(o_mask[27]), .B(n34863), .X(n26362) );
  inv_x1_sg U59881 ( .A(n26364), .X(n42522) );
  nand_x1_sg U59882 ( .A(n42521), .B(n31046), .X(n26366) );
  nand_x1_sg U59883 ( .A(o_mask[26]), .B(n30960), .X(n26365) );
  inv_x1_sg U59884 ( .A(n26367), .X(n42521) );
  nand_x1_sg U59885 ( .A(n42520), .B(n31249), .X(n26369) );
  nand_x1_sg U59886 ( .A(o_mask[25]), .B(n34866), .X(n26368) );
  inv_x1_sg U59887 ( .A(n26370), .X(n42520) );
  nand_x1_sg U59888 ( .A(n42519), .B(n30633), .X(n26372) );
  nand_x1_sg U59889 ( .A(o_mask[24]), .B(n30201), .X(n26371) );
  inv_x1_sg U59890 ( .A(n26373), .X(n42519) );
  nand_x1_sg U59891 ( .A(n42518), .B(n31252), .X(n26375) );
  nand_x1_sg U59892 ( .A(o_mask[23]), .B(n34865), .X(n26374) );
  inv_x1_sg U59893 ( .A(n26376), .X(n42518) );
  nand_x1_sg U59894 ( .A(n42517), .B(n34870), .X(n26378) );
  nand_x1_sg U59895 ( .A(o_mask[22]), .B(n33857), .X(n26377) );
  inv_x1_sg U59896 ( .A(n26379), .X(n42517) );
  nand_x1_sg U59897 ( .A(n42516), .B(n31252), .X(n26381) );
  nand_x1_sg U59898 ( .A(o_mask[21]), .B(n34864), .X(n26380) );
  inv_x1_sg U59899 ( .A(n26382), .X(n42516) );
  nand_x1_sg U59900 ( .A(n42515), .B(n31622), .X(n26384) );
  nand_x1_sg U59901 ( .A(o_mask[20]), .B(n30953), .X(n26383) );
  inv_x1_sg U59902 ( .A(n26385), .X(n42515) );
  nand_x1_sg U59903 ( .A(n42514), .B(n34873), .X(n26387) );
  nand_x1_sg U59904 ( .A(o_mask[19]), .B(n34864), .X(n26386) );
  inv_x1_sg U59905 ( .A(n26388), .X(n42514) );
  nand_x1_sg U59906 ( .A(n42513), .B(n34869), .X(n26390) );
  nand_x1_sg U59907 ( .A(o_mask[18]), .B(n33843), .X(n26389) );
  inv_x1_sg U59908 ( .A(n26391), .X(n42513) );
  nand_x1_sg U59909 ( .A(n42512), .B(n31748), .X(n26393) );
  nand_x1_sg U59910 ( .A(o_mask[17]), .B(n30961), .X(n26392) );
  inv_x1_sg U59911 ( .A(n26394), .X(n42512) );
  nand_x1_sg U59912 ( .A(n42511), .B(n34874), .X(n26396) );
  nand_x1_sg U59913 ( .A(o_mask[16]), .B(n30957), .X(n26395) );
  inv_x1_sg U59914 ( .A(n26397), .X(n42511) );
  nand_x1_sg U59915 ( .A(n42510), .B(n31251), .X(n26399) );
  nand_x1_sg U59916 ( .A(o_mask[15]), .B(n33855), .X(n26398) );
  inv_x1_sg U59917 ( .A(n26400), .X(n42510) );
  nand_x1_sg U59918 ( .A(n42509), .B(n31044), .X(n26402) );
  nand_x1_sg U59919 ( .A(o_mask[14]), .B(n33850), .X(n26401) );
  inv_x1_sg U59920 ( .A(n26403), .X(n42509) );
  nand_x1_sg U59921 ( .A(n42508), .B(n34875), .X(n26405) );
  nand_x1_sg U59922 ( .A(o_mask[13]), .B(n33846), .X(n26404) );
  inv_x1_sg U59923 ( .A(n26406), .X(n42508) );
  nand_x1_sg U59924 ( .A(n42507), .B(n30632), .X(n26408) );
  nand_x1_sg U59925 ( .A(o_mask[12]), .B(n33842), .X(n26407) );
  inv_x1_sg U59926 ( .A(n26409), .X(n42507) );
  nand_x1_sg U59927 ( .A(n42506), .B(n34872), .X(n26411) );
  nand_x1_sg U59928 ( .A(o_mask[11]), .B(n30957), .X(n26410) );
  inv_x1_sg U59929 ( .A(n26412), .X(n42506) );
  nand_x1_sg U59930 ( .A(n42505), .B(n31250), .X(n26414) );
  nand_x1_sg U59931 ( .A(o_mask[10]), .B(n33853), .X(n26413) );
  inv_x1_sg U59932 ( .A(n26415), .X(n42505) );
  nand_x1_sg U59933 ( .A(n42504), .B(n31045), .X(n26417) );
  nand_x1_sg U59934 ( .A(o_mask[9]), .B(n30956), .X(n26416) );
  inv_x1_sg U59935 ( .A(n26418), .X(n42504) );
  nand_x1_sg U59936 ( .A(n42503), .B(n30632), .X(n26420) );
  nand_x1_sg U59937 ( .A(o_mask[8]), .B(n33845), .X(n26419) );
  inv_x1_sg U59938 ( .A(n26421), .X(n42503) );
  nand_x1_sg U59939 ( .A(n42502), .B(n31746), .X(n26423) );
  nand_x1_sg U59940 ( .A(o_mask[7]), .B(n33851), .X(n26422) );
  inv_x1_sg U59941 ( .A(n26424), .X(n42502) );
  nand_x1_sg U59942 ( .A(n42501), .B(n34872), .X(n26426) );
  nand_x1_sg U59943 ( .A(o_mask[6]), .B(n33848), .X(n26425) );
  inv_x1_sg U59944 ( .A(n26427), .X(n42501) );
  nand_x1_sg U59945 ( .A(n42500), .B(n34874), .X(n26429) );
  nand_x1_sg U59946 ( .A(o_mask[5]), .B(n33852), .X(n26428) );
  inv_x1_sg U59947 ( .A(n26430), .X(n42500) );
  nand_x1_sg U59948 ( .A(n42499), .B(n34876), .X(n26432) );
  nand_x1_sg U59949 ( .A(o_mask[4]), .B(n33858), .X(n26431) );
  inv_x1_sg U59950 ( .A(n26433), .X(n42499) );
  nand_x1_sg U59951 ( .A(n42498), .B(n34870), .X(n26435) );
  nand_x1_sg U59952 ( .A(o_mask[3]), .B(n30952), .X(n26434) );
  inv_x1_sg U59953 ( .A(n26436), .X(n42498) );
  nand_x1_sg U59954 ( .A(n42497), .B(n31249), .X(n26438) );
  nand_x1_sg U59955 ( .A(o_mask[2]), .B(n30952), .X(n26437) );
  inv_x1_sg U59956 ( .A(n26439), .X(n42497) );
  nand_x1_sg U59957 ( .A(n42496), .B(n34876), .X(n26441) );
  nand_x1_sg U59958 ( .A(o_mask[1]), .B(n33847), .X(n26440) );
  inv_x1_sg U59959 ( .A(n26442), .X(n42496) );
  nand_x1_sg U59960 ( .A(n42495), .B(n31621), .X(n26444) );
  nand_x1_sg U59961 ( .A(o_mask[0]), .B(n30960), .X(n26443) );
  inv_x1_sg U59962 ( .A(n26445), .X(n42495) );
  nand_x1_sg U59963 ( .A(n32887), .B(\filter_0/n8242 ), .X(n28970) );
  nand_x1_sg U59964 ( .A(n31879), .B(n32210), .X(n28971) );
  nand_x1_sg U59965 ( .A(n34869), .B(\mask_0/reg_w_mask[31] ), .X(n26446) );
  nand_x1_sg U59966 ( .A(\mask_0/reg_ww_mask[31] ), .B(n30956), .X(n26447) );
  nand_x1_sg U59967 ( .A(n31252), .B(\mask_0/reg_w_mask[30] ), .X(n26448) );
  nand_x1_sg U59968 ( .A(\mask_0/reg_ww_mask[30] ), .B(n33845), .X(n26449) );
  nand_x1_sg U59969 ( .A(n31249), .B(\mask_0/reg_w_mask[29] ), .X(n26450) );
  nand_x1_sg U59970 ( .A(\mask_0/reg_ww_mask[29] ), .B(n33853), .X(n26451) );
  nand_x1_sg U59971 ( .A(n34871), .B(\mask_0/reg_w_mask[28] ), .X(n26452) );
  nand_x1_sg U59972 ( .A(\mask_0/reg_ww_mask[28] ), .B(n34866), .X(n26453) );
  nand_x1_sg U59973 ( .A(n31749), .B(\mask_0/reg_w_mask[27] ), .X(n26454) );
  nand_x1_sg U59974 ( .A(\mask_0/reg_ww_mask[27] ), .B(n33858), .X(n26455) );
  nand_x1_sg U59975 ( .A(n31746), .B(\mask_0/reg_w_mask[26] ), .X(n26456) );
  nand_x1_sg U59976 ( .A(\mask_0/reg_ww_mask[26] ), .B(n33848), .X(n26457) );
  nand_x1_sg U59977 ( .A(n31746), .B(\mask_0/reg_w_mask[25] ), .X(n26458) );
  nand_x1_sg U59978 ( .A(\mask_0/reg_ww_mask[25] ), .B(n33847), .X(n26459) );
  nand_x1_sg U59979 ( .A(n31749), .B(\mask_0/reg_w_mask[24] ), .X(n26460) );
  nand_x1_sg U59980 ( .A(\mask_0/reg_ww_mask[24] ), .B(n33856), .X(n26461) );
  nand_x1_sg U59981 ( .A(n34870), .B(\mask_0/reg_w_mask[23] ), .X(n26462) );
  nand_x1_sg U59982 ( .A(\mask_0/reg_ww_mask[23] ), .B(n30957), .X(n26463) );
  nand_x1_sg U59983 ( .A(n31748), .B(\mask_0/reg_w_mask[22] ), .X(n26464) );
  nand_x1_sg U59984 ( .A(\mask_0/reg_ww_mask[22] ), .B(n33852), .X(n26465) );
  nand_x1_sg U59985 ( .A(n34870), .B(\mask_0/reg_w_mask[21] ), .X(n26466) );
  nand_x1_sg U59986 ( .A(\mask_0/reg_ww_mask[21] ), .B(n30957), .X(n26467) );
  nand_x1_sg U59987 ( .A(n31749), .B(\mask_0/reg_w_mask[20] ), .X(n26468) );
  nand_x1_sg U59988 ( .A(\mask_0/reg_ww_mask[20] ), .B(n33847), .X(n26469) );
  nand_x1_sg U59989 ( .A(n31749), .B(\mask_0/reg_w_mask[19] ), .X(n26470) );
  nand_x1_sg U59990 ( .A(\mask_0/reg_ww_mask[19] ), .B(n34863), .X(n26471) );
  nand_x1_sg U59991 ( .A(n34875), .B(\mask_0/reg_w_mask[18] ), .X(n26472) );
  nand_x1_sg U59992 ( .A(\mask_0/reg_ww_mask[18] ), .B(n33853), .X(n26473) );
  nand_x1_sg U59993 ( .A(n34873), .B(\mask_0/reg_w_mask[17] ), .X(n26474) );
  nand_x1_sg U59994 ( .A(\mask_0/reg_ww_mask[17] ), .B(n33845), .X(n26475) );
  nand_x1_sg U59995 ( .A(n34874), .B(\mask_0/reg_w_mask[16] ), .X(n26476) );
  nand_x1_sg U59996 ( .A(\mask_0/reg_ww_mask[16] ), .B(n30201), .X(n26477) );
  nand_x1_sg U59997 ( .A(n30203), .B(\mask_0/reg_w_mask[15] ), .X(n26478) );
  nand_x1_sg U59998 ( .A(\mask_0/reg_ww_mask[15] ), .B(n30952), .X(n26479) );
  nand_x1_sg U59999 ( .A(n34871), .B(\mask_0/reg_w_mask[14] ), .X(n26480) );
  nand_x1_sg U60000 ( .A(\mask_0/reg_ww_mask[14] ), .B(n34864), .X(n26481) );
  nand_x1_sg U60001 ( .A(n34872), .B(\mask_0/reg_w_mask[13] ), .X(n26482) );
  nand_x1_sg U60002 ( .A(\mask_0/reg_ww_mask[13] ), .B(n30960), .X(n26483) );
  nand_x1_sg U60003 ( .A(n31045), .B(\mask_0/reg_w_mask[12] ), .X(n26484) );
  nand_x1_sg U60004 ( .A(\mask_0/reg_ww_mask[12] ), .B(n33858), .X(n26485) );
  nand_x1_sg U60005 ( .A(n34873), .B(\mask_0/reg_w_mask[11] ), .X(n26486) );
  nand_x1_sg U60006 ( .A(\mask_0/reg_ww_mask[11] ), .B(n30960), .X(n26487) );
  nand_x1_sg U60007 ( .A(n31046), .B(\mask_0/reg_w_mask[10] ), .X(n26488) );
  nand_x1_sg U60008 ( .A(\mask_0/reg_ww_mask[10] ), .B(n33850), .X(n26489) );
  nand_x1_sg U60009 ( .A(n34872), .B(\mask_0/reg_w_mask[9] ), .X(n26490) );
  nand_x1_sg U60010 ( .A(\mask_0/reg_ww_mask[9] ), .B(n30201), .X(n26491) );
  nand_x1_sg U60011 ( .A(n30203), .B(\mask_0/reg_w_mask[8] ), .X(n26492) );
  nand_x1_sg U60012 ( .A(\mask_0/reg_ww_mask[8] ), .B(n33853), .X(n26493) );
  nand_x1_sg U60013 ( .A(n30632), .B(\mask_0/reg_w_mask[7] ), .X(n26494) );
  nand_x1_sg U60014 ( .A(\mask_0/reg_ww_mask[7] ), .B(n33847), .X(n26495) );
  nand_x1_sg U60015 ( .A(n31621), .B(\mask_0/reg_w_mask[6] ), .X(n26496) );
  nand_x1_sg U60016 ( .A(\mask_0/reg_ww_mask[6] ), .B(n33846), .X(n26497) );
  nand_x1_sg U60017 ( .A(n34873), .B(\mask_0/reg_w_mask[5] ), .X(n26498) );
  nand_x1_sg U60018 ( .A(\mask_0/reg_ww_mask[5] ), .B(n33842), .X(n26499) );
  nand_x1_sg U60019 ( .A(n31250), .B(\mask_0/reg_w_mask[4] ), .X(n26500) );
  nand_x1_sg U60020 ( .A(\mask_0/reg_ww_mask[4] ), .B(n30953), .X(n26501) );
  nand_x1_sg U60021 ( .A(n34875), .B(\mask_0/reg_w_mask[3] ), .X(n26502) );
  nand_x1_sg U60022 ( .A(\mask_0/reg_ww_mask[3] ), .B(n30961), .X(n26503) );
  nand_x1_sg U60023 ( .A(n30633), .B(\mask_0/reg_w_mask[2] ), .X(n26504) );
  nand_x1_sg U60024 ( .A(\mask_0/reg_ww_mask[2] ), .B(n33855), .X(n26505) );
  nand_x1_sg U60025 ( .A(n31046), .B(\mask_0/reg_w_mask[1] ), .X(n26506) );
  nand_x1_sg U60026 ( .A(\mask_0/reg_ww_mask[1] ), .B(n34866), .X(n26507) );
  nand_x1_sg U60027 ( .A(n31621), .B(\mask_0/reg_w_mask[0] ), .X(n26508) );
  nand_x1_sg U60028 ( .A(\mask_0/reg_ww_mask[0] ), .B(n34865), .X(n26509) );
  nand_x1_sg U60029 ( .A(n31044), .B(\mask_0/reg_i_mask[31] ), .X(n26510) );
  nand_x1_sg U60030 ( .A(\mask_0/reg_ii_mask[31] ), .B(n30953), .X(n26511) );
  nand_x1_sg U60031 ( .A(n31621), .B(\mask_0/reg_i_mask[30] ), .X(n26512) );
  nand_x1_sg U60032 ( .A(\mask_0/reg_ii_mask[30] ), .B(n33858), .X(n26513) );
  nand_x1_sg U60033 ( .A(n30203), .B(\mask_0/reg_i_mask[29] ), .X(n26514) );
  nand_x1_sg U60034 ( .A(\mask_0/reg_ii_mask[29] ), .B(n33855), .X(n26515) );
  nand_x1_sg U60035 ( .A(n31252), .B(\mask_0/reg_i_mask[28] ), .X(n26516) );
  nand_x1_sg U60036 ( .A(\mask_0/reg_ii_mask[28] ), .B(n33852), .X(n26517) );
  nand_x1_sg U60037 ( .A(n31622), .B(\mask_0/reg_i_mask[27] ), .X(n26518) );
  nand_x1_sg U60038 ( .A(\mask_0/reg_ii_mask[27] ), .B(n33850), .X(n26519) );
  nand_x1_sg U60039 ( .A(n30203), .B(\mask_0/reg_i_mask[26] ), .X(n26520) );
  nand_x1_sg U60040 ( .A(\mask_0/reg_ii_mask[26] ), .B(n30956), .X(n26521) );
  nand_x1_sg U60041 ( .A(n34869), .B(\mask_0/reg_i_mask[25] ), .X(n26522) );
  nand_x1_sg U60042 ( .A(\mask_0/reg_ii_mask[25] ), .B(n33851), .X(n26523) );
  nand_x1_sg U60043 ( .A(n31046), .B(\mask_0/reg_i_mask[24] ), .X(n26524) );
  nand_x1_sg U60044 ( .A(\mask_0/reg_ii_mask[24] ), .B(n33852), .X(n26525) );
  nand_x1_sg U60045 ( .A(n31622), .B(\mask_0/reg_i_mask[23] ), .X(n26526) );
  nand_x1_sg U60046 ( .A(\mask_0/reg_ii_mask[23] ), .B(n33848), .X(n26527) );
  nand_x1_sg U60047 ( .A(n31622), .B(\mask_0/reg_i_mask[22] ), .X(n26528) );
  nand_x1_sg U60048 ( .A(\mask_0/reg_ii_mask[22] ), .B(n33857), .X(n26529) );
  nand_x1_sg U60049 ( .A(n31045), .B(\mask_0/reg_i_mask[21] ), .X(n26530) );
  nand_x1_sg U60050 ( .A(\mask_0/reg_ii_mask[21] ), .B(n34865), .X(n26531) );
  nand_x1_sg U60051 ( .A(n31251), .B(\mask_0/reg_i_mask[20] ), .X(n26532) );
  nand_x1_sg U60052 ( .A(\mask_0/reg_ii_mask[20] ), .B(n33855), .X(n26533) );
  nand_x1_sg U60053 ( .A(n30633), .B(\mask_0/reg_i_mask[19] ), .X(n26534) );
  nand_x1_sg U60054 ( .A(\mask_0/reg_ii_mask[19] ), .B(n30961), .X(n26535) );
  nand_x1_sg U60055 ( .A(n34871), .B(\mask_0/reg_i_mask[18] ), .X(n26536) );
  nand_x1_sg U60056 ( .A(\mask_0/reg_ii_mask[18] ), .B(n33846), .X(n26537) );
  nand_x1_sg U60057 ( .A(n31747), .B(\mask_0/reg_i_mask[17] ), .X(n26538) );
  nand_x1_sg U60058 ( .A(\mask_0/reg_ii_mask[17] ), .B(n33848), .X(n26539) );
  nand_x1_sg U60059 ( .A(n31747), .B(\mask_0/reg_i_mask[16] ), .X(n26540) );
  nand_x1_sg U60060 ( .A(\mask_0/reg_ii_mask[16] ), .B(n33843), .X(n26541) );
  nand_x1_sg U60061 ( .A(n31251), .B(\mask_0/reg_i_mask[15] ), .X(n26542) );
  nand_x1_sg U60062 ( .A(\mask_0/reg_ii_mask[15] ), .B(n33842), .X(n26543) );
  nand_x1_sg U60063 ( .A(n31747), .B(\mask_0/reg_i_mask[14] ), .X(n26544) );
  nand_x1_sg U60064 ( .A(\mask_0/reg_ii_mask[14] ), .B(n33843), .X(n26545) );
  nand_x1_sg U60065 ( .A(n34876), .B(\mask_0/reg_i_mask[13] ), .X(n26546) );
  nand_x1_sg U60066 ( .A(\mask_0/reg_ii_mask[13] ), .B(n33851), .X(n26547) );
  nand_x1_sg U60067 ( .A(n31748), .B(\mask_0/reg_i_mask[12] ), .X(n26548) );
  nand_x1_sg U60068 ( .A(\mask_0/reg_ii_mask[12] ), .B(n33856), .X(n26549) );
  nand_x1_sg U60069 ( .A(n31746), .B(\mask_0/reg_i_mask[11] ), .X(n26550) );
  nand_x1_sg U60070 ( .A(\mask_0/reg_ii_mask[11] ), .B(n33846), .X(n26551) );
  nand_x1_sg U60071 ( .A(n30633), .B(\mask_0/reg_i_mask[10] ), .X(n26552) );
  nand_x1_sg U60072 ( .A(\mask_0/reg_ii_mask[10] ), .B(n34864), .X(n26553) );
  nand_x1_sg U60073 ( .A(n31251), .B(\mask_0/reg_i_mask[9] ), .X(n26554) );
  nand_x1_sg U60074 ( .A(\mask_0/reg_ii_mask[9] ), .B(n34863), .X(n26555) );
  nand_x1_sg U60075 ( .A(n34876), .B(\mask_0/reg_i_mask[8] ), .X(n26556) );
  nand_x1_sg U60076 ( .A(\mask_0/reg_ii_mask[8] ), .B(n33857), .X(n26557) );
  nand_x1_sg U60077 ( .A(n31044), .B(\mask_0/reg_i_mask[7] ), .X(n26558) );
  nand_x1_sg U60078 ( .A(\mask_0/reg_ii_mask[7] ), .B(n33850), .X(n26559) );
  nand_x1_sg U60079 ( .A(n31748), .B(\mask_0/reg_i_mask[6] ), .X(n26560) );
  nand_x1_sg U60080 ( .A(\mask_0/reg_ii_mask[6] ), .B(n33843), .X(n26561) );
  nand_x1_sg U60081 ( .A(n34874), .B(\mask_0/reg_i_mask[5] ), .X(n26562) );
  nand_x1_sg U60082 ( .A(\mask_0/reg_ii_mask[5] ), .B(n33842), .X(n26563) );
  nand_x1_sg U60083 ( .A(n31249), .B(\mask_0/reg_i_mask[4] ), .X(n26564) );
  nand_x1_sg U60084 ( .A(\mask_0/reg_ii_mask[4] ), .B(n30952), .X(n26565) );
  nand_x1_sg U60085 ( .A(n31250), .B(\mask_0/reg_i_mask[3] ), .X(n26566) );
  nand_x1_sg U60086 ( .A(\mask_0/reg_ii_mask[3] ), .B(n33856), .X(n26567) );
  nand_x1_sg U60087 ( .A(n34875), .B(\mask_0/reg_i_mask[2] ), .X(n26568) );
  nand_x1_sg U60088 ( .A(\mask_0/reg_ii_mask[2] ), .B(n33845), .X(n26569) );
  nand_x1_sg U60089 ( .A(n30632), .B(\mask_0/reg_i_mask[1] ), .X(n26570) );
  nand_x1_sg U60090 ( .A(\mask_0/reg_ii_mask[1] ), .B(n33857), .X(n26571) );
  nand_x1_sg U60091 ( .A(n31045), .B(\mask_0/reg_i_mask[0] ), .X(n26572) );
  nand_x1_sg U60092 ( .A(\mask_0/reg_ii_mask[0] ), .B(n33851), .X(n26573) );
  nand_x1_sg U60093 ( .A(n32885), .B(\filter_0/n7917 ), .X(n28260) );
  nand_x1_sg U60094 ( .A(n30389), .B(n32211), .X(n28261) );
  nand_x1_sg U60095 ( .A(n32886), .B(\filter_0/n7914 ), .X(n28268) );
  nand_x1_sg U60096 ( .A(n31121), .B(n32212), .X(n28269) );
  nand_x1_sg U60097 ( .A(n32885), .B(\filter_0/n7912 ), .X(n28272) );
  nand_x1_sg U60098 ( .A(\filter_0/i_pointer[2] ), .B(n32212), .X(n28273) );
  nand_x1_sg U60099 ( .A(n32885), .B(\filter_0/n7916 ), .X(n28262) );
  nand_x1_sg U60100 ( .A(n31594), .B(n32212), .X(n28263) );
  nand_x1_sg U60101 ( .A(n32887), .B(\filter_0/n7913 ), .X(n28270) );
  nand_x1_sg U60102 ( .A(n31593), .B(n32210), .X(n28271) );
  nand_x1_sg U60103 ( .A(n32884), .B(\filter_0/n7919 ), .X(n28266) );
  nand_x1_sg U60104 ( .A(n31875), .B(n32211), .X(n28267) );
  nand_x1_sg U60105 ( .A(n32884), .B(\filter_0/n7918 ), .X(n28257) );
  nand_x1_sg U60106 ( .A(n31656), .B(n32211), .X(n28258) );
  nand_x1_sg U60107 ( .A(n32886), .B(\filter_0/n7915 ), .X(n28264) );
  nand_x1_sg U60108 ( .A(n32001), .B(n32210), .X(n28265) );
  nor_x1_sg U60109 ( .A(\filter_0/i_pointer[2] ), .B(n31118), .X(n28965) );
  nor_x1_sg U60110 ( .A(\filter_0/w_pointer[2] ), .B(n31123), .X(n29664) );
  nor_x1_sg U60111 ( .A(\filter_0/i_pointer[1] ), .B(n35257), .X(n28878) );
  nor_x1_sg U60112 ( .A(\shifter_0/reg_w_7[8] ), .B(\shifter_0/reg_w_7[9] ), 
        .X(n21138) );
  nor_x1_sg U60113 ( .A(\shifter_0/reg_w_7[6] ), .B(\shifter_0/reg_w_7[5] ), 
        .X(n21136) );
  nor_x1_sg U60114 ( .A(\shifter_0/reg_w_7[7] ), .B(n42715), .X(n21137) );
  nor_x1_sg U60115 ( .A(n31878), .B(n31657), .X(n29666) );
  nor_x1_sg U60116 ( .A(\shifter_0/reg_w_7[3] ), .B(\shifter_0/reg_w_7[4] ), 
        .X(n21135) );
  nor_x1_sg U60117 ( .A(\shifter_0/reg_w_7[17] ), .B(\shifter_0/reg_w_7[18] ), 
        .X(n21146) );
  nor_x1_sg U60118 ( .A(\shifter_0/reg_w_7[11] ), .B(n42716), .X(n21142) );
  nor_x1_sg U60119 ( .A(\shifter_0/reg_w_7[12] ), .B(\shifter_0/reg_w_7[13] ), 
        .X(n21143) );
  nor_x1_sg U60120 ( .A(\shifter_0/reg_w_7[1] ), .B(\shifter_0/reg_w_7[19] ), 
        .X(n21133) );
  nor_x1_sg U60121 ( .A(\shifter_0/reg_w_7[2] ), .B(n42714), .X(n21134) );
  nor_x1_sg U60122 ( .A(\shifter_0/reg_w_7[15] ), .B(\shifter_0/reg_w_7[14] ), 
        .X(n21144) );
  nor_x1_sg U60123 ( .A(\shifter_0/reg_w_7[16] ), .B(n42717), .X(n21145) );
  nor_x1_sg U60124 ( .A(n42412), .B(n31885), .X(n26578) );
  nor_x1_sg U60125 ( .A(n26583), .B(n26586), .X(n26585) );
  nor_x1_sg U60126 ( .A(filter_state[1]), .B(n42413), .X(n26586) );
  nand_x1_sg U60127 ( .A(n26578), .B(filter_state[0]), .X(n26580) );
  nand_x1_sg U60128 ( .A(n26582), .B(n32426), .X(n26581) );
  nor_x1_sg U60129 ( .A(n26578), .B(n26583), .X(n26582) );
  nor_x1_sg U60130 ( .A(\shifter_0/reg_i_7[8] ), .B(\shifter_0/reg_i_7[9] ), 
        .X(n21534) );
  nor_x1_sg U60131 ( .A(\shifter_0/reg_i_7[12] ), .B(\shifter_0/reg_i_7[13] ), 
        .X(n21539) );
  inv_x1_sg U60132 ( .A(\mask_0/state[1] ), .X(n42529) );
  nor_x1_sg U60133 ( .A(\shifter_0/reg_i_7[6] ), .B(\shifter_0/reg_i_7[5] ), 
        .X(n21532) );
  nor_x1_sg U60134 ( .A(\shifter_0/reg_i_7[7] ), .B(n42605), .X(n21533) );
  nor_x1_sg U60135 ( .A(\shifter_0/reg_i_7[10] ), .B(\shifter_0/reg_i_7[0] ), 
        .X(n21537) );
  nor_x1_sg U60136 ( .A(\shifter_0/reg_i_7[11] ), .B(n42606), .X(n21538) );
  nand_x1_sg U60137 ( .A(n35682), .B(reg_w_mask[31]), .X(n26345) );
  nand_x1_sg U60138 ( .A(\mask_0/reg_w_mask[31] ), .B(n34797), .X(n26346) );
  nand_x1_sg U60139 ( .A(n34391), .B(reg_w_mask[30]), .X(n26343) );
  nand_x1_sg U60140 ( .A(\mask_0/reg_w_mask[30] ), .B(n30644), .X(n26344) );
  nand_x1_sg U60141 ( .A(n34399), .B(reg_w_mask[29]), .X(n26341) );
  nand_x1_sg U60142 ( .A(\mask_0/reg_w_mask[29] ), .B(n32533), .X(n26342) );
  nand_x1_sg U60143 ( .A(n34400), .B(reg_w_mask[28]), .X(n26339) );
  nand_x1_sg U60144 ( .A(\mask_0/reg_w_mask[28] ), .B(n32533), .X(n26340) );
  nand_x1_sg U60145 ( .A(n34393), .B(reg_w_mask[27]), .X(n26337) );
  nand_x1_sg U60146 ( .A(\mask_0/reg_w_mask[27] ), .B(n32528), .X(n26338) );
  nand_x1_sg U60147 ( .A(n34399), .B(reg_w_mask[26]), .X(n26335) );
  nand_x1_sg U60148 ( .A(\mask_0/reg_w_mask[26] ), .B(n32534), .X(n26336) );
  nand_x1_sg U60149 ( .A(n34394), .B(reg_w_mask[25]), .X(n26333) );
  nand_x1_sg U60150 ( .A(\mask_0/reg_w_mask[25] ), .B(n32529), .X(n26334) );
  nand_x1_sg U60151 ( .A(n34399), .B(reg_w_mask[24]), .X(n26331) );
  nand_x1_sg U60152 ( .A(\mask_0/reg_w_mask[24] ), .B(n30645), .X(n26332) );
  nand_x1_sg U60153 ( .A(n34392), .B(reg_w_mask[23]), .X(n26329) );
  nand_x1_sg U60154 ( .A(\mask_0/reg_w_mask[23] ), .B(n34798), .X(n26330) );
  nand_x1_sg U60155 ( .A(n34394), .B(reg_w_mask[22]), .X(n26327) );
  nand_x1_sg U60156 ( .A(\mask_0/reg_w_mask[22] ), .B(n32534), .X(n26328) );
  nand_x1_sg U60157 ( .A(n33887), .B(reg_w_mask[21]), .X(n26325) );
  nand_x1_sg U60158 ( .A(\mask_0/reg_w_mask[21] ), .B(n32536), .X(n26326) );
  nand_x1_sg U60159 ( .A(n33885), .B(reg_w_mask[20]), .X(n26323) );
  nand_x1_sg U60160 ( .A(\mask_0/reg_w_mask[20] ), .B(n32537), .X(n26324) );
  nand_x1_sg U60161 ( .A(n33887), .B(reg_w_mask[19]), .X(n26321) );
  nand_x1_sg U60162 ( .A(\mask_0/reg_w_mask[19] ), .B(n32531), .X(n26322) );
  nand_x1_sg U60163 ( .A(n33888), .B(reg_w_mask[18]), .X(n26319) );
  nand_x1_sg U60164 ( .A(\mask_0/reg_w_mask[18] ), .B(n32534), .X(n26320) );
  nand_x1_sg U60165 ( .A(n33884), .B(reg_w_mask[17]), .X(n26317) );
  nand_x1_sg U60166 ( .A(\mask_0/reg_w_mask[17] ), .B(n34797), .X(n26318) );
  nand_x1_sg U60167 ( .A(n33885), .B(reg_w_mask[16]), .X(n26315) );
  nand_x1_sg U60168 ( .A(\mask_0/reg_w_mask[16] ), .B(n32538), .X(n26316) );
  nand_x1_sg U60169 ( .A(n34398), .B(reg_w_mask[15]), .X(n26313) );
  nand_x1_sg U60170 ( .A(\mask_0/reg_w_mask[15] ), .B(n30188), .X(n26314) );
  nand_x1_sg U60171 ( .A(n34401), .B(reg_w_mask[14]), .X(n26311) );
  nand_x1_sg U60172 ( .A(\mask_0/reg_w_mask[14] ), .B(n32532), .X(n26312) );
  nand_x1_sg U60173 ( .A(n33882), .B(reg_w_mask[13]), .X(n26309) );
  nand_x1_sg U60174 ( .A(\mask_0/reg_w_mask[13] ), .B(n34799), .X(n26310) );
  nand_x1_sg U60175 ( .A(n33882), .B(reg_w_mask[12]), .X(n26307) );
  nand_x1_sg U60176 ( .A(\mask_0/reg_w_mask[12] ), .B(n34796), .X(n26308) );
  nand_x1_sg U60177 ( .A(n33888), .B(reg_w_mask[11]), .X(n26305) );
  nand_x1_sg U60178 ( .A(\mask_0/reg_w_mask[11] ), .B(n32531), .X(n26306) );
  nand_x1_sg U60179 ( .A(n33882), .B(reg_w_mask[10]), .X(n26303) );
  nand_x1_sg U60180 ( .A(\mask_0/reg_w_mask[10] ), .B(n32533), .X(n26304) );
  nand_x1_sg U60181 ( .A(n34396), .B(reg_w_mask[9]), .X(n26301) );
  nand_x1_sg U60182 ( .A(\mask_0/reg_w_mask[9] ), .B(n32532), .X(n26302) );
  nand_x1_sg U60183 ( .A(n34392), .B(reg_w_mask[8]), .X(n26299) );
  nand_x1_sg U60184 ( .A(\mask_0/reg_w_mask[8] ), .B(n32534), .X(n26300) );
  nand_x1_sg U60185 ( .A(n34400), .B(reg_w_mask[7]), .X(n26297) );
  nand_x1_sg U60186 ( .A(\mask_0/reg_w_mask[7] ), .B(n34799), .X(n26298) );
  nand_x1_sg U60187 ( .A(n34396), .B(reg_w_mask[6]), .X(n26295) );
  nand_x1_sg U60188 ( .A(\mask_0/reg_w_mask[6] ), .B(n32538), .X(n26296) );
  nand_x1_sg U60189 ( .A(n34392), .B(reg_w_mask[5]), .X(n26293) );
  nand_x1_sg U60190 ( .A(\mask_0/reg_w_mask[5] ), .B(n34798), .X(n26294) );
  nand_x1_sg U60191 ( .A(n35682), .B(reg_w_mask[4]), .X(n26291) );
  nand_x1_sg U60192 ( .A(\mask_0/reg_w_mask[4] ), .B(n32539), .X(n26292) );
  nand_x1_sg U60193 ( .A(n34396), .B(reg_w_mask[3]), .X(n26289) );
  nand_x1_sg U60194 ( .A(\mask_0/reg_w_mask[3] ), .B(n34799), .X(n26290) );
  nand_x1_sg U60195 ( .A(n33881), .B(reg_w_mask[2]), .X(n26287) );
  nand_x1_sg U60196 ( .A(\mask_0/reg_w_mask[2] ), .B(n30188), .X(n26288) );
  nand_x1_sg U60197 ( .A(n33881), .B(reg_w_mask[1]), .X(n26285) );
  nand_x1_sg U60198 ( .A(\mask_0/reg_w_mask[1] ), .B(n32532), .X(n26286) );
  nand_x1_sg U60199 ( .A(n34397), .B(reg_w_mask[0]), .X(n26283) );
  nand_x1_sg U60200 ( .A(\mask_0/reg_w_mask[0] ), .B(n32536), .X(n26284) );
  nand_x1_sg U60201 ( .A(n34394), .B(reg_i_mask[31]), .X(n26281) );
  nand_x1_sg U60202 ( .A(\mask_0/reg_i_mask[31] ), .B(n30644), .X(n26282) );
  nand_x1_sg U60203 ( .A(n33879), .B(reg_i_mask[30]), .X(n26279) );
  nand_x1_sg U60204 ( .A(\mask_0/reg_i_mask[30] ), .B(n32537), .X(n26280) );
  nand_x1_sg U60205 ( .A(n35682), .B(reg_i_mask[29]), .X(n26277) );
  nand_x1_sg U60206 ( .A(\mask_0/reg_i_mask[29] ), .B(n32529), .X(n26278) );
  nand_x1_sg U60207 ( .A(n34394), .B(reg_i_mask[28]), .X(n26275) );
  nand_x1_sg U60208 ( .A(\mask_0/reg_i_mask[28] ), .B(n32539), .X(n26276) );
  nand_x1_sg U60209 ( .A(n34397), .B(reg_i_mask[27]), .X(n26273) );
  nand_x1_sg U60210 ( .A(\mask_0/reg_i_mask[27] ), .B(n32537), .X(n26274) );
  nand_x1_sg U60211 ( .A(n34392), .B(reg_i_mask[26]), .X(n26271) );
  nand_x1_sg U60212 ( .A(\mask_0/reg_i_mask[26] ), .B(n30645), .X(n26272) );
  nand_x1_sg U60213 ( .A(n34393), .B(reg_i_mask[25]), .X(n26269) );
  nand_x1_sg U60214 ( .A(\mask_0/reg_i_mask[25] ), .B(n32538), .X(n26270) );
  nand_x1_sg U60215 ( .A(n34391), .B(reg_i_mask[24]), .X(n26267) );
  nand_x1_sg U60216 ( .A(\mask_0/reg_i_mask[24] ), .B(n32531), .X(n26268) );
  nand_x1_sg U60217 ( .A(n34391), .B(reg_i_mask[23]), .X(n26265) );
  nand_x1_sg U60218 ( .A(\mask_0/reg_i_mask[23] ), .B(n32533), .X(n26266) );
  nand_x1_sg U60219 ( .A(n35682), .B(reg_i_mask[22]), .X(n26263) );
  nand_x1_sg U60220 ( .A(\mask_0/reg_i_mask[22] ), .B(n34798), .X(n26264) );
  nand_x1_sg U60221 ( .A(n34401), .B(reg_i_mask[21]), .X(n26261) );
  nand_x1_sg U60222 ( .A(\mask_0/reg_i_mask[21] ), .B(n34796), .X(n26262) );
  nand_x1_sg U60223 ( .A(n34398), .B(reg_i_mask[20]), .X(n26259) );
  nand_x1_sg U60224 ( .A(\mask_0/reg_i_mask[20] ), .B(n30645), .X(n26260) );
  nand_x1_sg U60225 ( .A(n34398), .B(reg_i_mask[19]), .X(n26257) );
  nand_x1_sg U60226 ( .A(\mask_0/reg_i_mask[19] ), .B(n32539), .X(n26258) );
  nand_x1_sg U60227 ( .A(n34398), .B(reg_i_mask[18]), .X(n26255) );
  nand_x1_sg U60228 ( .A(\mask_0/reg_i_mask[18] ), .B(n30644), .X(n26256) );
  nand_x1_sg U60229 ( .A(n34397), .B(reg_i_mask[17]), .X(n26253) );
  nand_x1_sg U60230 ( .A(\mask_0/reg_i_mask[17] ), .B(n32531), .X(n26254) );
  nand_x1_sg U60231 ( .A(n33881), .B(reg_i_mask[16]), .X(n26251) );
  nand_x1_sg U60232 ( .A(\mask_0/reg_i_mask[16] ), .B(n32536), .X(n26252) );
  nand_x1_sg U60233 ( .A(n34399), .B(reg_i_mask[15]), .X(n26249) );
  nand_x1_sg U60234 ( .A(\mask_0/reg_i_mask[15] ), .B(n34799), .X(n26250) );
  nand_x1_sg U60235 ( .A(n34393), .B(reg_i_mask[14]), .X(n26247) );
  nand_x1_sg U60236 ( .A(\mask_0/reg_i_mask[14] ), .B(n32528), .X(n26248) );
  nand_x1_sg U60237 ( .A(n34396), .B(reg_i_mask[13]), .X(n26245) );
  nand_x1_sg U60238 ( .A(\mask_0/reg_i_mask[13] ), .B(n32538), .X(n26246) );
  nand_x1_sg U60239 ( .A(n33879), .B(reg_i_mask[12]), .X(n26243) );
  nand_x1_sg U60240 ( .A(\mask_0/reg_i_mask[12] ), .B(n32529), .X(n26244) );
  nand_x1_sg U60241 ( .A(n34397), .B(reg_i_mask[11]), .X(n26241) );
  nand_x1_sg U60242 ( .A(\mask_0/reg_i_mask[11] ), .B(n32528), .X(n26242) );
  nand_x1_sg U60243 ( .A(n34391), .B(reg_i_mask[10]), .X(n26239) );
  nand_x1_sg U60244 ( .A(\mask_0/reg_i_mask[10] ), .B(n32532), .X(n26240) );
  nand_x1_sg U60245 ( .A(n33885), .B(reg_i_mask[9]), .X(n26237) );
  nand_x1_sg U60246 ( .A(\mask_0/reg_i_mask[9] ), .B(n32536), .X(n26238) );
  nand_x1_sg U60247 ( .A(n34389), .B(reg_i_mask[8]), .X(n26235) );
  nand_x1_sg U60248 ( .A(\mask_0/reg_i_mask[8] ), .B(n32537), .X(n26236) );
  nand_x1_sg U60249 ( .A(n34401), .B(reg_i_mask[7]), .X(n26233) );
  nand_x1_sg U60250 ( .A(\mask_0/reg_i_mask[7] ), .B(n30645), .X(n26234) );
  nand_x1_sg U60251 ( .A(n33887), .B(reg_i_mask[6]), .X(n26231) );
  nand_x1_sg U60252 ( .A(\mask_0/reg_i_mask[6] ), .B(n34796), .X(n26232) );
  nand_x1_sg U60253 ( .A(n33884), .B(reg_i_mask[5]), .X(n26229) );
  nand_x1_sg U60254 ( .A(\mask_0/reg_i_mask[5] ), .B(n32539), .X(n26230) );
  nand_x1_sg U60255 ( .A(n34400), .B(reg_i_mask[4]), .X(n26227) );
  nand_x1_sg U60256 ( .A(\mask_0/reg_i_mask[4] ), .B(n34796), .X(n26228) );
  nand_x1_sg U60257 ( .A(n33881), .B(reg_i_mask[3]), .X(n26225) );
  nand_x1_sg U60258 ( .A(\mask_0/reg_i_mask[3] ), .B(n30644), .X(n26226) );
  nand_x1_sg U60259 ( .A(n33882), .B(reg_i_mask[2]), .X(n26223) );
  nand_x1_sg U60260 ( .A(\mask_0/reg_i_mask[2] ), .B(n32528), .X(n26224) );
  nand_x1_sg U60261 ( .A(n33888), .B(reg_i_mask[1]), .X(n26221) );
  nand_x1_sg U60262 ( .A(\mask_0/reg_i_mask[1] ), .B(n32529), .X(n26222) );
  nand_x1_sg U60263 ( .A(n33884), .B(reg_i_mask[0]), .X(n26217) );
  nand_x1_sg U60264 ( .A(\mask_0/reg_i_mask[0] ), .B(n34798), .X(n26218) );
  nor_x1_sg U60265 ( .A(\shifter_0/reg_i_7[3] ), .B(\shifter_0/reg_i_7[4] ), 
        .X(n21531) );
  nor_x1_sg U60266 ( .A(\shifter_0/reg_i_7[1] ), .B(\shifter_0/reg_i_7[19] ), 
        .X(n21529) );
  nand_x1_sg U60267 ( .A(n35141), .B(n21531), .X(n21530) );
  nor_x1_sg U60268 ( .A(shifter_state[1]), .B(n35251), .X(n21744) );
  nand_x1_sg U60269 ( .A(\mask_0/state[0] ), .B(n42529), .X(n26206) );
  nor_x1_sg U60270 ( .A(\filter_0/i_pointer[1] ), .B(\filter_0/i_pointer[0] ), 
        .X(n28967) );
  nor_x1_sg U60271 ( .A(\shifter_0/reg_w_7[10] ), .B(\shifter_0/reg_w_7[0] ), 
        .X(n21141) );
  nand_x1_sg U60272 ( .A(n32884), .B(\filter_0/done ), .X(n26576) );
  nand_x1_sg U60273 ( .A(n26578), .B(filter_state[1]), .X(n26577) );
  nor_x1_sg U60274 ( .A(n31670), .B(\shifter_0/i_pointer[1] ), .X(n11637) );
  nor_x1_sg U60275 ( .A(\shifter_0/reg_w_8[8] ), .B(\shifter_0/reg_w_8[9] ), 
        .X(n21238) );
  nor_x1_sg U60276 ( .A(\shifter_0/reg_w_8[3] ), .B(\shifter_0/reg_w_8[4] ), 
        .X(n21235) );
  nor_x1_sg U60277 ( .A(\shifter_0/reg_w_8[17] ), .B(\shifter_0/reg_w_8[18] ), 
        .X(n21246) );
  nor_x1_sg U60278 ( .A(\shifter_0/reg_w_8[6] ), .B(\shifter_0/reg_w_8[5] ), 
        .X(n21236) );
  nor_x1_sg U60279 ( .A(\shifter_0/reg_w_8[7] ), .B(n42719), .X(n21237) );
  nor_x1_sg U60280 ( .A(\shifter_0/reg_w_8[1] ), .B(\shifter_0/reg_w_8[19] ), 
        .X(n21233) );
  nor_x1_sg U60281 ( .A(\shifter_0/reg_w_8[2] ), .B(n42718), .X(n21234) );
  nor_x1_sg U60282 ( .A(\shifter_0/reg_w_8[15] ), .B(\shifter_0/reg_w_8[14] ), 
        .X(n21244) );
  nor_x1_sg U60283 ( .A(\shifter_0/reg_w_8[16] ), .B(n42721), .X(n21245) );
  nor_x1_sg U60284 ( .A(\shifter_0/reg_i_8[8] ), .B(\shifter_0/reg_i_8[9] ), 
        .X(n21591) );
  nor_x1_sg U60285 ( .A(\shifter_0/reg_w_8[11] ), .B(n42720), .X(n21242) );
  nor_x1_sg U60286 ( .A(\shifter_0/reg_w_8[12] ), .B(\shifter_0/reg_w_8[13] ), 
        .X(n21243) );
  nor_x1_sg U60287 ( .A(\shifter_0/reg_i_8[6] ), .B(\shifter_0/reg_i_8[5] ), 
        .X(n21589) );
  nor_x1_sg U60288 ( .A(\shifter_0/reg_i_8[7] ), .B(n42608), .X(n21590) );
  nor_x1_sg U60289 ( .A(\shifter_0/reg_i_8[12] ), .B(\shifter_0/reg_i_8[13] ), 
        .X(n21596) );
  nor_x1_sg U60290 ( .A(\shifter_0/reg_i_8[10] ), .B(\shifter_0/reg_i_8[0] ), 
        .X(n21594) );
  nor_x1_sg U60291 ( .A(\shifter_0/reg_i_8[11] ), .B(n42609), .X(n21595) );
  nor_x1_sg U60292 ( .A(\shifter_0/reg_i_7[16] ), .B(n21542), .X(n21541) );
  nand_x1_sg U60293 ( .A(n35140), .B(n35139), .X(n21542) );
  nor_x1_sg U60294 ( .A(\shifter_0/reg_i_7[15] ), .B(\shifter_0/reg_i_7[14] ), 
        .X(n21540) );
  nor_x1_sg U60295 ( .A(\shifter_0/reg_i_8[3] ), .B(\shifter_0/reg_i_8[4] ), 
        .X(n21588) );
  nor_x1_sg U60296 ( .A(\shifter_0/reg_i_8[1] ), .B(\shifter_0/reg_i_8[19] ), 
        .X(n21586) );
  nor_x1_sg U60297 ( .A(\shifter_0/reg_i_8[2] ), .B(n42607), .X(n21587) );
  nor_x1_sg U60298 ( .A(\shifter_0/reg_i_14[3] ), .B(\shifter_0/reg_i_14[4] ), 
        .X(n21713) );
  nor_x1_sg U60299 ( .A(\shifter_0/reg_i_14[1] ), .B(\shifter_0/reg_i_14[19] ), 
        .X(n21711) );
  nor_x1_sg U60300 ( .A(\shifter_0/reg_i_14[2] ), .B(n42643), .X(n21712) );
  nor_x1_sg U60301 ( .A(\shifter_0/reg_i_8[16] ), .B(n42610), .X(n21598) );
  nor_x1_sg U60302 ( .A(\shifter_0/reg_i_8[17] ), .B(\shifter_0/reg_i_8[18] ), 
        .X(n21599) );
  nor_x1_sg U60303 ( .A(n26200), .B(\mask_0/state[0] ), .X(n26347) );
  nand_x1_sg U60304 ( .A(\filter_0/w_pointer[3] ), .B(n35256), .X(n29620) );
  nand_x1_sg U60305 ( .A(\filter_0/w_pointer[3] ), .B(\filter_0/w_pointer[2] ), 
        .X(n29444) );
  nand_x1_sg U60306 ( .A(\filter_0/i_pointer[3] ), .B(\filter_0/i_pointer[2] ), 
        .X(n28745) );
  nor_x1_sg U60307 ( .A(\shifter_0/reg_i_12[3] ), .B(\shifter_0/reg_i_12[4] ), 
        .X(n21695) );
  nor_x1_sg U60308 ( .A(\shifter_0/reg_i_12[1] ), .B(\shifter_0/reg_i_12[19] ), 
        .X(n21693) );
  nor_x1_sg U60309 ( .A(\shifter_0/reg_i_12[2] ), .B(n42629), .X(n21694) );
  nand_x1_sg U60310 ( .A(\filter_0/i_pointer[3] ), .B(n35258), .X(n28921) );
  nor_x1_sg U60311 ( .A(\shifter_0/reg_w_14[7] ), .B(n21216), .X(n21215) );
  nor_x1_sg U60312 ( .A(\shifter_0/reg_w_14[6] ), .B(\shifter_0/reg_w_14[5] ), 
        .X(n21214) );
  nand_x1_sg U60313 ( .A(n42760), .B(n42761), .X(n21216) );
  nor_x1_sg U60314 ( .A(\shifter_0/reg_w_14[2] ), .B(n21213), .X(n21212) );
  nor_x1_sg U60315 ( .A(\shifter_0/reg_w_14[1] ), .B(\shifter_0/reg_w_14[19] ), 
        .X(n21211) );
  nand_x1_sg U60316 ( .A(n42758), .B(n42759), .X(n21213) );
  nor_x1_sg U60317 ( .A(\shifter_0/reg_w_14[16] ), .B(n21224), .X(n21223) );
  nor_x1_sg U60318 ( .A(\shifter_0/reg_w_14[15] ), .B(\shifter_0/reg_w_14[14] ), .X(n21222) );
  nand_x1_sg U60319 ( .A(n42764), .B(n42765), .X(n21224) );
  nor_x1_sg U60320 ( .A(\shifter_0/reg_w_14[10] ), .B(\shifter_0/reg_w_14[0] ), 
        .X(n21219) );
  nor_x1_sg U60321 ( .A(\shifter_0/reg_w_14[11] ), .B(n21221), .X(n21220) );
  nand_x1_sg U60322 ( .A(n42762), .B(n42763), .X(n21221) );
  nor_x1_sg U60323 ( .A(n30460), .B(n21059), .X(n21058) );
  nor_x1_sg U60324 ( .A(n30459), .B(n30458), .X(n21057) );
  nand_x1_sg U60325 ( .A(n42684), .B(n42685), .X(n21059) );
  nor_x1_sg U60326 ( .A(n30461), .B(n30455), .X(n21062) );
  nor_x1_sg U60327 ( .A(n30462), .B(n21064), .X(n21063) );
  nand_x1_sg U60328 ( .A(n42686), .B(n42687), .X(n21064) );
  nor_x1_sg U60329 ( .A(n30457), .B(n21056), .X(n21055) );
  nor_x1_sg U60330 ( .A(n30456), .B(n30466), .X(n21054) );
  nand_x1_sg U60331 ( .A(n42682), .B(n42683), .X(n21056) );
  nor_x1_sg U60332 ( .A(n30465), .B(n21067), .X(n21066) );
  nor_x1_sg U60333 ( .A(n30464), .B(n30463), .X(n21065) );
  nand_x1_sg U60334 ( .A(n42688), .B(n42689), .X(n21067) );
  nor_x1_sg U60335 ( .A(\shifter_0/reg_w_12[7] ), .B(n21198), .X(n21197) );
  nor_x1_sg U60336 ( .A(\shifter_0/reg_w_12[6] ), .B(\shifter_0/reg_w_12[5] ), 
        .X(n21196) );
  nand_x1_sg U60337 ( .A(n42744), .B(n42745), .X(n21198) );
  nor_x1_sg U60338 ( .A(\shifter_0/reg_w_12[16] ), .B(n21206), .X(n21205) );
  nor_x1_sg U60339 ( .A(\shifter_0/reg_w_12[15] ), .B(\shifter_0/reg_w_12[14] ), .X(n21204) );
  nand_x1_sg U60340 ( .A(n42748), .B(n42749), .X(n21206) );
  nor_x1_sg U60341 ( .A(\shifter_0/reg_i_9[3] ), .B(\shifter_0/reg_i_9[4] ), 
        .X(n21644) );
  nor_x1_sg U60342 ( .A(\shifter_0/reg_w_12[10] ), .B(\shifter_0/reg_w_12[0] ), 
        .X(n21201) );
  nor_x1_sg U60343 ( .A(\shifter_0/reg_w_12[11] ), .B(n21203), .X(n21202) );
  nand_x1_sg U60344 ( .A(n42746), .B(n42747), .X(n21203) );
  nor_x1_sg U60345 ( .A(\shifter_0/reg_w_12[2] ), .B(n21195), .X(n21194) );
  nor_x1_sg U60346 ( .A(\shifter_0/reg_w_12[1] ), .B(\shifter_0/reg_w_12[19] ), 
        .X(n21193) );
  nand_x1_sg U60347 ( .A(n42742), .B(n42743), .X(n21195) );
  inv_x1_sg U60348 ( .A(\shifter_0/reg_w_3[4] ), .X(n42683) );
  inv_x1_sg U60349 ( .A(\shifter_0/reg_w_3[9] ), .X(n42685) );
  inv_x1_sg U60350 ( .A(\shifter_0/reg_w_3[18] ), .X(n42689) );
  nor_x1_sg U60351 ( .A(\shifter_0/reg_i_9[1] ), .B(\shifter_0/reg_i_9[19] ), 
        .X(n21642) );
  nor_x1_sg U60352 ( .A(\shifter_0/reg_i_9[2] ), .B(n42611), .X(n21643) );
  inv_x1_sg U60353 ( .A(\shifter_0/reg_w_3[3] ), .X(n42682) );
  inv_x1_sg U60354 ( .A(\shifter_0/reg_w_3[8] ), .X(n42684) );
  inv_x1_sg U60355 ( .A(\shifter_0/reg_w_3[12] ), .X(n42686) );
  inv_x1_sg U60356 ( .A(\shifter_0/reg_w_3[13] ), .X(n42687) );
  inv_x1_sg U60357 ( .A(\shifter_0/reg_w_3[17] ), .X(n42688) );
  nand_x1_sg U60358 ( .A(mask_input_ready), .B(n42529), .X(n26200) );
  inv_x1_sg U60359 ( .A(\shifter_0/reg_w_14[9] ), .X(n42761) );
  inv_x1_sg U60360 ( .A(\shifter_0/reg_w_14[8] ), .X(n42760) );
  inv_x1_sg U60361 ( .A(\shifter_0/reg_w_14[4] ), .X(n42759) );
  inv_x1_sg U60362 ( .A(\shifter_0/reg_w_14[3] ), .X(n42758) );
  inv_x1_sg U60363 ( .A(\shifter_0/reg_w_14[18] ), .X(n42765) );
  inv_x1_sg U60364 ( .A(\shifter_0/reg_w_14[17] ), .X(n42764) );
  inv_x1_sg U60365 ( .A(\shifter_0/reg_w_14[13] ), .X(n42763) );
  nor_x1_sg U60366 ( .A(\shifter_0/reg_i_14[17] ), .B(\shifter_0/reg_i_14[18] ), .X(n21724) );
  inv_x1_sg U60367 ( .A(\shifter_0/reg_w_14[12] ), .X(n42762) );
  nor_x1_sg U60368 ( .A(\shifter_0/reg_i_14[15] ), .B(\shifter_0/reg_i_14[14] ), .X(n21722) );
  nand_x1_sg U60369 ( .A(n42649), .B(n21724), .X(n21723) );
  nor_x1_sg U60370 ( .A(n31708), .B(\shifter_0/w_pointer[1] ), .X(n11612) );
  nor_x1_sg U60371 ( .A(\shifter_0/reg_i_11[3] ), .B(\shifter_0/reg_i_11[4] ), 
        .X(n21626) );
  nor_x1_sg U60372 ( .A(\shifter_0/reg_i_10[8] ), .B(\shifter_0/reg_i_10[9] ), 
        .X(n21609) );
  nor_x1_sg U60373 ( .A(\shifter_0/reg_i_11[1] ), .B(\shifter_0/reg_i_11[19] ), 
        .X(n21624) );
  nor_x1_sg U60374 ( .A(\shifter_0/reg_i_11[2] ), .B(n42622), .X(n21625) );
  nor_x1_sg U60375 ( .A(\shifter_0/reg_i_10[6] ), .B(\shifter_0/reg_i_10[5] ), 
        .X(n21607) );
  nor_x1_sg U60376 ( .A(\shifter_0/reg_i_10[7] ), .B(n42619), .X(n21608) );
  nor_x1_sg U60377 ( .A(\shifter_0/reg_i_10[12] ), .B(\shifter_0/reg_i_10[13] ), .X(n21614) );
  nor_x1_sg U60378 ( .A(\shifter_0/reg_i_10[10] ), .B(\shifter_0/reg_i_10[0] ), 
        .X(n21612) );
  nor_x1_sg U60379 ( .A(\shifter_0/reg_i_10[11] ), .B(n42620), .X(n21613) );
  inv_x1_sg U60380 ( .A(\shifter_0/reg_w_12[9] ), .X(n42745) );
  inv_x1_sg U60381 ( .A(\shifter_0/reg_w_12[8] ), .X(n42744) );
  inv_x1_sg U60382 ( .A(\shifter_0/reg_w_12[4] ), .X(n42743) );
  inv_x1_sg U60383 ( .A(\shifter_0/reg_w_12[18] ), .X(n42749) );
  nor_x1_sg U60384 ( .A(\shifter_0/reg_w_10[8] ), .B(\shifter_0/reg_w_10[9] ), 
        .X(n21256) );
  nor_x1_sg U60385 ( .A(\shifter_0/reg_w_10[17] ), .B(\shifter_0/reg_w_10[18] ), .X(n21264) );
  nor_x1_sg U60386 ( .A(\shifter_0/reg_i_10[3] ), .B(\shifter_0/reg_i_10[4] ), 
        .X(n21606) );
  nor_x1_sg U60387 ( .A(n30396), .B(n30390), .X(n21445) );
  nor_x1_sg U60388 ( .A(\shifter_0/reg_w_8[10] ), .B(\shifter_0/reg_w_8[0] ), 
        .X(n21241) );
  nor_x1_sg U60389 ( .A(\shifter_0/reg_i_8[15] ), .B(\shifter_0/reg_i_8[14] ), 
        .X(n21597) );
  nor_x1_sg U60390 ( .A(\shifter_0/reg_i_10[1] ), .B(\shifter_0/reg_i_10[19] ), 
        .X(n21604) );
  nor_x1_sg U60391 ( .A(\shifter_0/reg_i_10[2] ), .B(n42618), .X(n21605) );
  inv_x1_sg U60392 ( .A(\shifter_0/reg_w_12[3] ), .X(n42742) );
  inv_x1_sg U60393 ( .A(\shifter_0/reg_w_12[17] ), .X(n42748) );
  inv_x1_sg U60394 ( .A(\shifter_0/reg_w_12[13] ), .X(n42747) );
  inv_x1_sg U60395 ( .A(\shifter_0/reg_w_12[12] ), .X(n42746) );
  nor_x1_sg U60396 ( .A(n30395), .B(n21442), .X(n21441) );
  nor_x1_sg U60397 ( .A(n30394), .B(n30393), .X(n21440) );
  nand_x1_sg U60398 ( .A(n42574), .B(n42575), .X(n21442) );
  nor_x1_sg U60399 ( .A(n30392), .B(n21439), .X(n21438) );
  nor_x1_sg U60400 ( .A(n30391), .B(n30401), .X(n21437) );
  nand_x1_sg U60401 ( .A(n42572), .B(n42573), .X(n21439) );
  nor_x1_sg U60402 ( .A(n30400), .B(n21450), .X(n21449) );
  nor_x1_sg U60403 ( .A(n30399), .B(n30398), .X(n21448) );
  nand_x1_sg U60404 ( .A(n42578), .B(n42579), .X(n21450) );
  nor_x1_sg U60405 ( .A(\shifter_0/reg_w_10[6] ), .B(\shifter_0/reg_w_10[5] ), 
        .X(n21254) );
  nor_x1_sg U60406 ( .A(\shifter_0/reg_w_10[7] ), .B(n42731), .X(n21255) );
  nor_x1_sg U60407 ( .A(\shifter_0/reg_w_10[15] ), .B(\shifter_0/reg_w_10[14] ), .X(n21262) );
  nor_x1_sg U60408 ( .A(\shifter_0/reg_w_10[16] ), .B(n42733), .X(n21263) );
  nor_x1_sg U60409 ( .A(\shifter_0/reg_w_10[3] ), .B(\shifter_0/reg_w_10[4] ), 
        .X(n21253) );
  nor_x1_sg U60410 ( .A(n30397), .B(n21447), .X(n21446) );
  nand_x1_sg U60411 ( .A(n42576), .B(n42577), .X(n21447) );
  nor_x1_sg U60412 ( .A(\shifter_0/reg_w_10[11] ), .B(n42732), .X(n21260) );
  nor_x1_sg U60413 ( .A(\shifter_0/reg_w_10[12] ), .B(\shifter_0/reg_w_10[13] ), .X(n21261) );
  nor_x1_sg U60414 ( .A(\shifter_0/reg_i_12[17] ), .B(\shifter_0/reg_i_12[18] ), .X(n21706) );
  nor_x1_sg U60415 ( .A(\shifter_0/reg_i_12[15] ), .B(\shifter_0/reg_i_12[14] ), .X(n21704) );
  nand_x1_sg U60416 ( .A(n42635), .B(n21706), .X(n21705) );
  nor_x1_sg U60417 ( .A(\shifter_0/reg_w_10[1] ), .B(\shifter_0/reg_w_10[19] ), 
        .X(n21251) );
  nor_x1_sg U60418 ( .A(\shifter_0/reg_w_10[2] ), .B(n42730), .X(n21252) );
  nor_x1_sg U60419 ( .A(n42532), .B(n33964), .X(n26583) );
  inv_x1_sg U60420 ( .A(\filter_0/done ), .X(n42532) );
  nor_x1_sg U60421 ( .A(\shifter_0/reg_w_6[7] ), .B(n21118), .X(n21117) );
  nor_x1_sg U60422 ( .A(\shifter_0/reg_w_6[6] ), .B(\shifter_0/reg_w_6[5] ), 
        .X(n21116) );
  nand_x1_sg U60423 ( .A(n42708), .B(n42709), .X(n21118) );
  nor_x1_sg U60424 ( .A(\shifter_0/reg_i_14[10] ), .B(\shifter_0/reg_i_14[0] ), 
        .X(n21719) );
  nor_x1_sg U60425 ( .A(\shifter_0/reg_i_14[11] ), .B(n21721), .X(n21720) );
  nand_x1_sg U60426 ( .A(n42646), .B(n42647), .X(n21721) );
  nor_x1_sg U60427 ( .A(\shifter_0/reg_i_14[7] ), .B(n21716), .X(n21715) );
  nor_x1_sg U60428 ( .A(\shifter_0/reg_i_14[6] ), .B(\shifter_0/reg_i_14[5] ), 
        .X(n21714) );
  nand_x1_sg U60429 ( .A(n42644), .B(n42645), .X(n21716) );
  nor_x1_sg U60430 ( .A(\shifter_0/reg_i_10[16] ), .B(n42621), .X(n21616) );
  nor_x1_sg U60431 ( .A(\shifter_0/reg_i_10[17] ), .B(\shifter_0/reg_i_10[18] ), .X(n21617) );
  nor_x1_sg U60432 ( .A(\shifter_0/reg_w_6[10] ), .B(\shifter_0/reg_w_6[0] ), 
        .X(n21121) );
  nor_x1_sg U60433 ( .A(\shifter_0/reg_w_6[11] ), .B(n21123), .X(n21122) );
  nand_x1_sg U60434 ( .A(n42710), .B(n42711), .X(n21123) );
  inv_x1_sg U60435 ( .A(\shifter_0/reg_i_3[9] ), .X(n42575) );
  nor_x1_sg U60436 ( .A(\shifter_0/reg_w_6[2] ), .B(n21115), .X(n21114) );
  nor_x1_sg U60437 ( .A(\shifter_0/reg_w_6[1] ), .B(\shifter_0/reg_w_6[19] ), 
        .X(n21113) );
  nand_x1_sg U60438 ( .A(n42706), .B(n42707), .X(n21115) );
  nor_x1_sg U60439 ( .A(\shifter_0/reg_w_6[16] ), .B(n21126), .X(n21125) );
  nor_x1_sg U60440 ( .A(\shifter_0/reg_w_6[15] ), .B(\shifter_0/reg_w_6[14] ), 
        .X(n21124) );
  nand_x1_sg U60441 ( .A(n42712), .B(n42713), .X(n21126) );
  nor_x1_sg U60442 ( .A(\shifter_0/reg_w_5[7] ), .B(n21156), .X(n21155) );
  nor_x1_sg U60443 ( .A(\shifter_0/reg_w_5[6] ), .B(\shifter_0/reg_w_5[5] ), 
        .X(n21154) );
  nand_x1_sg U60444 ( .A(n42700), .B(n42701), .X(n21156) );
  inv_x1_sg U60445 ( .A(\shifter_0/reg_i_3[3] ), .X(n42572) );
  inv_x1_sg U60446 ( .A(\shifter_0/reg_i_3[4] ), .X(n42573) );
  inv_x1_sg U60447 ( .A(\shifter_0/reg_i_3[8] ), .X(n42574) );
  inv_x1_sg U60448 ( .A(\shifter_0/reg_i_3[13] ), .X(n42577) );
  inv_x1_sg U60449 ( .A(\shifter_0/reg_i_3[17] ), .X(n42578) );
  inv_x1_sg U60450 ( .A(\shifter_0/reg_i_3[18] ), .X(n42579) );
  nor_x1_sg U60451 ( .A(\shifter_0/reg_w_5[10] ), .B(\shifter_0/reg_w_5[0] ), 
        .X(n21159) );
  nor_x1_sg U60452 ( .A(\shifter_0/reg_w_5[11] ), .B(n21161), .X(n21160) );
  nand_x1_sg U60453 ( .A(n42702), .B(n42703), .X(n21161) );
  nor_x1_sg U60454 ( .A(\shifter_0/reg_w_5[2] ), .B(n21153), .X(n21152) );
  nor_x1_sg U60455 ( .A(\shifter_0/reg_w_5[1] ), .B(\shifter_0/reg_w_5[19] ), 
        .X(n21151) );
  nand_x1_sg U60456 ( .A(n42698), .B(n42699), .X(n21153) );
  nor_x1_sg U60457 ( .A(\shifter_0/reg_w_5[16] ), .B(n21164), .X(n21163) );
  nor_x1_sg U60458 ( .A(\shifter_0/reg_w_5[15] ), .B(\shifter_0/reg_w_5[14] ), 
        .X(n21162) );
  nand_x1_sg U60459 ( .A(n42704), .B(n42705), .X(n21164) );
  inv_x1_sg U60460 ( .A(\shifter_0/reg_i_3[12] ), .X(n42576) );
  nor_x1_sg U60461 ( .A(\shifter_0/reg_i_12[7] ), .B(n21698), .X(n21697) );
  nor_x1_sg U60462 ( .A(\shifter_0/reg_i_12[6] ), .B(\shifter_0/reg_i_12[5] ), 
        .X(n21696) );
  nand_x1_sg U60463 ( .A(n42630), .B(n42631), .X(n21698) );
  nand_x1_sg U60464 ( .A(\shifter_0/i_pointer[1] ), .B(n31669), .X(n19587) );
  nor_x1_sg U60465 ( .A(\shifter_0/reg_i_13[3] ), .B(\shifter_0/reg_i_13[4] ), 
        .X(n21674) );
  nor_x1_sg U60466 ( .A(\shifter_0/reg_i_12[10] ), .B(\shifter_0/reg_i_12[0] ), 
        .X(n21701) );
  nor_x1_sg U60467 ( .A(\shifter_0/reg_i_12[11] ), .B(n21703), .X(n21702) );
  nand_x1_sg U60468 ( .A(n42632), .B(n42633), .X(n21703) );
  nor_x1_sg U60469 ( .A(\shifter_0/reg_i_9[17] ), .B(\shifter_0/reg_i_9[18] ), 
        .X(n21655) );
  nor_x1_sg U60470 ( .A(\shifter_0/reg_i_13[1] ), .B(\shifter_0/reg_i_13[19] ), 
        .X(n21672) );
  nor_x1_sg U60471 ( .A(\shifter_0/reg_i_13[2] ), .B(n42636), .X(n21673) );
  inv_x1_sg U60472 ( .A(\shifter_0/reg_w_6[4] ), .X(n42707) );
  inv_x1_sg U60473 ( .A(\shifter_0/reg_w_6[8] ), .X(n42708) );
  inv_x1_sg U60474 ( .A(\shifter_0/reg_w_6[9] ), .X(n42709) );
  inv_x1_sg U60475 ( .A(\shifter_0/reg_w_6[18] ), .X(n42713) );
  inv_x1_sg U60476 ( .A(\shifter_0/reg_i_14[9] ), .X(n42645) );
  nor_x1_sg U60477 ( .A(\shifter_0/reg_i_9[15] ), .B(\shifter_0/reg_i_9[14] ), 
        .X(n21653) );
  nand_x1_sg U60478 ( .A(n42617), .B(n21655), .X(n21654) );
  inv_x1_sg U60479 ( .A(\shifter_0/reg_w_6[3] ), .X(n42706) );
  inv_x1_sg U60480 ( .A(\shifter_0/reg_w_6[12] ), .X(n42710) );
  inv_x1_sg U60481 ( .A(\shifter_0/reg_w_6[13] ), .X(n42711) );
  inv_x1_sg U60482 ( .A(\shifter_0/reg_w_6[17] ), .X(n42712) );
  inv_x1_sg U60483 ( .A(\shifter_0/reg_i_14[8] ), .X(n42644) );
  inv_x1_sg U60484 ( .A(\shifter_0/reg_i_14[13] ), .X(n42647) );
  inv_x1_sg U60485 ( .A(\shifter_0/reg_i_14[12] ), .X(n42646) );
  inv_x1_sg U60486 ( .A(\shifter_0/reg_w_5[4] ), .X(n42699) );
  inv_x1_sg U60487 ( .A(\shifter_0/reg_w_5[8] ), .X(n42700) );
  inv_x1_sg U60488 ( .A(\shifter_0/reg_w_5[9] ), .X(n42701) );
  inv_x1_sg U60489 ( .A(\shifter_0/reg_w_5[18] ), .X(n42705) );
  nor_x1_sg U60490 ( .A(\shifter_0/reg_w_2[2] ), .B(n21036), .X(n21035) );
  nor_x1_sg U60491 ( .A(\shifter_0/reg_w_2[1] ), .B(\shifter_0/reg_w_2[19] ), 
        .X(n21034) );
  nand_x1_sg U60492 ( .A(n42674), .B(n42675), .X(n21036) );
  nor_x1_sg U60493 ( .A(\shifter_0/reg_w_2[16] ), .B(n21047), .X(n21046) );
  nor_x1_sg U60494 ( .A(\shifter_0/reg_w_2[15] ), .B(\shifter_0/reg_w_2[14] ), 
        .X(n21045) );
  nand_x1_sg U60495 ( .A(n42680), .B(n42681), .X(n21047) );
  inv_x1_sg U60496 ( .A(\shifter_0/reg_w_5[3] ), .X(n42698) );
  inv_x1_sg U60497 ( .A(\shifter_0/reg_w_5[12] ), .X(n42702) );
  inv_x1_sg U60498 ( .A(\shifter_0/reg_w_5[13] ), .X(n42703) );
  inv_x1_sg U60499 ( .A(\shifter_0/reg_w_5[17] ), .X(n42704) );
  nor_x1_sg U60500 ( .A(\shifter_0/reg_w_2[7] ), .B(n21039), .X(n21038) );
  nor_x1_sg U60501 ( .A(\shifter_0/reg_w_2[6] ), .B(\shifter_0/reg_w_2[5] ), 
        .X(n21037) );
  nand_x1_sg U60502 ( .A(n42676), .B(n42677), .X(n21039) );
  nor_x1_sg U60503 ( .A(\shifter_0/reg_w_2[10] ), .B(\shifter_0/reg_w_2[0] ), 
        .X(n21042) );
  nor_x1_sg U60504 ( .A(\shifter_0/reg_w_2[11] ), .B(n21044), .X(n21043) );
  nand_x1_sg U60505 ( .A(n42678), .B(n42679), .X(n21044) );
  nor_x1_sg U60506 ( .A(\shifter_0/reg_i_11[17] ), .B(\shifter_0/reg_i_11[18] ), .X(n21637) );
  inv_x1_sg U60507 ( .A(\shifter_0/reg_i_12[9] ), .X(n42631) );
  nor_x1_sg U60508 ( .A(\shifter_0/reg_i_11[15] ), .B(\shifter_0/reg_i_11[14] ), .X(n21635) );
  nand_x1_sg U60509 ( .A(n42628), .B(n21637), .X(n21636) );
  nor_x1_sg U60510 ( .A(\shifter_0/reg_i_6[2] ), .B(n21511), .X(n21510) );
  nor_x1_sg U60511 ( .A(\shifter_0/reg_i_6[1] ), .B(\shifter_0/reg_i_6[19] ), 
        .X(n21509) );
  nand_x1_sg U60512 ( .A(n42596), .B(n42597), .X(n21511) );
  nor_x1_sg U60513 ( .A(\shifter_0/reg_i_6[16] ), .B(n21522), .X(n21521) );
  nor_x1_sg U60514 ( .A(\shifter_0/reg_i_6[15] ), .B(\shifter_0/reg_i_6[14] ), 
        .X(n21520) );
  nand_x1_sg U60515 ( .A(n42602), .B(n42603), .X(n21522) );
  inv_x1_sg U60516 ( .A(\shifter_0/reg_i_12[8] ), .X(n42630) );
  inv_x1_sg U60517 ( .A(\shifter_0/reg_i_12[13] ), .X(n42633) );
  nor_x1_sg U60518 ( .A(\shifter_0/reg_i_6[7] ), .B(n21514), .X(n21513) );
  nor_x1_sg U60519 ( .A(\shifter_0/reg_i_6[6] ), .B(\shifter_0/reg_i_6[5] ), 
        .X(n21512) );
  nand_x1_sg U60520 ( .A(n42598), .B(n42599), .X(n21514) );
  nor_x1_sg U60521 ( .A(\shifter_0/reg_i_6[10] ), .B(\shifter_0/reg_i_6[0] ), 
        .X(n21517) );
  nor_x1_sg U60522 ( .A(\shifter_0/reg_i_6[11] ), .B(n21519), .X(n21518) );
  nand_x1_sg U60523 ( .A(n42600), .B(n42601), .X(n21519) );
  nor_x1_sg U60524 ( .A(\shifter_0/reg_i_9[10] ), .B(\shifter_0/reg_i_9[0] ), 
        .X(n21650) );
  nor_x1_sg U60525 ( .A(\shifter_0/reg_i_9[11] ), .B(n21652), .X(n21651) );
  nand_x1_sg U60526 ( .A(n42614), .B(n42615), .X(n21652) );
  nor_x1_sg U60527 ( .A(\shifter_0/reg_i_9[7] ), .B(n21647), .X(n21646) );
  nor_x1_sg U60528 ( .A(\shifter_0/reg_i_9[6] ), .B(\shifter_0/reg_i_9[5] ), 
        .X(n21645) );
  nand_x1_sg U60529 ( .A(n42612), .B(n42613), .X(n21647) );
  inv_x1_sg U60530 ( .A(\shifter_0/reg_i_12[12] ), .X(n42632) );
  inv_x1_sg U60531 ( .A(\shifter_0/reg_i_14[16] ), .X(n42649) );
  nor_x1_sg U60532 ( .A(\shifter_0/reg_i_5[7] ), .B(n21552), .X(n21551) );
  nor_x1_sg U60533 ( .A(\shifter_0/reg_i_5[6] ), .B(\shifter_0/reg_i_5[5] ), 
        .X(n21550) );
  nand_x1_sg U60534 ( .A(n42590), .B(n42591), .X(n21552) );
  nor_x1_sg U60535 ( .A(\shifter_0/reg_i_5[2] ), .B(n21549), .X(n21548) );
  nor_x1_sg U60536 ( .A(\shifter_0/reg_i_5[1] ), .B(\shifter_0/reg_i_5[19] ), 
        .X(n21547) );
  nand_x1_sg U60537 ( .A(n42588), .B(n42589), .X(n21549) );
  nor_x1_sg U60538 ( .A(\shifter_0/reg_i_5[16] ), .B(n21560), .X(n21559) );
  nor_x1_sg U60539 ( .A(\shifter_0/reg_i_5[15] ), .B(\shifter_0/reg_i_5[14] ), 
        .X(n21558) );
  nand_x1_sg U60540 ( .A(n42594), .B(n42595), .X(n21560) );
  inv_x1_sg U60541 ( .A(\shifter_0/reg_w_2[9] ), .X(n42677) );
  nor_x1_sg U60542 ( .A(\shifter_0/reg_i_5[10] ), .B(\shifter_0/reg_i_5[0] ), 
        .X(n21555) );
  nor_x1_sg U60543 ( .A(\shifter_0/reg_i_5[11] ), .B(n21557), .X(n21556) );
  nand_x1_sg U60544 ( .A(n42592), .B(n42593), .X(n21557) );
  nor_x1_sg U60545 ( .A(\shifter_0/reg_w_9[7] ), .B(n21294), .X(n21293) );
  nor_x1_sg U60546 ( .A(\shifter_0/reg_w_9[6] ), .B(\shifter_0/reg_w_9[5] ), 
        .X(n21292) );
  nand_x1_sg U60547 ( .A(n42724), .B(n42725), .X(n21294) );
  inv_x1_sg U60548 ( .A(\shifter_0/reg_w_2[3] ), .X(n42674) );
  inv_x1_sg U60549 ( .A(\shifter_0/reg_w_2[4] ), .X(n42675) );
  inv_x1_sg U60550 ( .A(\shifter_0/reg_w_2[8] ), .X(n42676) );
  inv_x1_sg U60551 ( .A(\shifter_0/reg_w_2[13] ), .X(n42679) );
  inv_x1_sg U60552 ( .A(\shifter_0/reg_w_2[17] ), .X(n42680) );
  inv_x1_sg U60553 ( .A(\shifter_0/reg_w_2[18] ), .X(n42681) );
  nor_x1_sg U60554 ( .A(\shifter_0/reg_w_9[10] ), .B(\shifter_0/reg_w_9[0] ), 
        .X(n21297) );
  nor_x1_sg U60555 ( .A(\shifter_0/reg_w_9[11] ), .B(n21299), .X(n21298) );
  nand_x1_sg U60556 ( .A(n42726), .B(n42727), .X(n21299) );
  nor_x1_sg U60557 ( .A(\shifter_0/reg_i_11[7] ), .B(n21629), .X(n21628) );
  nor_x1_sg U60558 ( .A(\shifter_0/reg_i_11[6] ), .B(\shifter_0/reg_i_11[5] ), 
        .X(n21627) );
  nand_x1_sg U60559 ( .A(n42623), .B(n42624), .X(n21629) );
  nor_x1_sg U60560 ( .A(\shifter_0/reg_w_13[7] ), .B(n21177), .X(n21176) );
  nor_x1_sg U60561 ( .A(\shifter_0/reg_w_13[6] ), .B(\shifter_0/reg_w_13[5] ), 
        .X(n21175) );
  nand_x1_sg U60562 ( .A(n42752), .B(n42753), .X(n21177) );
  nor_x1_sg U60563 ( .A(\shifter_0/reg_w_13[2] ), .B(n21174), .X(n21173) );
  nor_x1_sg U60564 ( .A(\shifter_0/reg_w_13[1] ), .B(\shifter_0/reg_w_13[19] ), 
        .X(n21172) );
  nand_x1_sg U60565 ( .A(n42750), .B(n42751), .X(n21174) );
  nor_x1_sg U60566 ( .A(\shifter_0/reg_w_13[16] ), .B(n21185), .X(n21184) );
  nor_x1_sg U60567 ( .A(\shifter_0/reg_w_13[15] ), .B(\shifter_0/reg_w_13[14] ), .X(n21183) );
  nand_x1_sg U60568 ( .A(n42756), .B(n42757), .X(n21185) );
  nor_x1_sg U60569 ( .A(\shifter_0/reg_w_9[2] ), .B(n21291), .X(n21290) );
  nor_x1_sg U60570 ( .A(\shifter_0/reg_w_9[1] ), .B(\shifter_0/reg_w_9[19] ), 
        .X(n21289) );
  nand_x1_sg U60571 ( .A(n42722), .B(n42723), .X(n21291) );
  nor_x1_sg U60572 ( .A(\shifter_0/reg_w_9[16] ), .B(n21302), .X(n21301) );
  nor_x1_sg U60573 ( .A(\shifter_0/reg_w_9[15] ), .B(\shifter_0/reg_w_9[14] ), 
        .X(n21300) );
  nand_x1_sg U60574 ( .A(n42728), .B(n42729), .X(n21302) );
  inv_x1_sg U60575 ( .A(\shifter_0/reg_i_6[9] ), .X(n42599) );
  inv_x1_sg U60576 ( .A(\shifter_0/reg_w_2[12] ), .X(n42678) );
  nor_x1_sg U60577 ( .A(\shifter_0/reg_i_2[7] ), .B(n21422), .X(n21421) );
  nor_x1_sg U60578 ( .A(\shifter_0/reg_i_2[6] ), .B(\shifter_0/reg_i_2[5] ), 
        .X(n21420) );
  nand_x1_sg U60579 ( .A(n42566), .B(n42567), .X(n21422) );
  nor_x1_sg U60580 ( .A(\shifter_0/reg_i_11[10] ), .B(\shifter_0/reg_i_11[0] ), 
        .X(n21632) );
  nor_x1_sg U60581 ( .A(\shifter_0/reg_i_11[11] ), .B(n21634), .X(n21633) );
  nand_x1_sg U60582 ( .A(n42625), .B(n42626), .X(n21634) );
  nor_x1_sg U60583 ( .A(\shifter_0/reg_w_11[7] ), .B(n21276), .X(n21275) );
  nor_x1_sg U60584 ( .A(\shifter_0/reg_w_11[6] ), .B(\shifter_0/reg_w_11[5] ), 
        .X(n21274) );
  nand_x1_sg U60585 ( .A(n42736), .B(n42737), .X(n21276) );
  nor_x1_sg U60586 ( .A(\shifter_0/reg_w_11[2] ), .B(n21273), .X(n21272) );
  nor_x1_sg U60587 ( .A(\shifter_0/reg_w_11[1] ), .B(\shifter_0/reg_w_11[19] ), 
        .X(n21271) );
  nand_x1_sg U60588 ( .A(n42734), .B(n42735), .X(n21273) );
  nor_x1_sg U60589 ( .A(\shifter_0/reg_w_11[16] ), .B(n21284), .X(n21283) );
  nor_x1_sg U60590 ( .A(\shifter_0/reg_w_11[15] ), .B(\shifter_0/reg_w_11[14] ), .X(n21282) );
  nand_x1_sg U60591 ( .A(n42740), .B(n42741), .X(n21284) );
  nor_x1_sg U60592 ( .A(\shifter_0/reg_w_13[10] ), .B(\shifter_0/reg_w_13[0] ), 
        .X(n21180) );
  nor_x1_sg U60593 ( .A(\shifter_0/reg_w_13[11] ), .B(n21182), .X(n21181) );
  nand_x1_sg U60594 ( .A(n42754), .B(n42755), .X(n21182) );
  inv_x1_sg U60595 ( .A(\shifter_0/reg_i_6[3] ), .X(n42596) );
  inv_x1_sg U60596 ( .A(\shifter_0/reg_i_6[4] ), .X(n42597) );
  inv_x1_sg U60597 ( .A(\shifter_0/reg_i_6[8] ), .X(n42598) );
  inv_x1_sg U60598 ( .A(\shifter_0/reg_i_6[13] ), .X(n42601) );
  inv_x1_sg U60599 ( .A(\shifter_0/reg_i_6[17] ), .X(n42602) );
  inv_x1_sg U60600 ( .A(\shifter_0/reg_i_6[18] ), .X(n42603) );
  nor_x1_sg U60601 ( .A(\shifter_0/reg_i_2[2] ), .B(n21419), .X(n21418) );
  nor_x1_sg U60602 ( .A(\shifter_0/reg_i_2[1] ), .B(\shifter_0/reg_i_2[19] ), 
        .X(n21417) );
  nand_x1_sg U60603 ( .A(n42564), .B(n42565), .X(n21419) );
  nor_x1_sg U60604 ( .A(\shifter_0/reg_i_2[16] ), .B(n21430), .X(n21429) );
  nor_x1_sg U60605 ( .A(\shifter_0/reg_i_2[15] ), .B(\shifter_0/reg_i_2[14] ), 
        .X(n21428) );
  nand_x1_sg U60606 ( .A(n42570), .B(n42571), .X(n21430) );
  nor_x1_sg U60607 ( .A(\shifter_0/reg_i_2[10] ), .B(\shifter_0/reg_i_2[0] ), 
        .X(n21425) );
  nor_x1_sg U60608 ( .A(\shifter_0/reg_i_2[11] ), .B(n21427), .X(n21426) );
  nand_x1_sg U60609 ( .A(n42568), .B(n42569), .X(n21427) );
  nor_x1_sg U60610 ( .A(\shifter_0/reg_w_11[10] ), .B(\shifter_0/reg_w_11[0] ), 
        .X(n21279) );
  nor_x1_sg U60611 ( .A(\shifter_0/reg_w_11[11] ), .B(n21281), .X(n21280) );
  nand_x1_sg U60612 ( .A(n42738), .B(n42739), .X(n21281) );
  inv_x1_sg U60613 ( .A(\shifter_0/reg_i_6[12] ), .X(n42600) );
  inv_x1_sg U60614 ( .A(\shifter_0/reg_i_5[9] ), .X(n42591) );
  inv_x1_sg U60615 ( .A(\shifter_0/reg_w_1[4] ), .X(n42667) );
  inv_x1_sg U60616 ( .A(\shifter_0/reg_w_1[8] ), .X(n42668) );
  inv_x1_sg U60617 ( .A(\shifter_0/reg_w_1[9] ), .X(n42669) );
  inv_x1_sg U60618 ( .A(\shifter_0/reg_w_1[18] ), .X(n42673) );
  inv_x1_sg U60619 ( .A(\shifter_0/reg_i_12[16] ), .X(n42635) );
  inv_x1_sg U60620 ( .A(\shifter_0/reg_i_9[9] ), .X(n42613) );
  nor_x1_sg U60621 ( .A(\shifter_0/reg_w_1[6] ), .B(\shifter_0/reg_w_1[5] ), 
        .X(n21075) );
  nor_x1_sg U60622 ( .A(\shifter_0/reg_w_1[7] ), .B(n21077), .X(n21076) );
  nand_x1_sg U60623 ( .A(n42668), .B(n42669), .X(n21077) );
  nor_x1_sg U60624 ( .A(\shifter_0/reg_w_1[1] ), .B(\shifter_0/reg_w_1[19] ), 
        .X(n21072) );
  nor_x1_sg U60625 ( .A(\shifter_0/reg_w_1[2] ), .B(n21074), .X(n21073) );
  nand_x1_sg U60626 ( .A(n42666), .B(n42667), .X(n21074) );
  nor_x1_sg U60627 ( .A(\shifter_0/reg_w_1[15] ), .B(\shifter_0/reg_w_1[14] ), 
        .X(n21083) );
  nor_x1_sg U60628 ( .A(\shifter_0/reg_w_1[16] ), .B(n21085), .X(n21084) );
  nand_x1_sg U60629 ( .A(n42672), .B(n42673), .X(n21085) );
  nor_x1_sg U60630 ( .A(\shifter_0/reg_i_10[15] ), .B(\shifter_0/reg_i_10[14] ), .X(n21615) );
  nor_x1_sg U60631 ( .A(\shifter_0/reg_w_1[11] ), .B(n21082), .X(n21081) );
  nand_x1_sg U60632 ( .A(n42670), .B(n42671), .X(n21082) );
  inv_x1_sg U60633 ( .A(\shifter_0/reg_i_5[3] ), .X(n42588) );
  inv_x1_sg U60634 ( .A(\shifter_0/reg_i_5[4] ), .X(n42589) );
  inv_x1_sg U60635 ( .A(\shifter_0/reg_i_5[8] ), .X(n42590) );
  inv_x1_sg U60636 ( .A(\shifter_0/reg_i_5[13] ), .X(n42593) );
  inv_x1_sg U60637 ( .A(\shifter_0/reg_i_5[17] ), .X(n42594) );
  inv_x1_sg U60638 ( .A(\shifter_0/reg_i_5[18] ), .X(n42595) );
  inv_x1_sg U60639 ( .A(\shifter_0/reg_w_1[3] ), .X(n42666) );
  inv_x1_sg U60640 ( .A(\shifter_0/reg_w_1[12] ), .X(n42670) );
  inv_x1_sg U60641 ( .A(\shifter_0/reg_w_1[13] ), .X(n42671) );
  inv_x1_sg U60642 ( .A(\shifter_0/reg_w_1[17] ), .X(n42672) );
  inv_x1_sg U60643 ( .A(\shifter_0/reg_i_9[8] ), .X(n42612) );
  inv_x1_sg U60644 ( .A(\shifter_0/reg_i_9[13] ), .X(n42615) );
  inv_x1_sg U60645 ( .A(\shifter_0/reg_i_9[12] ), .X(n42614) );
  inv_x1_sg U60646 ( .A(\shifter_0/reg_i_5[12] ), .X(n42592) );
  nor_x1_sg U60647 ( .A(\shifter_0/reg_i_13[17] ), .B(\shifter_0/reg_i_13[18] ), .X(n21685) );
  inv_x1_sg U60648 ( .A(\shifter_0/reg_i_2[9] ), .X(n42567) );
  inv_x1_sg U60649 ( .A(\shifter_0/reg_w_9[18] ), .X(n42729) );
  inv_x1_sg U60650 ( .A(\shifter_0/reg_w_9[9] ), .X(n42725) );
  nor_x1_sg U60651 ( .A(\shifter_0/reg_i_13[15] ), .B(\shifter_0/reg_i_13[14] ), .X(n21683) );
  nand_x1_sg U60652 ( .A(n42642), .B(n21685), .X(n21684) );
  nor_x1_sg U60653 ( .A(\shifter_0/reg_w_10[10] ), .B(\shifter_0/reg_w_10[0] ), 
        .X(n21259) );
  nor_x1_sg U60654 ( .A(\shifter_0/reg_w_1[10] ), .B(\shifter_0/reg_w_1[0] ), 
        .X(n21080) );
  inv_x1_sg U60655 ( .A(\shifter_0/reg_i_2[3] ), .X(n42564) );
  inv_x1_sg U60656 ( .A(\shifter_0/reg_i_2[4] ), .X(n42565) );
  inv_x1_sg U60657 ( .A(\shifter_0/reg_i_2[8] ), .X(n42566) );
  inv_x1_sg U60658 ( .A(\shifter_0/reg_i_2[13] ), .X(n42569) );
  inv_x1_sg U60659 ( .A(\shifter_0/reg_i_2[17] ), .X(n42570) );
  inv_x1_sg U60660 ( .A(\shifter_0/reg_i_2[18] ), .X(n42571) );
  inv_x1_sg U60661 ( .A(\shifter_0/reg_i_11[9] ), .X(n42624) );
  inv_x1_sg U60662 ( .A(\shifter_0/reg_i_11[8] ), .X(n42623) );
  inv_x1_sg U60663 ( .A(\shifter_0/reg_w_13[9] ), .X(n42753) );
  inv_x1_sg U60664 ( .A(\shifter_0/reg_w_13[8] ), .X(n42752) );
  inv_x1_sg U60665 ( .A(\shifter_0/reg_w_13[4] ), .X(n42751) );
  inv_x1_sg U60666 ( .A(\shifter_0/reg_w_13[3] ), .X(n42750) );
  inv_x1_sg U60667 ( .A(\shifter_0/reg_w_13[18] ), .X(n42757) );
  inv_x1_sg U60668 ( .A(\shifter_0/reg_w_13[17] ), .X(n42756) );
  inv_x1_sg U60669 ( .A(\shifter_0/reg_w_13[13] ), .X(n42755) );
  inv_x1_sg U60670 ( .A(\shifter_0/reg_w_9[4] ), .X(n42723) );
  inv_x1_sg U60671 ( .A(\shifter_0/reg_w_9[3] ), .X(n42722) );
  inv_x1_sg U60672 ( .A(\shifter_0/reg_w_9[17] ), .X(n42728) );
  inv_x1_sg U60673 ( .A(\shifter_0/reg_w_9[8] ), .X(n42724) );
  inv_x1_sg U60674 ( .A(\shifter_0/reg_w_9[12] ), .X(n42726) );
  inv_x1_sg U60675 ( .A(\shifter_0/reg_w_9[13] ), .X(n42727) );
  inv_x1_sg U60676 ( .A(\shifter_0/reg_i_2[12] ), .X(n42568) );
  inv_x1_sg U60677 ( .A(\shifter_0/reg_w_11[9] ), .X(n42737) );
  inv_x1_sg U60678 ( .A(\shifter_0/reg_w_11[8] ), .X(n42736) );
  inv_x1_sg U60679 ( .A(\shifter_0/reg_w_11[4] ), .X(n42735) );
  inv_x1_sg U60680 ( .A(\shifter_0/reg_w_11[3] ), .X(n42734) );
  inv_x1_sg U60681 ( .A(\shifter_0/reg_w_11[18] ), .X(n42741) );
  inv_x1_sg U60682 ( .A(\shifter_0/reg_w_11[17] ), .X(n42740) );
  inv_x1_sg U60683 ( .A(\shifter_0/reg_w_11[13] ), .X(n42739) );
  inv_x1_sg U60684 ( .A(\shifter_0/reg_i_11[13] ), .X(n42626) );
  inv_x1_sg U60685 ( .A(\shifter_0/reg_i_11[12] ), .X(n42625) );
  inv_x1_sg U60686 ( .A(\shifter_0/reg_w_13[12] ), .X(n42754) );
  nor_x1_sg U60687 ( .A(\shifter_0/reg_i_1[11] ), .B(n21465), .X(n21464) );
  nand_x1_sg U60688 ( .A(n42560), .B(n42561), .X(n21465) );
  inv_x1_sg U60689 ( .A(\shifter_0/reg_i_1[4] ), .X(n42557) );
  inv_x1_sg U60690 ( .A(\shifter_0/reg_i_1[8] ), .X(n42558) );
  inv_x1_sg U60691 ( .A(\shifter_0/reg_i_1[9] ), .X(n42559) );
  inv_x1_sg U60692 ( .A(\shifter_0/reg_i_1[13] ), .X(n42561) );
  inv_x1_sg U60693 ( .A(\shifter_0/reg_i_1[17] ), .X(n42562) );
  inv_x1_sg U60694 ( .A(\shifter_0/reg_i_1[18] ), .X(n42563) );
  inv_x1_sg U60695 ( .A(\shifter_0/reg_w_11[12] ), .X(n42738) );
  inv_x1_sg U60696 ( .A(\shifter_0/reg_i_9[16] ), .X(n42617) );
  nor_x1_sg U60697 ( .A(\shifter_0/reg_i_1[6] ), .B(\shifter_0/reg_i_1[5] ), 
        .X(n21458) );
  nor_x1_sg U60698 ( .A(\shifter_0/reg_i_1[7] ), .B(n21460), .X(n21459) );
  nand_x1_sg U60699 ( .A(n42558), .B(n42559), .X(n21460) );
  nor_x1_sg U60700 ( .A(\shifter_0/reg_i_1[1] ), .B(\shifter_0/reg_i_1[19] ), 
        .X(n21455) );
  nor_x1_sg U60701 ( .A(\shifter_0/reg_i_1[2] ), .B(n21457), .X(n21456) );
  nand_x1_sg U60702 ( .A(n42556), .B(n42557), .X(n21457) );
  nor_x1_sg U60703 ( .A(\shifter_0/reg_i_1[15] ), .B(\shifter_0/reg_i_1[14] ), 
        .X(n21466) );
  nor_x1_sg U60704 ( .A(\shifter_0/reg_i_1[16] ), .B(n21468), .X(n21467) );
  nand_x1_sg U60705 ( .A(n42562), .B(n42563), .X(n21468) );
  nand_x1_sg U60706 ( .A(\shifter_0/w_pointer[1] ), .B(n31708), .X(n19586) );
  inv_x1_sg U60707 ( .A(\shifter_0/reg_i_1[3] ), .X(n42556) );
  inv_x1_sg U60708 ( .A(\shifter_0/reg_i_1[12] ), .X(n42560) );
  nor_x1_sg U60709 ( .A(\shifter_0/reg_i_13[10] ), .B(\shifter_0/reg_i_13[0] ), 
        .X(n21680) );
  nor_x1_sg U60710 ( .A(\shifter_0/reg_i_13[7] ), .B(n21677), .X(n21676) );
  nor_x1_sg U60711 ( .A(\shifter_0/reg_i_13[6] ), .B(\shifter_0/reg_i_13[5] ), 
        .X(n21675) );
  nand_x1_sg U60712 ( .A(n42637), .B(n42638), .X(n21677) );
  nor_x1_sg U60713 ( .A(\shifter_0/reg_i_13[11] ), .B(n21682), .X(n21681) );
  nand_x1_sg U60714 ( .A(n42639), .B(n42640), .X(n21682) );
  nor_x1_sg U60715 ( .A(\shifter_0/reg_i_1[10] ), .B(\shifter_0/reg_i_1[0] ), 
        .X(n21463) );
  inv_x1_sg U60716 ( .A(\shifter_0/reg_i_11[16] ), .X(n42628) );
  inv_x1_sg U60717 ( .A(\shifter_0/reg_i_13[9] ), .X(n42638) );
  inv_x1_sg U60718 ( .A(\shifter_0/reg_i_13[8] ), .X(n42637) );
  inv_x1_sg U60719 ( .A(\shifter_0/reg_i_13[13] ), .X(n42640) );
  nor_x1_sg U60720 ( .A(\shifter_0/reg_w_0[7] ), .B(n21021), .X(n21020) );
  nor_x1_sg U60721 ( .A(\shifter_0/reg_w_0[6] ), .B(\shifter_0/reg_w_0[5] ), 
        .X(n21019) );
  nand_x1_sg U60722 ( .A(n42660), .B(n42661), .X(n21021) );
  nor_x1_sg U60723 ( .A(\shifter_0/reg_w_0[16] ), .B(n21029), .X(n21028) );
  nor_x1_sg U60724 ( .A(\shifter_0/reg_w_0[15] ), .B(\shifter_0/reg_w_0[14] ), 
        .X(n21027) );
  nand_x1_sg U60725 ( .A(n42664), .B(n42665), .X(n21029) );
  inv_x1_sg U60726 ( .A(\shifter_0/reg_i_13[12] ), .X(n42639) );
  nor_x1_sg U60727 ( .A(\shifter_0/reg_w_0[10] ), .B(\shifter_0/reg_w_0[0] ), 
        .X(n21024) );
  nor_x1_sg U60728 ( .A(\shifter_0/reg_w_0[11] ), .B(n21026), .X(n21025) );
  nand_x1_sg U60729 ( .A(n42662), .B(n42663), .X(n21026) );
  nor_x1_sg U60730 ( .A(\shifter_0/reg_w_0[2] ), .B(n21018), .X(n21017) );
  nor_x1_sg U60731 ( .A(\shifter_0/reg_w_0[1] ), .B(\shifter_0/reg_w_0[19] ), 
        .X(n21016) );
  nand_x1_sg U60732 ( .A(n42658), .B(n42659), .X(n21018) );
  nor_x1_sg U60733 ( .A(\shifter_0/reg_i_15[4] ), .B(n21735), .X(n21732) );
  nand_x1_sg U60734 ( .A(n42651), .B(n42652), .X(n21735) );
  nor_x1_sg U60735 ( .A(n30446), .B(n21731), .X(n21730) );
  nor_x1_sg U60736 ( .A(n30454), .B(\shifter_0/reg_i_15[18] ), .X(n21729) );
  nand_x1_sg U60737 ( .A(n35136), .B(n42650), .X(n21731) );
  inv_x1_sg U60738 ( .A(\shifter_0/reg_w_4[3] ), .X(n42690) );
  inv_x1_sg U60739 ( .A(\shifter_0/reg_w_4[4] ), .X(n42691) );
  inv_x1_sg U60740 ( .A(\shifter_0/reg_w_4[8] ), .X(n42692) );
  inv_x1_sg U60741 ( .A(\shifter_0/reg_w_4[9] ), .X(n42693) );
  inv_x1_sg U60742 ( .A(\shifter_0/reg_w_4[13] ), .X(n42695) );
  inv_x1_sg U60743 ( .A(\shifter_0/reg_w_4[17] ), .X(n42696) );
  inv_x1_sg U60744 ( .A(\shifter_0/reg_w_4[18] ), .X(n42697) );
  nor_x1_sg U60745 ( .A(\shifter_0/reg_w_4[11] ), .B(n21105), .X(n21104) );
  nand_x1_sg U60746 ( .A(n42694), .B(n42695), .X(n21105) );
  nor_x1_sg U60747 ( .A(\shifter_0/reg_w_4[6] ), .B(\shifter_0/reg_w_4[5] ), 
        .X(n21098) );
  nor_x1_sg U60748 ( .A(\shifter_0/reg_w_4[7] ), .B(n21100), .X(n21099) );
  nand_x1_sg U60749 ( .A(n42692), .B(n42693), .X(n21100) );
  nor_x1_sg U60750 ( .A(\shifter_0/reg_w_4[1] ), .B(\shifter_0/reg_w_4[19] ), 
        .X(n21095) );
  nor_x1_sg U60751 ( .A(\shifter_0/reg_w_4[2] ), .B(n21097), .X(n21096) );
  nand_x1_sg U60752 ( .A(n42690), .B(n42691), .X(n21097) );
  nor_x1_sg U60753 ( .A(\shifter_0/reg_w_4[15] ), .B(\shifter_0/reg_w_4[14] ), 
        .X(n21106) );
  nor_x1_sg U60754 ( .A(\shifter_0/reg_w_4[16] ), .B(n21108), .X(n21107) );
  nand_x1_sg U60755 ( .A(n42696), .B(n42697), .X(n21108) );
  inv_x1_sg U60756 ( .A(\shifter_0/reg_w_4[12] ), .X(n42694) );
  nor_x1_sg U60757 ( .A(n30451), .B(n30450), .X(n21741) );
  nor_x1_sg U60758 ( .A(n30452), .B(n21743), .X(n21742) );
  nand_x1_sg U60759 ( .A(n42657), .B(n35130), .X(n21743) );
  inv_x1_sg U60760 ( .A(\shifter_0/reg_i_13[16] ), .X(n42642) );
  nor_x1_sg U60761 ( .A(n30509), .B(n21315), .X(n21312) );
  nor_x1_sg U60762 ( .A(n30510), .B(n21314), .X(n21313) );
  nand_x1_sg U60763 ( .A(n42768), .B(n42769), .X(n21315) );
  inv_x1_sg U60764 ( .A(\shifter_0/reg_w_15[9] ), .X(n42771) );
  nor_x1_sg U60765 ( .A(\shifter_0/reg_w_4[10] ), .B(\shifter_0/reg_w_4[0] ), 
        .X(n21103) );
  inv_x1_sg U60766 ( .A(\shifter_0/reg_w_0[4] ), .X(n42659) );
  inv_x1_sg U60767 ( .A(\shifter_0/reg_w_0[8] ), .X(n42660) );
  inv_x1_sg U60768 ( .A(\shifter_0/reg_w_0[9] ), .X(n42661) );
  inv_x1_sg U60769 ( .A(\shifter_0/reg_w_0[13] ), .X(n42663) );
  inv_x1_sg U60770 ( .A(\shifter_0/reg_w_0[17] ), .X(n42664) );
  inv_x1_sg U60771 ( .A(\shifter_0/reg_w_0[18] ), .X(n42665) );
  nor_x1_sg U60772 ( .A(n30513), .B(n30512), .X(n21321) );
  nor_x1_sg U60773 ( .A(n30514), .B(n21323), .X(n21322) );
  nand_x1_sg U60774 ( .A(n42774), .B(n42775), .X(n21323) );
  nor_x1_sg U60775 ( .A(n30516), .B(n30515), .X(n21309) );
  nor_x1_sg U60776 ( .A(n30508), .B(n21311), .X(n21310) );
  nand_x1_sg U60777 ( .A(n42766), .B(n42767), .X(n21311) );
  inv_x1_sg U60778 ( .A(\shifter_0/reg_w_15[8] ), .X(n42770) );
  inv_x1_sg U60779 ( .A(\shifter_0/reg_w_15[12] ), .X(n42773) );
  inv_x1_sg U60780 ( .A(\shifter_0/reg_w_15[17] ), .X(n42775) );
  inv_x1_sg U60781 ( .A(\shifter_0/reg_w_15[16] ), .X(n42774) );
  inv_x1_sg U60782 ( .A(\shifter_0/reg_w_15[6] ), .X(n42769) );
  inv_x1_sg U60783 ( .A(\shifter_0/reg_w_15[3] ), .X(n42767) );
  inv_x1_sg U60784 ( .A(\shifter_0/reg_w_0[3] ), .X(n42658) );
  inv_x1_sg U60785 ( .A(\shifter_0/reg_w_0[12] ), .X(n42662) );
  inv_x1_sg U60786 ( .A(\shifter_0/reg_w_15[11] ), .X(n42772) );
  inv_x1_sg U60787 ( .A(\shifter_0/reg_w_15[5] ), .X(n42768) );
  inv_x1_sg U60788 ( .A(\shifter_0/reg_w_15[2] ), .X(n42766) );
  nor_x1_sg U60789 ( .A(\shifter_0/reg_i_0[7] ), .B(n21404), .X(n21403) );
  nor_x1_sg U60790 ( .A(\shifter_0/reg_i_0[6] ), .B(\shifter_0/reg_i_0[5] ), 
        .X(n21402) );
  nand_x1_sg U60791 ( .A(n42550), .B(n42551), .X(n21404) );
  nor_x1_sg U60792 ( .A(\shifter_0/reg_i_0[10] ), .B(\shifter_0/reg_i_0[0] ), 
        .X(n21407) );
  nor_x1_sg U60793 ( .A(\shifter_0/reg_i_0[11] ), .B(n21409), .X(n21408) );
  nand_x1_sg U60794 ( .A(n42552), .B(n42553), .X(n21409) );
  nor_x1_sg U60795 ( .A(\shifter_0/reg_i_0[2] ), .B(n21401), .X(n21400) );
  nor_x1_sg U60796 ( .A(\shifter_0/reg_i_0[1] ), .B(\shifter_0/reg_i_0[19] ), 
        .X(n21399) );
  nand_x1_sg U60797 ( .A(n42548), .B(n42549), .X(n21401) );
  nor_x1_sg U60798 ( .A(\shifter_0/reg_i_0[16] ), .B(n21412), .X(n21411) );
  nor_x1_sg U60799 ( .A(\shifter_0/reg_i_0[15] ), .B(\shifter_0/reg_i_0[14] ), 
        .X(n21410) );
  nand_x1_sg U60800 ( .A(n42554), .B(n42555), .X(n21412) );
  inv_x1_sg U60801 ( .A(\shifter_0/reg_i_4[18] ), .X(n42587) );
  inv_x1_sg U60802 ( .A(\shifter_0/reg_i_4[9] ), .X(n42583) );
  nor_x1_sg U60803 ( .A(\shifter_0/reg_i_4[6] ), .B(\shifter_0/reg_i_4[5] ), 
        .X(n21494) );
  nor_x1_sg U60804 ( .A(\shifter_0/reg_i_4[7] ), .B(n21496), .X(n21495) );
  nand_x1_sg U60805 ( .A(n42582), .B(n42583), .X(n21496) );
  nor_x1_sg U60806 ( .A(\shifter_0/reg_i_4[15] ), .B(\shifter_0/reg_i_4[14] ), 
        .X(n21502) );
  nor_x1_sg U60807 ( .A(\shifter_0/reg_i_4[16] ), .B(n21504), .X(n21503) );
  nand_x1_sg U60808 ( .A(n42586), .B(n42587), .X(n21504) );
  inv_x1_sg U60809 ( .A(\shifter_0/reg_i_4[4] ), .X(n42581) );
  inv_x1_sg U60810 ( .A(\shifter_0/reg_i_4[17] ), .X(n42586) );
  inv_x1_sg U60811 ( .A(\shifter_0/reg_i_4[3] ), .X(n42580) );
  inv_x1_sg U60812 ( .A(\shifter_0/reg_i_4[8] ), .X(n42582) );
  inv_x1_sg U60813 ( .A(\shifter_0/reg_i_4[12] ), .X(n42584) );
  inv_x1_sg U60814 ( .A(\shifter_0/reg_i_4[13] ), .X(n42585) );
  nor_x1_sg U60815 ( .A(\shifter_0/reg_i_4[11] ), .B(n21501), .X(n21500) );
  nand_x1_sg U60816 ( .A(n42584), .B(n42585), .X(n21501) );
  nor_x1_sg U60817 ( .A(\shifter_0/reg_i_4[1] ), .B(\shifter_0/reg_i_4[19] ), 
        .X(n21491) );
  nor_x1_sg U60818 ( .A(\shifter_0/reg_i_4[2] ), .B(n21493), .X(n21492) );
  nand_x1_sg U60819 ( .A(n42580), .B(n42581), .X(n21493) );
  nor_x1_sg U60820 ( .A(\shifter_0/reg_i_4[10] ), .B(\shifter_0/reg_i_4[0] ), 
        .X(n21499) );
  inv_x1_sg U60821 ( .A(\shifter_0/reg_i_0[4] ), .X(n42549) );
  inv_x1_sg U60822 ( .A(\shifter_0/reg_i_0[8] ), .X(n42550) );
  inv_x1_sg U60823 ( .A(\shifter_0/reg_i_0[9] ), .X(n42551) );
  inv_x1_sg U60824 ( .A(\shifter_0/reg_i_0[18] ), .X(n42555) );
  nand_x1_sg U60825 ( .A(n26216), .B(n42528), .X(n26214) );
  nor_x1_sg U60826 ( .A(\mask_0/counter[1] ), .B(\mask_0/counter[0] ), .X(
        n26216) );
  nand_x1_sg U60827 ( .A(n26209), .B(\mask_0/state[0] ), .X(n26210) );
  nor_x1_sg U60828 ( .A(n26209), .B(n42527), .X(n26212) );
  inv_x1_sg U60829 ( .A(\shifter_0/reg_i_0[3] ), .X(n42548) );
  inv_x1_sg U60830 ( .A(\shifter_0/reg_i_0[12] ), .X(n42552) );
  inv_x1_sg U60831 ( .A(\shifter_0/reg_i_0[13] ), .X(n42553) );
  inv_x1_sg U60832 ( .A(\shifter_0/reg_i_0[17] ), .X(n42554) );
  nor_x1_sg U60833 ( .A(n30448), .B(n21734), .X(n21733) );
  nand_x1_sg U60834 ( .A(n42653), .B(n42654), .X(n21734) );
  inv_x1_sg U60835 ( .A(\shifter_0/reg_i_15[12] ), .X(n42656) );
  inv_x1_sg U60836 ( .A(\shifter_0/reg_i_15[3] ), .X(n42650) );
  inv_x1_sg U60837 ( .A(\shifter_0/reg_i_15[6] ), .X(n42652) );
  inv_x1_sg U60838 ( .A(\shifter_0/reg_i_15[9] ), .X(n42654) );
  inv_x1_sg U60839 ( .A(\shifter_0/reg_i_15[8] ), .X(n42653) );
  inv_x1_sg U60840 ( .A(\shifter_0/reg_i_15[11] ), .X(n42655) );
  inv_x1_sg U60841 ( .A(\shifter_0/reg_i_15[16] ), .X(n42657) );
  inv_x1_sg U60842 ( .A(\shifter_0/reg_i_15[5] ), .X(n42651) );
  nand_x1_sg U60843 ( .A(n42527), .B(n35418), .X(n26207) );
  nand_x1_sg U60844 ( .A(n26209), .B(\mask_0/state[1] ), .X(n26208) );
  nand_x1_sg U60845 ( .A(n26203), .B(n42528), .X(n26202) );
  nand_x1_sg U60846 ( .A(\mask_0/counter[1] ), .B(n26204), .X(n26201) );
  nor_x1_sg U60847 ( .A(\mask_0/counter[1] ), .B(n42530), .X(n26203) );
  nand_x1_sg U60848 ( .A(n26197), .B(n26198), .X(\mask_0/n774 ) );
  nand_x1_sg U60849 ( .A(n26199), .B(\mask_0/counter[0] ), .X(n26198) );
  nor_x1_sg U60850 ( .A(n42528), .B(n42411), .X(n26199) );
  inv_x1_sg U60851 ( .A(n26200), .X(n42411) );
  nor_x1_sg U60852 ( .A(n22219), .B(n22220), .X(n22214) );
  nand_x1_sg U60853 ( .A(n35251), .B(shifter_state[1]), .X(n22219) );
  inv_x1_sg U60854 ( .A(o_mask[30]), .X(n42494) );
  inv_x1_sg U60855 ( .A(o_mask[29]), .X(n42493) );
  nor_x1_sg U60856 ( .A(n35581), .B(\mask_0/reg_ww_mask[31] ), .X(n28254) );
  nor_x1_sg U60857 ( .A(n42494), .B(\mask_0/reg_ww_mask[30] ), .X(n28249) );
  nor_x1_sg U60858 ( .A(n42493), .B(\mask_0/reg_ww_mask[29] ), .X(n28244) );
  inv_x1_sg U60859 ( .A(o_mask[27]), .X(n42492) );
  inv_x1_sg U60860 ( .A(o_mask[26]), .X(n42491) );
  inv_x1_sg U60861 ( .A(o_mask[24]), .X(n42490) );
  inv_x1_sg U60862 ( .A(o_mask[22]), .X(n42489) );
  inv_x1_sg U60863 ( .A(o_mask[21]), .X(n42488) );
  inv_x1_sg U60864 ( .A(o_mask[17]), .X(n42487) );
  inv_x1_sg U60865 ( .A(o_mask[16]), .X(n42486) );
  inv_x1_sg U60866 ( .A(o_mask[14]), .X(n42485) );
  inv_x1_sg U60867 ( .A(o_mask[13]), .X(n42484) );
  inv_x1_sg U60868 ( .A(o_mask[11]), .X(n42483) );
  inv_x1_sg U60869 ( .A(o_mask[10]), .X(n42482) );
  inv_x1_sg U60870 ( .A(o_mask[5]), .X(n42481) );
  inv_x1_sg U60871 ( .A(o_mask[2]), .X(n42480) );
  inv_x1_sg U60872 ( .A(o_mask[1]), .X(n42479) );
  nor_x1_sg U60873 ( .A(n35580), .B(\mask_0/reg_ww_mask[28] ), .X(n28239) );
  nor_x1_sg U60874 ( .A(n42492), .B(\mask_0/reg_ww_mask[27] ), .X(n28234) );
  nor_x1_sg U60875 ( .A(n42491), .B(\mask_0/reg_ww_mask[26] ), .X(n28229) );
  nor_x1_sg U60876 ( .A(n35579), .B(\mask_0/reg_ww_mask[25] ), .X(n28224) );
  nor_x1_sg U60877 ( .A(n42490), .B(\mask_0/reg_ww_mask[24] ), .X(n28219) );
  nor_x1_sg U60878 ( .A(n35578), .B(\mask_0/reg_ww_mask[23] ), .X(n28214) );
  nor_x1_sg U60879 ( .A(n42489), .B(\mask_0/reg_ww_mask[22] ), .X(n28209) );
  nor_x1_sg U60880 ( .A(n42488), .B(\mask_0/reg_ww_mask[21] ), .X(n28204) );
  nor_x1_sg U60881 ( .A(n35577), .B(\mask_0/reg_ww_mask[20] ), .X(n28199) );
  nor_x1_sg U60882 ( .A(n35576), .B(\mask_0/reg_ww_mask[19] ), .X(n28194) );
  nor_x1_sg U60883 ( .A(n35575), .B(\mask_0/reg_ww_mask[18] ), .X(n28189) );
  nor_x1_sg U60884 ( .A(n42487), .B(\mask_0/reg_ww_mask[17] ), .X(n28184) );
  nor_x1_sg U60885 ( .A(n42486), .B(\mask_0/reg_ww_mask[16] ), .X(n28179) );
  nor_x1_sg U60886 ( .A(n35574), .B(\mask_0/reg_ww_mask[15] ), .X(n28174) );
  nor_x1_sg U60887 ( .A(n42485), .B(\mask_0/reg_ww_mask[14] ), .X(n28169) );
  nor_x1_sg U60888 ( .A(n42484), .B(\mask_0/reg_ww_mask[13] ), .X(n28164) );
  nor_x1_sg U60889 ( .A(n35573), .B(\mask_0/reg_ww_mask[12] ), .X(n28159) );
  nor_x1_sg U60890 ( .A(n42483), .B(\mask_0/reg_ww_mask[11] ), .X(n28154) );
  nor_x1_sg U60891 ( .A(n42482), .B(\mask_0/reg_ww_mask[10] ), .X(n28149) );
  nor_x1_sg U60892 ( .A(n35572), .B(\mask_0/reg_ww_mask[9] ), .X(n28144) );
  nor_x1_sg U60893 ( .A(n35571), .B(\mask_0/reg_ww_mask[8] ), .X(n28139) );
  nor_x1_sg U60894 ( .A(n35570), .B(\mask_0/reg_ww_mask[7] ), .X(n28134) );
  nor_x1_sg U60895 ( .A(n35569), .B(\mask_0/reg_ww_mask[6] ), .X(n28129) );
  nor_x1_sg U60896 ( .A(n42481), .B(\mask_0/reg_ww_mask[5] ), .X(n28124) );
  nor_x1_sg U60897 ( .A(n35568), .B(\mask_0/reg_ww_mask[4] ), .X(n28119) );
  nor_x1_sg U60898 ( .A(n35567), .B(\mask_0/reg_ww_mask[3] ), .X(n28114) );
  nor_x1_sg U60899 ( .A(n42480), .B(\mask_0/reg_ww_mask[2] ), .X(n28109) );
  nor_x1_sg U60900 ( .A(n42479), .B(\mask_0/reg_ww_mask[1] ), .X(n28104) );
  nor_x1_sg U60901 ( .A(n35566), .B(\mask_0/reg_ww_mask[0] ), .X(n28099) );
  nor_x1_sg U60902 ( .A(n35581), .B(\mask_0/reg_ii_mask[31] ), .X(n28094) );
  nor_x1_sg U60903 ( .A(n42494), .B(\mask_0/reg_ii_mask[30] ), .X(n28089) );
  nor_x1_sg U60904 ( .A(n42493), .B(\mask_0/reg_ii_mask[29] ), .X(n28084) );
  nor_x1_sg U60905 ( .A(n35580), .B(\mask_0/reg_ii_mask[28] ), .X(n28079) );
  nor_x1_sg U60906 ( .A(n42492), .B(\mask_0/reg_ii_mask[27] ), .X(n28074) );
  nor_x1_sg U60907 ( .A(n42491), .B(\mask_0/reg_ii_mask[26] ), .X(n28069) );
  nor_x1_sg U60908 ( .A(n35579), .B(\mask_0/reg_ii_mask[25] ), .X(n28064) );
  nor_x1_sg U60909 ( .A(n42490), .B(\mask_0/reg_ii_mask[24] ), .X(n28059) );
  nor_x1_sg U60910 ( .A(n35578), .B(\mask_0/reg_ii_mask[23] ), .X(n28054) );
  nor_x1_sg U60911 ( .A(n42489), .B(\mask_0/reg_ii_mask[22] ), .X(n28049) );
  nor_x1_sg U60912 ( .A(n42488), .B(\mask_0/reg_ii_mask[21] ), .X(n28044) );
  nor_x1_sg U60913 ( .A(n35577), .B(\mask_0/reg_ii_mask[20] ), .X(n28039) );
  nor_x1_sg U60914 ( .A(n35576), .B(\mask_0/reg_ii_mask[19] ), .X(n28034) );
  nor_x1_sg U60915 ( .A(n35575), .B(\mask_0/reg_ii_mask[18] ), .X(n28029) );
  nor_x1_sg U60916 ( .A(n42487), .B(\mask_0/reg_ii_mask[17] ), .X(n28024) );
  nor_x1_sg U60917 ( .A(n42486), .B(\mask_0/reg_ii_mask[16] ), .X(n28019) );
  nor_x1_sg U60918 ( .A(n35574), .B(\mask_0/reg_ii_mask[15] ), .X(n28014) );
  nor_x1_sg U60919 ( .A(n42485), .B(\mask_0/reg_ii_mask[14] ), .X(n28009) );
  nor_x1_sg U60920 ( .A(n42484), .B(\mask_0/reg_ii_mask[13] ), .X(n28004) );
  nor_x1_sg U60921 ( .A(n35573), .B(\mask_0/reg_ii_mask[12] ), .X(n27999) );
  nor_x1_sg U60922 ( .A(n42483), .B(\mask_0/reg_ii_mask[11] ), .X(n27994) );
  nor_x1_sg U60923 ( .A(n42482), .B(\mask_0/reg_ii_mask[10] ), .X(n27989) );
  nor_x1_sg U60924 ( .A(n35572), .B(\mask_0/reg_ii_mask[9] ), .X(n27984) );
  nor_x1_sg U60925 ( .A(n35571), .B(\mask_0/reg_ii_mask[8] ), .X(n27979) );
  nor_x1_sg U60926 ( .A(n35570), .B(\mask_0/reg_ii_mask[7] ), .X(n27974) );
  nor_x1_sg U60927 ( .A(n35569), .B(\mask_0/reg_ii_mask[6] ), .X(n27969) );
  nor_x1_sg U60928 ( .A(n42481), .B(\mask_0/reg_ii_mask[5] ), .X(n27964) );
  nor_x1_sg U60929 ( .A(n35568), .B(\mask_0/reg_ii_mask[4] ), .X(n27959) );
  nor_x1_sg U60930 ( .A(n35567), .B(\mask_0/reg_ii_mask[3] ), .X(n27954) );
  nor_x1_sg U60931 ( .A(n42480), .B(\mask_0/reg_ii_mask[2] ), .X(n27949) );
  nor_x1_sg U60932 ( .A(n42479), .B(\mask_0/reg_ii_mask[1] ), .X(n27944) );
  nor_x1_sg U60933 ( .A(n35566), .B(\mask_0/reg_ii_mask[0] ), .X(n27939) );
  nand_x1_sg U60934 ( .A(\mask_0/reg_ww_mask[31] ), .B(n35581), .X(n28253) );
  nand_x1_sg U60935 ( .A(\mask_0/reg_ww_mask[30] ), .B(n42494), .X(n28248) );
  nand_x1_sg U60936 ( .A(\mask_0/reg_ww_mask[29] ), .B(n42493), .X(n28243) );
  nand_x1_sg U60937 ( .A(\mask_0/reg_ww_mask[28] ), .B(n35580), .X(n28238) );
  nand_x1_sg U60938 ( .A(\mask_0/reg_ww_mask[27] ), .B(n42492), .X(n28233) );
  nand_x1_sg U60939 ( .A(\mask_0/reg_ww_mask[26] ), .B(n42491), .X(n28228) );
  nand_x1_sg U60940 ( .A(\mask_0/reg_ww_mask[25] ), .B(n35579), .X(n28223) );
  nand_x1_sg U60941 ( .A(\mask_0/reg_ww_mask[24] ), .B(n42490), .X(n28218) );
  nand_x1_sg U60942 ( .A(\mask_0/reg_ww_mask[23] ), .B(n35578), .X(n28213) );
  nand_x1_sg U60943 ( .A(\mask_0/reg_ww_mask[22] ), .B(n42489), .X(n28208) );
  nand_x1_sg U60944 ( .A(\mask_0/reg_ww_mask[21] ), .B(n42488), .X(n28203) );
  nand_x1_sg U60945 ( .A(\mask_0/reg_ww_mask[20] ), .B(n35577), .X(n28198) );
  nand_x1_sg U60946 ( .A(\mask_0/reg_ww_mask[19] ), .B(n35576), .X(n28193) );
  nand_x1_sg U60947 ( .A(\mask_0/reg_ww_mask[18] ), .B(n35575), .X(n28188) );
  nand_x1_sg U60948 ( .A(\mask_0/reg_ww_mask[17] ), .B(n42487), .X(n28183) );
  nand_x1_sg U60949 ( .A(\mask_0/reg_ww_mask[16] ), .B(n42486), .X(n28178) );
  nand_x1_sg U60950 ( .A(\mask_0/reg_ww_mask[15] ), .B(n35574), .X(n28173) );
  nand_x1_sg U60951 ( .A(\mask_0/reg_ww_mask[14] ), .B(n42485), .X(n28168) );
  nand_x1_sg U60952 ( .A(\mask_0/reg_ww_mask[13] ), .B(n42484), .X(n28163) );
  nand_x1_sg U60953 ( .A(\mask_0/reg_ww_mask[12] ), .B(n35573), .X(n28158) );
  nand_x1_sg U60954 ( .A(\mask_0/reg_ww_mask[11] ), .B(n42483), .X(n28153) );
  nand_x1_sg U60955 ( .A(\mask_0/reg_ww_mask[10] ), .B(n42482), .X(n28148) );
  nand_x1_sg U60956 ( .A(\mask_0/reg_ww_mask[9] ), .B(n35572), .X(n28143) );
  nand_x1_sg U60957 ( .A(\mask_0/reg_ww_mask[8] ), .B(n35571), .X(n28138) );
  nand_x1_sg U60958 ( .A(\mask_0/reg_ww_mask[7] ), .B(n35570), .X(n28133) );
  nand_x1_sg U60959 ( .A(\mask_0/reg_ww_mask[6] ), .B(n35569), .X(n28128) );
  nand_x1_sg U60960 ( .A(\mask_0/reg_ww_mask[5] ), .B(n42481), .X(n28123) );
  nand_x1_sg U60961 ( .A(\mask_0/reg_ww_mask[4] ), .B(n35568), .X(n28118) );
  nand_x1_sg U60962 ( .A(\mask_0/reg_ww_mask[3] ), .B(n35567), .X(n28113) );
  nand_x1_sg U60963 ( .A(\mask_0/reg_ww_mask[2] ), .B(n42480), .X(n28108) );
  nand_x1_sg U60964 ( .A(\mask_0/reg_ww_mask[1] ), .B(n42479), .X(n28103) );
  nand_x1_sg U60965 ( .A(\mask_0/reg_ww_mask[0] ), .B(n35566), .X(n28098) );
  nand_x1_sg U60966 ( .A(\mask_0/reg_ii_mask[31] ), .B(n35581), .X(n28093) );
  nand_x1_sg U60967 ( .A(\mask_0/reg_ii_mask[30] ), .B(n42494), .X(n28088) );
  nand_x1_sg U60968 ( .A(\mask_0/reg_ii_mask[29] ), .B(n42493), .X(n28083) );
  nand_x1_sg U60969 ( .A(\mask_0/reg_ii_mask[28] ), .B(n35580), .X(n28078) );
  nand_x1_sg U60970 ( .A(\mask_0/reg_ii_mask[27] ), .B(n42492), .X(n28073) );
  nand_x1_sg U60971 ( .A(\mask_0/reg_ii_mask[26] ), .B(n42491), .X(n28068) );
  nand_x1_sg U60972 ( .A(\mask_0/reg_ii_mask[25] ), .B(n35579), .X(n28063) );
  nand_x1_sg U60973 ( .A(\mask_0/reg_ii_mask[24] ), .B(n42490), .X(n28058) );
  nand_x1_sg U60974 ( .A(\mask_0/reg_ii_mask[23] ), .B(n35578), .X(n28053) );
  nand_x1_sg U60975 ( .A(\mask_0/reg_ii_mask[22] ), .B(n42489), .X(n28048) );
  nand_x1_sg U60976 ( .A(\mask_0/reg_ii_mask[21] ), .B(n42488), .X(n28043) );
  nand_x1_sg U60977 ( .A(\mask_0/reg_ii_mask[20] ), .B(n35577), .X(n28038) );
  nand_x1_sg U60978 ( .A(\mask_0/reg_ii_mask[19] ), .B(n35576), .X(n28033) );
  nand_x1_sg U60979 ( .A(\mask_0/reg_ii_mask[18] ), .B(n35575), .X(n28028) );
  nand_x1_sg U60980 ( .A(\mask_0/reg_ii_mask[17] ), .B(n42487), .X(n28023) );
  nand_x1_sg U60981 ( .A(\mask_0/reg_ii_mask[16] ), .B(n42486), .X(n28018) );
  nand_x1_sg U60982 ( .A(\mask_0/reg_ii_mask[15] ), .B(n35574), .X(n28013) );
  nand_x1_sg U60983 ( .A(\mask_0/reg_ii_mask[14] ), .B(n42485), .X(n28008) );
  nand_x1_sg U60984 ( .A(\mask_0/reg_ii_mask[13] ), .B(n42484), .X(n28003) );
  nand_x1_sg U60985 ( .A(\mask_0/reg_ii_mask[12] ), .B(n35573), .X(n27998) );
  nand_x1_sg U60986 ( .A(\mask_0/reg_ii_mask[11] ), .B(n42483), .X(n27993) );
  nand_x1_sg U60987 ( .A(\mask_0/reg_ii_mask[10] ), .B(n42482), .X(n27988) );
  nand_x1_sg U60988 ( .A(\mask_0/reg_ii_mask[9] ), .B(n35572), .X(n27983) );
  nand_x1_sg U60989 ( .A(\mask_0/reg_ii_mask[8] ), .B(n35571), .X(n27978) );
  nand_x1_sg U60990 ( .A(\mask_0/reg_ii_mask[7] ), .B(n35570), .X(n27973) );
  nand_x1_sg U60991 ( .A(\mask_0/reg_ii_mask[6] ), .B(n35569), .X(n27968) );
  nand_x1_sg U60992 ( .A(\mask_0/reg_ii_mask[5] ), .B(n42481), .X(n27963) );
  nand_x1_sg U60993 ( .A(\mask_0/reg_ii_mask[4] ), .B(n35568), .X(n27958) );
  nand_x1_sg U60994 ( .A(\mask_0/reg_ii_mask[3] ), .B(n35567), .X(n27953) );
  nand_x1_sg U60995 ( .A(\mask_0/reg_ii_mask[2] ), .B(n42480), .X(n27948) );
  nand_x1_sg U60996 ( .A(\mask_0/reg_ii_mask[1] ), .B(n42479), .X(n27943) );
  nand_x1_sg U60997 ( .A(\mask_0/reg_ii_mask[0] ), .B(n35566), .X(n27938) );
  inv_x1_sg U60998 ( .A(\mask_0/counter[0] ), .X(n42530) );
  nand_x1_sg U60999 ( .A(\mask_0/reg_i_mask[31] ), .B(\mask_0/reg_w_mask[31] ), 
        .X(n26351) );
  nand_x1_sg U61000 ( .A(\mask_0/reg_i_mask[30] ), .B(\mask_0/reg_w_mask[30] ), 
        .X(n26355) );
  nand_x1_sg U61001 ( .A(\mask_0/reg_i_mask[29] ), .B(\mask_0/reg_w_mask[29] ), 
        .X(n26358) );
  nand_x1_sg U61002 ( .A(\mask_0/reg_i_mask[28] ), .B(\mask_0/reg_w_mask[28] ), 
        .X(n26361) );
  nand_x1_sg U61003 ( .A(\mask_0/reg_i_mask[27] ), .B(\mask_0/reg_w_mask[27] ), 
        .X(n26364) );
  nand_x1_sg U61004 ( .A(\mask_0/reg_i_mask[26] ), .B(\mask_0/reg_w_mask[26] ), 
        .X(n26367) );
  nand_x1_sg U61005 ( .A(\mask_0/reg_i_mask[25] ), .B(\mask_0/reg_w_mask[25] ), 
        .X(n26370) );
  nand_x1_sg U61006 ( .A(\mask_0/reg_i_mask[24] ), .B(\mask_0/reg_w_mask[24] ), 
        .X(n26373) );
  nand_x1_sg U61007 ( .A(\mask_0/reg_i_mask[23] ), .B(\mask_0/reg_w_mask[23] ), 
        .X(n26376) );
  nand_x1_sg U61008 ( .A(\mask_0/reg_i_mask[22] ), .B(\mask_0/reg_w_mask[22] ), 
        .X(n26379) );
  nand_x1_sg U61009 ( .A(\mask_0/reg_i_mask[21] ), .B(\mask_0/reg_w_mask[21] ), 
        .X(n26382) );
  nand_x1_sg U61010 ( .A(\mask_0/reg_i_mask[20] ), .B(\mask_0/reg_w_mask[20] ), 
        .X(n26385) );
  nand_x1_sg U61011 ( .A(\mask_0/reg_i_mask[19] ), .B(\mask_0/reg_w_mask[19] ), 
        .X(n26388) );
  nand_x1_sg U61012 ( .A(\mask_0/reg_i_mask[18] ), .B(\mask_0/reg_w_mask[18] ), 
        .X(n26391) );
  nand_x1_sg U61013 ( .A(\mask_0/reg_i_mask[17] ), .B(\mask_0/reg_w_mask[17] ), 
        .X(n26394) );
  nand_x1_sg U61014 ( .A(\mask_0/reg_i_mask[16] ), .B(\mask_0/reg_w_mask[16] ), 
        .X(n26397) );
  nand_x1_sg U61015 ( .A(\mask_0/reg_i_mask[15] ), .B(\mask_0/reg_w_mask[15] ), 
        .X(n26400) );
  nand_x1_sg U61016 ( .A(\mask_0/reg_i_mask[14] ), .B(\mask_0/reg_w_mask[14] ), 
        .X(n26403) );
  nand_x1_sg U61017 ( .A(\mask_0/reg_i_mask[13] ), .B(\mask_0/reg_w_mask[13] ), 
        .X(n26406) );
  nand_x1_sg U61018 ( .A(\mask_0/reg_i_mask[12] ), .B(\mask_0/reg_w_mask[12] ), 
        .X(n26409) );
  nand_x1_sg U61019 ( .A(\mask_0/reg_i_mask[11] ), .B(\mask_0/reg_w_mask[11] ), 
        .X(n26412) );
  nand_x1_sg U61020 ( .A(\mask_0/reg_i_mask[10] ), .B(\mask_0/reg_w_mask[10] ), 
        .X(n26415) );
  nand_x1_sg U61021 ( .A(\mask_0/reg_i_mask[9] ), .B(\mask_0/reg_w_mask[9] ), 
        .X(n26418) );
  nand_x1_sg U61022 ( .A(\mask_0/reg_i_mask[8] ), .B(\mask_0/reg_w_mask[8] ), 
        .X(n26421) );
  nand_x1_sg U61023 ( .A(\mask_0/reg_i_mask[7] ), .B(\mask_0/reg_w_mask[7] ), 
        .X(n26424) );
  nand_x1_sg U61024 ( .A(\mask_0/reg_i_mask[6] ), .B(\mask_0/reg_w_mask[6] ), 
        .X(n26427) );
  nand_x1_sg U61025 ( .A(\mask_0/reg_i_mask[5] ), .B(\mask_0/reg_w_mask[5] ), 
        .X(n26430) );
  nand_x1_sg U61026 ( .A(\mask_0/reg_i_mask[4] ), .B(\mask_0/reg_w_mask[4] ), 
        .X(n26433) );
  nand_x1_sg U61027 ( .A(\mask_0/reg_i_mask[3] ), .B(\mask_0/reg_w_mask[3] ), 
        .X(n26436) );
  nand_x1_sg U61028 ( .A(\mask_0/reg_i_mask[2] ), .B(\mask_0/reg_w_mask[2] ), 
        .X(n26439) );
  nand_x1_sg U61029 ( .A(\mask_0/reg_i_mask[1] ), .B(\mask_0/reg_w_mask[1] ), 
        .X(n26442) );
  nand_x1_sg U61030 ( .A(\mask_0/reg_i_mask[0] ), .B(\mask_0/reg_w_mask[0] ), 
        .X(n26445) );
  nor_x1_sg U61031 ( .A(n31659), .B(n31707), .X(n11609) );
  nor_x1_sg U61032 ( .A(n31597), .B(n31595), .X(n11639) );
  nor_x1_sg U61033 ( .A(n31658), .B(n35305), .X(n15189) );
  nor_x1_sg U61034 ( .A(n35097), .B(n35257), .X(n15065) );
  nor_x1_sg U61035 ( .A(n31597), .B(n35102), .X(n13611) );
  nor_x1_sg U61036 ( .A(n41044), .B(n34545), .X(n12948) );
  nor_x1_sg U61037 ( .A(n14953), .B(n14954), .X(n14952) );
  nor_x1_sg U61038 ( .A(\shifter_0/reg_i_6[17] ), .B(n32894), .X(n14953) );
  nor_x1_sg U61039 ( .A(n40928), .B(n34544), .X(n12794) );
  nor_x1_sg U61040 ( .A(n14205), .B(n14206), .X(n14204) );
  nor_x1_sg U61041 ( .A(\shifter_0/reg_w_6[13] ), .B(n32893), .X(n14205) );
  nor_x1_sg U61042 ( .A(n40924), .B(n32054), .X(n12806) );
  nor_x1_sg U61043 ( .A(n14267), .B(n14268), .X(n14266) );
  nor_x1_sg U61044 ( .A(\shifter_0/reg_w_6[15] ), .B(n34855), .X(n14267) );
  nor_x1_sg U61045 ( .A(n40921), .B(n35416), .X(n12818) );
  nor_x1_sg U61046 ( .A(n14329), .B(n14330), .X(n14328) );
  nor_x1_sg U61047 ( .A(\shifter_0/reg_w_6[17] ), .B(n30200), .X(n14329) );
  nor_x1_sg U61048 ( .A(n40918), .B(n31302), .X(n12830) );
  nor_x1_sg U61049 ( .A(n14391), .B(n14392), .X(n14390) );
  nor_x1_sg U61050 ( .A(\shifter_0/reg_w_6[19] ), .B(n32899), .X(n14391) );
  nor_x1_sg U61051 ( .A(n41069), .B(n34545), .X(n12852) );
  nor_x1_sg U61052 ( .A(n14454), .B(n14455), .X(n14453) );
  nor_x1_sg U61053 ( .A(\shifter_0/reg_i_6[1] ), .B(n32899), .X(n14454) );
  nor_x1_sg U61054 ( .A(n41066), .B(n30137), .X(n12864) );
  nor_x1_sg U61055 ( .A(n14518), .B(n14519), .X(n14517) );
  nor_x1_sg U61056 ( .A(\shifter_0/reg_i_6[3] ), .B(n32897), .X(n14518) );
  nor_x1_sg U61057 ( .A(n41063), .B(n32058), .X(n12876) );
  nor_x1_sg U61058 ( .A(n14580), .B(n14581), .X(n14579) );
  nor_x1_sg U61059 ( .A(\shifter_0/reg_i_6[5] ), .B(n32929), .X(n14580) );
  nor_x1_sg U61060 ( .A(n41059), .B(n34546), .X(n12888) );
  nor_x1_sg U61061 ( .A(n14642), .B(n14643), .X(n14641) );
  nor_x1_sg U61062 ( .A(\shifter_0/reg_i_6[7] ), .B(n34854), .X(n14642) );
  nor_x1_sg U61063 ( .A(n41057), .B(n32056), .X(n12900) );
  nor_x1_sg U61064 ( .A(n14704), .B(n14705), .X(n14703) );
  nor_x1_sg U61065 ( .A(\shifter_0/reg_i_6[9] ), .B(n34856), .X(n14704) );
  nor_x1_sg U61066 ( .A(n41053), .B(n29750), .X(n12912) );
  nor_x1_sg U61067 ( .A(n14766), .B(n14767), .X(n14765) );
  nor_x1_sg U61068 ( .A(\shifter_0/reg_i_6[11] ), .B(n34858), .X(n14766) );
  nor_x1_sg U61069 ( .A(n41051), .B(n31302), .X(n12924) );
  nor_x1_sg U61070 ( .A(n14828), .B(n14829), .X(n14827) );
  nor_x1_sg U61071 ( .A(\shifter_0/reg_i_6[13] ), .B(n32899), .X(n14828) );
  nor_x1_sg U61072 ( .A(n41047), .B(n32054), .X(n12936) );
  nor_x1_sg U61073 ( .A(n14890), .B(n14891), .X(n14889) );
  nor_x1_sg U61074 ( .A(\shifter_0/reg_i_6[15] ), .B(n32898), .X(n14890) );
  nor_x1_sg U61075 ( .A(\shifter_0/reg_i_7[4] ), .B(n30967), .X(n14551) );
  nor_x1_sg U61076 ( .A(\shifter_0/reg_w_7[6] ), .B(n33836), .X(n13989) );
  nor_x1_sg U61077 ( .A(\shifter_0/reg_w_7[7] ), .B(n33833), .X(n14020) );
  nor_x1_sg U61078 ( .A(\shifter_0/reg_w_7[8] ), .B(n33833), .X(n14051) );
  nor_x1_sg U61079 ( .A(\shifter_0/reg_w_7[9] ), .B(n33837), .X(n14082) );
  nor_x1_sg U61080 ( .A(\shifter_0/reg_w_7[10] ), .B(n30963), .X(n14113) );
  nor_x1_sg U61081 ( .A(\shifter_0/reg_w_7[11] ), .B(n33837), .X(n14144) );
  nor_x1_sg U61082 ( .A(\shifter_0/reg_w_7[12] ), .B(n33832), .X(n14175) );
  nor_x1_sg U61083 ( .A(\shifter_0/reg_w_7[13] ), .B(n33837), .X(n14206) );
  nor_x1_sg U61084 ( .A(\shifter_0/reg_w_7[14] ), .B(n34808), .X(n14237) );
  nor_x1_sg U61085 ( .A(\shifter_0/reg_w_7[15] ), .B(n30638), .X(n14268) );
  nor_x1_sg U61086 ( .A(\shifter_0/reg_w_7[16] ), .B(n32925), .X(n14299) );
  nor_x1_sg U61087 ( .A(\shifter_0/reg_w_7[17] ), .B(n34861), .X(n14330) );
  nor_x1_sg U61088 ( .A(\shifter_0/reg_w_7[18] ), .B(n34861), .X(n14361) );
  nor_x1_sg U61089 ( .A(\shifter_0/reg_w_7[19] ), .B(n33834), .X(n14392) );
  nor_x1_sg U61090 ( .A(n31126), .B(n33832), .X(n14424) );
  nor_x1_sg U61091 ( .A(n31128), .B(n33831), .X(n14455) );
  nor_x1_sg U61092 ( .A(n31130), .B(n33834), .X(n14519) );
  nor_x1_sg U61093 ( .A(n31133), .B(n33838), .X(n14581) );
  nor_x1_sg U61094 ( .A(\shifter_0/reg_i_7[6] ), .B(n33832), .X(n14612) );
  nor_x1_sg U61095 ( .A(n31137), .B(n33831), .X(n14643) );
  nor_x1_sg U61096 ( .A(n31139), .B(n33832), .X(n14674) );
  nor_x1_sg U61097 ( .A(n31141), .B(n30964), .X(n14705) );
  nor_x1_sg U61098 ( .A(\shifter_0/reg_i_7[10] ), .B(n30964), .X(n14736) );
  nor_x1_sg U61099 ( .A(n31145), .B(n34806), .X(n14767) );
  nor_x1_sg U61100 ( .A(n31147), .B(n32926), .X(n14798) );
  nor_x1_sg U61101 ( .A(n31149), .B(n32925), .X(n14829) );
  nor_x1_sg U61102 ( .A(\shifter_0/reg_i_7[14] ), .B(n30963), .X(n14860) );
  nor_x1_sg U61103 ( .A(\shifter_0/reg_i_7[15] ), .B(n33838), .X(n14891) );
  nor_x1_sg U61104 ( .A(\shifter_0/reg_i_7[16] ), .B(n34859), .X(n14922) );
  nor_x1_sg U61105 ( .A(n31157), .B(n33829), .X(n15015) );
  nor_x1_sg U61106 ( .A(\shifter_0/reg_w_7[0] ), .B(n34808), .X(n13797) );
  nor_x1_sg U61107 ( .A(\shifter_0/reg_w_7[1] ), .B(n33839), .X(n13834) );
  nor_x1_sg U61108 ( .A(\shifter_0/reg_w_7[2] ), .B(n34860), .X(n13865) );
  nor_x1_sg U61109 ( .A(\shifter_0/reg_w_7[3] ), .B(n34861), .X(n13896) );
  nor_x1_sg U61110 ( .A(n31169), .B(n30965), .X(n13927) );
  nor_x1_sg U61111 ( .A(\shifter_0/reg_w_7[5] ), .B(n34808), .X(n13958) );
  nor_x1_sg U61112 ( .A(n31655), .B(n33966), .X(\filter_0/n6285 ) );
  nor_x1_sg U61113 ( .A(\shifter_0/reg_w_3[0] ), .B(n33837), .X(n13790) );
  nor_x1_sg U61114 ( .A(\shifter_0/reg_w_3[1] ), .B(n34807), .X(n13827) );
  nor_x1_sg U61115 ( .A(\shifter_0/reg_w_3[2] ), .B(n34807), .X(n13858) );
  nor_x1_sg U61116 ( .A(\shifter_0/reg_w_3[5] ), .B(n33833), .X(n13951) );
  nor_x1_sg U61117 ( .A(\shifter_0/reg_w_3[6] ), .B(n34860), .X(n13982) );
  nor_x1_sg U61118 ( .A(\shifter_0/reg_w_3[7] ), .B(n34806), .X(n14013) );
  nor_x1_sg U61119 ( .A(\shifter_0/reg_w_3[10] ), .B(n32926), .X(n14106) );
  nor_x1_sg U61120 ( .A(\shifter_0/reg_w_3[11] ), .B(n32925), .X(n14137) );
  nor_x1_sg U61121 ( .A(\shifter_0/reg_w_3[14] ), .B(n33831), .X(n14230) );
  nor_x1_sg U61122 ( .A(\shifter_0/reg_w_3[15] ), .B(n34859), .X(n14261) );
  nor_x1_sg U61123 ( .A(\shifter_0/reg_w_3[16] ), .B(n33836), .X(n14292) );
  nor_x1_sg U61124 ( .A(\shifter_0/reg_w_3[19] ), .B(n34808), .X(n14385) );
  nor_x1_sg U61125 ( .A(\shifter_0/reg_i_3[0] ), .B(n30967), .X(n14417) );
  nor_x1_sg U61126 ( .A(\shifter_0/reg_i_3[1] ), .B(n30199), .X(n14448) );
  nor_x1_sg U61127 ( .A(\shifter_0/reg_i_3[2] ), .B(n34807), .X(n14480) );
  nor_x1_sg U61128 ( .A(\shifter_0/reg_i_3[5] ), .B(n33834), .X(n14574) );
  nor_x1_sg U61129 ( .A(\shifter_0/reg_i_3[6] ), .B(n30638), .X(n14605) );
  nor_x1_sg U61130 ( .A(\shifter_0/reg_i_3[7] ), .B(n34806), .X(n14636) );
  nor_x1_sg U61131 ( .A(\shifter_0/reg_i_3[10] ), .B(n34860), .X(n14729) );
  nor_x1_sg U61132 ( .A(\shifter_0/reg_i_3[11] ), .B(n30638), .X(n14760) );
  nor_x1_sg U61133 ( .A(\shifter_0/reg_i_3[14] ), .B(n33836), .X(n14853) );
  nor_x1_sg U61134 ( .A(\shifter_0/reg_i_3[15] ), .B(n30963), .X(n14884) );
  nor_x1_sg U61135 ( .A(\shifter_0/reg_i_3[16] ), .B(n30638), .X(n14915) );
  nor_x1_sg U61136 ( .A(\shifter_0/reg_i_3[19] ), .B(n33828), .X(n15008) );
  nor_x1_sg U61137 ( .A(n30468), .B(n31694), .X(n13810) );
  nor_x1_sg U61138 ( .A(n30470), .B(n31049), .X(n13844) );
  nor_x1_sg U61139 ( .A(n30472), .B(n33991), .X(n13875) );
  nor_x1_sg U61140 ( .A(n30474), .B(n33990), .X(n13906) );
  nor_x1_sg U61141 ( .A(n30476), .B(n33990), .X(n13937) );
  nor_x1_sg U61142 ( .A(n30478), .B(n31694), .X(n13968) );
  nor_x1_sg U61143 ( .A(n30480), .B(n29704), .X(n13999) );
  nor_x1_sg U61144 ( .A(n30482), .B(n35414), .X(n14030) );
  nor_x1_sg U61145 ( .A(n30484), .B(n33991), .X(n14061) );
  nor_x1_sg U61146 ( .A(n30486), .B(n30021), .X(n14092) );
  nor_x1_sg U61147 ( .A(n30488), .B(n31048), .X(n14123) );
  nor_x1_sg U61148 ( .A(n30490), .B(n30021), .X(n14154) );
  nor_x1_sg U61149 ( .A(n30492), .B(n29704), .X(n14185) );
  nor_x1_sg U61150 ( .A(\shifter_0/reg_w_8[13] ), .B(n33989), .X(n14216) );
  nor_x1_sg U61151 ( .A(\shifter_0/reg_w_8[14] ), .B(n33991), .X(n14247) );
  nor_x1_sg U61152 ( .A(n30498), .B(n31049), .X(n14278) );
  nor_x1_sg U61153 ( .A(n30500), .B(n30530), .X(n14309) );
  nor_x1_sg U61154 ( .A(n30502), .B(n30530), .X(n14340) );
  nor_x1_sg U61155 ( .A(n30504), .B(n31048), .X(n14371) );
  nor_x1_sg U61156 ( .A(n30506), .B(n31694), .X(n14402) );
  nor_x1_sg U61157 ( .A(n30406), .B(n31048), .X(n14434) );
  nor_x1_sg U61158 ( .A(n30408), .B(n31049), .X(n14465) );
  nor_x1_sg U61159 ( .A(n30412), .B(n33989), .X(n14529) );
  nor_x1_sg U61160 ( .A(n30416), .B(n29704), .X(n14591) );
  nor_x1_sg U61161 ( .A(\shifter_0/reg_i_8[6] ), .B(n30530), .X(n14622) );
  nor_x1_sg U61162 ( .A(n30420), .B(n29704), .X(n14653) );
  nor_x1_sg U61163 ( .A(n30422), .B(n35414), .X(n14684) );
  nor_x1_sg U61164 ( .A(n30424), .B(n30021), .X(n14715) );
  nor_x1_sg U61165 ( .A(\shifter_0/reg_i_8[10] ), .B(n33990), .X(n14746) );
  nor_x1_sg U61166 ( .A(n30428), .B(n33991), .X(n14777) );
  nor_x1_sg U61167 ( .A(n30430), .B(n33989), .X(n14808) );
  nor_x1_sg U61168 ( .A(n30432), .B(n31694), .X(n14839) );
  nor_x1_sg U61169 ( .A(\shifter_0/reg_i_8[14] ), .B(n31048), .X(n14870) );
  nor_x1_sg U61170 ( .A(\shifter_0/reg_i_8[15] ), .B(n33989), .X(n14901) );
  nor_x1_sg U61171 ( .A(\shifter_0/reg_i_8[16] ), .B(n31049), .X(n14932) );
  nor_x1_sg U61172 ( .A(n30444), .B(n33990), .X(n15025) );
  nor_x1_sg U61173 ( .A(\shifter_0/reg_i_7[2] ), .B(n33838), .X(n14487) );
  nor_x1_sg U61174 ( .A(\shifter_0/reg_i_7[17] ), .B(n30968), .X(n14954) );
  nor_x1_sg U61175 ( .A(\shifter_0/reg_i_7[18] ), .B(n32926), .X(n14985) );
  nor_x1_sg U61176 ( .A(\shifter_0/reg_w_2[0] ), .B(n32929), .X(n13789) );
  nor_x1_sg U61177 ( .A(\shifter_0/reg_w_2[1] ), .B(n32896), .X(n13826) );
  nor_x1_sg U61178 ( .A(\shifter_0/reg_w_2[2] ), .B(n32897), .X(n13857) );
  nor_x1_sg U61179 ( .A(\shifter_0/reg_w_2[5] ), .B(n29771), .X(n13950) );
  nor_x1_sg U61180 ( .A(\shifter_0/reg_w_2[6] ), .B(n30200), .X(n13981) );
  nor_x1_sg U61181 ( .A(\shifter_0/reg_w_2[7] ), .B(n34854), .X(n14012) );
  nor_x1_sg U61182 ( .A(\shifter_0/reg_w_2[10] ), .B(n30636), .X(n14105) );
  nor_x1_sg U61183 ( .A(\shifter_0/reg_w_2[11] ), .B(n32896), .X(n14136) );
  nor_x1_sg U61184 ( .A(\shifter_0/reg_w_2[14] ), .B(n32931), .X(n14229) );
  nor_x1_sg U61185 ( .A(\shifter_0/reg_w_2[15] ), .B(n32891), .X(n14260) );
  nor_x1_sg U61186 ( .A(\shifter_0/reg_w_2[16] ), .B(n32930), .X(n14291) );
  nor_x1_sg U61187 ( .A(\shifter_0/reg_w_2[19] ), .B(n30636), .X(n14384) );
  nor_x1_sg U61188 ( .A(\shifter_0/reg_i_2[0] ), .B(n32892), .X(n14416) );
  nor_x1_sg U61189 ( .A(\shifter_0/reg_i_2[1] ), .B(n32888), .X(n14447) );
  nor_x1_sg U61190 ( .A(\shifter_0/reg_i_2[2] ), .B(n30635), .X(n14479) );
  nor_x1_sg U61191 ( .A(\shifter_0/reg_i_2[5] ), .B(n32930), .X(n14573) );
  nor_x1_sg U61192 ( .A(\shifter_0/reg_i_2[6] ), .B(n32889), .X(n14604) );
  nor_x1_sg U61193 ( .A(\shifter_0/reg_i_2[7] ), .B(n30200), .X(n14635) );
  nor_x1_sg U61194 ( .A(\shifter_0/reg_i_2[10] ), .B(n32931), .X(n14728) );
  nor_x1_sg U61195 ( .A(\shifter_0/reg_i_2[11] ), .B(n34857), .X(n14759) );
  nor_x1_sg U61196 ( .A(\shifter_0/reg_i_2[14] ), .B(n32891), .X(n14852) );
  nor_x1_sg U61197 ( .A(\shifter_0/reg_i_2[15] ), .B(n32892), .X(n14883) );
  nor_x1_sg U61198 ( .A(\shifter_0/reg_i_2[16] ), .B(n34855), .X(n14914) );
  nor_x1_sg U61199 ( .A(\shifter_0/reg_i_2[19] ), .B(n32892), .X(n15007) );
  nor_x1_sg U61200 ( .A(\shifter_0/reg_w_3[3] ), .B(n33839), .X(n13889) );
  nor_x1_sg U61201 ( .A(\shifter_0/reg_w_3[4] ), .B(n34859), .X(n13920) );
  nor_x1_sg U61202 ( .A(\shifter_0/reg_w_3[8] ), .B(n33839), .X(n14044) );
  nor_x1_sg U61203 ( .A(\shifter_0/reg_w_3[9] ), .B(n30968), .X(n14075) );
  nor_x1_sg U61204 ( .A(\shifter_0/reg_w_3[12] ), .B(n30964), .X(n14168) );
  nor_x1_sg U61205 ( .A(\shifter_0/reg_w_3[13] ), .B(n33838), .X(n14199) );
  nor_x1_sg U61206 ( .A(\shifter_0/reg_w_3[17] ), .B(n30963), .X(n14323) );
  nor_x1_sg U61207 ( .A(\shifter_0/reg_w_3[18] ), .B(n34807), .X(n14354) );
  nor_x1_sg U61208 ( .A(\shifter_0/reg_i_3[3] ), .B(n33834), .X(n14512) );
  nor_x1_sg U61209 ( .A(\shifter_0/reg_i_3[4] ), .B(n30967), .X(n14544) );
  nor_x1_sg U61210 ( .A(\shifter_0/reg_i_3[8] ), .B(n33829), .X(n14667) );
  nor_x1_sg U61211 ( .A(\shifter_0/reg_i_3[9] ), .B(n30967), .X(n14698) );
  nor_x1_sg U61212 ( .A(\shifter_0/reg_i_3[12] ), .B(n33831), .X(n14791) );
  nor_x1_sg U61213 ( .A(\shifter_0/reg_i_3[13] ), .B(n30968), .X(n14822) );
  nor_x1_sg U61214 ( .A(\shifter_0/reg_i_3[17] ), .B(n33829), .X(n14947) );
  nor_x1_sg U61215 ( .A(\shifter_0/reg_i_3[18] ), .B(n33828), .X(n14978) );
  nor_x1_sg U61216 ( .A(n41067), .B(n32057), .X(n12858) );
  nor_x1_sg U61217 ( .A(n14486), .B(n14487), .X(n14485) );
  nor_x1_sg U61218 ( .A(\shifter_0/reg_i_6[2] ), .B(n32898), .X(n14486) );
  nor_x1_sg U61219 ( .A(n41065), .B(n31303), .X(n12870) );
  nor_x1_sg U61220 ( .A(n14550), .B(n14551), .X(n14549) );
  nor_x1_sg U61221 ( .A(\shifter_0/reg_i_6[4] ), .B(n32930), .X(n14550) );
  nor_x1_sg U61222 ( .A(n41043), .B(n34546), .X(n12954) );
  nor_x1_sg U61223 ( .A(n14984), .B(n14985), .X(n14983) );
  nor_x1_sg U61224 ( .A(\shifter_0/reg_i_6[18] ), .B(n32897), .X(n14984) );
  nor_x1_sg U61225 ( .A(n40938), .B(n31302), .X(n12752) );
  nor_x1_sg U61226 ( .A(n13988), .B(n13989), .X(n13987) );
  nor_x1_sg U61227 ( .A(\shifter_0/reg_w_6[6] ), .B(n30962), .X(n13988) );
  nor_x1_sg U61228 ( .A(n40936), .B(n34544), .X(n12758) );
  nor_x1_sg U61229 ( .A(n14019), .B(n14020), .X(n14018) );
  nor_x1_sg U61230 ( .A(\shifter_0/reg_w_6[7] ), .B(n32898), .X(n14019) );
  nor_x1_sg U61231 ( .A(n40935), .B(n32053), .X(n12764) );
  nor_x1_sg U61232 ( .A(n14050), .B(n14051), .X(n14049) );
  nor_x1_sg U61233 ( .A(\shifter_0/reg_w_6[8] ), .B(n32893), .X(n14050) );
  nor_x1_sg U61234 ( .A(n40934), .B(n32057), .X(n12770) );
  nor_x1_sg U61235 ( .A(n14081), .B(n14082), .X(n14080) );
  nor_x1_sg U61236 ( .A(\shifter_0/reg_w_6[9] ), .B(n32894), .X(n14081) );
  nor_x1_sg U61237 ( .A(n40932), .B(n34544), .X(n12776) );
  nor_x1_sg U61238 ( .A(n14112), .B(n14113), .X(n14111) );
  nor_x1_sg U61239 ( .A(\shifter_0/reg_w_6[10] ), .B(n34856), .X(n14112) );
  nor_x1_sg U61240 ( .A(n40930), .B(n32057), .X(n12782) );
  nor_x1_sg U61241 ( .A(n14143), .B(n14144), .X(n14142) );
  nor_x1_sg U61242 ( .A(\shifter_0/reg_w_6[11] ), .B(n32897), .X(n14143) );
  nor_x1_sg U61243 ( .A(n40929), .B(n31302), .X(n12788) );
  nor_x1_sg U61244 ( .A(n14174), .B(n14175), .X(n14173) );
  nor_x1_sg U61245 ( .A(\shifter_0/reg_w_6[12] ), .B(n32928), .X(n14174) );
  nor_x1_sg U61246 ( .A(n40926), .B(n32053), .X(n12800) );
  nor_x1_sg U61247 ( .A(n14236), .B(n14237), .X(n14235) );
  nor_x1_sg U61248 ( .A(\shifter_0/reg_w_6[14] ), .B(n34856), .X(n14236) );
  nor_x1_sg U61249 ( .A(n40922), .B(n30137), .X(n12812) );
  nor_x1_sg U61250 ( .A(n14298), .B(n14299), .X(n14297) );
  nor_x1_sg U61251 ( .A(\shifter_0/reg_w_6[16] ), .B(n32928), .X(n14298) );
  nor_x1_sg U61252 ( .A(n40920), .B(n34546), .X(n12824) );
  nor_x1_sg U61253 ( .A(n14360), .B(n14361), .X(n14359) );
  nor_x1_sg U61254 ( .A(\shifter_0/reg_w_6[18] ), .B(n32888), .X(n14360) );
  nor_x1_sg U61255 ( .A(n41071), .B(n30137), .X(n12846) );
  nor_x1_sg U61256 ( .A(n14423), .B(n14424), .X(n14422) );
  nor_x1_sg U61257 ( .A(\shifter_0/reg_i_6[0] ), .B(n32930), .X(n14423) );
  nor_x1_sg U61258 ( .A(n41061), .B(n32058), .X(n12882) );
  nor_x1_sg U61259 ( .A(n14611), .B(n14612), .X(n14610) );
  nor_x1_sg U61260 ( .A(\shifter_0/reg_i_6[6] ), .B(n30636), .X(n14611) );
  nor_x1_sg U61261 ( .A(n41058), .B(n35416), .X(n12894) );
  nor_x1_sg U61262 ( .A(n14673), .B(n14674), .X(n14672) );
  nor_x1_sg U61263 ( .A(\shifter_0/reg_i_6[8] ), .B(n32931), .X(n14673) );
  nor_x1_sg U61264 ( .A(n41055), .B(n32056), .X(n12906) );
  nor_x1_sg U61265 ( .A(n14735), .B(n14736), .X(n14734) );
  nor_x1_sg U61266 ( .A(\shifter_0/reg_i_6[10] ), .B(n32929), .X(n14735) );
  nor_x1_sg U61267 ( .A(n41052), .B(n31303), .X(n12918) );
  nor_x1_sg U61268 ( .A(n14797), .B(n14798), .X(n14796) );
  nor_x1_sg U61269 ( .A(\shifter_0/reg_i_6[12] ), .B(n32898), .X(n14797) );
  nor_x1_sg U61270 ( .A(n41049), .B(n32054), .X(n12930) );
  nor_x1_sg U61271 ( .A(n14859), .B(n14860), .X(n14858) );
  nor_x1_sg U61272 ( .A(\shifter_0/reg_i_6[14] ), .B(n32888), .X(n14859) );
  nor_x1_sg U61273 ( .A(n41045), .B(n32058), .X(n12942) );
  nor_x1_sg U61274 ( .A(n14921), .B(n14922), .X(n14920) );
  nor_x1_sg U61275 ( .A(\shifter_0/reg_i_6[16] ), .B(n34857), .X(n14921) );
  nor_x1_sg U61276 ( .A(n41041), .B(n31303), .X(n12960) );
  nor_x1_sg U61277 ( .A(n15014), .B(n15015), .X(n15013) );
  nor_x1_sg U61278 ( .A(\shifter_0/reg_i_6[19] ), .B(n32892), .X(n15014) );
  nor_x1_sg U61279 ( .A(n40948), .B(n34544), .X(n12715) );
  nor_x1_sg U61280 ( .A(n13796), .B(n13797), .X(n13795) );
  nor_x1_sg U61281 ( .A(\shifter_0/reg_w_6[0] ), .B(n32928), .X(n13796) );
  nor_x1_sg U61282 ( .A(n40946), .B(n34545), .X(n12722) );
  nor_x1_sg U61283 ( .A(n13833), .B(n13834), .X(n13832) );
  nor_x1_sg U61284 ( .A(\shifter_0/reg_w_6[1] ), .B(n32928), .X(n13833) );
  nor_x1_sg U61285 ( .A(n40944), .B(n32053), .X(n12728) );
  nor_x1_sg U61286 ( .A(n13864), .B(n13865), .X(n13863) );
  nor_x1_sg U61287 ( .A(\shifter_0/reg_w_6[2] ), .B(n32888), .X(n13864) );
  nor_x1_sg U61288 ( .A(n40943), .B(n32056), .X(n12734) );
  nor_x1_sg U61289 ( .A(n13895), .B(n13896), .X(n13894) );
  nor_x1_sg U61290 ( .A(\shifter_0/reg_w_6[3] ), .B(n30639), .X(n13895) );
  nor_x1_sg U61291 ( .A(n40942), .B(n32057), .X(n12740) );
  nor_x1_sg U61292 ( .A(n13926), .B(n13927), .X(n13925) );
  nor_x1_sg U61293 ( .A(\shifter_0/reg_w_6[4] ), .B(n32894), .X(n13926) );
  nor_x1_sg U61294 ( .A(n40940), .B(n34546), .X(n12746) );
  nor_x1_sg U61295 ( .A(n13957), .B(n13958), .X(n13956) );
  nor_x1_sg U61296 ( .A(\shifter_0/reg_w_6[5] ), .B(n32931), .X(n13957) );
  nor_x1_sg U61297 ( .A(\shifter_0/reg_w_10[0] ), .B(n33993), .X(n13809) );
  nor_x1_sg U61298 ( .A(\shifter_0/reg_w_10[1] ), .B(n31051), .X(n13843) );
  nor_x1_sg U61299 ( .A(\shifter_0/reg_w_10[2] ), .B(n33993), .X(n13874) );
  nor_x1_sg U61300 ( .A(\shifter_0/reg_w_10[5] ), .B(n33993), .X(n13967) );
  nor_x1_sg U61301 ( .A(\shifter_0/reg_w_10[6] ), .B(n31051), .X(n13998) );
  nor_x1_sg U61302 ( .A(\shifter_0/reg_w_10[7] ), .B(n31052), .X(n14029) );
  nor_x1_sg U61303 ( .A(\shifter_0/reg_w_10[8] ), .B(n30022), .X(n14060) );
  nor_x1_sg U61304 ( .A(\shifter_0/reg_w_10[9] ), .B(n30532), .X(n14091) );
  nor_x1_sg U61305 ( .A(\shifter_0/reg_w_10[10] ), .B(n33993), .X(n14122) );
  nor_x1_sg U61306 ( .A(\shifter_0/reg_w_10[11] ), .B(n31693), .X(n14153) );
  nor_x1_sg U61307 ( .A(\shifter_0/reg_w_10[12] ), .B(n33994), .X(n14184) );
  nor_x1_sg U61308 ( .A(\shifter_0/reg_w_10[13] ), .B(n33994), .X(n14215) );
  nor_x1_sg U61309 ( .A(\shifter_0/reg_w_10[14] ), .B(n35413), .X(n14246) );
  nor_x1_sg U61310 ( .A(\shifter_0/reg_w_10[15] ), .B(n35413), .X(n14277) );
  nor_x1_sg U61311 ( .A(\shifter_0/reg_w_10[16] ), .B(n31693), .X(n14308) );
  nor_x1_sg U61312 ( .A(\shifter_0/reg_w_10[19] ), .B(n30532), .X(n14401) );
  nor_x1_sg U61313 ( .A(\shifter_0/reg_i_10[0] ), .B(n33995), .X(n14433) );
  nor_x1_sg U61314 ( .A(\shifter_0/reg_i_10[1] ), .B(n29703), .X(n14464) );
  nor_x1_sg U61315 ( .A(\shifter_0/reg_i_10[3] ), .B(n30022), .X(n14528) );
  nor_x1_sg U61316 ( .A(\shifter_0/reg_i_10[5] ), .B(n31051), .X(n14590) );
  nor_x1_sg U61317 ( .A(\shifter_0/reg_i_10[6] ), .B(n33995), .X(n14621) );
  nor_x1_sg U61318 ( .A(\shifter_0/reg_i_10[7] ), .B(n31051), .X(n14652) );
  nor_x1_sg U61319 ( .A(\shifter_0/reg_i_10[10] ), .B(n33995), .X(n14745) );
  nor_x1_sg U61320 ( .A(\shifter_0/reg_i_10[11] ), .B(n31693), .X(n14776) );
  nor_x1_sg U61321 ( .A(\shifter_0/reg_i_10[14] ), .B(n31052), .X(n14869) );
  nor_x1_sg U61322 ( .A(\shifter_0/reg_i_10[15] ), .B(n31693), .X(n14900) );
  nor_x1_sg U61323 ( .A(\shifter_0/reg_i_10[19] ), .B(n31052), .X(n15024) );
  nor_x1_sg U61324 ( .A(n11767), .B(n35302), .X(n11766) );
  nor_x1_sg U61325 ( .A(n11768), .B(n34520), .X(n11767) );
  nor_x1_sg U61326 ( .A(n41418), .B(n11770), .X(n11768) );
  nor_x1_sg U61327 ( .A(n13486), .B(n32222), .X(n13485) );
  nor_x1_sg U61328 ( .A(n31659), .B(n35252), .X(n13486) );
  nor_x1_sg U61329 ( .A(\shifter_0/reg_i_15[4] ), .B(n34287), .X(
        \shifter_0/n8937 ) );
  nor_x1_sg U61330 ( .A(\shifter_0/reg_i_15[18] ), .B(n34284), .X(
        \shifter_0/n8881 ) );
  nor_x1_sg U61331 ( .A(\shifter_0/reg_w_2[3] ), .B(n32891), .X(n13888) );
  nor_x1_sg U61332 ( .A(\shifter_0/reg_w_2[4] ), .B(n30966), .X(n13919) );
  nor_x1_sg U61333 ( .A(\shifter_0/reg_w_2[8] ), .B(n34857), .X(n14043) );
  nor_x1_sg U61334 ( .A(\shifter_0/reg_w_2[9] ), .B(n34855), .X(n14074) );
  nor_x1_sg U61335 ( .A(\shifter_0/reg_w_2[12] ), .B(n34858), .X(n14167) );
  nor_x1_sg U61336 ( .A(\shifter_0/reg_w_2[13] ), .B(n30635), .X(n14198) );
  nor_x1_sg U61337 ( .A(\shifter_0/reg_w_2[17] ), .B(n34858), .X(n14322) );
  nor_x1_sg U61338 ( .A(\shifter_0/reg_w_2[18] ), .B(n30636), .X(n14353) );
  nor_x1_sg U61339 ( .A(\shifter_0/reg_i_2[3] ), .B(n32889), .X(n14511) );
  nor_x1_sg U61340 ( .A(\shifter_0/reg_i_2[4] ), .B(n29771), .X(n14543) );
  nor_x1_sg U61341 ( .A(\shifter_0/reg_i_2[8] ), .B(n32893), .X(n14666) );
  nor_x1_sg U61342 ( .A(\shifter_0/reg_i_2[9] ), .B(n32894), .X(n14697) );
  nor_x1_sg U61343 ( .A(\shifter_0/reg_i_2[12] ), .B(n32893), .X(n14790) );
  nor_x1_sg U61344 ( .A(\shifter_0/reg_i_2[13] ), .B(n32889), .X(n14821) );
  nor_x1_sg U61345 ( .A(\shifter_0/reg_i_2[17] ), .B(n32899), .X(n14946) );
  nor_x1_sg U61346 ( .A(\shifter_0/reg_i_2[18] ), .B(n32891), .X(n14977) );
  nor_x1_sg U61347 ( .A(\shifter_0/reg_i_15[0] ), .B(n31793), .X(
        \shifter_0/n6393 ) );
  nor_x1_sg U61348 ( .A(\shifter_0/reg_i_15[1] ), .B(n34286), .X(
        \shifter_0/n8949 ) );
  nor_x1_sg U61349 ( .A(\shifter_0/reg_i_15[7] ), .B(n31794), .X(
        \shifter_0/n8925 ) );
  nor_x1_sg U61350 ( .A(\shifter_0/reg_i_15[10] ), .B(n34285), .X(
        \shifter_0/n8913 ) );
  nor_x1_sg U61351 ( .A(\shifter_0/reg_i_15[13] ), .B(n31365), .X(
        \shifter_0/n8901 ) );
  nor_x1_sg U61352 ( .A(\shifter_0/reg_i_15[14] ), .B(n34285), .X(
        \shifter_0/n8897 ) );
  nor_x1_sg U61353 ( .A(\shifter_0/reg_i_15[15] ), .B(n31793), .X(
        \shifter_0/n8893 ) );
  nor_x1_sg U61354 ( .A(\shifter_0/reg_i_15[19] ), .B(n31365), .X(
        \shifter_0/n8877 ) );
  nor_x1_sg U61355 ( .A(\shifter_0/reg_w_15[0] ), .B(n34380), .X(
        \shifter_0/n6473 ) );
  nor_x1_sg U61356 ( .A(\shifter_0/reg_w_15[1] ), .B(n31309), .X(
        \shifter_0/n6469 ) );
  nor_x1_sg U61357 ( .A(\shifter_0/reg_w_15[4] ), .B(n31309), .X(
        \shifter_0/n6457 ) );
  nor_x1_sg U61358 ( .A(\shifter_0/reg_w_15[7] ), .B(n34382), .X(
        \shifter_0/n6445 ) );
  nor_x1_sg U61359 ( .A(\shifter_0/reg_w_15[10] ), .B(n30362), .X(
        \shifter_0/n6433 ) );
  nor_x1_sg U61360 ( .A(\shifter_0/reg_w_15[13] ), .B(n30362), .X(
        \shifter_0/n6421 ) );
  nor_x1_sg U61361 ( .A(\shifter_0/reg_w_15[14] ), .B(n34379), .X(
        \shifter_0/n6417 ) );
  nor_x1_sg U61362 ( .A(\shifter_0/reg_w_15[15] ), .B(n31308), .X(
        \shifter_0/n6413 ) );
  nor_x1_sg U61363 ( .A(\shifter_0/reg_w_15[18] ), .B(n34380), .X(
        \shifter_0/n6401 ) );
  nor_x1_sg U61364 ( .A(\shifter_0/reg_w_15[19] ), .B(n31756), .X(
        \shifter_0/n6397 ) );
  nand_x1_sg U61365 ( .A(\shifter_0/reg_w_9[0] ), .B(n34447), .X(n11898) );
  nand_x1_sg U61366 ( .A(\shifter_0/reg_w_9[1] ), .B(n34447), .X(n11910) );
  nand_x1_sg U61367 ( .A(\shifter_0/reg_w_9[2] ), .B(n32188), .X(n11921) );
  nand_x1_sg U61368 ( .A(\shifter_0/reg_w_9[3] ), .B(n34448), .X(n11932) );
  nand_x1_sg U61369 ( .A(\shifter_0/reg_w_9[4] ), .B(n34448), .X(n11943) );
  nand_x1_sg U61370 ( .A(\shifter_0/reg_w_9[5] ), .B(n32191), .X(n11954) );
  nand_x1_sg U61371 ( .A(\shifter_0/reg_w_9[6] ), .B(n34450), .X(n11965) );
  nand_x1_sg U61372 ( .A(\shifter_0/reg_w_9[7] ), .B(n35653), .X(n11976) );
  nand_x1_sg U61373 ( .A(\shifter_0/reg_w_9[8] ), .B(n32190), .X(n11987) );
  nand_x1_sg U61374 ( .A(\shifter_0/reg_w_9[9] ), .B(n32191), .X(n11998) );
  nand_x1_sg U61375 ( .A(\shifter_0/reg_w_9[10] ), .B(n30835), .X(n12009) );
  nand_x1_sg U61376 ( .A(\shifter_0/reg_w_9[11] ), .B(n34449), .X(n12020) );
  nand_x1_sg U61377 ( .A(\shifter_0/reg_w_9[12] ), .B(n32189), .X(n12031) );
  nand_x1_sg U61378 ( .A(\shifter_0/reg_w_9[13] ), .B(n32190), .X(n12042) );
  nand_x1_sg U61379 ( .A(\shifter_0/reg_w_9[14] ), .B(n32186), .X(n12053) );
  nand_x1_sg U61380 ( .A(\shifter_0/reg_w_9[15] ), .B(n32191), .X(n12064) );
  nand_x1_sg U61381 ( .A(\shifter_0/reg_w_9[16] ), .B(n32188), .X(n12075) );
  nand_x1_sg U61382 ( .A(\shifter_0/reg_w_9[17] ), .B(n34447), .X(n12086) );
  nand_x1_sg U61383 ( .A(\shifter_0/reg_w_9[18] ), .B(n34450), .X(n12097) );
  nand_x1_sg U61384 ( .A(\shifter_0/reg_w_9[19] ), .B(n32189), .X(n12108) );
  nand_x1_sg U61385 ( .A(\shifter_0/reg_i_9[0] ), .B(n34450), .X(n12126) );
  nand_x1_sg U61386 ( .A(\shifter_0/reg_i_9[1] ), .B(n32186), .X(n12138) );
  nand_x1_sg U61387 ( .A(\shifter_0/reg_i_9[2] ), .B(n32190), .X(n12149) );
  nand_x1_sg U61388 ( .A(\shifter_0/reg_i_9[3] ), .B(n30834), .X(n12160) );
  nand_x1_sg U61389 ( .A(\shifter_0/reg_i_9[4] ), .B(n32191), .X(n12171) );
  nand_x1_sg U61390 ( .A(\shifter_0/reg_i_9[5] ), .B(n32189), .X(n12182) );
  nand_x1_sg U61391 ( .A(\shifter_0/reg_i_9[6] ), .B(n34449), .X(n12193) );
  nand_x1_sg U61392 ( .A(\shifter_0/reg_i_9[7] ), .B(n30835), .X(n12204) );
  nand_x1_sg U61393 ( .A(\shifter_0/reg_i_9[8] ), .B(n32189), .X(n12215) );
  nand_x1_sg U61394 ( .A(\shifter_0/reg_i_9[9] ), .B(n32188), .X(n12226) );
  nand_x1_sg U61395 ( .A(\shifter_0/reg_i_9[10] ), .B(n30834), .X(n12237) );
  nand_x1_sg U61396 ( .A(\shifter_0/reg_i_9[11] ), .B(n32186), .X(n12248) );
  nand_x1_sg U61397 ( .A(\shifter_0/reg_i_9[12] ), .B(n30834), .X(n12259) );
  nand_x1_sg U61398 ( .A(\shifter_0/reg_i_9[13] ), .B(n35653), .X(n12270) );
  nand_x1_sg U61399 ( .A(\shifter_0/reg_i_9[14] ), .B(n32190), .X(n12281) );
  nand_x1_sg U61400 ( .A(\shifter_0/reg_i_9[15] ), .B(n34449), .X(n12292) );
  nand_x1_sg U61401 ( .A(\shifter_0/reg_i_9[16] ), .B(n32188), .X(n12303) );
  nand_x1_sg U61402 ( .A(\shifter_0/reg_i_9[17] ), .B(n34448), .X(n12314) );
  nand_x1_sg U61403 ( .A(\shifter_0/reg_i_9[18] ), .B(n34448), .X(n12325) );
  nand_x1_sg U61404 ( .A(\shifter_0/reg_i_9[19] ), .B(n30835), .X(n12336) );
  nor_x1_sg U61405 ( .A(\shifter_0/reg_i_15[2] ), .B(n11535), .X(
        \shifter_0/n8945 ) );
  nor_x1_sg U61406 ( .A(\shifter_0/reg_i_15[17] ), .B(n34287), .X(
        \shifter_0/n8885 ) );
  nor_x1_sg U61407 ( .A(\filter_0/reg_xor_i_mask[18] ), .B(n32124), .X(n15135)
         );
  nor_x1_sg U61408 ( .A(\filter_0/reg_xor_i_mask[17] ), .B(n32118), .X(n15139)
         );
  nor_x1_sg U61409 ( .A(\filter_0/reg_xor_i_mask[19] ), .B(n32205), .X(n15130)
         );
  nor_x1_sg U61410 ( .A(\filter_0/reg_xor_i_mask[21] ), .B(n32115), .X(n15129)
         );
  nor_x1_sg U61411 ( .A(\filter_0/reg_xor_i_mask[23] ), .B(n32504), .X(n15132)
         );
  nor_x1_sg U61412 ( .A(\filter_0/reg_xor_i_mask[31] ), .B(n32503), .X(n15146)
         );
  nor_x1_sg U61413 ( .A(\filter_0/reg_xor_i_mask[30] ), .B(n32136), .X(n15145)
         );
  nor_x1_sg U61414 ( .A(\filter_0/reg_xor_i_mask[0] ), .B(n32127), .X(n15094)
         );
  nor_x1_sg U61415 ( .A(\filter_0/reg_xor_w_mask[18] ), .B(n32122), .X(n15264)
         );
  nor_x1_sg U61416 ( .A(\filter_0/reg_xor_w_mask[17] ), .B(n32120), .X(n15268)
         );
  nor_x1_sg U61417 ( .A(\filter_0/reg_xor_w_mask[19] ), .B(n32205), .X(n15259)
         );
  nor_x1_sg U61418 ( .A(\filter_0/reg_xor_w_mask[21] ), .B(n32114), .X(n15258)
         );
  nor_x1_sg U61419 ( .A(\filter_0/reg_xor_w_mask[23] ), .B(n29669), .X(n15261)
         );
  nor_x1_sg U61420 ( .A(\filter_0/reg_xor_w_mask[31] ), .B(n32503), .X(n15275)
         );
  nor_x1_sg U61421 ( .A(\filter_0/reg_xor_w_mask[30] ), .B(n32135), .X(n15274)
         );
  nor_x1_sg U61422 ( .A(\filter_0/reg_xor_w_mask[0] ), .B(n32127), .X(n15227)
         );
  nor_x1_sg U61423 ( .A(n32128), .B(\filter_0/reg_xor_i_mask[24] ), .X(n15152)
         );
  nor_x1_sg U61424 ( .A(n32123), .B(\filter_0/reg_xor_i_mask[26] ), .X(n15151)
         );
  nor_x1_sg U61425 ( .A(n32128), .B(\filter_0/reg_xor_i_mask[8] ), .X(n15119)
         );
  nor_x1_sg U61426 ( .A(n32124), .B(\filter_0/reg_xor_i_mask[10] ), .X(n15118)
         );
  nor_x1_sg U61427 ( .A(n32128), .B(\filter_0/reg_xor_w_mask[24] ), .X(n15281)
         );
  nor_x1_sg U61428 ( .A(n32122), .B(\filter_0/reg_xor_w_mask[26] ), .X(n15280)
         );
  nor_x1_sg U61429 ( .A(n32127), .B(\filter_0/reg_xor_w_mask[8] ), .X(n15248)
         );
  nor_x1_sg U61430 ( .A(n32124), .B(\filter_0/reg_xor_w_mask[10] ), .X(n15247)
         );
  nand_x1_sg U61431 ( .A(n32172), .B(n13847), .X(n13846) );
  nand_x1_sg U61432 ( .A(n31992), .B(n40904), .X(n13847) );
  inv_x1_sg U61433 ( .A(\shifter_0/reg_w_11[1] ), .X(n40904) );
  nand_x1_sg U61434 ( .A(n34550), .B(n13878), .X(n13877) );
  nand_x1_sg U61435 ( .A(n31751), .B(n40903), .X(n13878) );
  inv_x1_sg U61436 ( .A(\shifter_0/reg_w_11[2] ), .X(n40903) );
  nand_x1_sg U61437 ( .A(n32167), .B(n14002), .X(n14001) );
  nand_x1_sg U61438 ( .A(n31993), .B(n40901), .X(n14002) );
  inv_x1_sg U61439 ( .A(\shifter_0/reg_w_11[6] ), .X(n40901) );
  nand_x1_sg U61440 ( .A(n30784), .B(n14126), .X(n14125) );
  nand_x1_sg U61441 ( .A(n31994), .B(n40899), .X(n14126) );
  inv_x1_sg U61442 ( .A(\shifter_0/reg_w_11[10] ), .X(n40899) );
  nand_x1_sg U61443 ( .A(n34551), .B(n14157), .X(n14156) );
  nand_x1_sg U61444 ( .A(n30855), .B(n40898), .X(n14157) );
  inv_x1_sg U61445 ( .A(\shifter_0/reg_w_11[11] ), .X(n40898) );
  nand_x1_sg U61446 ( .A(n34549), .B(n14281), .X(n14280) );
  nand_x1_sg U61447 ( .A(n31992), .B(n40896), .X(n14281) );
  inv_x1_sg U61448 ( .A(\shifter_0/reg_w_11[15] ), .X(n40896) );
  nand_x1_sg U61449 ( .A(n34548), .B(n14405), .X(n14404) );
  nand_x1_sg U61450 ( .A(n34409), .B(n40894), .X(n14405) );
  inv_x1_sg U61451 ( .A(\shifter_0/reg_w_11[19] ), .X(n40894) );
  nand_x1_sg U61452 ( .A(n30138), .B(n14437), .X(n14436) );
  nand_x1_sg U61453 ( .A(n30855), .B(n41029), .X(n14437) );
  inv_x1_sg U61454 ( .A(\shifter_0/reg_i_11[0] ), .X(n41029) );
  nand_x1_sg U61455 ( .A(n31300), .B(n14625), .X(n14624) );
  nand_x1_sg U61456 ( .A(n31751), .B(n41025), .X(n14625) );
  inv_x1_sg U61457 ( .A(\shifter_0/reg_i_11[6] ), .X(n41025) );
  nand_x1_sg U61458 ( .A(n30784), .B(n14749), .X(n14748) );
  nand_x1_sg U61459 ( .A(n34411), .B(n41023), .X(n14749) );
  inv_x1_sg U61460 ( .A(\shifter_0/reg_i_11[10] ), .X(n41023) );
  nand_x1_sg U61461 ( .A(n31299), .B(n14780), .X(n14779) );
  nand_x1_sg U61462 ( .A(n31994), .B(n41022), .X(n14780) );
  inv_x1_sg U61463 ( .A(\shifter_0/reg_i_11[11] ), .X(n41022) );
  nand_x1_sg U61464 ( .A(n34550), .B(n14904), .X(n14903) );
  nand_x1_sg U61465 ( .A(n34410), .B(n41020), .X(n14904) );
  inv_x1_sg U61466 ( .A(\shifter_0/reg_i_11[15] ), .X(n41020) );
  nand_x1_sg U61467 ( .A(n31507), .B(\shifter_0/reg_w_1[1] ), .X(n13851) );
  nand_x1_sg U61468 ( .A(n33955), .B(\shifter_0/reg_w_1[5] ), .X(n13975) );
  nand_x1_sg U61469 ( .A(n33955), .B(\shifter_0/reg_w_1[7] ), .X(n14037) );
  nand_x1_sg U61470 ( .A(n33955), .B(\shifter_0/reg_w_1[11] ), .X(n14161) );
  nand_x1_sg U61471 ( .A(n30015), .B(\shifter_0/reg_w_1[15] ), .X(n14285) );
  nand_x1_sg U61472 ( .A(n33957), .B(\shifter_0/reg_w_1[19] ), .X(n14409) );
  nand_x1_sg U61473 ( .A(n33956), .B(\shifter_0/reg_i_1[1] ), .X(n14472) );
  nand_x1_sg U61474 ( .A(n30015), .B(\shifter_0/reg_i_1[5] ), .X(n14598) );
  nand_x1_sg U61475 ( .A(n33954), .B(\shifter_0/reg_i_1[7] ), .X(n14660) );
  nand_x1_sg U61476 ( .A(n31506), .B(\shifter_0/reg_i_1[11] ), .X(n14784) );
  nand_x1_sg U61477 ( .A(n31506), .B(\shifter_0/reg_i_1[15] ), .X(n14908) );
  nor_x1_sg U61478 ( .A(\shifter_0/reg_i_15[3] ), .B(n31794), .X(
        \shifter_0/n8941 ) );
  nor_x1_sg U61479 ( .A(\shifter_0/reg_i_15[5] ), .B(n31366), .X(
        \shifter_0/n8933 ) );
  nor_x1_sg U61480 ( .A(\shifter_0/reg_i_15[6] ), .B(n31793), .X(
        \shifter_0/n8929 ) );
  nor_x1_sg U61481 ( .A(\shifter_0/reg_i_15[8] ), .B(n34284), .X(
        \shifter_0/n8921 ) );
  nor_x1_sg U61482 ( .A(\shifter_0/reg_i_15[9] ), .B(n29725), .X(
        \shifter_0/n8917 ) );
  nor_x1_sg U61483 ( .A(\shifter_0/reg_i_15[11] ), .B(n31366), .X(
        \shifter_0/n8909 ) );
  nor_x1_sg U61484 ( .A(\shifter_0/reg_i_15[12] ), .B(n34285), .X(
        \shifter_0/n8905 ) );
  nor_x1_sg U61485 ( .A(\shifter_0/reg_i_15[16] ), .B(n30324), .X(
        \shifter_0/n8889 ) );
  nor_x1_sg U61486 ( .A(\shifter_0/reg_w_15[2] ), .B(n31756), .X(
        \shifter_0/n6465 ) );
  nor_x1_sg U61487 ( .A(\shifter_0/reg_w_15[3] ), .B(n31756), .X(
        \shifter_0/n6461 ) );
  nor_x1_sg U61488 ( .A(\shifter_0/reg_w_15[5] ), .B(n34381), .X(
        \shifter_0/n6453 ) );
  nor_x1_sg U61489 ( .A(\shifter_0/reg_w_15[6] ), .B(n31308), .X(
        \shifter_0/n6449 ) );
  nor_x1_sg U61490 ( .A(\shifter_0/reg_w_15[8] ), .B(n34382), .X(
        \shifter_0/n6441 ) );
  nor_x1_sg U61491 ( .A(\shifter_0/reg_w_15[9] ), .B(n35483), .X(
        \shifter_0/n6437 ) );
  nor_x1_sg U61492 ( .A(\shifter_0/reg_w_15[11] ), .B(n34381), .X(
        \shifter_0/n6429 ) );
  nor_x1_sg U61493 ( .A(\shifter_0/reg_w_15[12] ), .B(n34382), .X(
        \shifter_0/n6425 ) );
  nor_x1_sg U61494 ( .A(\shifter_0/reg_w_15[16] ), .B(n29706), .X(
        \shifter_0/n6409 ) );
  nor_x1_sg U61495 ( .A(\shifter_0/reg_w_15[17] ), .B(n31755), .X(
        \shifter_0/n6405 ) );
  nand_x1_sg U61496 ( .A(n34549), .B(n13813), .X(n13812) );
  nand_x1_sg U61497 ( .A(n31993), .B(n40905), .X(n13813) );
  inv_x1_sg U61498 ( .A(\shifter_0/reg_w_11[0] ), .X(n40905) );
  nand_x1_sg U61499 ( .A(n32170), .B(n13971), .X(n13970) );
  nand_x1_sg U61500 ( .A(n34410), .B(n40902), .X(n13971) );
  inv_x1_sg U61501 ( .A(\shifter_0/reg_w_11[5] ), .X(n40902) );
  nand_x1_sg U61502 ( .A(n34548), .B(n14250), .X(n14249) );
  nand_x1_sg U61503 ( .A(n34408), .B(n40897), .X(n14250) );
  inv_x1_sg U61504 ( .A(\shifter_0/reg_w_11[14] ), .X(n40897) );
  nand_x1_sg U61505 ( .A(n32171), .B(n14532), .X(n14531) );
  nand_x1_sg U61506 ( .A(n31751), .B(n41027), .X(n14532) );
  inv_x1_sg U61507 ( .A(\shifter_0/reg_i_11[3] ), .X(n41027) );
  nand_x1_sg U61508 ( .A(n32170), .B(n14594), .X(n14593) );
  nand_x1_sg U61509 ( .A(n31993), .B(n41026), .X(n14594) );
  inv_x1_sg U61510 ( .A(\shifter_0/reg_i_11[5] ), .X(n41026) );
  nand_x1_sg U61511 ( .A(n34549), .B(n14873), .X(n14872) );
  nand_x1_sg U61512 ( .A(n30855), .B(n41021), .X(n14873) );
  inv_x1_sg U61513 ( .A(\shifter_0/reg_i_11[14] ), .X(n41021) );
  nand_x1_sg U61514 ( .A(n33956), .B(\shifter_0/reg_w_1[0] ), .X(n13819) );
  nand_x1_sg U61515 ( .A(n33956), .B(\shifter_0/reg_w_1[2] ), .X(n13882) );
  nand_x1_sg U61516 ( .A(n33954), .B(\shifter_0/reg_w_1[6] ), .X(n14006) );
  nand_x1_sg U61517 ( .A(n33955), .B(\shifter_0/reg_w_1[10] ), .X(n14130) );
  nand_x1_sg U61518 ( .A(n33954), .B(\shifter_0/reg_w_1[14] ), .X(n14254) );
  nand_x1_sg U61519 ( .A(n31507), .B(\shifter_0/reg_w_1[16] ), .X(n14316) );
  nand_x1_sg U61520 ( .A(n31506), .B(\shifter_0/reg_i_1[0] ), .X(n14441) );
  nand_x1_sg U61521 ( .A(n33954), .B(\shifter_0/reg_i_1[2] ), .X(n14505) );
  nand_x1_sg U61522 ( .A(n30015), .B(\shifter_0/reg_i_1[6] ), .X(n14629) );
  nand_x1_sg U61523 ( .A(n33957), .B(\shifter_0/reg_i_1[10] ), .X(n14753) );
  nand_x1_sg U61524 ( .A(n33957), .B(\shifter_0/reg_i_1[14] ), .X(n14877) );
  nand_x1_sg U61525 ( .A(n30015), .B(\shifter_0/reg_i_1[16] ), .X(n14939) );
  nand_x1_sg U61526 ( .A(n31506), .B(\shifter_0/reg_i_1[19] ), .X(n15032) );
  nand_x1_sg U61527 ( .A(\shifter_0/reg_w_5[13] ), .B(n32064), .X(n14202) );
  nor_x1_sg U61528 ( .A(n12794), .B(n14203), .X(n14201) );
  nor_x1_sg U61529 ( .A(n30016), .B(n42695), .X(n14203) );
  nor_x1_sg U61530 ( .A(n12806), .B(n41125), .X(n14263) );
  nand_x1_sg U61531 ( .A(\shifter_0/reg_w_5[15] ), .B(n31022), .X(n14264) );
  inv_x1_sg U61532 ( .A(n14265), .X(n41125) );
  nand_x1_sg U61533 ( .A(\shifter_0/reg_w_5[17] ), .B(n32064), .X(n14326) );
  nor_x1_sg U61534 ( .A(n12818), .B(n14327), .X(n14325) );
  nor_x1_sg U61535 ( .A(n29688), .B(n42696), .X(n14327) );
  nor_x1_sg U61536 ( .A(n12830), .B(n41123), .X(n14387) );
  nand_x1_sg U61537 ( .A(\shifter_0/reg_w_5[19] ), .B(n30135), .X(n14388) );
  inv_x1_sg U61538 ( .A(n14389), .X(n41123) );
  nor_x1_sg U61539 ( .A(n12852), .B(n41121), .X(n14450) );
  nand_x1_sg U61540 ( .A(\shifter_0/reg_i_5[1] ), .B(n34541), .X(n14451) );
  inv_x1_sg U61541 ( .A(n14452), .X(n41121) );
  nand_x1_sg U61542 ( .A(\shifter_0/reg_i_5[3] ), .B(n32059), .X(n14515) );
  nor_x1_sg U61543 ( .A(n12864), .B(n14516), .X(n14514) );
  nor_x1_sg U61544 ( .A(n31652), .B(n42580), .X(n14516) );
  nor_x1_sg U61545 ( .A(n12876), .B(n41119), .X(n14576) );
  nand_x1_sg U61546 ( .A(\shifter_0/reg_i_5[5] ), .B(n32062), .X(n14577) );
  inv_x1_sg U61547 ( .A(n14578), .X(n41119) );
  nor_x1_sg U61548 ( .A(n12888), .B(n41117), .X(n14638) );
  nand_x1_sg U61549 ( .A(\shifter_0/reg_i_5[7] ), .B(n32063), .X(n14639) );
  inv_x1_sg U61550 ( .A(n14640), .X(n41117) );
  nand_x1_sg U61551 ( .A(\shifter_0/reg_i_5[9] ), .B(n32063), .X(n14701) );
  nor_x1_sg U61552 ( .A(n12900), .B(n14702), .X(n14700) );
  nor_x1_sg U61553 ( .A(n31653), .B(n42583), .X(n14702) );
  nor_x1_sg U61554 ( .A(n12912), .B(n41115), .X(n14762) );
  nand_x1_sg U61555 ( .A(\shifter_0/reg_i_5[11] ), .B(n34540), .X(n14763) );
  inv_x1_sg U61556 ( .A(n14764), .X(n41115) );
  nand_x1_sg U61557 ( .A(\shifter_0/reg_i_5[13] ), .B(n31023), .X(n14825) );
  nor_x1_sg U61558 ( .A(n12924), .B(n14826), .X(n14824) );
  nor_x1_sg U61559 ( .A(n33961), .B(n42585), .X(n14826) );
  nor_x1_sg U61560 ( .A(n12936), .B(n41113), .X(n14886) );
  nand_x1_sg U61561 ( .A(\shifter_0/reg_i_5[15] ), .B(n34539), .X(n14887) );
  inv_x1_sg U61562 ( .A(n14888), .X(n41113) );
  nor_x1_sg U61563 ( .A(n12715), .B(n41134), .X(n13792) );
  nand_x1_sg U61564 ( .A(\shifter_0/reg_w_5[0] ), .B(n34542), .X(n13793) );
  inv_x1_sg U61565 ( .A(n13794), .X(n41134) );
  nor_x1_sg U61566 ( .A(n12722), .B(n41133), .X(n13829) );
  nand_x1_sg U61567 ( .A(\shifter_0/reg_w_5[1] ), .B(n32062), .X(n13830) );
  inv_x1_sg U61568 ( .A(n13831), .X(n41133) );
  nor_x1_sg U61569 ( .A(n12728), .B(n41132), .X(n13860) );
  nand_x1_sg U61570 ( .A(\shifter_0/reg_w_5[2] ), .B(n34542), .X(n13861) );
  inv_x1_sg U61571 ( .A(n13862), .X(n41132) );
  nor_x1_sg U61572 ( .A(n12734), .B(n13893), .X(n13891) );
  nand_x1_sg U61573 ( .A(\shifter_0/reg_w_5[3] ), .B(n34541), .X(n13892) );
  nor_x1_sg U61574 ( .A(n33959), .B(n42690), .X(n13893) );
  nor_x1_sg U61575 ( .A(n12740), .B(n13924), .X(n13922) );
  nand_x1_sg U61576 ( .A(\shifter_0/reg_w_5[4] ), .B(n30135), .X(n13923) );
  nor_x1_sg U61577 ( .A(n33960), .B(n42691), .X(n13924) );
  nor_x1_sg U61578 ( .A(n12746), .B(n41131), .X(n13953) );
  nand_x1_sg U61579 ( .A(\shifter_0/reg_w_5[5] ), .B(n32060), .X(n13954) );
  inv_x1_sg U61580 ( .A(n13955), .X(n41131) );
  nor_x1_sg U61581 ( .A(n12752), .B(n41130), .X(n13984) );
  nand_x1_sg U61582 ( .A(\shifter_0/reg_w_5[6] ), .B(n34539), .X(n13985) );
  inv_x1_sg U61583 ( .A(n13986), .X(n41130) );
  nor_x1_sg U61584 ( .A(n12758), .B(n41129), .X(n14015) );
  nand_x1_sg U61585 ( .A(\shifter_0/reg_w_5[7] ), .B(n32063), .X(n14016) );
  inv_x1_sg U61586 ( .A(n14017), .X(n41129) );
  nor_x1_sg U61587 ( .A(n12764), .B(n14048), .X(n14046) );
  nand_x1_sg U61588 ( .A(\shifter_0/reg_w_5[8] ), .B(n32059), .X(n14047) );
  nor_x1_sg U61589 ( .A(n31653), .B(n42692), .X(n14048) );
  nor_x1_sg U61590 ( .A(n12770), .B(n14079), .X(n14077) );
  nand_x1_sg U61591 ( .A(\shifter_0/reg_w_5[9] ), .B(n34540), .X(n14078) );
  nor_x1_sg U61592 ( .A(n33961), .B(n42693), .X(n14079) );
  nor_x1_sg U61593 ( .A(n12776), .B(n41128), .X(n14108) );
  nand_x1_sg U61594 ( .A(\shifter_0/reg_w_5[10] ), .B(n32064), .X(n14109) );
  inv_x1_sg U61595 ( .A(n14110), .X(n41128) );
  nor_x1_sg U61596 ( .A(n12782), .B(n41127), .X(n14139) );
  nand_x1_sg U61597 ( .A(\shifter_0/reg_w_5[11] ), .B(n32060), .X(n14140) );
  inv_x1_sg U61598 ( .A(n14141), .X(n41127) );
  nor_x1_sg U61599 ( .A(n12788), .B(n14172), .X(n14170) );
  nand_x1_sg U61600 ( .A(\shifter_0/reg_w_5[12] ), .B(n34542), .X(n14171) );
  nor_x1_sg U61601 ( .A(n33959), .B(n42694), .X(n14172) );
  nor_x1_sg U61602 ( .A(n12800), .B(n41126), .X(n14232) );
  nand_x1_sg U61603 ( .A(\shifter_0/reg_w_5[14] ), .B(n31023), .X(n14233) );
  inv_x1_sg U61604 ( .A(n14234), .X(n41126) );
  nor_x1_sg U61605 ( .A(n12812), .B(n41124), .X(n14294) );
  nand_x1_sg U61606 ( .A(\shifter_0/reg_w_5[16] ), .B(n31022), .X(n14295) );
  inv_x1_sg U61607 ( .A(n14296), .X(n41124) );
  nor_x1_sg U61608 ( .A(n12824), .B(n14358), .X(n14356) );
  nand_x1_sg U61609 ( .A(\shifter_0/reg_w_5[18] ), .B(n30135), .X(n14357) );
  nor_x1_sg U61610 ( .A(n33961), .B(n42697), .X(n14358) );
  nor_x1_sg U61611 ( .A(n12846), .B(n41122), .X(n14419) );
  nand_x1_sg U61612 ( .A(\shifter_0/reg_i_5[0] ), .B(n34541), .X(n14420) );
  inv_x1_sg U61613 ( .A(n14421), .X(n41122) );
  nor_x1_sg U61614 ( .A(n12882), .B(n41118), .X(n14607) );
  nand_x1_sg U61615 ( .A(\shifter_0/reg_i_5[6] ), .B(n34540), .X(n14608) );
  inv_x1_sg U61616 ( .A(n14609), .X(n41118) );
  nor_x1_sg U61617 ( .A(n12894), .B(n14671), .X(n14669) );
  nand_x1_sg U61618 ( .A(\shifter_0/reg_i_5[8] ), .B(n31023), .X(n14670) );
  nor_x1_sg U61619 ( .A(n33962), .B(n42582), .X(n14671) );
  nor_x1_sg U61620 ( .A(n12906), .B(n41116), .X(n14731) );
  nand_x1_sg U61621 ( .A(\shifter_0/reg_i_5[10] ), .B(n32060), .X(n14732) );
  inv_x1_sg U61622 ( .A(n14733), .X(n41116) );
  nor_x1_sg U61623 ( .A(n12918), .B(n14795), .X(n14793) );
  nand_x1_sg U61624 ( .A(\shifter_0/reg_i_5[12] ), .B(n31023), .X(n14794) );
  nor_x1_sg U61625 ( .A(n30016), .B(n42584), .X(n14795) );
  nor_x1_sg U61626 ( .A(n12930), .B(n41114), .X(n14855) );
  nand_x1_sg U61627 ( .A(\shifter_0/reg_i_5[14] ), .B(n32059), .X(n14856) );
  inv_x1_sg U61628 ( .A(n14857), .X(n41114) );
  nor_x1_sg U61629 ( .A(n12942), .B(n41112), .X(n14917) );
  nand_x1_sg U61630 ( .A(\shifter_0/reg_i_5[16] ), .B(n34542), .X(n14918) );
  inv_x1_sg U61631 ( .A(n14919), .X(n41112) );
  nor_x1_sg U61632 ( .A(n12960), .B(n41111), .X(n15010) );
  nand_x1_sg U61633 ( .A(\shifter_0/reg_i_5[19] ), .B(n34539), .X(n15011) );
  inv_x1_sg U61634 ( .A(n15012), .X(n41111) );
  inv_x1_sg U61635 ( .A(\shifter_0/reg_w_6[0] ), .X(n40949) );
  inv_x1_sg U61636 ( .A(\shifter_0/reg_w_6[1] ), .X(n40947) );
  inv_x1_sg U61637 ( .A(\shifter_0/reg_w_6[2] ), .X(n40945) );
  inv_x1_sg U61638 ( .A(\shifter_0/reg_w_6[5] ), .X(n40941) );
  inv_x1_sg U61639 ( .A(\shifter_0/reg_w_6[6] ), .X(n40939) );
  inv_x1_sg U61640 ( .A(\shifter_0/reg_w_6[7] ), .X(n40937) );
  inv_x1_sg U61641 ( .A(\shifter_0/reg_w_6[10] ), .X(n40933) );
  inv_x1_sg U61642 ( .A(\shifter_0/reg_w_6[11] ), .X(n40931) );
  inv_x1_sg U61643 ( .A(\shifter_0/reg_w_6[14] ), .X(n40927) );
  inv_x1_sg U61644 ( .A(\shifter_0/reg_w_6[15] ), .X(n40925) );
  inv_x1_sg U61645 ( .A(\shifter_0/reg_w_6[16] ), .X(n40923) );
  inv_x1_sg U61646 ( .A(\shifter_0/reg_w_6[19] ), .X(n40919) );
  inv_x1_sg U61647 ( .A(\shifter_0/reg_i_6[0] ), .X(n41072) );
  inv_x1_sg U61648 ( .A(\shifter_0/reg_i_6[1] ), .X(n41070) );
  inv_x1_sg U61649 ( .A(\shifter_0/reg_i_6[2] ), .X(n41068) );
  inv_x1_sg U61650 ( .A(\shifter_0/reg_i_6[5] ), .X(n41064) );
  inv_x1_sg U61651 ( .A(\shifter_0/reg_i_6[6] ), .X(n41062) );
  inv_x1_sg U61652 ( .A(\shifter_0/reg_i_6[7] ), .X(n41060) );
  inv_x1_sg U61653 ( .A(\shifter_0/reg_i_6[10] ), .X(n41056) );
  inv_x1_sg U61654 ( .A(\shifter_0/reg_i_6[11] ), .X(n41054) );
  inv_x1_sg U61655 ( .A(\shifter_0/reg_i_6[14] ), .X(n41050) );
  inv_x1_sg U61656 ( .A(\shifter_0/reg_i_6[15] ), .X(n41048) );
  inv_x1_sg U61657 ( .A(\shifter_0/reg_i_6[16] ), .X(n41046) );
  inv_x1_sg U61658 ( .A(\shifter_0/reg_i_6[19] ), .X(n41042) );
  inv_x1_sg U61659 ( .A(\shifter_0/reg_w_2[0] ), .X(n40973) );
  inv_x1_sg U61660 ( .A(\shifter_0/reg_w_2[1] ), .X(n40972) );
  inv_x1_sg U61661 ( .A(\shifter_0/reg_w_2[2] ), .X(n40971) );
  inv_x1_sg U61662 ( .A(\shifter_0/reg_w_2[5] ), .X(n40970) );
  inv_x1_sg U61663 ( .A(\shifter_0/reg_w_2[6] ), .X(n40969) );
  inv_x1_sg U61664 ( .A(\shifter_0/reg_w_2[7] ), .X(n40968) );
  inv_x1_sg U61665 ( .A(\shifter_0/reg_w_2[10] ), .X(n40967) );
  inv_x1_sg U61666 ( .A(\shifter_0/reg_w_2[11] ), .X(n40966) );
  inv_x1_sg U61667 ( .A(\shifter_0/reg_w_2[14] ), .X(n40965) );
  inv_x1_sg U61668 ( .A(\shifter_0/reg_w_2[15] ), .X(n40964) );
  inv_x1_sg U61669 ( .A(\shifter_0/reg_w_2[16] ), .X(n40963) );
  inv_x1_sg U61670 ( .A(\shifter_0/reg_w_2[19] ), .X(n40962) );
  inv_x1_sg U61671 ( .A(\shifter_0/reg_i_2[0] ), .X(n41096) );
  inv_x1_sg U61672 ( .A(\shifter_0/reg_i_2[1] ), .X(n41095) );
  inv_x1_sg U61673 ( .A(\shifter_0/reg_i_2[2] ), .X(n41094) );
  inv_x1_sg U61674 ( .A(\shifter_0/reg_i_2[5] ), .X(n41093) );
  inv_x1_sg U61675 ( .A(\shifter_0/reg_i_2[6] ), .X(n41092) );
  inv_x1_sg U61676 ( .A(\shifter_0/reg_i_2[7] ), .X(n41091) );
  inv_x1_sg U61677 ( .A(\shifter_0/reg_i_2[10] ), .X(n41090) );
  inv_x1_sg U61678 ( .A(\shifter_0/reg_i_2[11] ), .X(n41089) );
  inv_x1_sg U61679 ( .A(\shifter_0/reg_i_2[14] ), .X(n41088) );
  inv_x1_sg U61680 ( .A(\shifter_0/reg_i_2[15] ), .X(n41087) );
  inv_x1_sg U61681 ( .A(\shifter_0/reg_i_2[16] ), .X(n41086) );
  inv_x1_sg U61682 ( .A(\shifter_0/reg_i_2[19] ), .X(n41085) );
  nor_x1_sg U61683 ( .A(n15113), .B(n31203), .X(n15109) );
  nor_x1_sg U61684 ( .A(\filter_0/reg_xor_i_mask[15] ), .B(n32505), .X(n15113)
         );
  nor_x1_sg U61685 ( .A(n15242), .B(n35306), .X(n15238) );
  nor_x1_sg U61686 ( .A(\filter_0/reg_xor_w_mask[15] ), .B(n29669), .X(n15242)
         );
  nand_x1_sg U61687 ( .A(n30389), .B(n31204), .X(n15164) );
  nand_x1_sg U61688 ( .A(n31656), .B(n35154), .X(n15163) );
  nand_x1_sg U61689 ( .A(n13301), .B(n13302), .X(n13300) );
  nand_x1_sg U61690 ( .A(\shifter_0/reg_i_3[2] ), .B(n32069), .X(n13302) );
  nand_x1_sg U61691 ( .A(n13308), .B(n13309), .X(n13307) );
  nand_x1_sg U61692 ( .A(\shifter_0/reg_i_3[4] ), .B(n31019), .X(n13309) );
  nand_x1_sg U61693 ( .A(n13348), .B(n13349), .X(n13347) );
  nand_x1_sg U61694 ( .A(\shifter_0/reg_i_3[17] ), .B(n32065), .X(n13349) );
  nand_x1_sg U61695 ( .A(n13352), .B(n13353), .X(n13351) );
  nand_x1_sg U61696 ( .A(\shifter_0/reg_i_3[18] ), .B(n34534), .X(n13353) );
  nand_x1_sg U61697 ( .A(n35096), .B(n30584), .X(n15213) );
  nand_x1_sg U61698 ( .A(n31658), .B(n30543), .X(n15214) );
  inv_x1_sg U61699 ( .A(\shifter_0/reg_w_5[0] ), .X(n40961) );
  inv_x1_sg U61700 ( .A(\shifter_0/reg_w_5[1] ), .X(n40960) );
  inv_x1_sg U61701 ( .A(\shifter_0/reg_w_5[2] ), .X(n40959) );
  inv_x1_sg U61702 ( .A(\shifter_0/reg_w_5[5] ), .X(n40958) );
  inv_x1_sg U61703 ( .A(\shifter_0/reg_w_5[6] ), .X(n40957) );
  inv_x1_sg U61704 ( .A(\shifter_0/reg_w_5[7] ), .X(n40956) );
  inv_x1_sg U61705 ( .A(\shifter_0/reg_w_5[10] ), .X(n40955) );
  inv_x1_sg U61706 ( .A(\shifter_0/reg_w_5[11] ), .X(n40954) );
  inv_x1_sg U61707 ( .A(\shifter_0/reg_w_5[14] ), .X(n40953) );
  inv_x1_sg U61708 ( .A(\shifter_0/reg_w_5[15] ), .X(n40952) );
  inv_x1_sg U61709 ( .A(\shifter_0/reg_w_5[16] ), .X(n40951) );
  inv_x1_sg U61710 ( .A(\shifter_0/reg_w_5[19] ), .X(n40950) );
  inv_x1_sg U61711 ( .A(\shifter_0/reg_i_5[0] ), .X(n41084) );
  inv_x1_sg U61712 ( .A(\shifter_0/reg_i_5[1] ), .X(n41083) );
  inv_x1_sg U61713 ( .A(\shifter_0/reg_i_5[2] ), .X(n41082) );
  inv_x1_sg U61714 ( .A(\shifter_0/reg_i_5[5] ), .X(n41081) );
  inv_x1_sg U61715 ( .A(\shifter_0/reg_i_5[6] ), .X(n41080) );
  inv_x1_sg U61716 ( .A(\shifter_0/reg_i_5[7] ), .X(n41079) );
  inv_x1_sg U61717 ( .A(\shifter_0/reg_i_5[10] ), .X(n41078) );
  inv_x1_sg U61718 ( .A(\shifter_0/reg_i_5[11] ), .X(n41077) );
  inv_x1_sg U61719 ( .A(\shifter_0/reg_i_5[14] ), .X(n41076) );
  inv_x1_sg U61720 ( .A(\shifter_0/reg_i_5[15] ), .X(n41075) );
  inv_x1_sg U61721 ( .A(\shifter_0/reg_i_5[16] ), .X(n41074) );
  inv_x1_sg U61722 ( .A(\shifter_0/reg_i_5[19] ), .X(n41073) );
  nor_x1_sg U61723 ( .A(n15161), .B(n42371), .X(n15159) );
  nand_x1_sg U61724 ( .A(n31594), .B(n31204), .X(n15160) );
  inv_x1_sg U61725 ( .A(n32205), .X(n42371) );
  nand_x1_sg U61726 ( .A(\shifter_0/reg_i_14[4] ), .B(n34442), .X(n12177) );
  nand_x1_sg U61727 ( .A(n31158), .B(n34440), .X(n12176) );
  nand_x1_sg U61728 ( .A(\shifter_0/reg_i_14[18] ), .B(n11561), .X(n12331) );
  nand_x1_sg U61729 ( .A(n31159), .B(n30839), .X(n12330) );
  nor_x1_sg U61730 ( .A(n30254), .B(n15061), .X(n15058) );
  nand_x1_sg U61731 ( .A(n31118), .B(n35565), .X(n15059) );
  nor_x1_sg U61732 ( .A(n35103), .B(n35565), .X(n15061) );
  nor_x1_sg U61733 ( .A(n30253), .B(n15197), .X(n15194) );
  nand_x1_sg U61734 ( .A(n31123), .B(n35564), .X(n15195) );
  nor_x1_sg U61735 ( .A(n35104), .B(n35564), .X(n15197) );
  nor_x1_sg U61736 ( .A(\filter_0/reg_i_8[19] ), .B(n34312), .X(
        \filter_0/n4980 ) );
  nor_x1_sg U61737 ( .A(\filter_0/reg_i_8[18] ), .B(n35599), .X(
        \filter_0/n7588 ) );
  nor_x1_sg U61738 ( .A(\filter_0/reg_i_8[17] ), .B(n31350), .X(
        \filter_0/n7584 ) );
  nor_x1_sg U61739 ( .A(\filter_0/reg_i_8[16] ), .B(n31783), .X(
        \filter_0/n7580 ) );
  nor_x1_sg U61740 ( .A(\filter_0/reg_i_8[15] ), .B(n34309), .X(
        \filter_0/n7576 ) );
  nor_x1_sg U61741 ( .A(\filter_0/reg_i_8[14] ), .B(n30097), .X(
        \filter_0/n7572 ) );
  nor_x1_sg U61742 ( .A(\filter_0/reg_i_8[13] ), .B(n30097), .X(
        \filter_0/n7568 ) );
  nor_x1_sg U61743 ( .A(\filter_0/reg_i_8[12] ), .B(n34310), .X(
        \filter_0/n7564 ) );
  nor_x1_sg U61744 ( .A(\filter_0/reg_i_8[11] ), .B(n34310), .X(
        \filter_0/n7560 ) );
  nor_x1_sg U61745 ( .A(\filter_0/reg_i_8[10] ), .B(n34309), .X(
        \filter_0/n7556 ) );
  nor_x1_sg U61746 ( .A(\filter_0/reg_i_8[9] ), .B(n31784), .X(
        \filter_0/n7552 ) );
  nor_x1_sg U61747 ( .A(\filter_0/reg_i_8[8] ), .B(n31783), .X(
        \filter_0/n7548 ) );
  nor_x1_sg U61748 ( .A(\filter_0/reg_i_8[7] ), .B(n29720), .X(
        \filter_0/n7544 ) );
  nor_x1_sg U61749 ( .A(\filter_0/reg_i_8[6] ), .B(n31350), .X(
        \filter_0/n7540 ) );
  nor_x1_sg U61750 ( .A(\filter_0/reg_i_8[5] ), .B(n31351), .X(
        \filter_0/n7536 ) );
  nor_x1_sg U61751 ( .A(\filter_0/reg_i_8[4] ), .B(n31783), .X(
        \filter_0/n7532 ) );
  nor_x1_sg U61752 ( .A(\filter_0/reg_i_8[3] ), .B(n34309), .X(
        \filter_0/n7528 ) );
  nor_x1_sg U61753 ( .A(\filter_0/reg_i_8[2] ), .B(n31783), .X(
        \filter_0/n7524 ) );
  nor_x1_sg U61754 ( .A(\filter_0/reg_i_8[1] ), .B(n30334), .X(
        \filter_0/n7520 ) );
  nor_x1_sg U61755 ( .A(\filter_0/reg_i_8[0] ), .B(n31350), .X(
        \filter_0/n7516 ) );
  nor_x1_sg U61756 ( .A(\filter_0/reg_i_9[19] ), .B(n31820), .X(
        \filter_0/n7512 ) );
  nor_x1_sg U61757 ( .A(\filter_0/reg_i_9[18] ), .B(n31417), .X(
        \filter_0/n7508 ) );
  nor_x1_sg U61758 ( .A(\filter_0/reg_i_9[17] ), .B(n34201), .X(
        \filter_0/n7504 ) );
  nor_x1_sg U61759 ( .A(\filter_0/reg_i_9[16] ), .B(n34202), .X(
        \filter_0/n7500 ) );
  nor_x1_sg U61760 ( .A(\filter_0/reg_i_9[15] ), .B(n15037), .X(
        \filter_0/n7496 ) );
  nor_x1_sg U61761 ( .A(\filter_0/reg_i_9[14] ), .B(n30283), .X(
        \filter_0/n7492 ) );
  nor_x1_sg U61762 ( .A(\filter_0/reg_i_9[13] ), .B(n31417), .X(
        \filter_0/n7488 ) );
  nor_x1_sg U61763 ( .A(\filter_0/reg_i_9[12] ), .B(n31417), .X(
        \filter_0/n7484 ) );
  nor_x1_sg U61764 ( .A(\filter_0/reg_i_9[11] ), .B(n31416), .X(
        \filter_0/n7480 ) );
  nor_x1_sg U61765 ( .A(\filter_0/reg_i_9[10] ), .B(n30075), .X(
        \filter_0/n7476 ) );
  nor_x1_sg U61766 ( .A(\filter_0/reg_i_9[9] ), .B(n34202), .X(
        \filter_0/n7472 ) );
  nor_x1_sg U61767 ( .A(\filter_0/reg_i_9[8] ), .B(n31821), .X(
        \filter_0/n7468 ) );
  nor_x1_sg U61768 ( .A(\filter_0/reg_i_9[7] ), .B(n31416), .X(
        \filter_0/n7464 ) );
  nor_x1_sg U61769 ( .A(\filter_0/reg_i_9[6] ), .B(n30283), .X(
        \filter_0/n7460 ) );
  nor_x1_sg U61770 ( .A(\filter_0/reg_i_9[5] ), .B(n30283), .X(
        \filter_0/n7456 ) );
  nor_x1_sg U61771 ( .A(\filter_0/reg_i_9[4] ), .B(n34200), .X(
        \filter_0/n7452 ) );
  nor_x1_sg U61772 ( .A(\filter_0/reg_i_9[3] ), .B(n31820), .X(
        \filter_0/n7448 ) );
  nor_x1_sg U61773 ( .A(\filter_0/reg_i_9[2] ), .B(n30075), .X(
        \filter_0/n7444 ) );
  nor_x1_sg U61774 ( .A(\filter_0/reg_i_9[1] ), .B(n34200), .X(
        \filter_0/n7440 ) );
  nor_x1_sg U61775 ( .A(\filter_0/reg_i_9[0] ), .B(n34200), .X(
        \filter_0/n7436 ) );
  nor_x1_sg U61776 ( .A(\filter_0/reg_i_10[19] ), .B(n29736), .X(
        \filter_0/n7432 ) );
  nor_x1_sg U61777 ( .A(\filter_0/reg_i_10[18] ), .B(n31823), .X(
        \filter_0/n7428 ) );
  nor_x1_sg U61778 ( .A(\filter_0/reg_i_10[17] ), .B(n34194), .X(
        \filter_0/n7424 ) );
  nor_x1_sg U61779 ( .A(\filter_0/reg_i_10[16] ), .B(n34195), .X(
        \filter_0/n7420 ) );
  nor_x1_sg U61780 ( .A(\filter_0/reg_i_10[15] ), .B(n30281), .X(
        \filter_0/n7416 ) );
  nor_x1_sg U61781 ( .A(\filter_0/reg_i_10[14] ), .B(n34197), .X(
        \filter_0/n7412 ) );
  nor_x1_sg U61782 ( .A(\filter_0/reg_i_10[13] ), .B(n34196), .X(
        \filter_0/n7408 ) );
  nor_x1_sg U61783 ( .A(\filter_0/reg_i_10[12] ), .B(n34195), .X(
        \filter_0/n7404 ) );
  nor_x1_sg U61784 ( .A(\filter_0/reg_i_10[11] ), .B(n31822), .X(
        \filter_0/n7400 ) );
  nor_x1_sg U61785 ( .A(\filter_0/reg_i_10[10] ), .B(n34197), .X(
        \filter_0/n7396 ) );
  nor_x1_sg U61786 ( .A(\filter_0/reg_i_10[9] ), .B(n31823), .X(
        \filter_0/n7392 ) );
  nor_x1_sg U61787 ( .A(\filter_0/reg_i_10[8] ), .B(n31822), .X(
        \filter_0/n7388 ) );
  nor_x1_sg U61788 ( .A(\filter_0/reg_i_10[7] ), .B(n30074), .X(
        \filter_0/n7384 ) );
  nor_x1_sg U61789 ( .A(\filter_0/reg_i_10[6] ), .B(n15038), .X(
        \filter_0/n7380 ) );
  nor_x1_sg U61790 ( .A(\filter_0/reg_i_10[5] ), .B(n31419), .X(
        \filter_0/n7376 ) );
  nor_x1_sg U61791 ( .A(\filter_0/reg_i_10[4] ), .B(n34194), .X(
        \filter_0/n7372 ) );
  nor_x1_sg U61792 ( .A(\filter_0/reg_i_10[3] ), .B(n31420), .X(
        \filter_0/n7368 ) );
  nor_x1_sg U61793 ( .A(\filter_0/reg_i_10[2] ), .B(n34195), .X(
        \filter_0/n7364 ) );
  nor_x1_sg U61794 ( .A(\filter_0/reg_i_10[1] ), .B(n31420), .X(
        \filter_0/n7360 ) );
  nor_x1_sg U61795 ( .A(\filter_0/reg_i_10[0] ), .B(n30281), .X(
        \filter_0/n7356 ) );
  nor_x1_sg U61796 ( .A(\filter_0/reg_i_11[19] ), .B(n34191), .X(
        \filter_0/n7352 ) );
  nor_x1_sg U61797 ( .A(\filter_0/reg_i_11[18] ), .B(n31422), .X(
        \filter_0/n7348 ) );
  nor_x1_sg U61798 ( .A(\filter_0/reg_i_11[17] ), .B(n31825), .X(
        \filter_0/n7344 ) );
  nor_x1_sg U61799 ( .A(\filter_0/reg_i_11[16] ), .B(n30073), .X(
        \filter_0/n7340 ) );
  nor_x1_sg U61800 ( .A(\filter_0/reg_i_11[15] ), .B(n31825), .X(
        \filter_0/n7336 ) );
  nor_x1_sg U61801 ( .A(\filter_0/reg_i_11[14] ), .B(n34192), .X(
        \filter_0/n7332 ) );
  nor_x1_sg U61802 ( .A(\filter_0/reg_i_11[13] ), .B(n34189), .X(
        \filter_0/n7328 ) );
  nor_x1_sg U61803 ( .A(\filter_0/reg_i_11[12] ), .B(n34190), .X(
        \filter_0/n7324 ) );
  nor_x1_sg U61804 ( .A(\filter_0/reg_i_11[11] ), .B(n34191), .X(
        \filter_0/n7320 ) );
  nor_x1_sg U61805 ( .A(\filter_0/reg_i_11[10] ), .B(n31422), .X(
        \filter_0/n7316 ) );
  nor_x1_sg U61806 ( .A(\filter_0/reg_i_11[9] ), .B(n29737), .X(
        \filter_0/n7312 ) );
  nor_x1_sg U61807 ( .A(\filter_0/reg_i_11[8] ), .B(n34190), .X(
        \filter_0/n7308 ) );
  nor_x1_sg U61808 ( .A(\filter_0/reg_i_11[7] ), .B(n29737), .X(
        \filter_0/n7304 ) );
  nor_x1_sg U61809 ( .A(\filter_0/reg_i_11[6] ), .B(n31824), .X(
        \filter_0/n7300 ) );
  nor_x1_sg U61810 ( .A(\filter_0/reg_i_11[5] ), .B(n31824), .X(
        \filter_0/n7296 ) );
  nor_x1_sg U61811 ( .A(\filter_0/reg_i_11[4] ), .B(n31824), .X(
        \filter_0/n7292 ) );
  nor_x1_sg U61812 ( .A(\filter_0/reg_i_11[3] ), .B(n30279), .X(
        \filter_0/n7288 ) );
  nor_x1_sg U61813 ( .A(\filter_0/reg_i_11[2] ), .B(n34192), .X(
        \filter_0/n7284 ) );
  nor_x1_sg U61814 ( .A(\filter_0/reg_i_11[1] ), .B(n34192), .X(
        \filter_0/n7280 ) );
  nor_x1_sg U61815 ( .A(\filter_0/reg_i_11[0] ), .B(n34190), .X(
        \filter_0/n7276 ) );
  nor_x1_sg U61816 ( .A(\filter_0/reg_i_15[19] ), .B(n34232), .X(
        \filter_0/n7272 ) );
  nor_x1_sg U61817 ( .A(\filter_0/reg_i_15[18] ), .B(n31399), .X(
        \filter_0/n7268 ) );
  nor_x1_sg U61818 ( .A(\filter_0/reg_i_15[17] ), .B(n30298), .X(
        \filter_0/n7264 ) );
  nor_x1_sg U61819 ( .A(\filter_0/reg_i_15[16] ), .B(n30081), .X(
        \filter_0/n7260 ) );
  nor_x1_sg U61820 ( .A(\filter_0/reg_i_15[15] ), .B(n31812), .X(
        \filter_0/n7256 ) );
  nor_x1_sg U61821 ( .A(\filter_0/reg_i_15[14] ), .B(n34230), .X(
        \filter_0/n7252 ) );
  nor_x1_sg U61822 ( .A(\filter_0/reg_i_15[13] ), .B(n34229), .X(
        \filter_0/n7248 ) );
  nor_x1_sg U61823 ( .A(\filter_0/reg_i_15[12] ), .B(n30081), .X(
        \filter_0/n7244 ) );
  nor_x1_sg U61824 ( .A(\filter_0/reg_i_15[11] ), .B(n34229), .X(
        \filter_0/n7240 ) );
  nor_x1_sg U61825 ( .A(\filter_0/reg_i_15[10] ), .B(n34229), .X(
        \filter_0/n7236 ) );
  nor_x1_sg U61826 ( .A(\filter_0/reg_i_15[9] ), .B(n31811), .X(
        \filter_0/n7232 ) );
  nor_x1_sg U61827 ( .A(\filter_0/reg_i_15[8] ), .B(n35633), .X(
        \filter_0/n7228 ) );
  nor_x1_sg U61828 ( .A(\filter_0/reg_i_15[7] ), .B(n34230), .X(
        \filter_0/n7224 ) );
  nor_x1_sg U61829 ( .A(\filter_0/reg_i_15[6] ), .B(n34231), .X(
        \filter_0/n7220 ) );
  nor_x1_sg U61830 ( .A(\filter_0/reg_i_15[5] ), .B(n31812), .X(
        \filter_0/n7216 ) );
  nor_x1_sg U61831 ( .A(\filter_0/reg_i_15[4] ), .B(n34231), .X(
        \filter_0/n7212 ) );
  nor_x1_sg U61832 ( .A(\filter_0/reg_i_15[3] ), .B(n34230), .X(
        \filter_0/n7208 ) );
  nor_x1_sg U61833 ( .A(\filter_0/reg_i_15[2] ), .B(n31399), .X(
        \filter_0/n7204 ) );
  nor_x1_sg U61834 ( .A(\filter_0/reg_i_15[1] ), .B(n29732), .X(
        \filter_0/n7200 ) );
  nor_x1_sg U61835 ( .A(\filter_0/reg_i_15[0] ), .B(n31812), .X(
        \filter_0/n7196 ) );
  nor_x1_sg U61836 ( .A(\filter_0/reg_i_12[19] ), .B(n31347), .X(
        \filter_0/n7192 ) );
  nor_x1_sg U61837 ( .A(\filter_0/reg_i_12[18] ), .B(n30336), .X(
        \filter_0/n7188 ) );
  nor_x1_sg U61838 ( .A(\filter_0/reg_i_12[17] ), .B(n31347), .X(
        \filter_0/n7184 ) );
  nor_x1_sg U61839 ( .A(\filter_0/reg_i_12[16] ), .B(n31782), .X(
        \filter_0/n7180 ) );
  nor_x1_sg U61840 ( .A(\filter_0/reg_i_12[15] ), .B(n34317), .X(
        \filter_0/n7176 ) );
  nor_x1_sg U61841 ( .A(\filter_0/reg_i_12[14] ), .B(n31348), .X(
        \filter_0/n7172 ) );
  nor_x1_sg U61842 ( .A(\filter_0/reg_i_12[13] ), .B(n35598), .X(
        \filter_0/n7168 ) );
  nor_x1_sg U61843 ( .A(\filter_0/reg_i_12[12] ), .B(n31781), .X(
        \filter_0/n7164 ) );
  nor_x1_sg U61844 ( .A(\filter_0/reg_i_12[11] ), .B(n30098), .X(
        \filter_0/n7160 ) );
  nor_x1_sg U61845 ( .A(\filter_0/reg_i_12[10] ), .B(n34315), .X(
        \filter_0/n7156 ) );
  nor_x1_sg U61846 ( .A(\filter_0/reg_i_12[9] ), .B(n34316), .X(
        \filter_0/n7152 ) );
  nor_x1_sg U61847 ( .A(\filter_0/reg_i_12[8] ), .B(n31348), .X(
        \filter_0/n7148 ) );
  nor_x1_sg U61848 ( .A(\filter_0/reg_i_12[7] ), .B(n34316), .X(
        \filter_0/n7144 ) );
  nor_x1_sg U61849 ( .A(\filter_0/reg_i_12[6] ), .B(n31782), .X(
        \filter_0/n7140 ) );
  nor_x1_sg U61850 ( .A(\filter_0/reg_i_12[5] ), .B(n31782), .X(
        \filter_0/n7136 ) );
  nor_x1_sg U61851 ( .A(\filter_0/reg_i_12[4] ), .B(n31348), .X(
        \filter_0/n7132 ) );
  nor_x1_sg U61852 ( .A(\filter_0/reg_i_12[3] ), .B(n34315), .X(
        \filter_0/n7128 ) );
  nor_x1_sg U61853 ( .A(\filter_0/reg_i_12[2] ), .B(n34314), .X(
        \filter_0/n7124 ) );
  nor_x1_sg U61854 ( .A(\filter_0/reg_i_12[1] ), .B(n34317), .X(
        \filter_0/n7120 ) );
  nor_x1_sg U61855 ( .A(\filter_0/reg_i_12[0] ), .B(n34315), .X(
        \filter_0/n7116 ) );
  nor_x1_sg U61856 ( .A(\filter_0/reg_i_13[19] ), .B(n31386), .X(
        \filter_0/n7112 ) );
  nor_x1_sg U61857 ( .A(\filter_0/reg_i_13[18] ), .B(n34250), .X(
        \filter_0/n7108 ) );
  nor_x1_sg U61858 ( .A(\filter_0/reg_i_13[17] ), .B(n34250), .X(
        \filter_0/n7104 ) );
  nor_x1_sg U61859 ( .A(\filter_0/reg_i_13[16] ), .B(n29728), .X(
        \filter_0/n7100 ) );
  nor_x1_sg U61860 ( .A(\filter_0/reg_i_13[15] ), .B(n31387), .X(
        \filter_0/n7096 ) );
  nor_x1_sg U61861 ( .A(\filter_0/reg_i_13[14] ), .B(n35632), .X(
        \filter_0/n7092 ) );
  nor_x1_sg U61862 ( .A(\filter_0/reg_i_13[13] ), .B(n34252), .X(
        \filter_0/n7088 ) );
  nor_x1_sg U61863 ( .A(\filter_0/reg_i_13[12] ), .B(n30306), .X(
        \filter_0/n7084 ) );
  nor_x1_sg U61864 ( .A(\filter_0/reg_i_13[11] ), .B(n34252), .X(
        \filter_0/n7080 ) );
  nor_x1_sg U61865 ( .A(\filter_0/reg_i_13[10] ), .B(n30085), .X(
        \filter_0/n7076 ) );
  nor_x1_sg U61866 ( .A(\filter_0/reg_i_13[9] ), .B(n34252), .X(
        \filter_0/n7072 ) );
  nor_x1_sg U61867 ( .A(\filter_0/reg_i_13[8] ), .B(n34249), .X(
        \filter_0/n7068 ) );
  nor_x1_sg U61868 ( .A(\filter_0/reg_i_13[7] ), .B(n31386), .X(
        \filter_0/n7064 ) );
  nor_x1_sg U61869 ( .A(\filter_0/reg_i_13[6] ), .B(n31803), .X(
        \filter_0/n7060 ) );
  nor_x1_sg U61870 ( .A(\filter_0/reg_i_13[5] ), .B(n31387), .X(
        \filter_0/n7056 ) );
  nor_x1_sg U61871 ( .A(\filter_0/reg_i_13[4] ), .B(n34249), .X(
        \filter_0/n7052 ) );
  nor_x1_sg U61872 ( .A(\filter_0/reg_i_13[3] ), .B(n31386), .X(
        \filter_0/n7048 ) );
  nor_x1_sg U61873 ( .A(\filter_0/reg_i_13[2] ), .B(n30306), .X(
        \filter_0/n7044 ) );
  nor_x1_sg U61874 ( .A(\filter_0/reg_i_13[1] ), .B(n34249), .X(
        \filter_0/n7040 ) );
  nor_x1_sg U61875 ( .A(\filter_0/reg_i_13[0] ), .B(n31804), .X(
        \filter_0/n7036 ) );
  nor_x1_sg U61876 ( .A(\filter_0/reg_i_14[19] ), .B(n31768), .X(
        \filter_0/n7032 ) );
  nor_x1_sg U61877 ( .A(\filter_0/reg_i_14[18] ), .B(n34351), .X(
        \filter_0/n7028 ) );
  nor_x1_sg U61878 ( .A(\filter_0/reg_i_14[17] ), .B(n34350), .X(
        \filter_0/n7024 ) );
  nor_x1_sg U61879 ( .A(\filter_0/reg_i_14[16] ), .B(n31326), .X(
        \filter_0/n7020 ) );
  nor_x1_sg U61880 ( .A(\filter_0/reg_i_14[15] ), .B(n31327), .X(
        \filter_0/n7016 ) );
  nor_x1_sg U61881 ( .A(\filter_0/reg_i_14[14] ), .B(n31767), .X(
        \filter_0/n7012 ) );
  nor_x1_sg U61882 ( .A(\filter_0/reg_i_14[13] ), .B(n31767), .X(
        \filter_0/n7008 ) );
  nor_x1_sg U61883 ( .A(\filter_0/reg_i_14[12] ), .B(n34352), .X(
        \filter_0/n7004 ) );
  nor_x1_sg U61884 ( .A(\filter_0/reg_i_14[11] ), .B(n29712), .X(
        \filter_0/n7000 ) );
  nor_x1_sg U61885 ( .A(\filter_0/reg_i_14[10] ), .B(n34352), .X(
        \filter_0/n6996 ) );
  nor_x1_sg U61886 ( .A(\filter_0/reg_i_14[9] ), .B(n31768), .X(
        \filter_0/n6992 ) );
  nor_x1_sg U61887 ( .A(\filter_0/reg_i_14[8] ), .B(n31327), .X(
        \filter_0/n6988 ) );
  nor_x1_sg U61888 ( .A(\filter_0/reg_i_14[7] ), .B(n30105), .X(
        \filter_0/n6984 ) );
  nor_x1_sg U61889 ( .A(\filter_0/reg_i_14[6] ), .B(n30350), .X(
        \filter_0/n6980 ) );
  nor_x1_sg U61890 ( .A(\filter_0/reg_i_14[5] ), .B(n34352), .X(
        \filter_0/n6976 ) );
  nor_x1_sg U61891 ( .A(\filter_0/reg_i_14[4] ), .B(n30105), .X(
        \filter_0/n6972 ) );
  nor_x1_sg U61892 ( .A(\filter_0/reg_i_14[3] ), .B(n34350), .X(
        \filter_0/n6968 ) );
  nor_x1_sg U61893 ( .A(\filter_0/reg_i_14[2] ), .B(n34352), .X(
        \filter_0/n6964 ) );
  nor_x1_sg U61894 ( .A(\filter_0/reg_i_14[1] ), .B(n30105), .X(
        \filter_0/n6960 ) );
  nor_x1_sg U61895 ( .A(\filter_0/reg_i_14[0] ), .B(n34350), .X(
        \filter_0/n6956 ) );
  nor_x1_sg U61896 ( .A(\filter_0/reg_i_4[19] ), .B(n31444), .X(
        \filter_0/n6952 ) );
  nor_x1_sg U61897 ( .A(\filter_0/reg_i_4[18] ), .B(n31838), .X(
        \filter_0/n6948 ) );
  nor_x1_sg U61898 ( .A(\filter_0/reg_i_4[17] ), .B(n31443), .X(
        \filter_0/n6944 ) );
  nor_x1_sg U61899 ( .A(\filter_0/reg_i_4[16] ), .B(n34154), .X(
        \filter_0/n6940 ) );
  nor_x1_sg U61900 ( .A(\filter_0/reg_i_4[15] ), .B(n31443), .X(
        \filter_0/n6936 ) );
  nor_x1_sg U61901 ( .A(\filter_0/reg_i_4[14] ), .B(n30066), .X(
        \filter_0/n6932 ) );
  nor_x1_sg U61902 ( .A(\filter_0/reg_i_4[13] ), .B(n34157), .X(
        \filter_0/n6928 ) );
  nor_x1_sg U61903 ( .A(\filter_0/reg_i_4[12] ), .B(n30265), .X(
        \filter_0/n6924 ) );
  nor_x1_sg U61904 ( .A(\filter_0/reg_i_4[11] ), .B(n34155), .X(
        \filter_0/n6920 ) );
  nor_x1_sg U61905 ( .A(\filter_0/reg_i_4[10] ), .B(n31838), .X(
        \filter_0/n6916 ) );
  nor_x1_sg U61906 ( .A(\filter_0/reg_i_4[9] ), .B(n29744), .X(
        \filter_0/n6912 ) );
  nor_x1_sg U61907 ( .A(\filter_0/reg_i_4[8] ), .B(n34155), .X(
        \filter_0/n6908 ) );
  nor_x1_sg U61908 ( .A(\filter_0/reg_i_4[7] ), .B(n34156), .X(
        \filter_0/n6904 ) );
  nor_x1_sg U61909 ( .A(\filter_0/reg_i_4[6] ), .B(n31839), .X(
        \filter_0/n6900 ) );
  nor_x1_sg U61910 ( .A(\filter_0/reg_i_4[5] ), .B(n31839), .X(
        \filter_0/n6896 ) );
  nor_x1_sg U61911 ( .A(\filter_0/reg_i_4[4] ), .B(n31839), .X(
        \filter_0/n6892 ) );
  nor_x1_sg U61912 ( .A(\filter_0/reg_i_4[3] ), .B(n34154), .X(
        \filter_0/n6888 ) );
  nor_x1_sg U61913 ( .A(\filter_0/reg_i_4[2] ), .B(n34156), .X(
        \filter_0/n6884 ) );
  nor_x1_sg U61914 ( .A(\filter_0/reg_i_4[1] ), .B(n31443), .X(
        \filter_0/n6880 ) );
  nor_x1_sg U61915 ( .A(\filter_0/reg_i_4[0] ), .B(n30265), .X(
        \filter_0/n6876 ) );
  nor_x1_sg U61916 ( .A(\filter_0/reg_i_5[19] ), .B(n31786), .X(
        \filter_0/n6872 ) );
  nor_x1_sg U61917 ( .A(\filter_0/reg_i_5[18] ), .B(n34305), .X(
        \filter_0/n6868 ) );
  nor_x1_sg U61918 ( .A(\filter_0/reg_i_5[17] ), .B(n31353), .X(
        \filter_0/n6864 ) );
  nor_x1_sg U61919 ( .A(\filter_0/reg_i_5[16] ), .B(n34306), .X(
        \filter_0/n6860 ) );
  nor_x1_sg U61920 ( .A(\filter_0/reg_i_5[15] ), .B(n34307), .X(
        \filter_0/n6856 ) );
  nor_x1_sg U61921 ( .A(\filter_0/reg_i_5[14] ), .B(n31785), .X(
        \filter_0/n6852 ) );
  nor_x1_sg U61922 ( .A(\filter_0/reg_i_5[13] ), .B(n30332), .X(
        \filter_0/n6848 ) );
  nor_x1_sg U61923 ( .A(\filter_0/reg_i_5[12] ), .B(n31786), .X(
        \filter_0/n6844 ) );
  nor_x1_sg U61924 ( .A(\filter_0/reg_i_5[11] ), .B(n31353), .X(
        \filter_0/n6840 ) );
  nor_x1_sg U61925 ( .A(\filter_0/reg_i_5[10] ), .B(n31785), .X(
        \filter_0/n6836 ) );
  nor_x1_sg U61926 ( .A(\filter_0/reg_i_5[9] ), .B(n34307), .X(
        \filter_0/n6832 ) );
  nor_x1_sg U61927 ( .A(\filter_0/reg_i_5[8] ), .B(n15046), .X(
        \filter_0/n6828 ) );
  nor_x1_sg U61928 ( .A(\filter_0/reg_i_5[7] ), .B(n34307), .X(
        \filter_0/n6824 ) );
  nor_x1_sg U61929 ( .A(\filter_0/reg_i_5[6] ), .B(n31353), .X(
        \filter_0/n6820 ) );
  nor_x1_sg U61930 ( .A(\filter_0/reg_i_5[5] ), .B(n30096), .X(
        \filter_0/n6816 ) );
  nor_x1_sg U61931 ( .A(\filter_0/reg_i_5[4] ), .B(n31354), .X(
        \filter_0/n6812 ) );
  nor_x1_sg U61932 ( .A(\filter_0/reg_i_5[3] ), .B(n31354), .X(
        \filter_0/n6808 ) );
  nor_x1_sg U61933 ( .A(\filter_0/reg_i_5[2] ), .B(n34304), .X(
        \filter_0/n6804 ) );
  nor_x1_sg U61934 ( .A(\filter_0/reg_i_5[1] ), .B(n34305), .X(
        \filter_0/n6800 ) );
  nor_x1_sg U61935 ( .A(\filter_0/reg_i_5[0] ), .B(n31353), .X(
        \filter_0/n6796 ) );
  nor_x1_sg U61936 ( .A(\filter_0/reg_i_6[19] ), .B(n31335), .X(
        \filter_0/n6792 ) );
  nor_x1_sg U61937 ( .A(\filter_0/reg_i_6[18] ), .B(n31336), .X(
        \filter_0/n6788 ) );
  nor_x1_sg U61938 ( .A(\filter_0/reg_i_6[17] ), .B(n34336), .X(
        \filter_0/n6784 ) );
  nor_x1_sg U61939 ( .A(\filter_0/reg_i_6[16] ), .B(n30344), .X(
        \filter_0/n6780 ) );
  nor_x1_sg U61940 ( .A(\filter_0/reg_i_6[15] ), .B(n31774), .X(
        \filter_0/n6776 ) );
  nor_x1_sg U61941 ( .A(\filter_0/reg_i_6[14] ), .B(n30102), .X(
        \filter_0/n6772 ) );
  nor_x1_sg U61942 ( .A(\filter_0/reg_i_6[13] ), .B(n30344), .X(
        \filter_0/n6768 ) );
  nor_x1_sg U61943 ( .A(\filter_0/reg_i_6[12] ), .B(n34334), .X(
        \filter_0/n6764 ) );
  nor_x1_sg U61944 ( .A(\filter_0/reg_i_6[11] ), .B(n34337), .X(
        \filter_0/n6760 ) );
  nor_x1_sg U61945 ( .A(\filter_0/reg_i_6[10] ), .B(n31774), .X(
        \filter_0/n6756 ) );
  nor_x1_sg U61946 ( .A(\filter_0/reg_i_6[9] ), .B(n34337), .X(
        \filter_0/n6752 ) );
  nor_x1_sg U61947 ( .A(\filter_0/reg_i_6[8] ), .B(n29715), .X(
        \filter_0/n6748 ) );
  nor_x1_sg U61948 ( .A(\filter_0/reg_i_6[7] ), .B(n34336), .X(
        \filter_0/n6744 ) );
  nor_x1_sg U61949 ( .A(\filter_0/reg_i_6[6] ), .B(n30102), .X(
        \filter_0/n6740 ) );
  nor_x1_sg U61950 ( .A(\filter_0/reg_i_6[5] ), .B(n34337), .X(
        \filter_0/n6736 ) );
  nor_x1_sg U61951 ( .A(\filter_0/reg_i_6[4] ), .B(n31773), .X(
        \filter_0/n6732 ) );
  nor_x1_sg U61952 ( .A(\filter_0/reg_i_6[3] ), .B(n34336), .X(
        \filter_0/n6728 ) );
  nor_x1_sg U61953 ( .A(\filter_0/reg_i_6[2] ), .B(n34337), .X(
        \filter_0/n6724 ) );
  nor_x1_sg U61954 ( .A(\filter_0/reg_i_6[1] ), .B(n34335), .X(
        \filter_0/n6720 ) );
  nor_x1_sg U61955 ( .A(\filter_0/reg_i_6[0] ), .B(n31774), .X(
        \filter_0/n6716 ) );
  nor_x1_sg U61956 ( .A(\filter_0/reg_i_7[19] ), .B(n31446), .X(
        \filter_0/n6712 ) );
  nor_x1_sg U61957 ( .A(\filter_0/reg_i_7[18] ), .B(n31446), .X(
        \filter_0/n6708 ) );
  nor_x1_sg U61958 ( .A(\filter_0/reg_i_7[17] ), .B(n31840), .X(
        \filter_0/n6704 ) );
  nor_x1_sg U61959 ( .A(\filter_0/reg_i_7[16] ), .B(n34149), .X(
        \filter_0/n6700 ) );
  nor_x1_sg U61960 ( .A(\filter_0/reg_i_7[15] ), .B(n31841), .X(
        \filter_0/n6696 ) );
  nor_x1_sg U61961 ( .A(\filter_0/reg_i_7[14] ), .B(n15048), .X(
        \filter_0/n6692 ) );
  nor_x1_sg U61962 ( .A(\filter_0/reg_i_7[13] ), .B(n34151), .X(
        \filter_0/n6688 ) );
  nor_x1_sg U61963 ( .A(\filter_0/reg_i_7[12] ), .B(n34152), .X(
        \filter_0/n6684 ) );
  nor_x1_sg U61964 ( .A(\filter_0/reg_i_7[11] ), .B(n34151), .X(
        \filter_0/n6680 ) );
  nor_x1_sg U61965 ( .A(\filter_0/reg_i_7[10] ), .B(n34152), .X(
        \filter_0/n6676 ) );
  nor_x1_sg U61966 ( .A(\filter_0/reg_i_7[9] ), .B(n31447), .X(
        \filter_0/n6672 ) );
  nor_x1_sg U61967 ( .A(\filter_0/reg_i_7[8] ), .B(n34151), .X(
        \filter_0/n6668 ) );
  nor_x1_sg U61968 ( .A(\filter_0/reg_i_7[7] ), .B(n34150), .X(
        \filter_0/n6664 ) );
  nor_x1_sg U61969 ( .A(\filter_0/reg_i_7[6] ), .B(n34149), .X(
        \filter_0/n6660 ) );
  nor_x1_sg U61970 ( .A(\filter_0/reg_i_7[5] ), .B(n31840), .X(
        \filter_0/n6656 ) );
  nor_x1_sg U61971 ( .A(\filter_0/reg_i_7[4] ), .B(n31841), .X(
        \filter_0/n6652 ) );
  nor_x1_sg U61972 ( .A(\filter_0/reg_i_7[3] ), .B(n31840), .X(
        \filter_0/n6648 ) );
  nor_x1_sg U61973 ( .A(\filter_0/reg_i_7[2] ), .B(n34152), .X(
        \filter_0/n6644 ) );
  nor_x1_sg U61974 ( .A(\filter_0/reg_i_7[1] ), .B(n30263), .X(
        \filter_0/n6640 ) );
  nor_x1_sg U61975 ( .A(\filter_0/reg_i_7[0] ), .B(n34150), .X(
        \filter_0/n6636 ) );
  nor_x1_sg U61976 ( .A(\filter_0/reg_i_0[19] ), .B(n34176), .X(
        \filter_0/n6632 ) );
  nor_x1_sg U61977 ( .A(\filter_0/reg_i_0[18] ), .B(n31431), .X(
        \filter_0/n6628 ) );
  nor_x1_sg U61978 ( .A(\filter_0/reg_i_0[17] ), .B(n31431), .X(
        \filter_0/n6624 ) );
  nor_x1_sg U61979 ( .A(\filter_0/reg_i_0[16] ), .B(n31431), .X(
        \filter_0/n6620 ) );
  nor_x1_sg U61980 ( .A(\filter_0/reg_i_0[15] ), .B(n15049), .X(
        \filter_0/n6616 ) );
  nor_x1_sg U61981 ( .A(\filter_0/reg_i_0[14] ), .B(n34175), .X(
        \filter_0/n6612 ) );
  nor_x1_sg U61982 ( .A(\filter_0/reg_i_0[13] ), .B(n30273), .X(
        \filter_0/n6608 ) );
  nor_x1_sg U61983 ( .A(\filter_0/reg_i_0[12] ), .B(n34174), .X(
        \filter_0/n6604 ) );
  nor_x1_sg U61984 ( .A(\filter_0/reg_i_0[11] ), .B(n34176), .X(
        \filter_0/n6600 ) );
  nor_x1_sg U61985 ( .A(\filter_0/reg_i_0[10] ), .B(n31831), .X(
        \filter_0/n6596 ) );
  nor_x1_sg U61986 ( .A(\filter_0/reg_i_0[9] ), .B(n30273), .X(
        \filter_0/n6592 ) );
  nor_x1_sg U61987 ( .A(\filter_0/reg_i_0[8] ), .B(n34175), .X(
        \filter_0/n6588 ) );
  nor_x1_sg U61988 ( .A(\filter_0/reg_i_0[7] ), .B(n31830), .X(
        \filter_0/n6584 ) );
  nor_x1_sg U61989 ( .A(\filter_0/reg_i_0[6] ), .B(n31831), .X(
        \filter_0/n6580 ) );
  nor_x1_sg U61990 ( .A(\filter_0/reg_i_0[5] ), .B(n34174), .X(
        \filter_0/n6576 ) );
  nor_x1_sg U61991 ( .A(\filter_0/reg_i_0[4] ), .B(n31432), .X(
        \filter_0/n6572 ) );
  nor_x1_sg U61992 ( .A(\filter_0/reg_i_0[3] ), .B(n34176), .X(
        \filter_0/n6568 ) );
  nor_x1_sg U61993 ( .A(\filter_0/reg_i_0[2] ), .B(n34177), .X(
        \filter_0/n6564 ) );
  nor_x1_sg U61994 ( .A(\filter_0/reg_i_0[1] ), .B(n31431), .X(
        \filter_0/n6560 ) );
  nor_x1_sg U61995 ( .A(\filter_0/reg_i_0[0] ), .B(n34175), .X(
        \filter_0/n6556 ) );
  nor_x1_sg U61996 ( .A(\filter_0/reg_i_1[19] ), .B(n31787), .X(
        \filter_0/n6552 ) );
  nor_x1_sg U61997 ( .A(\filter_0/reg_i_1[18] ), .B(n30095), .X(
        \filter_0/n6548 ) );
  nor_x1_sg U61998 ( .A(\filter_0/reg_i_1[17] ), .B(n34301), .X(
        \filter_0/n6544 ) );
  nor_x1_sg U61999 ( .A(\filter_0/reg_i_1[16] ), .B(n31788), .X(
        \filter_0/n6540 ) );
  nor_x1_sg U62000 ( .A(\filter_0/reg_i_1[15] ), .B(n31788), .X(
        \filter_0/n6536 ) );
  nor_x1_sg U62001 ( .A(\filter_0/reg_i_1[14] ), .B(n15050), .X(
        \filter_0/n6532 ) );
  nor_x1_sg U62002 ( .A(\filter_0/reg_i_1[13] ), .B(n31356), .X(
        \filter_0/n6528 ) );
  nor_x1_sg U62003 ( .A(\filter_0/reg_i_1[12] ), .B(n29722), .X(
        \filter_0/n6524 ) );
  nor_x1_sg U62004 ( .A(\filter_0/reg_i_1[11] ), .B(n31357), .X(
        \filter_0/n6520 ) );
  nor_x1_sg U62005 ( .A(\filter_0/reg_i_1[10] ), .B(n34300), .X(
        \filter_0/n6516 ) );
  nor_x1_sg U62006 ( .A(\filter_0/reg_i_1[9] ), .B(n31787), .X(
        \filter_0/n6512 ) );
  nor_x1_sg U62007 ( .A(\filter_0/reg_i_1[8] ), .B(n30095), .X(
        \filter_0/n6508 ) );
  nor_x1_sg U62008 ( .A(\filter_0/reg_i_1[7] ), .B(n34300), .X(
        \filter_0/n6504 ) );
  nor_x1_sg U62009 ( .A(\filter_0/reg_i_1[6] ), .B(n31787), .X(
        \filter_0/n6500 ) );
  nor_x1_sg U62010 ( .A(\filter_0/reg_i_1[5] ), .B(n34299), .X(
        \filter_0/n6496 ) );
  nor_x1_sg U62011 ( .A(\filter_0/reg_i_1[4] ), .B(n31356), .X(
        \filter_0/n6492 ) );
  nor_x1_sg U62012 ( .A(\filter_0/reg_i_1[3] ), .B(n31356), .X(
        \filter_0/n6488 ) );
  nor_x1_sg U62013 ( .A(\filter_0/reg_i_1[2] ), .B(n31357), .X(
        \filter_0/n6484 ) );
  nor_x1_sg U62014 ( .A(\filter_0/reg_i_1[1] ), .B(n34302), .X(
        \filter_0/n6480 ) );
  nor_x1_sg U62015 ( .A(\filter_0/reg_i_1[0] ), .B(n31787), .X(
        \filter_0/n6476 ) );
  nor_x1_sg U62016 ( .A(\filter_0/reg_i_2[19] ), .B(n29705), .X(
        \filter_0/n6472 ) );
  nor_x1_sg U62017 ( .A(\filter_0/reg_i_2[18] ), .B(n31306), .X(
        \filter_0/n6468 ) );
  nor_x1_sg U62018 ( .A(\filter_0/reg_i_2[17] ), .B(n31753), .X(
        \filter_0/n6464 ) );
  nor_x1_sg U62019 ( .A(\filter_0/reg_i_2[16] ), .B(n31754), .X(
        \filter_0/n6460 ) );
  nor_x1_sg U62020 ( .A(\filter_0/reg_i_2[15] ), .B(n34384), .X(
        \filter_0/n6456 ) );
  nor_x1_sg U62021 ( .A(\filter_0/reg_i_2[14] ), .B(n31753), .X(
        \filter_0/n6452 ) );
  nor_x1_sg U62022 ( .A(\filter_0/reg_i_2[13] ), .B(n30364), .X(
        \filter_0/n6448 ) );
  nor_x1_sg U62023 ( .A(\filter_0/reg_i_2[12] ), .B(n31305), .X(
        \filter_0/n6444 ) );
  nor_x1_sg U62024 ( .A(\filter_0/reg_i_2[11] ), .B(n30112), .X(
        \filter_0/n6440 ) );
  nor_x1_sg U62025 ( .A(\filter_0/reg_i_2[10] ), .B(n15053), .X(
        \filter_0/n6436 ) );
  nor_x1_sg U62026 ( .A(\filter_0/reg_i_2[9] ), .B(n29705), .X(
        \filter_0/n6432 ) );
  nor_x1_sg U62027 ( .A(\filter_0/reg_i_2[8] ), .B(n34386), .X(
        \filter_0/n6428 ) );
  nor_x1_sg U62028 ( .A(\filter_0/reg_i_2[7] ), .B(n31306), .X(
        \filter_0/n6424 ) );
  nor_x1_sg U62029 ( .A(\filter_0/reg_i_2[6] ), .B(n34387), .X(
        \filter_0/n6420 ) );
  nor_x1_sg U62030 ( .A(\filter_0/reg_i_2[5] ), .B(n31753), .X(
        \filter_0/n6416 ) );
  nor_x1_sg U62031 ( .A(\filter_0/reg_i_2[4] ), .B(n34385), .X(
        \filter_0/n6412 ) );
  nor_x1_sg U62032 ( .A(\filter_0/reg_i_2[3] ), .B(n31754), .X(
        \filter_0/n6408 ) );
  nor_x1_sg U62033 ( .A(\filter_0/reg_i_2[2] ), .B(n34387), .X(
        \filter_0/n6404 ) );
  nor_x1_sg U62034 ( .A(\filter_0/reg_i_2[1] ), .B(n34384), .X(
        \filter_0/n6400 ) );
  nor_x1_sg U62035 ( .A(\filter_0/reg_i_2[0] ), .B(n34385), .X(
        \filter_0/n6396 ) );
  nor_x1_sg U62036 ( .A(\filter_0/reg_i_3[19] ), .B(n34170), .X(
        \filter_0/n6392 ) );
  nor_x1_sg U62037 ( .A(\filter_0/reg_i_3[18] ), .B(n34169), .X(
        \filter_0/n6388 ) );
  nor_x1_sg U62038 ( .A(\filter_0/reg_i_3[17] ), .B(n30271), .X(
        \filter_0/n6384 ) );
  nor_x1_sg U62039 ( .A(\filter_0/reg_i_3[16] ), .B(n34170), .X(
        \filter_0/n6380 ) );
  nor_x1_sg U62040 ( .A(\filter_0/reg_i_3[15] ), .B(n31832), .X(
        \filter_0/n6376 ) );
  nor_x1_sg U62041 ( .A(\filter_0/reg_i_3[14] ), .B(n34170), .X(
        \filter_0/n6372 ) );
  nor_x1_sg U62042 ( .A(\filter_0/reg_i_3[13] ), .B(n31832), .X(
        \filter_0/n6368 ) );
  nor_x1_sg U62043 ( .A(\filter_0/reg_i_3[12] ), .B(n34170), .X(
        \filter_0/n6364 ) );
  nor_x1_sg U62044 ( .A(\filter_0/reg_i_3[11] ), .B(n31832), .X(
        \filter_0/n6360 ) );
  nor_x1_sg U62045 ( .A(\filter_0/reg_i_3[10] ), .B(n34172), .X(
        \filter_0/n6356 ) );
  nor_x1_sg U62046 ( .A(\filter_0/reg_i_3[9] ), .B(n31434), .X(
        \filter_0/n6352 ) );
  nor_x1_sg U62047 ( .A(\filter_0/reg_i_3[8] ), .B(n31435), .X(
        \filter_0/n6348 ) );
  nor_x1_sg U62048 ( .A(\filter_0/reg_i_3[7] ), .B(n15055), .X(
        \filter_0/n6344 ) );
  nor_x1_sg U62049 ( .A(\filter_0/reg_i_3[6] ), .B(n31434), .X(
        \filter_0/n6340 ) );
  nor_x1_sg U62050 ( .A(\filter_0/reg_i_3[5] ), .B(n34169), .X(
        \filter_0/n6336 ) );
  nor_x1_sg U62051 ( .A(\filter_0/reg_i_3[4] ), .B(n30271), .X(
        \filter_0/n6332 ) );
  nor_x1_sg U62052 ( .A(\filter_0/reg_i_3[3] ), .B(n34172), .X(
        \filter_0/n6328 ) );
  nor_x1_sg U62053 ( .A(\filter_0/reg_i_3[2] ), .B(n31832), .X(
        \filter_0/n6324 ) );
  nor_x1_sg U62054 ( .A(\filter_0/reg_i_3[1] ), .B(n34171), .X(
        \filter_0/n6320 ) );
  nor_x1_sg U62055 ( .A(\filter_0/reg_i_3[0] ), .B(n34172), .X(
        \filter_0/n6316 ) );
  nor_x1_sg U62056 ( .A(\filter_0/reg_w_8[19] ), .B(n34322), .X(
        \filter_0/n6276 ) );
  nor_x1_sg U62057 ( .A(\filter_0/reg_w_8[18] ), .B(n31780), .X(
        \filter_0/n6272 ) );
  nor_x1_sg U62058 ( .A(\filter_0/reg_w_8[17] ), .B(n31780), .X(
        \filter_0/n6268 ) );
  nor_x1_sg U62059 ( .A(\filter_0/reg_w_8[16] ), .B(n34320), .X(
        \filter_0/n6264 ) );
  nor_x1_sg U62060 ( .A(\filter_0/reg_w_8[15] ), .B(n31779), .X(
        \filter_0/n6260 ) );
  nor_x1_sg U62061 ( .A(\filter_0/reg_w_8[14] ), .B(n30099), .X(
        \filter_0/n6256 ) );
  nor_x1_sg U62062 ( .A(\filter_0/reg_w_8[13] ), .B(n34322), .X(
        \filter_0/n6252 ) );
  nor_x1_sg U62063 ( .A(\filter_0/reg_w_8[12] ), .B(n34320), .X(
        \filter_0/n6248 ) );
  nor_x1_sg U62064 ( .A(\filter_0/reg_w_8[11] ), .B(n31780), .X(
        \filter_0/n6244 ) );
  nor_x1_sg U62065 ( .A(\filter_0/reg_w_8[10] ), .B(n31779), .X(
        \filter_0/n6240 ) );
  nor_x1_sg U62066 ( .A(\filter_0/reg_w_8[9] ), .B(n34321), .X(
        \filter_0/n6236 ) );
  nor_x1_sg U62067 ( .A(\filter_0/reg_w_8[8] ), .B(n31344), .X(
        \filter_0/n6232 ) );
  nor_x1_sg U62068 ( .A(\filter_0/reg_w_8[7] ), .B(n31344), .X(
        \filter_0/n6228 ) );
  nor_x1_sg U62069 ( .A(\filter_0/reg_w_8[6] ), .B(n31345), .X(
        \filter_0/n6224 ) );
  nor_x1_sg U62070 ( .A(\filter_0/reg_w_8[5] ), .B(n29718), .X(
        \filter_0/n6220 ) );
  nor_x1_sg U62071 ( .A(\filter_0/reg_w_8[4] ), .B(n34319), .X(
        \filter_0/n6216 ) );
  nor_x1_sg U62072 ( .A(\filter_0/reg_w_8[3] ), .B(n34319), .X(
        \filter_0/n6212 ) );
  nor_x1_sg U62073 ( .A(\filter_0/reg_w_8[2] ), .B(n34320), .X(
        \filter_0/n6208 ) );
  nor_x1_sg U62074 ( .A(\filter_0/reg_w_8[1] ), .B(n29718), .X(
        \filter_0/n6204 ) );
  nor_x1_sg U62075 ( .A(\filter_0/reg_w_8[0] ), .B(n34321), .X(
        \filter_0/n6200 ) );
  nor_x1_sg U62076 ( .A(\filter_0/reg_w_9[19] ), .B(n34187), .X(
        \filter_0/n6196 ) );
  nor_x1_sg U62077 ( .A(\filter_0/reg_w_9[18] ), .B(n15170), .X(
        \filter_0/n6192 ) );
  nor_x1_sg U62078 ( .A(\filter_0/reg_w_9[17] ), .B(n31426), .X(
        \filter_0/n6188 ) );
  nor_x1_sg U62079 ( .A(\filter_0/reg_w_9[16] ), .B(n34184), .X(
        \filter_0/n6184 ) );
  nor_x1_sg U62080 ( .A(\filter_0/reg_w_9[15] ), .B(n29738), .X(
        \filter_0/n6180 ) );
  nor_x1_sg U62081 ( .A(\filter_0/reg_w_9[14] ), .B(n34186), .X(
        \filter_0/n6176 ) );
  nor_x1_sg U62082 ( .A(\filter_0/reg_w_9[13] ), .B(n34187), .X(
        \filter_0/n6172 ) );
  nor_x1_sg U62083 ( .A(\filter_0/reg_w_9[12] ), .B(n34187), .X(
        \filter_0/n6168 ) );
  nor_x1_sg U62084 ( .A(\filter_0/reg_w_9[11] ), .B(n30277), .X(
        \filter_0/n6164 ) );
  nor_x1_sg U62085 ( .A(\filter_0/reg_w_9[10] ), .B(n34184), .X(
        \filter_0/n6160 ) );
  nor_x1_sg U62086 ( .A(\filter_0/reg_w_9[9] ), .B(n30277), .X(
        \filter_0/n6156 ) );
  nor_x1_sg U62087 ( .A(\filter_0/reg_w_9[8] ), .B(n31425), .X(
        \filter_0/n6152 ) );
  nor_x1_sg U62088 ( .A(\filter_0/reg_w_9[7] ), .B(n31425), .X(
        \filter_0/n6148 ) );
  nor_x1_sg U62089 ( .A(\filter_0/reg_w_9[6] ), .B(n34185), .X(
        \filter_0/n6144 ) );
  nor_x1_sg U62090 ( .A(\filter_0/reg_w_9[5] ), .B(n31425), .X(
        \filter_0/n6140 ) );
  nor_x1_sg U62091 ( .A(\filter_0/reg_w_9[4] ), .B(n34187), .X(
        \filter_0/n6136 ) );
  nor_x1_sg U62092 ( .A(\filter_0/reg_w_9[3] ), .B(n34185), .X(
        \filter_0/n6132 ) );
  nor_x1_sg U62093 ( .A(\filter_0/reg_w_9[2] ), .B(n31826), .X(
        \filter_0/n6128 ) );
  nor_x1_sg U62094 ( .A(\filter_0/reg_w_9[1] ), .B(n31827), .X(
        \filter_0/n6124 ) );
  nor_x1_sg U62095 ( .A(\filter_0/reg_w_9[0] ), .B(n34185), .X(
        \filter_0/n6120 ) );
  nor_x1_sg U62096 ( .A(\filter_0/reg_w_10[19] ), .B(n34132), .X(
        \filter_0/n6116 ) );
  nor_x1_sg U62097 ( .A(\filter_0/reg_w_10[18] ), .B(n31848), .X(
        \filter_0/n6112 ) );
  nor_x1_sg U62098 ( .A(\filter_0/reg_w_10[17] ), .B(n30060), .X(
        \filter_0/n6108 ) );
  nor_x1_sg U62099 ( .A(\filter_0/reg_w_10[16] ), .B(n30060), .X(
        \filter_0/n6104 ) );
  nor_x1_sg U62100 ( .A(\filter_0/reg_w_10[15] ), .B(n34132), .X(
        \filter_0/n6100 ) );
  nor_x1_sg U62101 ( .A(\filter_0/reg_w_10[14] ), .B(n31848), .X(
        \filter_0/n6096 ) );
  nor_x1_sg U62102 ( .A(\filter_0/reg_w_10[13] ), .B(n31849), .X(
        \filter_0/n6092 ) );
  nor_x1_sg U62103 ( .A(\filter_0/reg_w_10[12] ), .B(n31849), .X(
        \filter_0/n6088 ) );
  nor_x1_sg U62104 ( .A(\filter_0/reg_w_10[11] ), .B(n34129), .X(
        \filter_0/n6084 ) );
  nor_x1_sg U62105 ( .A(\filter_0/reg_w_10[10] ), .B(n34130), .X(
        \filter_0/n6080 ) );
  nor_x1_sg U62106 ( .A(\filter_0/reg_w_10[9] ), .B(n31459), .X(
        \filter_0/n6076 ) );
  nor_x1_sg U62107 ( .A(\filter_0/reg_w_10[8] ), .B(n31848), .X(
        \filter_0/n6072 ) );
  nor_x1_sg U62108 ( .A(\filter_0/reg_w_10[7] ), .B(n31459), .X(
        \filter_0/n6068 ) );
  nor_x1_sg U62109 ( .A(\filter_0/reg_w_10[6] ), .B(n34132), .X(
        \filter_0/n6064 ) );
  nor_x1_sg U62110 ( .A(\filter_0/reg_w_10[5] ), .B(n34131), .X(
        \filter_0/n6060 ) );
  nor_x1_sg U62111 ( .A(\filter_0/reg_w_10[4] ), .B(n31459), .X(
        \filter_0/n6056 ) );
  nor_x1_sg U62112 ( .A(\filter_0/reg_w_10[3] ), .B(n34129), .X(
        \filter_0/n6052 ) );
  nor_x1_sg U62113 ( .A(\filter_0/reg_w_10[2] ), .B(n31458), .X(
        \filter_0/n6048 ) );
  nor_x1_sg U62114 ( .A(\filter_0/reg_w_10[1] ), .B(n34131), .X(
        \filter_0/n6044 ) );
  nor_x1_sg U62115 ( .A(\filter_0/reg_w_10[0] ), .B(n34129), .X(
        \filter_0/n6040 ) );
  nor_x1_sg U62116 ( .A(\filter_0/reg_w_11[19] ), .B(n34179), .X(
        \filter_0/n6036 ) );
  nor_x1_sg U62117 ( .A(\filter_0/reg_w_11[18] ), .B(n31428), .X(
        \filter_0/n6032 ) );
  nor_x1_sg U62118 ( .A(\filter_0/reg_w_11[17] ), .B(n34182), .X(
        \filter_0/n6028 ) );
  nor_x1_sg U62119 ( .A(\filter_0/reg_w_11[16] ), .B(n31828), .X(
        \filter_0/n6024 ) );
  nor_x1_sg U62120 ( .A(\filter_0/reg_w_11[15] ), .B(n31428), .X(
        \filter_0/n6020 ) );
  nor_x1_sg U62121 ( .A(\filter_0/reg_w_11[14] ), .B(n34181), .X(
        \filter_0/n6016 ) );
  nor_x1_sg U62122 ( .A(\filter_0/reg_w_11[13] ), .B(n34180), .X(
        \filter_0/n6012 ) );
  nor_x1_sg U62123 ( .A(\filter_0/reg_w_11[12] ), .B(n31428), .X(
        \filter_0/n6008 ) );
  nor_x1_sg U62124 ( .A(\filter_0/reg_w_11[11] ), .B(n30071), .X(
        \filter_0/n6004 ) );
  nor_x1_sg U62125 ( .A(\filter_0/reg_w_11[10] ), .B(n31428), .X(
        \filter_0/n6000 ) );
  nor_x1_sg U62126 ( .A(\filter_0/reg_w_11[9] ), .B(n29739), .X(
        \filter_0/n5996 ) );
  nor_x1_sg U62127 ( .A(\filter_0/reg_w_11[8] ), .B(n34181), .X(
        \filter_0/n5992 ) );
  nor_x1_sg U62128 ( .A(\filter_0/reg_w_11[7] ), .B(n31828), .X(
        \filter_0/n5988 ) );
  nor_x1_sg U62129 ( .A(\filter_0/reg_w_11[6] ), .B(n31828), .X(
        \filter_0/n5984 ) );
  nor_x1_sg U62130 ( .A(\filter_0/reg_w_11[5] ), .B(n31829), .X(
        \filter_0/n5980 ) );
  nor_x1_sg U62131 ( .A(\filter_0/reg_w_11[4] ), .B(n30275), .X(
        \filter_0/n5976 ) );
  nor_x1_sg U62132 ( .A(\filter_0/reg_w_11[3] ), .B(n34179), .X(
        \filter_0/n5972 ) );
  nor_x1_sg U62133 ( .A(\filter_0/reg_w_11[2] ), .B(n31429), .X(
        \filter_0/n5968 ) );
  nor_x1_sg U62134 ( .A(\filter_0/reg_w_11[1] ), .B(n31829), .X(
        \filter_0/n5964 ) );
  nor_x1_sg U62135 ( .A(\filter_0/reg_w_11[0] ), .B(n34180), .X(
        \filter_0/n5960 ) );
  nor_x1_sg U62136 ( .A(\filter_0/reg_w_15[19] ), .B(n35630), .X(
        \filter_0/n5956 ) );
  nor_x1_sg U62137 ( .A(\filter_0/reg_w_15[18] ), .B(n34245), .X(
        \filter_0/n5952 ) );
  nor_x1_sg U62138 ( .A(\filter_0/reg_w_15[17] ), .B(n34246), .X(
        \filter_0/n5948 ) );
  nor_x1_sg U62139 ( .A(\filter_0/reg_w_15[16] ), .B(n34247), .X(
        \filter_0/n5944 ) );
  nor_x1_sg U62140 ( .A(\filter_0/reg_w_15[15] ), .B(n31389), .X(
        \filter_0/n5940 ) );
  nor_x1_sg U62141 ( .A(\filter_0/reg_w_15[14] ), .B(n34246), .X(
        \filter_0/n5936 ) );
  nor_x1_sg U62142 ( .A(\filter_0/reg_w_15[13] ), .B(n34246), .X(
        \filter_0/n5932 ) );
  nor_x1_sg U62143 ( .A(\filter_0/reg_w_15[12] ), .B(n34247), .X(
        \filter_0/n5928 ) );
  nor_x1_sg U62144 ( .A(\filter_0/reg_w_15[11] ), .B(n34245), .X(
        \filter_0/n5924 ) );
  nor_x1_sg U62145 ( .A(\filter_0/reg_w_15[10] ), .B(n31806), .X(
        \filter_0/n5920 ) );
  nor_x1_sg U62146 ( .A(\filter_0/reg_w_15[9] ), .B(n34244), .X(
        \filter_0/n5916 ) );
  nor_x1_sg U62147 ( .A(\filter_0/reg_w_15[8] ), .B(n31806), .X(
        \filter_0/n5912 ) );
  nor_x1_sg U62148 ( .A(\filter_0/reg_w_15[7] ), .B(n34247), .X(
        \filter_0/n5908 ) );
  nor_x1_sg U62149 ( .A(\filter_0/reg_w_15[6] ), .B(n34245), .X(
        \filter_0/n5904 ) );
  nor_x1_sg U62150 ( .A(\filter_0/reg_w_15[5] ), .B(n34245), .X(
        \filter_0/n5900 ) );
  nor_x1_sg U62151 ( .A(\filter_0/reg_w_15[4] ), .B(n31805), .X(
        \filter_0/n5896 ) );
  nor_x1_sg U62152 ( .A(\filter_0/reg_w_15[3] ), .B(n30304), .X(
        \filter_0/n5892 ) );
  nor_x1_sg U62153 ( .A(\filter_0/reg_w_15[2] ), .B(n30304), .X(
        \filter_0/n5888 ) );
  nor_x1_sg U62154 ( .A(\filter_0/reg_w_15[1] ), .B(n30084), .X(
        \filter_0/n5884 ) );
  nor_x1_sg U62155 ( .A(\filter_0/reg_w_15[0] ), .B(n34244), .X(
        \filter_0/n5880 ) );
  nor_x1_sg U62156 ( .A(\filter_0/reg_w_12[19] ), .B(n34240), .X(
        \filter_0/n5876 ) );
  nor_x1_sg U62157 ( .A(\filter_0/reg_w_12[18] ), .B(n34240), .X(
        \filter_0/n5872 ) );
  nor_x1_sg U62158 ( .A(\filter_0/reg_w_12[17] ), .B(n31807), .X(
        \filter_0/n5868 ) );
  nor_x1_sg U62159 ( .A(\filter_0/reg_w_12[16] ), .B(n31392), .X(
        \filter_0/n5864 ) );
  nor_x1_sg U62160 ( .A(\filter_0/reg_w_12[15] ), .B(n34239), .X(
        \filter_0/n5860 ) );
  nor_x1_sg U62161 ( .A(\filter_0/reg_w_12[14] ), .B(n31393), .X(
        \filter_0/n5856 ) );
  nor_x1_sg U62162 ( .A(\filter_0/reg_w_12[13] ), .B(n30083), .X(
        \filter_0/n5852 ) );
  nor_x1_sg U62163 ( .A(\filter_0/reg_w_12[12] ), .B(n34242), .X(
        \filter_0/n5848 ) );
  nor_x1_sg U62164 ( .A(\filter_0/reg_w_12[11] ), .B(n31393), .X(
        \filter_0/n5844 ) );
  nor_x1_sg U62165 ( .A(\filter_0/reg_w_12[10] ), .B(n31392), .X(
        \filter_0/n5840 ) );
  nor_x1_sg U62166 ( .A(\filter_0/reg_w_12[9] ), .B(n31807), .X(
        \filter_0/n5836 ) );
  nor_x1_sg U62167 ( .A(\filter_0/reg_w_12[8] ), .B(n34242), .X(
        \filter_0/n5832 ) );
  nor_x1_sg U62168 ( .A(\filter_0/reg_w_12[7] ), .B(n30083), .X(
        \filter_0/n5828 ) );
  nor_x1_sg U62169 ( .A(\filter_0/reg_w_12[6] ), .B(n30302), .X(
        \filter_0/n5824 ) );
  nor_x1_sg U62170 ( .A(\filter_0/reg_w_12[5] ), .B(n31808), .X(
        \filter_0/n5820 ) );
  nor_x1_sg U62171 ( .A(\filter_0/reg_w_12[4] ), .B(n34239), .X(
        \filter_0/n5816 ) );
  nor_x1_sg U62172 ( .A(\filter_0/reg_w_12[3] ), .B(n34239), .X(
        \filter_0/n5812 ) );
  nor_x1_sg U62173 ( .A(\filter_0/reg_w_12[2] ), .B(n31393), .X(
        \filter_0/n5808 ) );
  nor_x1_sg U62174 ( .A(\filter_0/reg_w_12[1] ), .B(n29730), .X(
        \filter_0/n5804 ) );
  nor_x1_sg U62175 ( .A(\filter_0/reg_w_12[0] ), .B(n31807), .X(
        \filter_0/n5800 ) );
  nor_x1_sg U62176 ( .A(\filter_0/reg_w_13[19] ), .B(n31342), .X(
        \filter_0/n5796 ) );
  nor_x1_sg U62177 ( .A(\filter_0/reg_w_13[18] ), .B(n34325), .X(
        \filter_0/n5792 ) );
  nor_x1_sg U62178 ( .A(\filter_0/reg_w_13[17] ), .B(n30340), .X(
        \filter_0/n5788 ) );
  nor_x1_sg U62179 ( .A(\filter_0/reg_w_13[16] ), .B(n34325), .X(
        \filter_0/n5784 ) );
  nor_x1_sg U62180 ( .A(\filter_0/reg_w_13[15] ), .B(n35596), .X(
        \filter_0/n5780 ) );
  nor_x1_sg U62181 ( .A(\filter_0/reg_w_13[14] ), .B(n34325), .X(
        \filter_0/n5776 ) );
  nor_x1_sg U62182 ( .A(\filter_0/reg_w_13[13] ), .B(n31778), .X(
        \filter_0/n5772 ) );
  nor_x1_sg U62183 ( .A(\filter_0/reg_w_13[12] ), .B(n30100), .X(
        \filter_0/n5768 ) );
  nor_x1_sg U62184 ( .A(\filter_0/reg_w_13[11] ), .B(n31777), .X(
        \filter_0/n5764 ) );
  nor_x1_sg U62185 ( .A(\filter_0/reg_w_13[10] ), .B(n31341), .X(
        \filter_0/n5760 ) );
  nor_x1_sg U62186 ( .A(\filter_0/reg_w_13[9] ), .B(n34326), .X(
        \filter_0/n5756 ) );
  nor_x1_sg U62187 ( .A(\filter_0/reg_w_13[8] ), .B(n34324), .X(
        \filter_0/n5752 ) );
  nor_x1_sg U62188 ( .A(\filter_0/reg_w_13[7] ), .B(n34324), .X(
        \filter_0/n5748 ) );
  nor_x1_sg U62189 ( .A(\filter_0/reg_w_13[6] ), .B(n29717), .X(
        \filter_0/n5744 ) );
  nor_x1_sg U62190 ( .A(\filter_0/reg_w_13[5] ), .B(n31778), .X(
        \filter_0/n5740 ) );
  nor_x1_sg U62191 ( .A(\filter_0/reg_w_13[4] ), .B(n31777), .X(
        \filter_0/n5736 ) );
  nor_x1_sg U62192 ( .A(\filter_0/reg_w_13[3] ), .B(n31341), .X(
        \filter_0/n5732 ) );
  nor_x1_sg U62193 ( .A(\filter_0/reg_w_13[2] ), .B(n31342), .X(
        \filter_0/n5728 ) );
  nor_x1_sg U62194 ( .A(\filter_0/reg_w_13[1] ), .B(n34327), .X(
        \filter_0/n5724 ) );
  nor_x1_sg U62195 ( .A(\filter_0/reg_w_13[0] ), .B(n34327), .X(
        \filter_0/n5720 ) );
  nor_x1_sg U62196 ( .A(\filter_0/reg_w_14[19] ), .B(n31339), .X(
        \filter_0/n5716 ) );
  nor_x1_sg U62197 ( .A(\filter_0/reg_w_14[18] ), .B(n30101), .X(
        \filter_0/n5712 ) );
  nor_x1_sg U62198 ( .A(\filter_0/reg_w_14[17] ), .B(n34330), .X(
        \filter_0/n5708 ) );
  nor_x1_sg U62199 ( .A(\filter_0/reg_w_14[16] ), .B(n31338), .X(
        \filter_0/n5704 ) );
  nor_x1_sg U62200 ( .A(\filter_0/reg_w_14[15] ), .B(n34330), .X(
        \filter_0/n5700 ) );
  nor_x1_sg U62201 ( .A(\filter_0/reg_w_14[14] ), .B(n35595), .X(
        \filter_0/n5696 ) );
  nor_x1_sg U62202 ( .A(\filter_0/reg_w_14[13] ), .B(n31338), .X(
        \filter_0/n5692 ) );
  nor_x1_sg U62203 ( .A(\filter_0/reg_w_14[12] ), .B(n34331), .X(
        \filter_0/n5688 ) );
  nor_x1_sg U62204 ( .A(\filter_0/reg_w_14[11] ), .B(n31775), .X(
        \filter_0/n5684 ) );
  nor_x1_sg U62205 ( .A(\filter_0/reg_w_14[10] ), .B(n30342), .X(
        \filter_0/n5680 ) );
  nor_x1_sg U62206 ( .A(\filter_0/reg_w_14[9] ), .B(n31775), .X(
        \filter_0/n5676 ) );
  nor_x1_sg U62207 ( .A(\filter_0/reg_w_14[8] ), .B(n31776), .X(
        \filter_0/n5672 ) );
  nor_x1_sg U62208 ( .A(\filter_0/reg_w_14[7] ), .B(n30101), .X(
        \filter_0/n5668 ) );
  nor_x1_sg U62209 ( .A(\filter_0/reg_w_14[6] ), .B(n31338), .X(
        \filter_0/n5664 ) );
  nor_x1_sg U62210 ( .A(\filter_0/reg_w_14[5] ), .B(n31775), .X(
        \filter_0/n5660 ) );
  nor_x1_sg U62211 ( .A(\filter_0/reg_w_14[4] ), .B(n34329), .X(
        \filter_0/n5656 ) );
  nor_x1_sg U62212 ( .A(\filter_0/reg_w_14[3] ), .B(n31776), .X(
        \filter_0/n5652 ) );
  nor_x1_sg U62213 ( .A(\filter_0/reg_w_14[2] ), .B(n34332), .X(
        \filter_0/n5648 ) );
  nor_x1_sg U62214 ( .A(\filter_0/reg_w_14[1] ), .B(n31338), .X(
        \filter_0/n5644 ) );
  nor_x1_sg U62215 ( .A(\filter_0/reg_w_14[0] ), .B(n34329), .X(
        \filter_0/n5640 ) );
  nor_x1_sg U62216 ( .A(\filter_0/reg_w_4[19] ), .B(n34144), .X(
        \filter_0/n5636 ) );
  nor_x1_sg U62217 ( .A(\filter_0/reg_w_4[18] ), .B(n31843), .X(
        \filter_0/n5632 ) );
  nor_x1_sg U62218 ( .A(\filter_0/reg_w_4[17] ), .B(n34146), .X(
        \filter_0/n5628 ) );
  nor_x1_sg U62219 ( .A(\filter_0/reg_w_4[16] ), .B(n34145), .X(
        \filter_0/n5624 ) );
  nor_x1_sg U62220 ( .A(\filter_0/reg_w_4[15] ), .B(n31450), .X(
        \filter_0/n5620 ) );
  nor_x1_sg U62221 ( .A(\filter_0/reg_w_4[14] ), .B(n29746), .X(
        \filter_0/n5616 ) );
  nor_x1_sg U62222 ( .A(\filter_0/reg_w_4[13] ), .B(n31842), .X(
        \filter_0/n5612 ) );
  nor_x1_sg U62223 ( .A(\filter_0/reg_w_4[12] ), .B(n30064), .X(
        \filter_0/n5608 ) );
  nor_x1_sg U62224 ( .A(\filter_0/reg_w_4[11] ), .B(n31842), .X(
        \filter_0/n5604 ) );
  nor_x1_sg U62225 ( .A(\filter_0/reg_w_4[10] ), .B(n34147), .X(
        \filter_0/n5600 ) );
  nor_x1_sg U62226 ( .A(\filter_0/reg_w_4[9] ), .B(n34146), .X(
        \filter_0/n5596 ) );
  nor_x1_sg U62227 ( .A(\filter_0/reg_w_4[8] ), .B(n31842), .X(
        \filter_0/n5592 ) );
  nor_x1_sg U62228 ( .A(\filter_0/reg_w_4[7] ), .B(n31842), .X(
        \filter_0/n5588 ) );
  nor_x1_sg U62229 ( .A(\filter_0/reg_w_4[6] ), .B(n31449), .X(
        \filter_0/n5584 ) );
  nor_x1_sg U62230 ( .A(\filter_0/reg_w_4[5] ), .B(n34147), .X(
        \filter_0/n5580 ) );
  nor_x1_sg U62231 ( .A(\filter_0/reg_w_4[4] ), .B(n34144), .X(
        \filter_0/n5576 ) );
  nor_x1_sg U62232 ( .A(\filter_0/reg_w_4[3] ), .B(n15177), .X(
        \filter_0/n5572 ) );
  nor_x1_sg U62233 ( .A(\filter_0/reg_w_4[2] ), .B(n34147), .X(
        \filter_0/n5568 ) );
  nor_x1_sg U62234 ( .A(\filter_0/reg_w_4[1] ), .B(n29746), .X(
        \filter_0/n5564 ) );
  nor_x1_sg U62235 ( .A(\filter_0/reg_w_4[0] ), .B(n31450), .X(
        \filter_0/n5560 ) );
  nor_x1_sg U62236 ( .A(\filter_0/reg_w_5[19] ), .B(n31359), .X(
        \filter_0/n5556 ) );
  nor_x1_sg U62237 ( .A(\filter_0/reg_w_5[18] ), .B(n34294), .X(
        \filter_0/n5552 ) );
  nor_x1_sg U62238 ( .A(\filter_0/reg_w_5[17] ), .B(n34294), .X(
        \filter_0/n5548 ) );
  nor_x1_sg U62239 ( .A(\filter_0/reg_w_5[16] ), .B(n30328), .X(
        \filter_0/n5544 ) );
  nor_x1_sg U62240 ( .A(\filter_0/reg_w_5[15] ), .B(n34295), .X(
        \filter_0/n5540 ) );
  nor_x1_sg U62241 ( .A(\filter_0/reg_w_5[14] ), .B(n30328), .X(
        \filter_0/n5536 ) );
  nor_x1_sg U62242 ( .A(\filter_0/reg_w_5[13] ), .B(n15179), .X(
        \filter_0/n5532 ) );
  nor_x1_sg U62243 ( .A(\filter_0/reg_w_5[12] ), .B(n31359), .X(
        \filter_0/n5528 ) );
  nor_x1_sg U62244 ( .A(\filter_0/reg_w_5[11] ), .B(n31359), .X(
        \filter_0/n5524 ) );
  nor_x1_sg U62245 ( .A(\filter_0/reg_w_5[10] ), .B(n31789), .X(
        \filter_0/n5520 ) );
  nor_x1_sg U62246 ( .A(\filter_0/reg_w_5[9] ), .B(n34297), .X(
        \filter_0/n5516 ) );
  nor_x1_sg U62247 ( .A(\filter_0/reg_w_5[8] ), .B(n34297), .X(
        \filter_0/n5512 ) );
  nor_x1_sg U62248 ( .A(\filter_0/reg_w_5[7] ), .B(n31789), .X(
        \filter_0/n5508 ) );
  nor_x1_sg U62249 ( .A(\filter_0/reg_w_5[6] ), .B(n31790), .X(
        \filter_0/n5504 ) );
  nor_x1_sg U62250 ( .A(\filter_0/reg_w_5[5] ), .B(n34295), .X(
        \filter_0/n5500 ) );
  nor_x1_sg U62251 ( .A(\filter_0/reg_w_5[4] ), .B(n34297), .X(
        \filter_0/n5496 ) );
  nor_x1_sg U62252 ( .A(\filter_0/reg_w_5[3] ), .B(n31360), .X(
        \filter_0/n5492 ) );
  nor_x1_sg U62253 ( .A(\filter_0/reg_w_5[2] ), .B(n34296), .X(
        \filter_0/n5488 ) );
  nor_x1_sg U62254 ( .A(\filter_0/reg_w_5[1] ), .B(n31789), .X(
        \filter_0/n5484 ) );
  nor_x1_sg U62255 ( .A(\filter_0/reg_w_5[0] ), .B(n34295), .X(
        \filter_0/n5480 ) );
  nor_x1_sg U62256 ( .A(\filter_0/reg_w_6[19] ), .B(n29747), .X(
        \filter_0/n5476 ) );
  nor_x1_sg U62257 ( .A(\filter_0/reg_w_6[18] ), .B(n31453), .X(
        \filter_0/n5472 ) );
  nor_x1_sg U62258 ( .A(\filter_0/reg_w_6[17] ), .B(n34142), .X(
        \filter_0/n5468 ) );
  nor_x1_sg U62259 ( .A(\filter_0/reg_w_6[16] ), .B(n30259), .X(
        \filter_0/n5464 ) );
  nor_x1_sg U62260 ( .A(\filter_0/reg_w_6[15] ), .B(n31845), .X(
        \filter_0/n5460 ) );
  nor_x1_sg U62261 ( .A(\filter_0/reg_w_6[14] ), .B(n31844), .X(
        \filter_0/n5456 ) );
  nor_x1_sg U62262 ( .A(\filter_0/reg_w_6[13] ), .B(n30259), .X(
        \filter_0/n5452 ) );
  nor_x1_sg U62263 ( .A(\filter_0/reg_w_6[12] ), .B(n34139), .X(
        \filter_0/n5448 ) );
  nor_x1_sg U62264 ( .A(\filter_0/reg_w_6[11] ), .B(n34139), .X(
        \filter_0/n5444 ) );
  nor_x1_sg U62265 ( .A(\filter_0/reg_w_6[10] ), .B(n34142), .X(
        \filter_0/n5440 ) );
  nor_x1_sg U62266 ( .A(\filter_0/reg_w_6[9] ), .B(n30259), .X(
        \filter_0/n5436 ) );
  nor_x1_sg U62267 ( .A(\filter_0/reg_w_6[8] ), .B(n34142), .X(
        \filter_0/n5432 ) );
  nor_x1_sg U62268 ( .A(\filter_0/reg_w_6[7] ), .B(n31453), .X(
        \filter_0/n5428 ) );
  nor_x1_sg U62269 ( .A(\filter_0/reg_w_6[6] ), .B(n15180), .X(
        \filter_0/n5424 ) );
  nor_x1_sg U62270 ( .A(\filter_0/reg_w_6[5] ), .B(n34141), .X(
        \filter_0/n5420 ) );
  nor_x1_sg U62271 ( .A(\filter_0/reg_w_6[4] ), .B(n31844), .X(
        \filter_0/n5416 ) );
  nor_x1_sg U62272 ( .A(\filter_0/reg_w_6[3] ), .B(n31844), .X(
        \filter_0/n5412 ) );
  nor_x1_sg U62273 ( .A(\filter_0/reg_w_6[2] ), .B(n34142), .X(
        \filter_0/n5408 ) );
  nor_x1_sg U62274 ( .A(\filter_0/reg_w_6[1] ), .B(n34140), .X(
        \filter_0/n5404 ) );
  nor_x1_sg U62275 ( .A(\filter_0/reg_w_6[0] ), .B(n31845), .X(
        \filter_0/n5400 ) );
  nor_x1_sg U62276 ( .A(\filter_0/reg_w_7[19] ), .B(n31455), .X(
        \filter_0/n5396 ) );
  nor_x1_sg U62277 ( .A(\filter_0/reg_w_7[18] ), .B(n31455), .X(
        \filter_0/n5392 ) );
  nor_x1_sg U62278 ( .A(\filter_0/reg_w_7[17] ), .B(n30257), .X(
        \filter_0/n5388 ) );
  nor_x1_sg U62279 ( .A(\filter_0/reg_w_7[16] ), .B(n31456), .X(
        \filter_0/n5384 ) );
  nor_x1_sg U62280 ( .A(\filter_0/reg_w_7[15] ), .B(n31847), .X(
        \filter_0/n5380 ) );
  nor_x1_sg U62281 ( .A(\filter_0/reg_w_7[14] ), .B(n31455), .X(
        \filter_0/n5376 ) );
  nor_x1_sg U62282 ( .A(\filter_0/reg_w_7[13] ), .B(n30257), .X(
        \filter_0/n5372 ) );
  nor_x1_sg U62283 ( .A(\filter_0/reg_w_7[12] ), .B(n34134), .X(
        \filter_0/n5368 ) );
  nor_x1_sg U62284 ( .A(\filter_0/reg_w_7[11] ), .B(n31456), .X(
        \filter_0/n5364 ) );
  nor_x1_sg U62285 ( .A(\filter_0/reg_w_7[10] ), .B(n34137), .X(
        \filter_0/n5360 ) );
  nor_x1_sg U62286 ( .A(\filter_0/reg_w_7[9] ), .B(n31456), .X(
        \filter_0/n5356 ) );
  nor_x1_sg U62287 ( .A(\filter_0/reg_w_7[8] ), .B(n31456), .X(
        \filter_0/n5352 ) );
  nor_x1_sg U62288 ( .A(\filter_0/reg_w_7[7] ), .B(n15181), .X(
        \filter_0/n5348 ) );
  nor_x1_sg U62289 ( .A(\filter_0/reg_w_7[6] ), .B(n34134), .X(
        \filter_0/n5344 ) );
  nor_x1_sg U62290 ( .A(\filter_0/reg_w_7[5] ), .B(n30062), .X(
        \filter_0/n5340 ) );
  nor_x1_sg U62291 ( .A(\filter_0/reg_w_7[4] ), .B(n31846), .X(
        \filter_0/n5336 ) );
  nor_x1_sg U62292 ( .A(\filter_0/reg_w_7[3] ), .B(n31846), .X(
        \filter_0/n5332 ) );
  nor_x1_sg U62293 ( .A(\filter_0/reg_w_7[2] ), .B(n34137), .X(
        \filter_0/n5328 ) );
  nor_x1_sg U62294 ( .A(\filter_0/reg_w_7[1] ), .B(n34135), .X(
        \filter_0/n5324 ) );
  nor_x1_sg U62295 ( .A(\filter_0/reg_w_7[0] ), .B(n31847), .X(
        \filter_0/n5320 ) );
  nor_x1_sg U62296 ( .A(\filter_0/reg_w_0[19] ), .B(n29742), .X(
        \filter_0/n5316 ) );
  nor_x1_sg U62297 ( .A(\filter_0/reg_w_0[18] ), .B(n31437), .X(
        \filter_0/n5312 ) );
  nor_x1_sg U62298 ( .A(\filter_0/reg_w_0[17] ), .B(n31834), .X(
        \filter_0/n5308 ) );
  nor_x1_sg U62299 ( .A(\filter_0/reg_w_0[16] ), .B(n34164), .X(
        \filter_0/n5304 ) );
  nor_x1_sg U62300 ( .A(\filter_0/reg_w_0[15] ), .B(n30068), .X(
        \filter_0/n5300 ) );
  nor_x1_sg U62301 ( .A(\filter_0/reg_w_0[14] ), .B(n34167), .X(
        \filter_0/n5296 ) );
  nor_x1_sg U62302 ( .A(\filter_0/reg_w_0[13] ), .B(n34165), .X(
        \filter_0/n5292 ) );
  nor_x1_sg U62303 ( .A(\filter_0/reg_w_0[12] ), .B(n31438), .X(
        \filter_0/n5288 ) );
  nor_x1_sg U62304 ( .A(\filter_0/reg_w_0[11] ), .B(n34166), .X(
        \filter_0/n5284 ) );
  nor_x1_sg U62305 ( .A(\filter_0/reg_w_0[10] ), .B(n31834), .X(
        \filter_0/n5280 ) );
  nor_x1_sg U62306 ( .A(\filter_0/reg_w_0[9] ), .B(n34165), .X(
        \filter_0/n5276 ) );
  nor_x1_sg U62307 ( .A(\filter_0/reg_w_0[8] ), .B(n31835), .X(
        \filter_0/n5272 ) );
  nor_x1_sg U62308 ( .A(\filter_0/reg_w_0[7] ), .B(n29742), .X(
        \filter_0/n5268 ) );
  nor_x1_sg U62309 ( .A(\filter_0/reg_w_0[6] ), .B(n30269), .X(
        \filter_0/n5264 ) );
  nor_x1_sg U62310 ( .A(\filter_0/reg_w_0[5] ), .B(n34164), .X(
        \filter_0/n5260 ) );
  nor_x1_sg U62311 ( .A(\filter_0/reg_w_0[4] ), .B(n31438), .X(
        \filter_0/n5256 ) );
  nor_x1_sg U62312 ( .A(\filter_0/reg_w_0[3] ), .B(n34166), .X(
        \filter_0/n5252 ) );
  nor_x1_sg U62313 ( .A(\filter_0/reg_w_0[2] ), .B(n31438), .X(
        \filter_0/n5248 ) );
  nor_x1_sg U62314 ( .A(\filter_0/reg_w_0[1] ), .B(n34164), .X(
        \filter_0/n5244 ) );
  nor_x1_sg U62315 ( .A(\filter_0/reg_w_0[0] ), .B(n15182), .X(
        \filter_0/n5240 ) );
  nor_x1_sg U62316 ( .A(\filter_0/reg_w_1[19] ), .B(n34291), .X(
        \filter_0/n5236 ) );
  nor_x1_sg U62317 ( .A(\filter_0/reg_w_1[18] ), .B(n31792), .X(
        \filter_0/n5232 ) );
  nor_x1_sg U62318 ( .A(\filter_0/reg_w_1[17] ), .B(n31363), .X(
        \filter_0/n5228 ) );
  nor_x1_sg U62319 ( .A(\filter_0/reg_w_1[16] ), .B(n34291), .X(
        \filter_0/n5224 ) );
  nor_x1_sg U62320 ( .A(\filter_0/reg_w_1[15] ), .B(n34292), .X(
        \filter_0/n5220 ) );
  nor_x1_sg U62321 ( .A(\filter_0/reg_w_1[14] ), .B(n31362), .X(
        \filter_0/n5216 ) );
  nor_x1_sg U62322 ( .A(\filter_0/reg_w_1[13] ), .B(n34290), .X(
        \filter_0/n5212 ) );
  nor_x1_sg U62323 ( .A(\filter_0/reg_w_1[12] ), .B(n31362), .X(
        \filter_0/n5208 ) );
  nor_x1_sg U62324 ( .A(\filter_0/reg_w_1[11] ), .B(n34290), .X(
        \filter_0/n5204 ) );
  nor_x1_sg U62325 ( .A(\filter_0/reg_w_1[10] ), .B(n31363), .X(
        \filter_0/n5200 ) );
  nor_x1_sg U62326 ( .A(\filter_0/reg_w_1[9] ), .B(n30326), .X(
        \filter_0/n5196 ) );
  nor_x1_sg U62327 ( .A(\filter_0/reg_w_1[8] ), .B(n31362), .X(
        \filter_0/n5192 ) );
  nor_x1_sg U62328 ( .A(\filter_0/reg_w_1[7] ), .B(n34289), .X(
        \filter_0/n5188 ) );
  nor_x1_sg U62329 ( .A(\filter_0/reg_w_1[6] ), .B(n31362), .X(
        \filter_0/n5184 ) );
  nor_x1_sg U62330 ( .A(\filter_0/reg_w_1[5] ), .B(n15184), .X(
        \filter_0/n5180 ) );
  nor_x1_sg U62331 ( .A(\filter_0/reg_w_1[4] ), .B(n34290), .X(
        \filter_0/n5176 ) );
  nor_x1_sg U62332 ( .A(\filter_0/reg_w_1[3] ), .B(n30326), .X(
        \filter_0/n5172 ) );
  nor_x1_sg U62333 ( .A(\filter_0/reg_w_1[2] ), .B(n34289), .X(
        \filter_0/n5168 ) );
  nor_x1_sg U62334 ( .A(\filter_0/reg_w_1[1] ), .B(n31792), .X(
        \filter_0/n5164 ) );
  nor_x1_sg U62335 ( .A(\filter_0/reg_w_1[0] ), .B(n31792), .X(
        \filter_0/n5160 ) );
  nor_x1_sg U62336 ( .A(\filter_0/reg_w_2[19] ), .B(n34340), .X(
        \filter_0/n5156 ) );
  nor_x1_sg U62337 ( .A(\filter_0/reg_w_2[18] ), .B(n34339), .X(
        \filter_0/n5152 ) );
  nor_x1_sg U62338 ( .A(\filter_0/reg_w_2[17] ), .B(n30346), .X(
        \filter_0/n5148 ) );
  nor_x1_sg U62339 ( .A(\filter_0/reg_w_2[16] ), .B(n34340), .X(
        \filter_0/n5144 ) );
  nor_x1_sg U62340 ( .A(\filter_0/reg_w_2[15] ), .B(n31771), .X(
        \filter_0/n5140 ) );
  nor_x1_sg U62341 ( .A(\filter_0/reg_w_2[14] ), .B(n34340), .X(
        \filter_0/n5136 ) );
  nor_x1_sg U62342 ( .A(\filter_0/reg_w_2[13] ), .B(n31771), .X(
        \filter_0/n5132 ) );
  nor_x1_sg U62343 ( .A(\filter_0/reg_w_2[12] ), .B(n34340), .X(
        \filter_0/n5128 ) );
  nor_x1_sg U62344 ( .A(\filter_0/reg_w_2[11] ), .B(n31771), .X(
        \filter_0/n5124 ) );
  nor_x1_sg U62345 ( .A(\filter_0/reg_w_2[10] ), .B(n34342), .X(
        \filter_0/n5120 ) );
  nor_x1_sg U62346 ( .A(\filter_0/reg_w_2[9] ), .B(n31332), .X(
        \filter_0/n5116 ) );
  nor_x1_sg U62347 ( .A(\filter_0/reg_w_2[8] ), .B(n31333), .X(
        \filter_0/n5112 ) );
  nor_x1_sg U62348 ( .A(\filter_0/reg_w_2[7] ), .B(n15187), .X(
        \filter_0/n5108 ) );
  nor_x1_sg U62349 ( .A(\filter_0/reg_w_2[6] ), .B(n31332), .X(
        \filter_0/n5104 ) );
  nor_x1_sg U62350 ( .A(\filter_0/reg_w_2[5] ), .B(n34339), .X(
        \filter_0/n5100 ) );
  nor_x1_sg U62351 ( .A(\filter_0/reg_w_2[4] ), .B(n30346), .X(
        \filter_0/n5096 ) );
  nor_x1_sg U62352 ( .A(\filter_0/reg_w_2[3] ), .B(n34342), .X(
        \filter_0/n5092 ) );
  nor_x1_sg U62353 ( .A(\filter_0/reg_w_2[2] ), .B(n31771), .X(
        \filter_0/n5088 ) );
  nor_x1_sg U62354 ( .A(\filter_0/reg_w_2[1] ), .B(n34341), .X(
        \filter_0/n5084 ) );
  nor_x1_sg U62355 ( .A(\filter_0/reg_w_2[0] ), .B(n34342), .X(
        \filter_0/n5080 ) );
  nor_x1_sg U62356 ( .A(\filter_0/reg_w_3[19] ), .B(n31440), .X(
        \filter_0/n5076 ) );
  nor_x1_sg U62357 ( .A(\filter_0/reg_w_3[18] ), .B(n31440), .X(
        \filter_0/n5072 ) );
  nor_x1_sg U62358 ( .A(\filter_0/reg_w_3[17] ), .B(n34159), .X(
        \filter_0/n5068 ) );
  nor_x1_sg U62359 ( .A(\filter_0/reg_w_3[16] ), .B(n31836), .X(
        \filter_0/n5064 ) );
  nor_x1_sg U62360 ( .A(\filter_0/reg_w_3[15] ), .B(n31441), .X(
        \filter_0/n5060 ) );
  nor_x1_sg U62361 ( .A(\filter_0/reg_w_3[14] ), .B(n31837), .X(
        \filter_0/n5056 ) );
  nor_x1_sg U62362 ( .A(\filter_0/reg_w_3[13] ), .B(n34161), .X(
        \filter_0/n5052 ) );
  nor_x1_sg U62363 ( .A(\filter_0/reg_w_3[12] ), .B(n34159), .X(
        \filter_0/n5048 ) );
  nor_x1_sg U62364 ( .A(\filter_0/reg_w_3[11] ), .B(n29743), .X(
        \filter_0/n5044 ) );
  nor_x1_sg U62365 ( .A(\filter_0/reg_w_3[10] ), .B(n31440), .X(
        \filter_0/n5040 ) );
  nor_x1_sg U62366 ( .A(\filter_0/reg_w_3[9] ), .B(n34162), .X(
        \filter_0/n5036 ) );
  nor_x1_sg U62367 ( .A(\filter_0/reg_w_3[8] ), .B(n34162), .X(
        \filter_0/n5032 ) );
  nor_x1_sg U62368 ( .A(\filter_0/reg_w_3[7] ), .B(n31837), .X(
        \filter_0/n5028 ) );
  nor_x1_sg U62369 ( .A(\filter_0/reg_w_3[6] ), .B(n30067), .X(
        \filter_0/n5024 ) );
  nor_x1_sg U62370 ( .A(\filter_0/reg_w_3[5] ), .B(n34161), .X(
        \filter_0/n5020 ) );
  nor_x1_sg U62371 ( .A(\filter_0/reg_w_3[4] ), .B(n15190), .X(
        \filter_0/n5016 ) );
  nor_x1_sg U62372 ( .A(\filter_0/reg_w_3[3] ), .B(n34162), .X(
        \filter_0/n5012 ) );
  nor_x1_sg U62373 ( .A(\filter_0/reg_w_3[2] ), .B(n34159), .X(
        \filter_0/n5008 ) );
  nor_x1_sg U62374 ( .A(\filter_0/reg_w_3[1] ), .B(n34161), .X(
        \filter_0/n5004 ) );
  nor_x1_sg U62375 ( .A(\filter_0/reg_w_3[0] ), .B(n30267), .X(
        \filter_0/n5000 ) );
  nand_x1_sg U62376 ( .A(\shifter_0/reg_w_14[0] ), .B(n32194), .X(n11904) );
  nand_x1_sg U62377 ( .A(\shifter_0/reg_w_15[0] ), .B(n34438), .X(n11903) );
  nand_x1_sg U62378 ( .A(\shifter_0/reg_w_14[1] ), .B(n34442), .X(n11916) );
  nand_x1_sg U62379 ( .A(\shifter_0/reg_w_15[1] ), .B(n34439), .X(n11915) );
  nand_x1_sg U62380 ( .A(\shifter_0/reg_w_14[4] ), .B(n34443), .X(n11949) );
  nand_x1_sg U62381 ( .A(\shifter_0/reg_w_15[4] ), .B(n30839), .X(n11948) );
  nand_x1_sg U62382 ( .A(\shifter_0/reg_w_14[7] ), .B(n34444), .X(n11982) );
  nand_x1_sg U62383 ( .A(\shifter_0/reg_w_15[7] ), .B(n31976), .X(n11981) );
  nand_x1_sg U62384 ( .A(\shifter_0/reg_w_14[10] ), .B(n32195), .X(n12015) );
  nand_x1_sg U62385 ( .A(\shifter_0/reg_w_15[10] ), .B(n30840), .X(n12014) );
  nand_x1_sg U62386 ( .A(\shifter_0/reg_w_14[13] ), .B(n32194), .X(n12048) );
  nand_x1_sg U62387 ( .A(\shifter_0/reg_w_15[13] ), .B(n31978), .X(n12047) );
  nand_x1_sg U62388 ( .A(\shifter_0/reg_w_14[14] ), .B(n30837), .X(n12059) );
  nand_x1_sg U62389 ( .A(\shifter_0/reg_w_15[14] ), .B(n34438), .X(n12058) );
  nand_x1_sg U62390 ( .A(\shifter_0/reg_w_14[15] ), .B(n34443), .X(n12070) );
  nand_x1_sg U62391 ( .A(\shifter_0/reg_w_15[15] ), .B(n34440), .X(n12069) );
  nand_x1_sg U62392 ( .A(\shifter_0/reg_w_14[18] ), .B(n30838), .X(n12103) );
  nand_x1_sg U62393 ( .A(\shifter_0/reg_w_15[18] ), .B(n31975), .X(n12102) );
  nand_x1_sg U62394 ( .A(\shifter_0/reg_w_14[19] ), .B(n32197), .X(n12114) );
  nand_x1_sg U62395 ( .A(\shifter_0/reg_w_15[19] ), .B(n34439), .X(n12113) );
  nand_x1_sg U62396 ( .A(\shifter_0/reg_i_14[0] ), .B(n32192), .X(n12132) );
  nand_x1_sg U62397 ( .A(\shifter_0/reg_i_15[0] ), .B(n34438), .X(n12131) );
  nand_x1_sg U62398 ( .A(\shifter_0/reg_i_14[1] ), .B(n30837), .X(n12144) );
  nand_x1_sg U62399 ( .A(\shifter_0/reg_i_15[1] ), .B(n34439), .X(n12143) );
  nand_x1_sg U62400 ( .A(\shifter_0/reg_i_14[7] ), .B(n34442), .X(n12210) );
  nand_x1_sg U62401 ( .A(\shifter_0/reg_i_15[7] ), .B(n31975), .X(n12209) );
  nand_x1_sg U62402 ( .A(\shifter_0/reg_i_14[10] ), .B(n32192), .X(n12243) );
  nand_x1_sg U62403 ( .A(\shifter_0/reg_i_15[10] ), .B(n30840), .X(n12242) );
  nand_x1_sg U62404 ( .A(\shifter_0/reg_i_14[13] ), .B(n34443), .X(n12276) );
  nand_x1_sg U62405 ( .A(\shifter_0/reg_i_15[13] ), .B(n31976), .X(n12275) );
  nand_x1_sg U62406 ( .A(\shifter_0/reg_i_14[14] ), .B(n32196), .X(n12287) );
  nand_x1_sg U62407 ( .A(\shifter_0/reg_i_15[14] ), .B(n34437), .X(n12286) );
  nand_x1_sg U62408 ( .A(\shifter_0/reg_i_14[15] ), .B(n30838), .X(n12298) );
  nand_x1_sg U62409 ( .A(\shifter_0/reg_i_15[15] ), .B(n31980), .X(n12297) );
  nand_x1_sg U62410 ( .A(\shifter_0/reg_i_14[19] ), .B(n34444), .X(n12342) );
  nand_x1_sg U62411 ( .A(\shifter_0/reg_i_15[19] ), .B(n30839), .X(n12341) );
  nand_x1_sg U62412 ( .A(n31119), .B(n35565), .X(n15063) );
  nor_x1_sg U62413 ( .A(n35565), .B(n31119), .X(n15064) );
  nand_x1_sg U62414 ( .A(n31124), .B(n35564), .X(n15199) );
  nor_x1_sg U62415 ( .A(n35564), .B(n31124), .X(n15200) );
  nand_x1_sg U62416 ( .A(n35097), .B(n35257), .X(n15077) );
  nand_x1_sg U62417 ( .A(n31121), .B(n15068), .X(n15078) );
  nand_x1_sg U62418 ( .A(n34225), .B(\shifter_0/reg_i_7[2] ), .X(n12629) );
  nor_x1_sg U62419 ( .A(n12630), .B(n12631), .X(n12628) );
  nor_x1_sg U62420 ( .A(n31810), .B(n41068), .X(n12631) );
  nor_x1_sg U62421 ( .A(n12639), .B(n12640), .X(n12637) );
  nand_x1_sg U62422 ( .A(n30080), .B(n31131), .X(n12638) );
  nor_x1_sg U62423 ( .A(n31810), .B(n42597), .X(n12640) );
  nand_x1_sg U62424 ( .A(n34226), .B(\shifter_0/reg_i_7[17] ), .X(n12691) );
  nor_x1_sg U62425 ( .A(n12692), .B(n12693), .X(n12690) );
  nor_x1_sg U62426 ( .A(n31809), .B(n42602), .X(n12693) );
  nand_x1_sg U62427 ( .A(n34225), .B(\shifter_0/reg_i_7[18] ), .X(n12696) );
  nor_x1_sg U62428 ( .A(n12697), .B(n12698), .X(n12695) );
  nor_x1_sg U62429 ( .A(n34235), .B(n42603), .X(n12698) );
  nand_x1_sg U62430 ( .A(\shifter_0/reg_i_14[2] ), .B(n32196), .X(n12155) );
  nand_x1_sg U62431 ( .A(\shifter_0/reg_i_15[2] ), .B(n34440), .X(n12154) );
  nand_x1_sg U62432 ( .A(\shifter_0/reg_i_14[17] ), .B(n32196), .X(n12320) );
  nand_x1_sg U62433 ( .A(\shifter_0/reg_i_15[17] ), .B(n34437), .X(n12319) );
  nor_x1_sg U62434 ( .A(n15099), .B(n15100), .X(n15098) );
  nor_x1_sg U62435 ( .A(n32505), .B(\filter_0/reg_xor_i_mask[7] ), .X(n15099)
         );
  nor_x1_sg U62436 ( .A(n32136), .B(\filter_0/reg_xor_i_mask[6] ), .X(n15100)
         );
  nor_x1_sg U62437 ( .A(n15102), .B(n15103), .X(n15097) );
  nor_x1_sg U62438 ( .A(n32206), .B(\filter_0/reg_xor_i_mask[3] ), .X(n15102)
         );
  nor_x1_sg U62439 ( .A(n32116), .B(\filter_0/reg_xor_i_mask[5] ), .X(n15103)
         );
  nor_x1_sg U62440 ( .A(n15231), .B(n15232), .X(n15230) );
  nor_x1_sg U62441 ( .A(n32504), .B(\filter_0/reg_xor_w_mask[7] ), .X(n15231)
         );
  nor_x1_sg U62442 ( .A(n32136), .B(\filter_0/reg_xor_w_mask[6] ), .X(n15232)
         );
  nor_x1_sg U62443 ( .A(n15233), .B(n15234), .X(n15229) );
  nor_x1_sg U62444 ( .A(n32207), .B(\filter_0/reg_xor_w_mask[3] ), .X(n15233)
         );
  nor_x1_sg U62445 ( .A(n32114), .B(\filter_0/reg_xor_w_mask[5] ), .X(n15234)
         );
  nand_x1_sg U62446 ( .A(n32172), .B(n14033), .X(n14032) );
  nand_x1_sg U62447 ( .A(n34411), .B(n40900), .X(n14033) );
  inv_x1_sg U62448 ( .A(\shifter_0/reg_w_11[7] ), .X(n40900) );
  nand_x1_sg U62449 ( .A(n31300), .B(n14312), .X(n14311) );
  nand_x1_sg U62450 ( .A(n30114), .B(n40895), .X(n14312) );
  inv_x1_sg U62451 ( .A(\shifter_0/reg_w_11[16] ), .X(n40895) );
  nand_x1_sg U62452 ( .A(n34550), .B(n14468), .X(n14467) );
  nand_x1_sg U62453 ( .A(n30855), .B(n41028), .X(n14468) );
  inv_x1_sg U62454 ( .A(\shifter_0/reg_i_11[1] ), .X(n41028) );
  nand_x1_sg U62455 ( .A(n31299), .B(n14656), .X(n14655) );
  nand_x1_sg U62456 ( .A(n30114), .B(n41024), .X(n14656) );
  inv_x1_sg U62457 ( .A(\shifter_0/reg_i_11[7] ), .X(n41024) );
  nand_x1_sg U62458 ( .A(n34548), .B(n15028), .X(n15027) );
  nand_x1_sg U62459 ( .A(n31992), .B(n41019), .X(n15028) );
  inv_x1_sg U62460 ( .A(\shifter_0/reg_i_11[19] ), .X(n41019) );
  nor_x1_sg U62461 ( .A(n15149), .B(n42373), .X(n15148) );
  nor_x1_sg U62462 ( .A(\filter_0/reg_xor_i_mask[28] ), .B(n32131), .X(n15149)
         );
  nor_x1_sg U62463 ( .A(n15151), .B(n15152), .X(n15150) );
  nor_x1_sg U62464 ( .A(n15116), .B(n42372), .X(n15115) );
  nor_x1_sg U62465 ( .A(\filter_0/reg_xor_i_mask[12] ), .B(n32131), .X(n15116)
         );
  nor_x1_sg U62466 ( .A(n15118), .B(n15119), .X(n15117) );
  nor_x1_sg U62467 ( .A(n15278), .B(n42375), .X(n15277) );
  nor_x1_sg U62468 ( .A(\filter_0/reg_xor_w_mask[28] ), .B(n32131), .X(n15278)
         );
  nor_x1_sg U62469 ( .A(n15280), .B(n15281), .X(n15279) );
  nor_x1_sg U62470 ( .A(n15245), .B(n42374), .X(n15244) );
  nor_x1_sg U62471 ( .A(\filter_0/reg_xor_w_mask[12] ), .B(n32132), .X(n15245)
         );
  nor_x1_sg U62472 ( .A(n15247), .B(n15248), .X(n15246) );
  nor_x1_sg U62473 ( .A(n15153), .B(n15154), .X(n15147) );
  nor_x1_sg U62474 ( .A(\filter_0/reg_xor_i_mask[25] ), .B(n32118), .X(n15153)
         );
  nor_x1_sg U62475 ( .A(\filter_0/reg_xor_i_mask[29] ), .B(n32115), .X(n15154)
         );
  nor_x1_sg U62476 ( .A(n15111), .B(n15112), .X(n15110) );
  nor_x1_sg U62477 ( .A(\filter_0/reg_xor_i_mask[11] ), .B(n32208), .X(n15111)
         );
  nor_x1_sg U62478 ( .A(\filter_0/reg_xor_i_mask[14] ), .B(n32134), .X(n15112)
         );
  nor_x1_sg U62479 ( .A(n15120), .B(n15121), .X(n15114) );
  nor_x1_sg U62480 ( .A(\filter_0/reg_xor_i_mask[9] ), .B(n32119), .X(n15120)
         );
  nor_x1_sg U62481 ( .A(\filter_0/reg_xor_i_mask[13] ), .B(n32116), .X(n15121)
         );
  nor_x1_sg U62482 ( .A(n15282), .B(n15283), .X(n15276) );
  nor_x1_sg U62483 ( .A(\filter_0/reg_xor_w_mask[25] ), .B(n32119), .X(n15282)
         );
  nor_x1_sg U62484 ( .A(\filter_0/reg_xor_w_mask[29] ), .B(n32115), .X(n15283)
         );
  nor_x1_sg U62485 ( .A(n15240), .B(n15241), .X(n15239) );
  nor_x1_sg U62486 ( .A(\filter_0/reg_xor_w_mask[11] ), .B(n32208), .X(n15240)
         );
  nor_x1_sg U62487 ( .A(\filter_0/reg_xor_w_mask[14] ), .B(n32135), .X(n15241)
         );
  nor_x1_sg U62488 ( .A(n15249), .B(n15250), .X(n15243) );
  nor_x1_sg U62489 ( .A(\filter_0/reg_xor_w_mask[9] ), .B(n32119), .X(n15249)
         );
  nor_x1_sg U62490 ( .A(\filter_0/reg_xor_w_mask[13] ), .B(n32116), .X(n15250)
         );
  nand_x1_sg U62491 ( .A(n31880), .B(n30584), .X(n15211) );
  nand_x1_sg U62492 ( .A(n31657), .B(n35305), .X(n15210) );
  inv_x1_sg U62493 ( .A(\shifter_0/reg_w_14[0] ), .X(n40869) );
  inv_x1_sg U62494 ( .A(\shifter_0/reg_w_14[1] ), .X(n40868) );
  inv_x1_sg U62495 ( .A(\shifter_0/reg_w_14[2] ), .X(n40867) );
  inv_x1_sg U62496 ( .A(\shifter_0/reg_w_14[5] ), .X(n40866) );
  inv_x1_sg U62497 ( .A(\shifter_0/reg_w_14[6] ), .X(n40865) );
  inv_x1_sg U62498 ( .A(\shifter_0/reg_w_14[7] ), .X(n40864) );
  inv_x1_sg U62499 ( .A(\shifter_0/reg_w_14[10] ), .X(n40863) );
  inv_x1_sg U62500 ( .A(\shifter_0/reg_w_14[11] ), .X(n40862) );
  inv_x1_sg U62501 ( .A(\shifter_0/reg_w_14[14] ), .X(n40861) );
  inv_x1_sg U62502 ( .A(\shifter_0/reg_w_14[15] ), .X(n40860) );
  inv_x1_sg U62503 ( .A(\shifter_0/reg_w_14[16] ), .X(n40859) );
  inv_x1_sg U62504 ( .A(\shifter_0/reg_w_14[19] ), .X(n40858) );
  inv_x1_sg U62505 ( .A(\shifter_0/reg_i_14[0] ), .X(n40996) );
  inv_x1_sg U62506 ( .A(\shifter_0/reg_i_14[1] ), .X(n40995) );
  inv_x1_sg U62507 ( .A(\shifter_0/reg_i_14[3] ), .X(n40994) );
  inv_x1_sg U62508 ( .A(\shifter_0/reg_i_14[5] ), .X(n40993) );
  inv_x1_sg U62509 ( .A(\shifter_0/reg_i_14[6] ), .X(n40992) );
  inv_x1_sg U62510 ( .A(\shifter_0/reg_i_14[7] ), .X(n40991) );
  inv_x1_sg U62511 ( .A(\shifter_0/reg_i_14[10] ), .X(n40990) );
  inv_x1_sg U62512 ( .A(\shifter_0/reg_i_14[11] ), .X(n40989) );
  inv_x1_sg U62513 ( .A(\shifter_0/reg_i_14[14] ), .X(n40988) );
  inv_x1_sg U62514 ( .A(\shifter_0/reg_i_14[15] ), .X(n40987) );
  inv_x1_sg U62515 ( .A(\shifter_0/reg_i_14[19] ), .X(n40986) );
  nor_x1_sg U62516 ( .A(n35614), .B(n12532), .X(n12529) );
  nand_x1_sg U62517 ( .A(n34227), .B(n31161), .X(n12530) );
  nor_x1_sg U62518 ( .A(n34236), .B(n40949), .X(n12532) );
  nor_x1_sg U62519 ( .A(n35561), .B(n12537), .X(n12535) );
  nand_x1_sg U62520 ( .A(n34227), .B(n31163), .X(n12536) );
  nor_x1_sg U62521 ( .A(n34234), .B(n40947), .X(n12537) );
  nor_x1_sg U62522 ( .A(n35613), .B(n12541), .X(n12539) );
  nand_x1_sg U62523 ( .A(n34226), .B(n31165), .X(n12540) );
  nor_x1_sg U62524 ( .A(n31395), .B(n40945), .X(n12541) );
  nor_x1_sg U62525 ( .A(n35509), .B(n12545), .X(n12543) );
  nand_x1_sg U62526 ( .A(n31813), .B(n31167), .X(n12544) );
  nor_x1_sg U62527 ( .A(n34237), .B(n42706), .X(n12545) );
  nor_x1_sg U62528 ( .A(n35604), .B(n12549), .X(n12547) );
  nand_x1_sg U62529 ( .A(n30297), .B(n31169), .X(n12548) );
  nor_x1_sg U62530 ( .A(n30300), .B(n42707), .X(n12549) );
  nor_x1_sg U62531 ( .A(n35619), .B(n12553), .X(n12551) );
  nand_x1_sg U62532 ( .A(n31402), .B(n31171), .X(n12552) );
  nor_x1_sg U62533 ( .A(n34234), .B(n40941), .X(n12553) );
  nor_x1_sg U62534 ( .A(n35514), .B(n12557), .X(n12555) );
  nand_x1_sg U62535 ( .A(n34224), .B(n31173), .X(n12556) );
  nor_x1_sg U62536 ( .A(n34235), .B(n40939), .X(n12557) );
  nor_x1_sg U62537 ( .A(n35618), .B(n12561), .X(n12559) );
  nand_x1_sg U62538 ( .A(n31401), .B(n31175), .X(n12560) );
  nor_x1_sg U62539 ( .A(n31809), .B(n40937), .X(n12561) );
  nor_x1_sg U62540 ( .A(n35612), .B(n12565), .X(n12563) );
  nand_x1_sg U62541 ( .A(n34224), .B(n31177), .X(n12564) );
  nor_x1_sg U62542 ( .A(n12533), .B(n42708), .X(n12565) );
  nor_x1_sg U62543 ( .A(n35617), .B(n12569), .X(n12567) );
  nand_x1_sg U62544 ( .A(n30295), .B(n31179), .X(n12568) );
  nor_x1_sg U62545 ( .A(n29731), .B(n42709), .X(n12569) );
  nor_x1_sg U62546 ( .A(n35602), .B(n12573), .X(n12571) );
  nand_x1_sg U62547 ( .A(n31401), .B(n31181), .X(n12572) );
  nor_x1_sg U62548 ( .A(n30082), .B(n40933), .X(n12573) );
  nor_x1_sg U62549 ( .A(n35616), .B(n12577), .X(n12575) );
  nand_x1_sg U62550 ( .A(n30295), .B(n31183), .X(n12576) );
  nor_x1_sg U62551 ( .A(n31809), .B(n40931), .X(n12577) );
  nor_x1_sg U62552 ( .A(n35611), .B(n12581), .X(n12579) );
  nand_x1_sg U62553 ( .A(n34227), .B(n31185), .X(n12580) );
  nor_x1_sg U62554 ( .A(n30082), .B(n42710), .X(n12581) );
  nor_x1_sg U62555 ( .A(n35615), .B(n12585), .X(n12583) );
  nand_x1_sg U62556 ( .A(n30295), .B(n31187), .X(n12584) );
  nor_x1_sg U62557 ( .A(n34237), .B(n42711), .X(n12585) );
  nor_x1_sg U62558 ( .A(n35610), .B(n12589), .X(n12587) );
  nand_x1_sg U62559 ( .A(n30080), .B(n31189), .X(n12588) );
  nor_x1_sg U62560 ( .A(n31395), .B(n40927), .X(n12589) );
  nor_x1_sg U62561 ( .A(n35609), .B(n12593), .X(n12591) );
  nand_x1_sg U62562 ( .A(n31401), .B(n31191), .X(n12592) );
  nor_x1_sg U62563 ( .A(n30300), .B(n40925), .X(n12593) );
  nor_x1_sg U62564 ( .A(n35601), .B(n12597), .X(n12595) );
  nand_x1_sg U62565 ( .A(n34225), .B(n31193), .X(n12596) );
  nor_x1_sg U62566 ( .A(n31396), .B(n40923), .X(n12597) );
  nor_x1_sg U62567 ( .A(n35608), .B(n12601), .X(n12599) );
  nand_x1_sg U62568 ( .A(n30080), .B(n31195), .X(n12600) );
  nor_x1_sg U62569 ( .A(n31396), .B(n42712), .X(n12601) );
  nor_x1_sg U62570 ( .A(n35607), .B(n12605), .X(n12603) );
  nand_x1_sg U62571 ( .A(n30295), .B(n31197), .X(n12604) );
  nor_x1_sg U62572 ( .A(n34234), .B(n42713), .X(n12605) );
  nor_x1_sg U62573 ( .A(n35603), .B(n12609), .X(n12607) );
  nand_x1_sg U62574 ( .A(n34226), .B(n31199), .X(n12608) );
  nor_x1_sg U62575 ( .A(n29731), .B(n40919), .X(n12609) );
  nor_x1_sg U62576 ( .A(n35503), .B(n12622), .X(n12620) );
  nand_x1_sg U62577 ( .A(n34224), .B(n31126), .X(n12621) );
  nor_x1_sg U62578 ( .A(n31810), .B(n41072), .X(n12622) );
  nor_x1_sg U62579 ( .A(n35593), .B(n12626), .X(n12624) );
  nand_x1_sg U62580 ( .A(n31402), .B(n31128), .X(n12625) );
  nor_x1_sg U62581 ( .A(n34235), .B(n41070), .X(n12626) );
  nor_x1_sg U62582 ( .A(n35592), .B(n12635), .X(n12633) );
  nand_x1_sg U62583 ( .A(n34224), .B(n31130), .X(n12634) );
  nor_x1_sg U62584 ( .A(n34235), .B(n42596), .X(n12635) );
  nor_x1_sg U62585 ( .A(n35591), .B(n12644), .X(n12642) );
  nand_x1_sg U62586 ( .A(n31402), .B(n31133), .X(n12643) );
  nor_x1_sg U62587 ( .A(n31809), .B(n41064), .X(n12644) );
  nor_x1_sg U62588 ( .A(n35590), .B(n12648), .X(n12646) );
  nand_x1_sg U62589 ( .A(n34226), .B(n31135), .X(n12647) );
  nor_x1_sg U62590 ( .A(n31396), .B(n41062), .X(n12648) );
  nor_x1_sg U62591 ( .A(n35506), .B(n12652), .X(n12650) );
  nand_x1_sg U62592 ( .A(n30297), .B(n31137), .X(n12651) );
  nor_x1_sg U62593 ( .A(n34236), .B(n41060), .X(n12652) );
  nor_x1_sg U62594 ( .A(n35589), .B(n12656), .X(n12654) );
  nand_x1_sg U62595 ( .A(n30297), .B(n31139), .X(n12655) );
  nor_x1_sg U62596 ( .A(n31395), .B(n42598), .X(n12656) );
  nor_x1_sg U62597 ( .A(n35588), .B(n12660), .X(n12658) );
  nand_x1_sg U62598 ( .A(n31401), .B(n31141), .X(n12659) );
  nor_x1_sg U62599 ( .A(n30300), .B(n42599), .X(n12660) );
  nor_x1_sg U62600 ( .A(n35513), .B(n12664), .X(n12662) );
  nand_x1_sg U62601 ( .A(n30297), .B(n31143), .X(n12663) );
  nor_x1_sg U62602 ( .A(n30082), .B(n41056), .X(n12664) );
  nor_x1_sg U62603 ( .A(n35587), .B(n12668), .X(n12666) );
  nand_x1_sg U62604 ( .A(n34227), .B(n31145), .X(n12667) );
  nor_x1_sg U62605 ( .A(n34236), .B(n41054), .X(n12668) );
  nor_x1_sg U62606 ( .A(n35586), .B(n12672), .X(n12670) );
  nand_x1_sg U62607 ( .A(n31813), .B(n31147), .X(n12671) );
  nor_x1_sg U62608 ( .A(n31395), .B(n42600), .X(n12672) );
  nor_x1_sg U62609 ( .A(n35505), .B(n12676), .X(n12674) );
  nand_x1_sg U62610 ( .A(n31402), .B(n31149), .X(n12675) );
  nor_x1_sg U62611 ( .A(n31396), .B(n42601), .X(n12676) );
  nor_x1_sg U62612 ( .A(n35585), .B(n12680), .X(n12678) );
  nand_x1_sg U62613 ( .A(n31813), .B(n31151), .X(n12679) );
  nor_x1_sg U62614 ( .A(n34237), .B(n41050), .X(n12680) );
  nor_x1_sg U62615 ( .A(n35584), .B(n12684), .X(n12682) );
  nand_x1_sg U62616 ( .A(n34225), .B(n31153), .X(n12683) );
  nor_x1_sg U62617 ( .A(n34237), .B(n41048), .X(n12684) );
  nor_x1_sg U62618 ( .A(n35512), .B(n12688), .X(n12686) );
  nand_x1_sg U62619 ( .A(n30080), .B(n31155), .X(n12687) );
  nor_x1_sg U62620 ( .A(n34234), .B(n41046), .X(n12688) );
  nor_x1_sg U62621 ( .A(n35583), .B(n12702), .X(n12700) );
  nand_x1_sg U62622 ( .A(n31813), .B(n31157), .X(n12701) );
  nor_x1_sg U62623 ( .A(n31810), .B(n41042), .X(n12702) );
  nand_x1_sg U62624 ( .A(\shifter_0/reg_w_15[2] ), .B(n34438), .X(n11926) );
  nand_x1_sg U62625 ( .A(\shifter_0/reg_w_14[2] ), .B(n32192), .X(n11927) );
  nand_x1_sg U62626 ( .A(\shifter_0/reg_w_14[3] ), .B(n32194), .X(n11938) );
  nand_x1_sg U62627 ( .A(\shifter_0/reg_w_15[3] ), .B(n30840), .X(n11937) );
  nand_x1_sg U62628 ( .A(\shifter_0/reg_w_15[5] ), .B(n31979), .X(n11959) );
  nand_x1_sg U62629 ( .A(\shifter_0/reg_w_14[5] ), .B(n32197), .X(n11960) );
  nand_x1_sg U62630 ( .A(\shifter_0/reg_w_15[6] ), .B(n31979), .X(n11970) );
  nand_x1_sg U62631 ( .A(\shifter_0/reg_w_14[6] ), .B(n34444), .X(n11971) );
  nand_x1_sg U62632 ( .A(\shifter_0/reg_w_14[8] ), .B(n32195), .X(n11993) );
  nand_x1_sg U62633 ( .A(\shifter_0/reg_w_15[8] ), .B(n31978), .X(n11992) );
  nand_x1_sg U62634 ( .A(\shifter_0/reg_w_14[9] ), .B(n34445), .X(n12004) );
  nand_x1_sg U62635 ( .A(\shifter_0/reg_w_15[9] ), .B(n31980), .X(n12003) );
  nand_x1_sg U62636 ( .A(\shifter_0/reg_w_15[11] ), .B(n31976), .X(n12025) );
  nand_x1_sg U62637 ( .A(\shifter_0/reg_w_14[11] ), .B(n32197), .X(n12026) );
  nand_x1_sg U62638 ( .A(\shifter_0/reg_w_14[12] ), .B(n32197), .X(n12037) );
  nand_x1_sg U62639 ( .A(\shifter_0/reg_w_15[12] ), .B(n31976), .X(n12036) );
  nand_x1_sg U62640 ( .A(\shifter_0/reg_w_15[16] ), .B(n31975), .X(n12080) );
  nand_x1_sg U62641 ( .A(\shifter_0/reg_w_14[16] ), .B(n30837), .X(n12081) );
  nand_x1_sg U62642 ( .A(\shifter_0/reg_w_14[17] ), .B(n32194), .X(n12092) );
  nand_x1_sg U62643 ( .A(\shifter_0/reg_w_15[17] ), .B(n31979), .X(n12091) );
  nand_x1_sg U62644 ( .A(\shifter_0/reg_i_15[3] ), .B(n34437), .X(n12165) );
  nand_x1_sg U62645 ( .A(\shifter_0/reg_i_14[3] ), .B(n34445), .X(n12166) );
  nand_x1_sg U62646 ( .A(\shifter_0/reg_i_15[5] ), .B(n31979), .X(n12187) );
  nand_x1_sg U62647 ( .A(\shifter_0/reg_i_14[5] ), .B(n34442), .X(n12188) );
  nand_x1_sg U62648 ( .A(\shifter_0/reg_i_15[6] ), .B(n31978), .X(n12198) );
  nand_x1_sg U62649 ( .A(\shifter_0/reg_i_14[6] ), .B(n11561), .X(n12199) );
  nand_x1_sg U62650 ( .A(\shifter_0/reg_i_14[8] ), .B(n32196), .X(n12221) );
  nand_x1_sg U62651 ( .A(\shifter_0/reg_i_15[8] ), .B(n34439), .X(n12220) );
  nand_x1_sg U62652 ( .A(\shifter_0/reg_i_14[9] ), .B(n34445), .X(n12232) );
  nand_x1_sg U62653 ( .A(\shifter_0/reg_i_15[9] ), .B(n30839), .X(n12231) );
  nand_x1_sg U62654 ( .A(\shifter_0/reg_i_15[11] ), .B(n30840), .X(n12253) );
  nand_x1_sg U62655 ( .A(\shifter_0/reg_i_14[11] ), .B(n32195), .X(n12254) );
  nand_x1_sg U62656 ( .A(\shifter_0/reg_i_14[12] ), .B(n30838), .X(n12265) );
  nand_x1_sg U62657 ( .A(\shifter_0/reg_i_15[12] ), .B(n31980), .X(n12264) );
  nand_x1_sg U62658 ( .A(\shifter_0/reg_i_14[16] ), .B(n32195), .X(n12309) );
  nand_x1_sg U62659 ( .A(\shifter_0/reg_i_15[16] ), .B(n31975), .X(n12308) );
  nand_x1_sg U62660 ( .A(\shifter_0/reg_w_1[0] ), .B(n32105), .X(n13618) );
  nand_x1_sg U62661 ( .A(\shifter_0/reg_w_1[1] ), .B(n34428), .X(n13623) );
  nand_x1_sg U62662 ( .A(\shifter_0/reg_w_1[2] ), .B(n34428), .X(n13627) );
  nand_x1_sg U62663 ( .A(\shifter_0/reg_w_1[3] ), .B(n30117), .X(n13631) );
  nand_x1_sg U62664 ( .A(\shifter_0/reg_w_1[4] ), .B(n34429), .X(n13635) );
  nand_x1_sg U62665 ( .A(\shifter_0/reg_w_1[5] ), .B(n32101), .X(n13639) );
  nand_x1_sg U62666 ( .A(\shifter_0/reg_w_1[6] ), .B(n32102), .X(n13643) );
  nand_x1_sg U62667 ( .A(\shifter_0/reg_w_1[7] ), .B(n32104), .X(n13647) );
  nand_x1_sg U62668 ( .A(\shifter_0/reg_w_1[8] ), .B(n32106), .X(n13651) );
  nand_x1_sg U62669 ( .A(\shifter_0/reg_w_1[9] ), .B(n32104), .X(n13655) );
  nand_x1_sg U62670 ( .A(\shifter_0/reg_w_1[10] ), .B(n34430), .X(n13659) );
  nand_x1_sg U62671 ( .A(\shifter_0/reg_w_1[11] ), .B(n34427), .X(n13663) );
  nand_x1_sg U62672 ( .A(\shifter_0/reg_w_1[12] ), .B(n34427), .X(n13667) );
  nand_x1_sg U62673 ( .A(\shifter_0/reg_w_1[13] ), .B(n30845), .X(n13671) );
  nand_x1_sg U62674 ( .A(\shifter_0/reg_w_1[14] ), .B(n32104), .X(n13675) );
  nand_x1_sg U62675 ( .A(\shifter_0/reg_w_1[15] ), .B(n32106), .X(n13679) );
  nand_x1_sg U62676 ( .A(\shifter_0/reg_w_1[16] ), .B(n34429), .X(n13683) );
  nand_x1_sg U62677 ( .A(\shifter_0/reg_w_1[17] ), .B(n32101), .X(n13687) );
  nand_x1_sg U62678 ( .A(\shifter_0/reg_w_1[18] ), .B(n32101), .X(n13691) );
  nand_x1_sg U62679 ( .A(\shifter_0/reg_w_1[19] ), .B(n34429), .X(n13695) );
  nand_x1_sg U62680 ( .A(\shifter_0/reg_i_1[0] ), .B(n34427), .X(n13705) );
  nand_x1_sg U62681 ( .A(\shifter_0/reg_i_1[1] ), .B(n32106), .X(n13709) );
  nand_x1_sg U62682 ( .A(\shifter_0/reg_i_1[3] ), .B(n30845), .X(n13716) );
  nand_x1_sg U62683 ( .A(\shifter_0/reg_i_1[5] ), .B(n30845), .X(n13723) );
  nand_x1_sg U62684 ( .A(\shifter_0/reg_i_1[6] ), .B(n30117), .X(n13727) );
  nand_x1_sg U62685 ( .A(\shifter_0/reg_i_1[7] ), .B(n34430), .X(n13731) );
  nand_x1_sg U62686 ( .A(\shifter_0/reg_i_1[8] ), .B(n34428), .X(n13735) );
  nand_x1_sg U62687 ( .A(\shifter_0/reg_i_1[9] ), .B(n30845), .X(n13739) );
  nand_x1_sg U62688 ( .A(\shifter_0/reg_i_1[10] ), .B(n32102), .X(n13743) );
  nand_x1_sg U62689 ( .A(\shifter_0/reg_i_1[11] ), .B(n32102), .X(n13747) );
  nand_x1_sg U62690 ( .A(\shifter_0/reg_i_1[12] ), .B(n34428), .X(n13751) );
  nand_x1_sg U62691 ( .A(\shifter_0/reg_i_1[13] ), .B(n32105), .X(n13755) );
  nand_x1_sg U62692 ( .A(\shifter_0/reg_i_1[14] ), .B(n32104), .X(n13759) );
  nand_x1_sg U62693 ( .A(\shifter_0/reg_i_1[15] ), .B(n32101), .X(n13763) );
  nand_x1_sg U62694 ( .A(\shifter_0/reg_i_1[16] ), .B(n32106), .X(n13767) );
  nand_x1_sg U62695 ( .A(\shifter_0/reg_i_1[19] ), .B(n34427), .X(n13777) );
  nand_x1_sg U62696 ( .A(\shifter_0/reg_w_13[0] ), .B(n34425), .X(n11902) );
  nand_x1_sg U62697 ( .A(\shifter_0/reg_w_13[1] ), .B(n32110), .X(n11914) );
  nand_x1_sg U62698 ( .A(\shifter_0/reg_w_13[2] ), .B(n30116), .X(n11925) );
  nand_x1_sg U62699 ( .A(\shifter_0/reg_w_13[5] ), .B(n32108), .X(n11958) );
  nand_x1_sg U62700 ( .A(\shifter_0/reg_w_13[6] ), .B(n30847), .X(n11969) );
  nand_x1_sg U62701 ( .A(\shifter_0/reg_w_13[7] ), .B(n32112), .X(n11980) );
  nand_x1_sg U62702 ( .A(\shifter_0/reg_w_13[10] ), .B(n32111), .X(n12013) );
  nand_x1_sg U62703 ( .A(\shifter_0/reg_w_13[11] ), .B(n30847), .X(n12024) );
  nand_x1_sg U62704 ( .A(\shifter_0/reg_w_13[14] ), .B(n34425), .X(n12057) );
  nand_x1_sg U62705 ( .A(\shifter_0/reg_w_13[15] ), .B(n32110), .X(n12068) );
  nand_x1_sg U62706 ( .A(\shifter_0/reg_w_13[16] ), .B(n30116), .X(n12079) );
  nand_x1_sg U62707 ( .A(\shifter_0/reg_w_13[19] ), .B(n32107), .X(n12112) );
  nand_x1_sg U62708 ( .A(\shifter_0/reg_i_13[0] ), .B(n32108), .X(n12130) );
  nand_x1_sg U62709 ( .A(\shifter_0/reg_i_13[1] ), .B(n32110), .X(n12142) );
  nand_x1_sg U62710 ( .A(\shifter_0/reg_i_13[3] ), .B(n34422), .X(n12164) );
  nand_x1_sg U62711 ( .A(\shifter_0/reg_i_13[5] ), .B(n30847), .X(n12186) );
  nand_x1_sg U62712 ( .A(\shifter_0/reg_i_13[6] ), .B(n34422), .X(n12197) );
  nand_x1_sg U62713 ( .A(\shifter_0/reg_i_13[7] ), .B(n34424), .X(n12208) );
  nand_x1_sg U62714 ( .A(\shifter_0/reg_i_13[10] ), .B(n32111), .X(n12241) );
  nand_x1_sg U62715 ( .A(\shifter_0/reg_i_13[11] ), .B(n34423), .X(n12252) );
  nand_x1_sg U62716 ( .A(\shifter_0/reg_i_13[14] ), .B(n34422), .X(n12285) );
  nand_x1_sg U62717 ( .A(\shifter_0/reg_i_13[15] ), .B(n30847), .X(n12296) );
  nand_x1_sg U62718 ( .A(\shifter_0/reg_i_13[19] ), .B(n34423), .X(n12340) );
  nand_x1_sg U62719 ( .A(\shifter_0/reg_w_12[0] ), .B(n32203), .X(n11901) );
  nand_x1_sg U62720 ( .A(\shifter_0/reg_w_12[1] ), .B(n32202), .X(n11913) );
  nand_x1_sg U62721 ( .A(\shifter_0/reg_w_12[2] ), .B(n34432), .X(n11924) );
  nand_x1_sg U62722 ( .A(\shifter_0/reg_w_12[5] ), .B(n30843), .X(n11957) );
  nand_x1_sg U62723 ( .A(\shifter_0/reg_w_12[6] ), .B(n34434), .X(n11968) );
  nand_x1_sg U62724 ( .A(\shifter_0/reg_w_12[7] ), .B(n32203), .X(n11979) );
  nand_x1_sg U62725 ( .A(\shifter_0/reg_w_12[10] ), .B(n32200), .X(n12012) );
  nand_x1_sg U62726 ( .A(\shifter_0/reg_w_12[11] ), .B(n32201), .X(n12023) );
  nand_x1_sg U62727 ( .A(\shifter_0/reg_w_12[14] ), .B(n34433), .X(n12056) );
  nand_x1_sg U62728 ( .A(\shifter_0/reg_w_12[15] ), .B(n32202), .X(n12067) );
  nand_x1_sg U62729 ( .A(\shifter_0/reg_w_12[16] ), .B(n32198), .X(n12078) );
  nand_x1_sg U62730 ( .A(\shifter_0/reg_w_12[19] ), .B(n32203), .X(n12111) );
  nand_x1_sg U62731 ( .A(\shifter_0/reg_i_12[0] ), .B(n30844), .X(n12129) );
  nand_x1_sg U62732 ( .A(\shifter_0/reg_i_12[1] ), .B(n30844), .X(n12141) );
  nand_x1_sg U62733 ( .A(\shifter_0/reg_i_12[3] ), .B(n34434), .X(n12163) );
  nand_x1_sg U62734 ( .A(\shifter_0/reg_i_12[5] ), .B(n34433), .X(n12185) );
  nand_x1_sg U62735 ( .A(\shifter_0/reg_i_12[6] ), .B(n32202), .X(n12196) );
  nand_x1_sg U62736 ( .A(\shifter_0/reg_i_12[7] ), .B(n30844), .X(n12207) );
  nand_x1_sg U62737 ( .A(\shifter_0/reg_i_12[10] ), .B(n34435), .X(n12240) );
  nand_x1_sg U62738 ( .A(\shifter_0/reg_i_12[11] ), .B(n34435), .X(n12251) );
  nand_x1_sg U62739 ( .A(\shifter_0/reg_i_12[14] ), .B(n32201), .X(n12284) );
  nand_x1_sg U62740 ( .A(\shifter_0/reg_i_12[15] ), .B(n34434), .X(n12295) );
  nand_x1_sg U62741 ( .A(\shifter_0/reg_i_12[19] ), .B(n32200), .X(n12339) );
  nand_x1_sg U62742 ( .A(\shifter_0/reg_w_11[0] ), .B(n34513), .X(n11900) );
  nand_x1_sg U62743 ( .A(\shifter_0/reg_w_11[1] ), .B(n32177), .X(n11912) );
  nand_x1_sg U62744 ( .A(\shifter_0/reg_w_11[2] ), .B(n32178), .X(n11923) );
  nand_x1_sg U62745 ( .A(\shifter_0/reg_w_11[5] ), .B(n32421), .X(n11956) );
  nand_x1_sg U62746 ( .A(\shifter_0/reg_w_11[6] ), .B(n34515), .X(n11967) );
  nand_x1_sg U62747 ( .A(\shifter_0/reg_w_11[7] ), .B(n34514), .X(n11978) );
  nand_x1_sg U62748 ( .A(\shifter_0/reg_w_11[10] ), .B(n32419), .X(n12011) );
  nand_x1_sg U62749 ( .A(\shifter_0/reg_w_11[11] ), .B(n32177), .X(n12022) );
  nand_x1_sg U62750 ( .A(\shifter_0/reg_w_11[14] ), .B(n32419), .X(n12055) );
  nand_x1_sg U62751 ( .A(\shifter_0/reg_w_11[15] ), .B(n32422), .X(n12066) );
  nand_x1_sg U62752 ( .A(\shifter_0/reg_w_11[16] ), .B(n30785), .X(n12077) );
  nand_x1_sg U62753 ( .A(\shifter_0/reg_w_11[19] ), .B(n32419), .X(n12110) );
  nand_x1_sg U62754 ( .A(\shifter_0/reg_i_11[0] ), .B(n34516), .X(n12128) );
  nand_x1_sg U62755 ( .A(\shifter_0/reg_i_11[1] ), .B(n30786), .X(n12140) );
  nand_x1_sg U62756 ( .A(\shifter_0/reg_i_11[3] ), .B(n34516), .X(n12162) );
  nand_x1_sg U62757 ( .A(\shifter_0/reg_i_11[5] ), .B(n34514), .X(n12184) );
  nand_x1_sg U62758 ( .A(\shifter_0/reg_i_11[6] ), .B(n32422), .X(n12195) );
  nand_x1_sg U62759 ( .A(\shifter_0/reg_i_11[7] ), .B(n32177), .X(n12206) );
  nand_x1_sg U62760 ( .A(\shifter_0/reg_i_11[10] ), .B(n30785), .X(n12239) );
  nand_x1_sg U62761 ( .A(\shifter_0/reg_i_11[11] ), .B(n34515), .X(n12250) );
  nand_x1_sg U62762 ( .A(\shifter_0/reg_i_11[14] ), .B(n32422), .X(n12283) );
  nand_x1_sg U62763 ( .A(\shifter_0/reg_i_11[15] ), .B(n32178), .X(n12294) );
  nand_x1_sg U62764 ( .A(\shifter_0/reg_i_11[19] ), .B(n34513), .X(n12338) );
  nand_x1_sg U62765 ( .A(n31377), .B(\shifter_0/reg_i_12[2] ), .X(n14503) );
  nand_x1_sg U62766 ( .A(n34262), .B(\shifter_0/reg_i_13[2] ), .X(n14502) );
  nand_x1_sg U62767 ( .A(n31377), .B(\shifter_0/reg_i_12[4] ), .X(n14565) );
  nand_x1_sg U62768 ( .A(n31380), .B(\shifter_0/reg_i_13[4] ), .X(n14564) );
  nand_x1_sg U62769 ( .A(n34265), .B(\shifter_0/reg_i_12[17] ), .X(n14968) );
  nand_x1_sg U62770 ( .A(n31380), .B(\shifter_0/reg_i_13[17] ), .X(n14967) );
  nand_x1_sg U62771 ( .A(n34264), .B(\shifter_0/reg_i_12[18] ), .X(n14999) );
  nand_x1_sg U62772 ( .A(n31801), .B(\shifter_0/reg_i_13[18] ), .X(n14998) );
  nand_x1_sg U62773 ( .A(n33987), .B(\shifter_0/reg_i_4[2] ), .X(n14484) );
  nand_x1_sg U62774 ( .A(n30909), .B(\shifter_0/reg_w_4[0] ), .X(n13794) );
  nand_x1_sg U62775 ( .A(n31696), .B(\shifter_0/reg_w_4[1] ), .X(n13831) );
  nand_x1_sg U62776 ( .A(n30908), .B(\shifter_0/reg_w_4[2] ), .X(n13862) );
  nand_x1_sg U62777 ( .A(n33985), .B(\shifter_0/reg_w_4[5] ), .X(n13955) );
  nand_x1_sg U62778 ( .A(n30909), .B(\shifter_0/reg_w_4[6] ), .X(n13986) );
  nand_x1_sg U62779 ( .A(n30909), .B(\shifter_0/reg_w_4[7] ), .X(n14017) );
  nand_x1_sg U62780 ( .A(n33985), .B(\shifter_0/reg_w_4[10] ), .X(n14110) );
  nand_x1_sg U62781 ( .A(n33986), .B(\shifter_0/reg_w_4[11] ), .X(n14141) );
  nand_x1_sg U62782 ( .A(n33984), .B(\shifter_0/reg_w_4[14] ), .X(n14234) );
  nand_x1_sg U62783 ( .A(n31695), .B(\shifter_0/reg_w_4[15] ), .X(n14265) );
  nand_x1_sg U62784 ( .A(n33984), .B(\shifter_0/reg_w_4[16] ), .X(n14296) );
  nand_x1_sg U62785 ( .A(n31695), .B(\shifter_0/reg_w_4[19] ), .X(n14389) );
  nand_x1_sg U62786 ( .A(n33985), .B(\shifter_0/reg_i_4[0] ), .X(n14421) );
  nand_x1_sg U62787 ( .A(n31696), .B(\shifter_0/reg_i_4[1] ), .X(n14452) );
  nand_x1_sg U62788 ( .A(n30020), .B(\shifter_0/reg_i_4[5] ), .X(n14578) );
  nand_x1_sg U62789 ( .A(n30908), .B(\shifter_0/reg_i_4[6] ), .X(n14609) );
  nand_x1_sg U62790 ( .A(n33984), .B(\shifter_0/reg_i_4[7] ), .X(n14640) );
  nand_x1_sg U62791 ( .A(n33987), .B(\shifter_0/reg_i_4[10] ), .X(n14733) );
  nand_x1_sg U62792 ( .A(n31695), .B(\shifter_0/reg_i_4[11] ), .X(n14764) );
  nand_x1_sg U62793 ( .A(n33987), .B(\shifter_0/reg_i_4[14] ), .X(n14857) );
  nand_x1_sg U62794 ( .A(n30908), .B(\shifter_0/reg_i_4[15] ), .X(n14888) );
  nand_x1_sg U62795 ( .A(n33986), .B(\shifter_0/reg_i_4[16] ), .X(n14919) );
  nand_x1_sg U62796 ( .A(n30020), .B(\shifter_0/reg_i_4[19] ), .X(n15012) );
  nand_x1_sg U62797 ( .A(n31121), .B(n35269), .X(n15074) );
  nand_x1_sg U62798 ( .A(n31593), .B(n35257), .X(n15075) );
  nand_x1_sg U62799 ( .A(\shifter_0/reg_w_10[0] ), .B(n34518), .X(n11899) );
  nand_x1_sg U62800 ( .A(\shifter_0/reg_w_10[1] ), .B(n32415), .X(n11911) );
  nand_x1_sg U62801 ( .A(\shifter_0/reg_w_10[2] ), .B(n32412), .X(n11922) );
  nand_x1_sg U62802 ( .A(\shifter_0/reg_w_10[3] ), .B(n32176), .X(n11933) );
  nand_x1_sg U62803 ( .A(\shifter_0/reg_w_10[4] ), .B(n32414), .X(n11944) );
  nand_x1_sg U62804 ( .A(\shifter_0/reg_w_10[5] ), .B(n32174), .X(n11955) );
  nand_x1_sg U62805 ( .A(\shifter_0/reg_w_10[6] ), .B(n32175), .X(n11966) );
  nand_x1_sg U62806 ( .A(\shifter_0/reg_w_10[7] ), .B(n32176), .X(n11977) );
  nand_x1_sg U62807 ( .A(\shifter_0/reg_w_10[8] ), .B(n32417), .X(n11988) );
  nand_x1_sg U62808 ( .A(\shifter_0/reg_w_10[9] ), .B(n32176), .X(n11999) );
  nand_x1_sg U62809 ( .A(\shifter_0/reg_w_10[10] ), .B(n32411), .X(n12010) );
  nand_x1_sg U62810 ( .A(\shifter_0/reg_w_10[11] ), .B(n32415), .X(n12021) );
  nand_x1_sg U62811 ( .A(\shifter_0/reg_w_10[12] ), .B(n32174), .X(n12032) );
  nand_x1_sg U62812 ( .A(\shifter_0/reg_w_10[13] ), .B(n32412), .X(n12043) );
  nand_x1_sg U62813 ( .A(\shifter_0/reg_w_10[14] ), .B(n32412), .X(n12054) );
  nand_x1_sg U62814 ( .A(\shifter_0/reg_w_10[15] ), .B(n32410), .X(n12065) );
  nand_x1_sg U62815 ( .A(\shifter_0/reg_w_10[16] ), .B(n32175), .X(n12076) );
  nand_x1_sg U62816 ( .A(\shifter_0/reg_w_10[17] ), .B(n32417), .X(n12087) );
  nand_x1_sg U62817 ( .A(\shifter_0/reg_w_10[18] ), .B(n32414), .X(n12098) );
  nand_x1_sg U62818 ( .A(\shifter_0/reg_w_10[19] ), .B(n32411), .X(n12109) );
  nand_x1_sg U62819 ( .A(\shifter_0/reg_i_10[0] ), .B(n32175), .X(n12127) );
  nand_x1_sg U62820 ( .A(\shifter_0/reg_i_10[1] ), .B(n32411), .X(n12139) );
  nand_x1_sg U62821 ( .A(\shifter_0/reg_i_10[3] ), .B(n32410), .X(n12161) );
  nand_x1_sg U62822 ( .A(\shifter_0/reg_i_10[5] ), .B(n32416), .X(n12183) );
  nand_x1_sg U62823 ( .A(\shifter_0/reg_i_10[6] ), .B(n34518), .X(n12194) );
  nand_x1_sg U62824 ( .A(\shifter_0/reg_i_10[7] ), .B(n32417), .X(n12205) );
  nand_x1_sg U62825 ( .A(\shifter_0/reg_i_10[8] ), .B(n32412), .X(n12216) );
  nand_x1_sg U62826 ( .A(\shifter_0/reg_i_10[9] ), .B(n32415), .X(n12227) );
  nand_x1_sg U62827 ( .A(\shifter_0/reg_i_10[10] ), .B(n32410), .X(n12238) );
  nand_x1_sg U62828 ( .A(\shifter_0/reg_i_10[11] ), .B(n32415), .X(n12249) );
  nand_x1_sg U62829 ( .A(\shifter_0/reg_i_10[12] ), .B(n32416), .X(n12260) );
  nand_x1_sg U62830 ( .A(\shifter_0/reg_i_10[13] ), .B(n32416), .X(n12271) );
  nand_x1_sg U62831 ( .A(\shifter_0/reg_i_10[14] ), .B(n32416), .X(n12282) );
  nand_x1_sg U62832 ( .A(\shifter_0/reg_i_10[15] ), .B(n32174), .X(n12293) );
  nand_x1_sg U62833 ( .A(\shifter_0/reg_i_10[16] ), .B(n32414), .X(n12304) );
  nand_x1_sg U62834 ( .A(\shifter_0/reg_i_10[19] ), .B(n32414), .X(n12337) );
  nand_x1_sg U62835 ( .A(\shifter_0/reg_i_13[4] ), .B(n32111), .X(n12175) );
  nand_x1_sg U62836 ( .A(\shifter_0/reg_i_13[18] ), .B(n32112), .X(n12329) );
  nand_x1_sg U62837 ( .A(\shifter_0/reg_w_13[4] ), .B(n32111), .X(n11947) );
  nand_x1_sg U62838 ( .A(\shifter_0/reg_w_13[13] ), .B(n32112), .X(n12046) );
  nand_x1_sg U62839 ( .A(\shifter_0/reg_w_13[18] ), .B(n34425), .X(n12101) );
  nand_x1_sg U62840 ( .A(\shifter_0/reg_i_13[13] ), .B(n32112), .X(n12274) );
  nand_x1_sg U62841 ( .A(\shifter_0/reg_i_13[2] ), .B(n32110), .X(n12153) );
  nand_x1_sg U62842 ( .A(\shifter_0/reg_i_13[17] ), .B(n30116), .X(n12318) );
  nand_x1_sg U62843 ( .A(\shifter_0/reg_w_13[3] ), .B(n34424), .X(n11936) );
  nand_x1_sg U62844 ( .A(\shifter_0/reg_w_13[8] ), .B(n32108), .X(n11991) );
  nand_x1_sg U62845 ( .A(\shifter_0/reg_w_13[9] ), .B(n34422), .X(n12002) );
  nand_x1_sg U62846 ( .A(\shifter_0/reg_w_13[12] ), .B(n34423), .X(n12035) );
  nand_x1_sg U62847 ( .A(\shifter_0/reg_w_13[17] ), .B(n34423), .X(n12090) );
  nand_x1_sg U62848 ( .A(\shifter_0/reg_i_13[8] ), .B(n32107), .X(n12219) );
  nand_x1_sg U62849 ( .A(\shifter_0/reg_i_13[9] ), .B(n32107), .X(n12230) );
  nand_x1_sg U62850 ( .A(\shifter_0/reg_i_13[12] ), .B(n34424), .X(n12263) );
  nand_x1_sg U62851 ( .A(\shifter_0/reg_i_13[16] ), .B(n32107), .X(n12307) );
  nand_x1_sg U62852 ( .A(\shifter_0/reg_w_12[3] ), .B(n30843), .X(n11935) );
  nand_x1_sg U62853 ( .A(\shifter_0/reg_w_12[4] ), .B(n34432), .X(n11946) );
  nand_x1_sg U62854 ( .A(\shifter_0/reg_w_12[8] ), .B(n30843), .X(n11990) );
  nand_x1_sg U62855 ( .A(\shifter_0/reg_w_12[9] ), .B(n32201), .X(n12001) );
  nand_x1_sg U62856 ( .A(\shifter_0/reg_w_12[12] ), .B(n32202), .X(n12034) );
  nand_x1_sg U62857 ( .A(\shifter_0/reg_w_12[13] ), .B(n32201), .X(n12045) );
  nand_x1_sg U62858 ( .A(\shifter_0/reg_w_12[17] ), .B(n32203), .X(n12089) );
  nand_x1_sg U62859 ( .A(\shifter_0/reg_w_12[18] ), .B(n34432), .X(n12100) );
  nand_x1_sg U62860 ( .A(\shifter_0/reg_i_12[2] ), .B(n32198), .X(n12152) );
  nand_x1_sg U62861 ( .A(\shifter_0/reg_i_12[4] ), .B(n32200), .X(n12174) );
  nand_x1_sg U62862 ( .A(\shifter_0/reg_i_12[8] ), .B(n32200), .X(n12218) );
  nand_x1_sg U62863 ( .A(\shifter_0/reg_i_12[9] ), .B(n34435), .X(n12229) );
  nand_x1_sg U62864 ( .A(\shifter_0/reg_i_12[12] ), .B(n35657), .X(n12262) );
  nand_x1_sg U62865 ( .A(\shifter_0/reg_i_12[13] ), .B(n34432), .X(n12273) );
  nand_x1_sg U62866 ( .A(\shifter_0/reg_i_12[16] ), .B(n34433), .X(n12306) );
  nand_x1_sg U62867 ( .A(\shifter_0/reg_i_12[17] ), .B(n32198), .X(n12317) );
  nand_x1_sg U62868 ( .A(\shifter_0/reg_i_12[18] ), .B(n35657), .X(n12328) );
  nand_x1_sg U62869 ( .A(\shifter_0/reg_w_11[3] ), .B(n30785), .X(n11934) );
  nand_x1_sg U62870 ( .A(\shifter_0/reg_w_11[4] ), .B(n30786), .X(n11945) );
  nand_x1_sg U62871 ( .A(\shifter_0/reg_w_11[8] ), .B(n32420), .X(n11989) );
  nand_x1_sg U62872 ( .A(\shifter_0/reg_w_11[9] ), .B(n34514), .X(n12000) );
  nand_x1_sg U62873 ( .A(\shifter_0/reg_w_11[12] ), .B(n32421), .X(n12033) );
  nand_x1_sg U62874 ( .A(\shifter_0/reg_w_11[13] ), .B(n30786), .X(n12044) );
  nand_x1_sg U62875 ( .A(\shifter_0/reg_w_11[17] ), .B(n32178), .X(n12088) );
  nand_x1_sg U62876 ( .A(\shifter_0/reg_w_11[18] ), .B(n32421), .X(n12099) );
  nand_x1_sg U62877 ( .A(\shifter_0/reg_i_11[2] ), .B(n34514), .X(n12151) );
  nand_x1_sg U62878 ( .A(\shifter_0/reg_i_11[4] ), .B(n32419), .X(n12173) );
  nand_x1_sg U62879 ( .A(\shifter_0/reg_i_11[8] ), .B(n32177), .X(n12217) );
  nand_x1_sg U62880 ( .A(\shifter_0/reg_i_11[9] ), .B(n34513), .X(n12228) );
  nand_x1_sg U62881 ( .A(\shifter_0/reg_i_11[12] ), .B(n30786), .X(n12261) );
  nand_x1_sg U62882 ( .A(\shifter_0/reg_i_11[13] ), .B(n32420), .X(n12272) );
  nand_x1_sg U62883 ( .A(\shifter_0/reg_i_11[16] ), .B(n32420), .X(n12305) );
  nand_x1_sg U62884 ( .A(\shifter_0/reg_i_11[17] ), .B(n34515), .X(n12316) );
  nand_x1_sg U62885 ( .A(\shifter_0/reg_i_11[18] ), .B(n30785), .X(n12327) );
  nand_x1_sg U62886 ( .A(\shifter_0/reg_i_10[2] ), .B(n32417), .X(n12150) );
  nand_x1_sg U62887 ( .A(\shifter_0/reg_i_10[4] ), .B(n32174), .X(n12172) );
  nand_x1_sg U62888 ( .A(\shifter_0/reg_i_10[17] ), .B(n32176), .X(n12315) );
  nand_x1_sg U62889 ( .A(\shifter_0/reg_i_10[18] ), .B(n32411), .X(n12326) );
  nand_x1_sg U62890 ( .A(\shifter_0/reg_i_5[17] ), .B(n31022), .X(n14950) );
  nor_x1_sg U62891 ( .A(n12948), .B(n14951), .X(n14949) );
  nor_x1_sg U62892 ( .A(n29688), .B(n42586), .X(n14951) );
  nor_x1_sg U62893 ( .A(n12858), .B(n41120), .X(n14482) );
  nand_x1_sg U62894 ( .A(\shifter_0/reg_i_5[2] ), .B(n34539), .X(n14483) );
  nor_x1_sg U62895 ( .A(n12870), .B(n14548), .X(n14546) );
  nand_x1_sg U62896 ( .A(\shifter_0/reg_i_5[4] ), .B(n32062), .X(n14547) );
  nor_x1_sg U62897 ( .A(n33960), .B(n42581), .X(n14548) );
  nor_x1_sg U62898 ( .A(n12954), .B(n14982), .X(n14980) );
  nand_x1_sg U62899 ( .A(\shifter_0/reg_i_5[18] ), .B(n32064), .X(n14981) );
  nor_x1_sg U62900 ( .A(n31653), .B(n42587), .X(n14982) );
  inv_x1_sg U62901 ( .A(\shifter_0/reg_w_0[0] ), .X(n40985) );
  inv_x1_sg U62902 ( .A(\shifter_0/reg_w_0[1] ), .X(n40984) );
  inv_x1_sg U62903 ( .A(\shifter_0/reg_w_0[2] ), .X(n40983) );
  inv_x1_sg U62904 ( .A(\shifter_0/reg_w_0[5] ), .X(n40982) );
  inv_x1_sg U62905 ( .A(\shifter_0/reg_w_0[6] ), .X(n40981) );
  inv_x1_sg U62906 ( .A(\shifter_0/reg_w_0[7] ), .X(n40980) );
  inv_x1_sg U62907 ( .A(\shifter_0/reg_w_0[10] ), .X(n40979) );
  inv_x1_sg U62908 ( .A(\shifter_0/reg_w_0[11] ), .X(n40978) );
  inv_x1_sg U62909 ( .A(\shifter_0/reg_w_0[14] ), .X(n40977) );
  inv_x1_sg U62910 ( .A(\shifter_0/reg_w_0[15] ), .X(n40976) );
  inv_x1_sg U62911 ( .A(\shifter_0/reg_w_0[16] ), .X(n40975) );
  inv_x1_sg U62912 ( .A(\shifter_0/reg_w_0[19] ), .X(n40974) );
  inv_x1_sg U62913 ( .A(\shifter_0/reg_i_0[0] ), .X(n41108) );
  inv_x1_sg U62914 ( .A(\shifter_0/reg_i_0[1] ), .X(n41107) );
  inv_x1_sg U62915 ( .A(\shifter_0/reg_i_0[2] ), .X(n41106) );
  inv_x1_sg U62916 ( .A(\shifter_0/reg_i_0[5] ), .X(n41105) );
  inv_x1_sg U62917 ( .A(\shifter_0/reg_i_0[6] ), .X(n41104) );
  inv_x1_sg U62918 ( .A(\shifter_0/reg_i_0[7] ), .X(n41103) );
  inv_x1_sg U62919 ( .A(\shifter_0/reg_i_0[10] ), .X(n41102) );
  inv_x1_sg U62920 ( .A(\shifter_0/reg_i_0[11] ), .X(n41101) );
  inv_x1_sg U62921 ( .A(\shifter_0/reg_i_0[14] ), .X(n41100) );
  inv_x1_sg U62922 ( .A(\shifter_0/reg_i_0[15] ), .X(n41099) );
  inv_x1_sg U62923 ( .A(\shifter_0/reg_i_0[16] ), .X(n41098) );
  inv_x1_sg U62924 ( .A(\shifter_0/reg_i_0[19] ), .X(n41097) );
  nand_x1_sg U62925 ( .A(\shifter_0/reg_w_3[0] ), .B(n31020), .X(n13229) );
  nand_x1_sg U62926 ( .A(\shifter_0/reg_w_3[1] ), .B(n32068), .X(n13232) );
  nand_x1_sg U62927 ( .A(\shifter_0/reg_w_3[2] ), .B(n32069), .X(n13235) );
  nand_x1_sg U62928 ( .A(\shifter_0/reg_w_3[5] ), .B(n30134), .X(n13244) );
  nand_x1_sg U62929 ( .A(\shifter_0/reg_w_3[6] ), .B(n32070), .X(n13247) );
  nand_x1_sg U62930 ( .A(\shifter_0/reg_w_3[7] ), .B(n32068), .X(n13250) );
  nand_x1_sg U62931 ( .A(\shifter_0/reg_w_3[10] ), .B(n32066), .X(n13259) );
  nand_x1_sg U62932 ( .A(\shifter_0/reg_w_3[11] ), .B(n34535), .X(n13262) );
  nand_x1_sg U62933 ( .A(\shifter_0/reg_w_3[14] ), .B(n34535), .X(n13271) );
  nand_x1_sg U62934 ( .A(\shifter_0/reg_w_3[15] ), .B(n34536), .X(n13274) );
  nand_x1_sg U62935 ( .A(\shifter_0/reg_w_3[16] ), .B(n34537), .X(n13277) );
  nand_x1_sg U62936 ( .A(\shifter_0/reg_w_3[19] ), .B(n32066), .X(n13286) );
  nand_x1_sg U62937 ( .A(\shifter_0/reg_i_3[0] ), .B(n34535), .X(n13295) );
  nand_x1_sg U62938 ( .A(\shifter_0/reg_i_3[1] ), .B(n34535), .X(n13298) );
  nand_x1_sg U62939 ( .A(\shifter_0/reg_i_3[5] ), .B(n31019), .X(n13312) );
  nand_x1_sg U62940 ( .A(\shifter_0/reg_i_3[6] ), .B(n32068), .X(n13315) );
  nand_x1_sg U62941 ( .A(\shifter_0/reg_i_3[7] ), .B(n32069), .X(n13318) );
  nand_x1_sg U62942 ( .A(\shifter_0/reg_i_3[10] ), .B(n32065), .X(n13327) );
  nand_x1_sg U62943 ( .A(\shifter_0/reg_i_3[11] ), .B(n34536), .X(n13330) );
  nand_x1_sg U62944 ( .A(\shifter_0/reg_i_3[14] ), .B(n34534), .X(n13339) );
  nand_x1_sg U62945 ( .A(\shifter_0/reg_i_3[15] ), .B(n34537), .X(n13342) );
  nand_x1_sg U62946 ( .A(\shifter_0/reg_i_3[16] ), .B(n32069), .X(n13345) );
  nand_x1_sg U62947 ( .A(\shifter_0/reg_i_3[19] ), .B(n34534), .X(n13356) );
  nand_x1_sg U62948 ( .A(\shifter_0/reg_w_3[3] ), .B(n32065), .X(n13238) );
  nand_x1_sg U62949 ( .A(\shifter_0/reg_w_3[4] ), .B(n32066), .X(n13241) );
  nand_x1_sg U62950 ( .A(\shifter_0/reg_w_3[8] ), .B(n32065), .X(n13253) );
  nand_x1_sg U62951 ( .A(\shifter_0/reg_w_3[9] ), .B(n32066), .X(n13256) );
  nand_x1_sg U62952 ( .A(\shifter_0/reg_w_3[12] ), .B(n31020), .X(n13265) );
  nand_x1_sg U62953 ( .A(\shifter_0/reg_w_3[13] ), .B(n32070), .X(n13268) );
  nand_x1_sg U62954 ( .A(\shifter_0/reg_w_3[17] ), .B(n34536), .X(n13280) );
  nand_x1_sg U62955 ( .A(\shifter_0/reg_w_3[18] ), .B(n31020), .X(n13283) );
  nand_x1_sg U62956 ( .A(\shifter_0/reg_i_3[3] ), .B(n34536), .X(n13305) );
  nand_x1_sg U62957 ( .A(\shifter_0/reg_i_3[8] ), .B(n32070), .X(n13321) );
  nand_x1_sg U62958 ( .A(\shifter_0/reg_i_3[9] ), .B(n31019), .X(n13324) );
  nand_x1_sg U62959 ( .A(\shifter_0/reg_i_3[12] ), .B(n31020), .X(n13333) );
  nand_x1_sg U62960 ( .A(\shifter_0/reg_i_3[13] ), .B(n32070), .X(n13336) );
  nand_x1_sg U62961 ( .A(\shifter_0/reg_i_1[2] ), .B(n34430), .X(n13712) );
  nand_x1_sg U62962 ( .A(\shifter_0/reg_i_1[4] ), .B(n32105), .X(n13719) );
  nand_x1_sg U62963 ( .A(\shifter_0/reg_i_1[17] ), .B(n30117), .X(n13770) );
  nand_x1_sg U62964 ( .A(\shifter_0/reg_i_1[18] ), .B(n32105), .X(n13773) );
  nand_x1_sg U62965 ( .A(n34259), .B(n40881), .X(n13815) );
  inv_x1_sg U62966 ( .A(\shifter_0/reg_w_13[0] ), .X(n40881) );
  nand_x1_sg U62967 ( .A(n31801), .B(n40880), .X(n13849) );
  inv_x1_sg U62968 ( .A(\shifter_0/reg_w_13[1] ), .X(n40880) );
  nand_x1_sg U62969 ( .A(n34259), .B(n40879), .X(n13880) );
  inv_x1_sg U62970 ( .A(\shifter_0/reg_w_13[2] ), .X(n40879) );
  nand_x1_sg U62971 ( .A(n31381), .B(n40878), .X(n13973) );
  inv_x1_sg U62972 ( .A(\shifter_0/reg_w_13[5] ), .X(n40878) );
  nand_x1_sg U62973 ( .A(n34259), .B(n40877), .X(n14004) );
  inv_x1_sg U62974 ( .A(\shifter_0/reg_w_13[6] ), .X(n40877) );
  nand_x1_sg U62975 ( .A(n34261), .B(n40876), .X(n14035) );
  inv_x1_sg U62976 ( .A(\shifter_0/reg_w_13[7] ), .X(n40876) );
  nand_x1_sg U62977 ( .A(n30087), .B(n40875), .X(n14128) );
  inv_x1_sg U62978 ( .A(\shifter_0/reg_w_13[10] ), .X(n40875) );
  nand_x1_sg U62979 ( .A(n34259), .B(n40874), .X(n14159) );
  inv_x1_sg U62980 ( .A(\shifter_0/reg_w_13[11] ), .X(n40874) );
  nand_x1_sg U62981 ( .A(n34260), .B(n40873), .X(n14252) );
  inv_x1_sg U62982 ( .A(\shifter_0/reg_w_13[14] ), .X(n40873) );
  nand_x1_sg U62983 ( .A(n30087), .B(n40872), .X(n14283) );
  inv_x1_sg U62984 ( .A(\shifter_0/reg_w_13[15] ), .X(n40872) );
  nand_x1_sg U62985 ( .A(n31801), .B(n40871), .X(n14314) );
  inv_x1_sg U62986 ( .A(\shifter_0/reg_w_13[16] ), .X(n40871) );
  nand_x1_sg U62987 ( .A(n30313), .B(n40870), .X(n14407) );
  inv_x1_sg U62988 ( .A(\shifter_0/reg_w_13[19] ), .X(n40870) );
  nand_x1_sg U62989 ( .A(n34262), .B(n41007), .X(n14439) );
  inv_x1_sg U62990 ( .A(\shifter_0/reg_i_13[0] ), .X(n41007) );
  nand_x1_sg U62991 ( .A(n31801), .B(n41006), .X(n14470) );
  inv_x1_sg U62992 ( .A(\shifter_0/reg_i_13[1] ), .X(n41006) );
  nand_x1_sg U62993 ( .A(n31381), .B(n41005), .X(n14534) );
  inv_x1_sg U62994 ( .A(\shifter_0/reg_i_13[3] ), .X(n41005) );
  nand_x1_sg U62995 ( .A(n31380), .B(n41004), .X(n14596) );
  inv_x1_sg U62996 ( .A(\shifter_0/reg_i_13[5] ), .X(n41004) );
  nand_x1_sg U62997 ( .A(n30311), .B(n41003), .X(n14627) );
  inv_x1_sg U62998 ( .A(\shifter_0/reg_i_13[6] ), .X(n41003) );
  nand_x1_sg U62999 ( .A(n30087), .B(n41002), .X(n14658) );
  inv_x1_sg U63000 ( .A(\shifter_0/reg_i_13[7] ), .X(n41002) );
  nand_x1_sg U63001 ( .A(n30311), .B(n41001), .X(n14751) );
  inv_x1_sg U63002 ( .A(\shifter_0/reg_i_13[10] ), .X(n41001) );
  nand_x1_sg U63003 ( .A(n34260), .B(n41000), .X(n14782) );
  inv_x1_sg U63004 ( .A(\shifter_0/reg_i_13[11] ), .X(n41000) );
  nand_x1_sg U63005 ( .A(n34262), .B(n40999), .X(n14875) );
  inv_x1_sg U63006 ( .A(\shifter_0/reg_i_13[14] ), .X(n40999) );
  nand_x1_sg U63007 ( .A(n30313), .B(n40998), .X(n14906) );
  inv_x1_sg U63008 ( .A(\shifter_0/reg_i_13[15] ), .X(n40998) );
  nand_x1_sg U63009 ( .A(n34261), .B(n40997), .X(n15030) );
  inv_x1_sg U63010 ( .A(\shifter_0/reg_i_13[19] ), .X(n40997) );
  nand_x1_sg U63011 ( .A(n14496), .B(\shifter_0/reg_i_10[2] ), .X(n14495) );
  nand_x1_sg U63012 ( .A(n14497), .B(n30410), .X(n14494) );
  nand_x1_sg U63013 ( .A(n30533), .B(\shifter_0/reg_i_10[4] ), .X(n14559) );
  nand_x1_sg U63014 ( .A(n30531), .B(n30414), .X(n14558) );
  nand_x1_sg U63015 ( .A(n14496), .B(\shifter_0/reg_i_10[17] ), .X(n14962) );
  nand_x1_sg U63016 ( .A(n14497), .B(n30440), .X(n14961) );
  nand_x1_sg U63017 ( .A(n30533), .B(\shifter_0/reg_i_10[18] ), .X(n14993) );
  nand_x1_sg U63018 ( .A(n30531), .B(n30442), .X(n14992) );
  nand_x1_sg U63019 ( .A(n30076), .B(n40917), .X(n13807) );
  nor_x1_sg U63020 ( .A(n13809), .B(n13810), .X(n13806) );
  inv_x1_sg U63021 ( .A(\shifter_0/reg_w_9[0] ), .X(n40917) );
  nand_x1_sg U63022 ( .A(n31413), .B(n40916), .X(n13842) );
  nor_x1_sg U63023 ( .A(n13843), .B(n13844), .X(n13841) );
  inv_x1_sg U63024 ( .A(\shifter_0/reg_w_9[1] ), .X(n40916) );
  nand_x1_sg U63025 ( .A(n34204), .B(n40915), .X(n13873) );
  nor_x1_sg U63026 ( .A(n13874), .B(n13875), .X(n13872) );
  inv_x1_sg U63027 ( .A(\shifter_0/reg_w_9[2] ), .X(n40915) );
  nand_x1_sg U63028 ( .A(n31414), .B(n42722), .X(n13904) );
  nor_x1_sg U63029 ( .A(n13905), .B(n13906), .X(n13903) );
  nor_x1_sg U63030 ( .A(\shifter_0/reg_w_10[3] ), .B(n33994), .X(n13905) );
  nand_x1_sg U63031 ( .A(n34206), .B(n42723), .X(n13935) );
  nor_x1_sg U63032 ( .A(n13936), .B(n13937), .X(n13934) );
  nor_x1_sg U63033 ( .A(\shifter_0/reg_w_10[4] ), .B(n29703), .X(n13936) );
  nand_x1_sg U63034 ( .A(n31819), .B(n40914), .X(n13966) );
  nor_x1_sg U63035 ( .A(n13967), .B(n13968), .X(n13965) );
  inv_x1_sg U63036 ( .A(\shifter_0/reg_w_9[5] ), .X(n40914) );
  nand_x1_sg U63037 ( .A(n34205), .B(n40913), .X(n13997) );
  nor_x1_sg U63038 ( .A(n13998), .B(n13999), .X(n13996) );
  inv_x1_sg U63039 ( .A(\shifter_0/reg_w_9[6] ), .X(n40913) );
  nand_x1_sg U63040 ( .A(n30076), .B(n40912), .X(n14028) );
  nor_x1_sg U63041 ( .A(n14029), .B(n14030), .X(n14027) );
  inv_x1_sg U63042 ( .A(\shifter_0/reg_w_9[7] ), .X(n40912) );
  nor_x1_sg U63043 ( .A(n14122), .B(n14123), .X(n14120) );
  inv_x1_sg U63044 ( .A(\shifter_0/reg_w_9[10] ), .X(n40911) );
  nor_x1_sg U63045 ( .A(n14153), .B(n14154), .X(n14151) );
  inv_x1_sg U63046 ( .A(\shifter_0/reg_w_9[11] ), .X(n40910) );
  nor_x1_sg U63047 ( .A(n14246), .B(n14247), .X(n14244) );
  inv_x1_sg U63048 ( .A(\shifter_0/reg_w_9[14] ), .X(n40909) );
  nor_x1_sg U63049 ( .A(n14277), .B(n14278), .X(n14275) );
  inv_x1_sg U63050 ( .A(\shifter_0/reg_w_9[15] ), .X(n40908) );
  nand_x1_sg U63051 ( .A(n34206), .B(n40907), .X(n14307) );
  nor_x1_sg U63052 ( .A(n14308), .B(n14309), .X(n14306) );
  inv_x1_sg U63053 ( .A(\shifter_0/reg_w_9[16] ), .X(n40907) );
  nand_x1_sg U63054 ( .A(n34204), .B(n42728), .X(n14338) );
  nor_x1_sg U63055 ( .A(n14339), .B(n14340), .X(n14337) );
  nor_x1_sg U63056 ( .A(\shifter_0/reg_w_10[17] ), .B(n29703), .X(n14339) );
  nand_x1_sg U63057 ( .A(n30287), .B(n42729), .X(n14369) );
  nor_x1_sg U63058 ( .A(n14370), .B(n14371), .X(n14368) );
  nor_x1_sg U63059 ( .A(\shifter_0/reg_w_10[18] ), .B(n29703), .X(n14370) );
  nand_x1_sg U63060 ( .A(n30285), .B(n40906), .X(n14400) );
  nor_x1_sg U63061 ( .A(n14401), .B(n14402), .X(n14399) );
  inv_x1_sg U63062 ( .A(\shifter_0/reg_w_9[19] ), .X(n40906) );
  nand_x1_sg U63063 ( .A(n34205), .B(n41040), .X(n14432) );
  nor_x1_sg U63064 ( .A(n14433), .B(n14434), .X(n14431) );
  inv_x1_sg U63065 ( .A(\shifter_0/reg_i_9[0] ), .X(n41040) );
  nand_x1_sg U63066 ( .A(n30076), .B(n41039), .X(n14463) );
  nor_x1_sg U63067 ( .A(n14464), .B(n14465), .X(n14462) );
  inv_x1_sg U63068 ( .A(\shifter_0/reg_i_9[1] ), .X(n41039) );
  nand_x1_sg U63069 ( .A(n34207), .B(n41038), .X(n14527) );
  nor_x1_sg U63070 ( .A(n14528), .B(n14529), .X(n14526) );
  inv_x1_sg U63071 ( .A(\shifter_0/reg_i_9[3] ), .X(n41038) );
  nand_x1_sg U63072 ( .A(n34205), .B(n41037), .X(n14589) );
  nor_x1_sg U63073 ( .A(n14590), .B(n14591), .X(n14588) );
  inv_x1_sg U63074 ( .A(\shifter_0/reg_i_9[5] ), .X(n41037) );
  nand_x1_sg U63075 ( .A(n31414), .B(n41036), .X(n14620) );
  nor_x1_sg U63076 ( .A(n14621), .B(n14622), .X(n14619) );
  inv_x1_sg U63077 ( .A(\shifter_0/reg_i_9[6] ), .X(n41036) );
  nand_x1_sg U63078 ( .A(n30287), .B(n41035), .X(n14651) );
  nor_x1_sg U63079 ( .A(n14652), .B(n14653), .X(n14650) );
  inv_x1_sg U63080 ( .A(\shifter_0/reg_i_9[7] ), .X(n41035) );
  nand_x1_sg U63081 ( .A(n30287), .B(n42612), .X(n14682) );
  nor_x1_sg U63082 ( .A(n14683), .B(n14684), .X(n14681) );
  nor_x1_sg U63083 ( .A(\shifter_0/reg_i_10[8] ), .B(n31052), .X(n14683) );
  nand_x1_sg U63084 ( .A(n34207), .B(n42613), .X(n14713) );
  nor_x1_sg U63085 ( .A(n14714), .B(n14715), .X(n14712) );
  nor_x1_sg U63086 ( .A(\shifter_0/reg_i_10[9] ), .B(n30532), .X(n14714) );
  nand_x1_sg U63087 ( .A(n30285), .B(n41034), .X(n14744) );
  nor_x1_sg U63088 ( .A(n14745), .B(n14746), .X(n14743) );
  inv_x1_sg U63089 ( .A(\shifter_0/reg_i_9[10] ), .X(n41034) );
  nand_x1_sg U63090 ( .A(n34206), .B(n41033), .X(n14775) );
  nor_x1_sg U63091 ( .A(n14776), .B(n14777), .X(n14774) );
  inv_x1_sg U63092 ( .A(\shifter_0/reg_i_9[11] ), .X(n41033) );
  nand_x1_sg U63093 ( .A(n34207), .B(n42614), .X(n14806) );
  nor_x1_sg U63094 ( .A(n14807), .B(n14808), .X(n14805) );
  nor_x1_sg U63095 ( .A(\shifter_0/reg_i_10[12] ), .B(n30022), .X(n14807) );
  nand_x1_sg U63096 ( .A(n34207), .B(n42615), .X(n14837) );
  nor_x1_sg U63097 ( .A(n14838), .B(n14839), .X(n14836) );
  nor_x1_sg U63098 ( .A(\shifter_0/reg_i_10[13] ), .B(n33995), .X(n14838) );
  nand_x1_sg U63099 ( .A(n34205), .B(n41032), .X(n14868) );
  nor_x1_sg U63100 ( .A(n14869), .B(n14870), .X(n14867) );
  inv_x1_sg U63101 ( .A(\shifter_0/reg_i_9[14] ), .X(n41032) );
  nand_x1_sg U63102 ( .A(n31414), .B(n41031), .X(n14899) );
  nor_x1_sg U63103 ( .A(n14900), .B(n14901), .X(n14898) );
  inv_x1_sg U63104 ( .A(\shifter_0/reg_i_9[15] ), .X(n41031) );
  nand_x1_sg U63105 ( .A(n31819), .B(n42617), .X(n14930) );
  nor_x1_sg U63106 ( .A(n14931), .B(n14932), .X(n14929) );
  nor_x1_sg U63107 ( .A(\shifter_0/reg_i_10[16] ), .B(n33994), .X(n14931) );
  nand_x1_sg U63108 ( .A(n30285), .B(n41030), .X(n15023) );
  nor_x1_sg U63109 ( .A(n15024), .B(n15025), .X(n15022) );
  inv_x1_sg U63110 ( .A(\shifter_0/reg_i_9[19] ), .X(n41030) );
  nor_x1_sg U63111 ( .A(n15138), .B(n15139), .X(n15133) );
  nor_x1_sg U63112 ( .A(n15135), .B(n42392), .X(n15134) );
  nor_x1_sg U63113 ( .A(\filter_0/reg_xor_i_mask[20] ), .B(n32130), .X(n15138)
         );
  nor_x1_sg U63114 ( .A(n15267), .B(n15268), .X(n15262) );
  nor_x1_sg U63115 ( .A(n15264), .B(n42389), .X(n15263) );
  nor_x1_sg U63116 ( .A(\filter_0/reg_xor_w_mask[20] ), .B(n32130), .X(n15267)
         );
  nor_x1_sg U63117 ( .A(n15131), .B(n15132), .X(n15127) );
  nor_x1_sg U63118 ( .A(n15129), .B(n15130), .X(n15128) );
  nor_x1_sg U63119 ( .A(\filter_0/reg_xor_i_mask[22] ), .B(n32135), .X(n15131)
         );
  nor_x1_sg U63120 ( .A(n15144), .B(n15145), .X(n15143) );
  nor_x1_sg U63121 ( .A(n15146), .B(n31203), .X(n15142) );
  nor_x1_sg U63122 ( .A(\filter_0/reg_xor_i_mask[27] ), .B(n32206), .X(n15144)
         );
  nor_x1_sg U63123 ( .A(n15260), .B(n15261), .X(n15256) );
  nor_x1_sg U63124 ( .A(n15258), .B(n15259), .X(n15257) );
  nor_x1_sg U63125 ( .A(\filter_0/reg_xor_w_mask[22] ), .B(n32134), .X(n15260)
         );
  nor_x1_sg U63126 ( .A(n15273), .B(n15274), .X(n15272) );
  nor_x1_sg U63127 ( .A(n15275), .B(n35306), .X(n15271) );
  nor_x1_sg U63128 ( .A(\filter_0/reg_xor_w_mask[27] ), .B(n32207), .X(n15273)
         );
  nor_x1_sg U63129 ( .A(n35614), .B(n12351), .X(\shifter_0/n7753 ) );
  nor_x1_sg U63130 ( .A(n12352), .B(n33292), .X(n12351) );
  nor_x1_sg U63131 ( .A(n31161), .B(n33809), .X(n12352) );
  nor_x1_sg U63132 ( .A(n35561), .B(n12356), .X(\shifter_0/n7749 ) );
  nor_x1_sg U63133 ( .A(n12357), .B(n33293), .X(n12356) );
  nor_x1_sg U63134 ( .A(n31163), .B(n33812), .X(n12357) );
  nor_x1_sg U63135 ( .A(n35613), .B(n12360), .X(\shifter_0/n7745 ) );
  nor_x1_sg U63136 ( .A(n12361), .B(n33292), .X(n12360) );
  nor_x1_sg U63137 ( .A(n31165), .B(n33809), .X(n12361) );
  nor_x1_sg U63138 ( .A(n35509), .B(n12364), .X(\shifter_0/n7741 ) );
  nor_x1_sg U63139 ( .A(n12365), .B(n33291), .X(n12364) );
  nor_x1_sg U63140 ( .A(n31167), .B(n33812), .X(n12365) );
  nor_x1_sg U63141 ( .A(n35604), .B(n12368), .X(\shifter_0/n7737 ) );
  nor_x1_sg U63142 ( .A(n12369), .B(n33293), .X(n12368) );
  nor_x1_sg U63143 ( .A(\shifter_0/reg_w_7[4] ), .B(n30980), .X(n12369) );
  nor_x1_sg U63144 ( .A(n35619), .B(n12372), .X(\shifter_0/n7733 ) );
  nor_x1_sg U63145 ( .A(n12373), .B(n33293), .X(n12372) );
  nor_x1_sg U63146 ( .A(n31171), .B(n33810), .X(n12373) );
  nor_x1_sg U63147 ( .A(n35514), .B(n12376), .X(\shifter_0/n7729 ) );
  nor_x1_sg U63148 ( .A(n12377), .B(n33290), .X(n12376) );
  nor_x1_sg U63149 ( .A(n31173), .B(n33811), .X(n12377) );
  nor_x1_sg U63150 ( .A(n35618), .B(n12380), .X(\shifter_0/n7725 ) );
  nor_x1_sg U63151 ( .A(n12381), .B(n33292), .X(n12380) );
  nor_x1_sg U63152 ( .A(n31175), .B(n33810), .X(n12381) );
  nor_x1_sg U63153 ( .A(n35612), .B(n12384), .X(\shifter_0/n7721 ) );
  nor_x1_sg U63154 ( .A(n12385), .B(n29915), .X(n12384) );
  nor_x1_sg U63155 ( .A(n31177), .B(n33812), .X(n12385) );
  nor_x1_sg U63156 ( .A(n35617), .B(n12388), .X(\shifter_0/n7717 ) );
  nor_x1_sg U63157 ( .A(n12389), .B(n33290), .X(n12388) );
  nor_x1_sg U63158 ( .A(n31179), .B(n30980), .X(n12389) );
  nor_x1_sg U63159 ( .A(n35602), .B(n12392), .X(\shifter_0/n7713 ) );
  nor_x1_sg U63160 ( .A(n12393), .B(n33290), .X(n12392) );
  nor_x1_sg U63161 ( .A(n31181), .B(n33812), .X(n12393) );
  nor_x1_sg U63162 ( .A(n35616), .B(n12396), .X(\shifter_0/n7709 ) );
  nor_x1_sg U63163 ( .A(n12397), .B(n33293), .X(n12396) );
  nor_x1_sg U63164 ( .A(n31183), .B(n30980), .X(n12397) );
  nor_x1_sg U63165 ( .A(n35611), .B(n12400), .X(\shifter_0/n7705 ) );
  nor_x1_sg U63166 ( .A(n12401), .B(n33291), .X(n12400) );
  nor_x1_sg U63167 ( .A(n31185), .B(n30979), .X(n12401) );
  nor_x1_sg U63168 ( .A(n35615), .B(n12404), .X(\shifter_0/n7701 ) );
  nor_x1_sg U63169 ( .A(n12405), .B(n29915), .X(n12404) );
  nor_x1_sg U63170 ( .A(n31187), .B(n33811), .X(n12405) );
  nor_x1_sg U63171 ( .A(n35610), .B(n12408), .X(\shifter_0/n7697 ) );
  nor_x1_sg U63172 ( .A(n12409), .B(n33292), .X(n12408) );
  nor_x1_sg U63173 ( .A(n31189), .B(n33811), .X(n12409) );
  nor_x1_sg U63174 ( .A(n35609), .B(n12412), .X(\shifter_0/n7693 ) );
  nor_x1_sg U63175 ( .A(n12413), .B(n33290), .X(n12412) );
  nor_x1_sg U63176 ( .A(n31191), .B(n33810), .X(n12413) );
  nor_x1_sg U63177 ( .A(n35601), .B(n12416), .X(\shifter_0/n7689 ) );
  nor_x1_sg U63178 ( .A(n12417), .B(n33291), .X(n12416) );
  nor_x1_sg U63179 ( .A(n31193), .B(n33810), .X(n12417) );
  nor_x1_sg U63180 ( .A(n35608), .B(n12420), .X(\shifter_0/n7685 ) );
  nor_x1_sg U63181 ( .A(n12421), .B(n33291), .X(n12420) );
  nor_x1_sg U63182 ( .A(n31195), .B(n33811), .X(n12421) );
  nor_x1_sg U63183 ( .A(n35607), .B(n12424), .X(\shifter_0/n7681 ) );
  nor_x1_sg U63184 ( .A(n12425), .B(n29915), .X(n12424) );
  nor_x1_sg U63185 ( .A(n31197), .B(n30979), .X(n12425) );
  nor_x1_sg U63186 ( .A(n35603), .B(n12428), .X(\shifter_0/n7677 ) );
  nor_x1_sg U63187 ( .A(n12429), .B(n29915), .X(n12428) );
  nor_x1_sg U63188 ( .A(n31199), .B(n33809), .X(n12429) );
  nor_x1_sg U63189 ( .A(n35503), .B(n12439), .X(\shifter_0/n7673 ) );
  nor_x1_sg U63190 ( .A(n12440), .B(n33878), .X(n12439) );
  nor_x1_sg U63191 ( .A(\shifter_0/reg_i_7[0] ), .B(n32923), .X(n12440) );
  nor_x1_sg U63192 ( .A(n35593), .B(n12444), .X(\shifter_0/n7669 ) );
  nor_x1_sg U63193 ( .A(n12445), .B(n33875), .X(n12444) );
  nor_x1_sg U63194 ( .A(\shifter_0/reg_i_7[1] ), .B(n32921), .X(n12445) );
  nor_x1_sg U63195 ( .A(n35592), .B(n12453), .X(\shifter_0/n7661 ) );
  nor_x1_sg U63196 ( .A(n12454), .B(n30941), .X(n12453) );
  nor_x1_sg U63197 ( .A(\shifter_0/reg_i_7[3] ), .B(n32924), .X(n12454) );
  nor_x1_sg U63198 ( .A(n35591), .B(n12462), .X(\shifter_0/n7653 ) );
  nor_x1_sg U63199 ( .A(n12463), .B(n30940), .X(n12462) );
  nor_x1_sg U63200 ( .A(\shifter_0/reg_i_7[5] ), .B(n32924), .X(n12463) );
  nor_x1_sg U63201 ( .A(n35590), .B(n12466), .X(\shifter_0/n7649 ) );
  nor_x1_sg U63202 ( .A(n12467), .B(n33877), .X(n12466) );
  nor_x1_sg U63203 ( .A(n31135), .B(n32924), .X(n12467) );
  nor_x1_sg U63204 ( .A(n35506), .B(n12470), .X(\shifter_0/n7645 ) );
  nor_x1_sg U63205 ( .A(n12471), .B(n33878), .X(n12470) );
  nor_x1_sg U63206 ( .A(\shifter_0/reg_i_7[7] ), .B(n29776), .X(n12471) );
  nor_x1_sg U63207 ( .A(n35589), .B(n12474), .X(\shifter_0/n7641 ) );
  nor_x1_sg U63208 ( .A(n12475), .B(n33876), .X(n12474) );
  nor_x1_sg U63209 ( .A(\shifter_0/reg_i_7[8] ), .B(n32923), .X(n12475) );
  nor_x1_sg U63210 ( .A(n35588), .B(n12478), .X(\shifter_0/n7637 ) );
  nor_x1_sg U63211 ( .A(n12479), .B(n33876), .X(n12478) );
  nor_x1_sg U63212 ( .A(\shifter_0/reg_i_7[9] ), .B(n32923), .X(n12479) );
  nor_x1_sg U63213 ( .A(n35513), .B(n12482), .X(\shifter_0/n7633 ) );
  nor_x1_sg U63214 ( .A(n12483), .B(n30941), .X(n12482) );
  nor_x1_sg U63215 ( .A(n31143), .B(n32921), .X(n12483) );
  nor_x1_sg U63216 ( .A(n35587), .B(n12486), .X(\shifter_0/n7629 ) );
  nor_x1_sg U63217 ( .A(n12487), .B(n33877), .X(n12486) );
  nor_x1_sg U63218 ( .A(\shifter_0/reg_i_7[11] ), .B(n32922), .X(n12487) );
  nor_x1_sg U63219 ( .A(n35586), .B(n12490), .X(\shifter_0/n7625 ) );
  nor_x1_sg U63220 ( .A(n12491), .B(n33875), .X(n12490) );
  nor_x1_sg U63221 ( .A(\shifter_0/reg_i_7[12] ), .B(n29776), .X(n12491) );
  nor_x1_sg U63222 ( .A(n35505), .B(n12494), .X(\shifter_0/n7621 ) );
  nor_x1_sg U63223 ( .A(n12495), .B(n33876), .X(n12494) );
  nor_x1_sg U63224 ( .A(\shifter_0/reg_i_7[13] ), .B(n32921), .X(n12495) );
  nor_x1_sg U63225 ( .A(n35585), .B(n12498), .X(\shifter_0/n7617 ) );
  nor_x1_sg U63226 ( .A(n12499), .B(n30940), .X(n12498) );
  nor_x1_sg U63227 ( .A(n31151), .B(n32922), .X(n12499) );
  nor_x1_sg U63228 ( .A(n35584), .B(n12502), .X(\shifter_0/n7613 ) );
  nor_x1_sg U63229 ( .A(n12503), .B(n33875), .X(n12502) );
  nor_x1_sg U63230 ( .A(n31153), .B(n32923), .X(n12503) );
  nor_x1_sg U63231 ( .A(n35512), .B(n12506), .X(\shifter_0/n7609 ) );
  nor_x1_sg U63232 ( .A(n12507), .B(n33878), .X(n12506) );
  nor_x1_sg U63233 ( .A(n31155), .B(n29776), .X(n12507) );
  nor_x1_sg U63234 ( .A(n35583), .B(n12520), .X(\shifter_0/n7597 ) );
  nor_x1_sg U63235 ( .A(n12521), .B(n33877), .X(n12520) );
  nor_x1_sg U63236 ( .A(\shifter_0/reg_i_7[19] ), .B(n32924), .X(n12521) );
  nand_x1_sg U63237 ( .A(n31993), .B(\shifter_0/reg_i_11[4] ), .X(n14562) );
  nand_x1_sg U63238 ( .A(n34255), .B(n31158), .X(n14563) );
  nand_x1_sg U63239 ( .A(n31994), .B(\shifter_0/reg_i_11[18] ), .X(n14996) );
  nand_x1_sg U63240 ( .A(n31384), .B(n31159), .X(n14997) );
  nor_x1_sg U63241 ( .A(n32001), .B(n15094), .X(n15091) );
  nor_x1_sg U63242 ( .A(n32123), .B(\filter_0/reg_xor_i_mask[2] ), .X(n15092)
         );
  nor_x1_sg U63243 ( .A(n32002), .B(n15227), .X(n15225) );
  nor_x1_sg U63244 ( .A(n32123), .B(\filter_0/reg_xor_w_mask[2] ), .X(n15226)
         );
  nand_x1_sg U63245 ( .A(n30319), .B(\shifter_0/reg_i_14[2] ), .X(n14492) );
  nand_x1_sg U63246 ( .A(n31413), .B(\shifter_0/reg_i_9[2] ), .X(n14493) );
  nand_x1_sg U63247 ( .A(n34409), .B(\shifter_0/reg_i_11[2] ), .X(n14500) );
  nand_x1_sg U63248 ( .A(n30310), .B(\shifter_0/reg_i_15[2] ), .X(n14501) );
  nand_x1_sg U63249 ( .A(n31375), .B(\shifter_0/reg_i_14[4] ), .X(n14556) );
  nand_x1_sg U63250 ( .A(n31819), .B(\shifter_0/reg_i_9[4] ), .X(n14557) );
  nand_x1_sg U63251 ( .A(n30319), .B(\shifter_0/reg_i_14[17] ), .X(n14959) );
  nand_x1_sg U63252 ( .A(n31413), .B(\shifter_0/reg_i_9[17] ), .X(n14960) );
  nand_x1_sg U63253 ( .A(n34409), .B(\shifter_0/reg_i_11[17] ), .X(n14965) );
  nand_x1_sg U63254 ( .A(n30086), .B(\shifter_0/reg_i_15[17] ), .X(n14966) );
  nand_x1_sg U63255 ( .A(n30317), .B(\shifter_0/reg_i_14[18] ), .X(n14990) );
  nand_x1_sg U63256 ( .A(n31819), .B(\shifter_0/reg_i_9[18] ), .X(n14991) );
  nand_x1_sg U63257 ( .A(n34264), .B(n40893), .X(n13802) );
  nand_x1_sg U63258 ( .A(n30317), .B(n40869), .X(n13803) );
  inv_x1_sg U63259 ( .A(\shifter_0/reg_w_12[0] ), .X(n40893) );
  nand_x1_sg U63260 ( .A(n31800), .B(n40892), .X(n13839) );
  nand_x1_sg U63261 ( .A(n34272), .B(n40868), .X(n13840) );
  inv_x1_sg U63262 ( .A(\shifter_0/reg_w_12[1] ), .X(n40892) );
  nand_x1_sg U63263 ( .A(n34265), .B(n40891), .X(n13870) );
  nand_x1_sg U63264 ( .A(n34272), .B(n40867), .X(n13871) );
  inv_x1_sg U63265 ( .A(\shifter_0/reg_w_12[2] ), .X(n40891) );
  nand_x1_sg U63266 ( .A(n31378), .B(n40890), .X(n13963) );
  nand_x1_sg U63267 ( .A(n34269), .B(n40866), .X(n13964) );
  inv_x1_sg U63268 ( .A(\shifter_0/reg_w_12[5] ), .X(n40890) );
  nand_x1_sg U63269 ( .A(n31800), .B(n40889), .X(n13994) );
  nand_x1_sg U63270 ( .A(n31374), .B(n40865), .X(n13995) );
  inv_x1_sg U63271 ( .A(\shifter_0/reg_w_12[6] ), .X(n40889) );
  nand_x1_sg U63272 ( .A(n34266), .B(n40888), .X(n14025) );
  nand_x1_sg U63273 ( .A(n34269), .B(n40864), .X(n14026) );
  inv_x1_sg U63274 ( .A(\shifter_0/reg_w_12[7] ), .X(n40888) );
  nand_x1_sg U63275 ( .A(n30316), .B(n40887), .X(n14118) );
  nand_x1_sg U63276 ( .A(n30317), .B(n40863), .X(n14119) );
  inv_x1_sg U63277 ( .A(\shifter_0/reg_w_12[10] ), .X(n40887) );
  nand_x1_sg U63278 ( .A(n34267), .B(n40886), .X(n14149) );
  nand_x1_sg U63279 ( .A(n31375), .B(n40862), .X(n14150) );
  inv_x1_sg U63280 ( .A(\shifter_0/reg_w_12[11] ), .X(n40886) );
  nand_x1_sg U63281 ( .A(n30314), .B(n40885), .X(n14242) );
  nand_x1_sg U63282 ( .A(n30089), .B(n40861), .X(n14243) );
  inv_x1_sg U63283 ( .A(\shifter_0/reg_w_12[14] ), .X(n40885) );
  nand_x1_sg U63284 ( .A(n30088), .B(n40884), .X(n14273) );
  nand_x1_sg U63285 ( .A(n30319), .B(n40860), .X(n14274) );
  inv_x1_sg U63286 ( .A(\shifter_0/reg_w_12[15] ), .X(n40884) );
  nand_x1_sg U63287 ( .A(n31378), .B(n40883), .X(n14304) );
  nand_x1_sg U63288 ( .A(n31374), .B(n40859), .X(n14305) );
  inv_x1_sg U63289 ( .A(\shifter_0/reg_w_12[16] ), .X(n40883) );
  nand_x1_sg U63290 ( .A(n30314), .B(n40882), .X(n14397) );
  nand_x1_sg U63291 ( .A(n34271), .B(n40858), .X(n14398) );
  inv_x1_sg U63292 ( .A(\shifter_0/reg_w_12[19] ), .X(n40882) );
  nand_x1_sg U63293 ( .A(n34266), .B(n41018), .X(n14429) );
  nand_x1_sg U63294 ( .A(n30089), .B(n40996), .X(n14430) );
  inv_x1_sg U63295 ( .A(\shifter_0/reg_i_12[0] ), .X(n41018) );
  nand_x1_sg U63296 ( .A(n31800), .B(n41017), .X(n14460) );
  nand_x1_sg U63297 ( .A(n31374), .B(n40995), .X(n14461) );
  inv_x1_sg U63298 ( .A(\shifter_0/reg_i_12[1] ), .X(n41017) );
  nand_x1_sg U63299 ( .A(n34264), .B(n41016), .X(n14524) );
  nand_x1_sg U63300 ( .A(n34270), .B(n40994), .X(n14525) );
  inv_x1_sg U63301 ( .A(\shifter_0/reg_i_12[3] ), .X(n41016) );
  nand_x1_sg U63302 ( .A(n31377), .B(n41015), .X(n14586) );
  nand_x1_sg U63303 ( .A(n31799), .B(n40993), .X(n14587) );
  inv_x1_sg U63304 ( .A(\shifter_0/reg_i_12[5] ), .X(n41015) );
  nand_x1_sg U63305 ( .A(n30088), .B(n41014), .X(n14617) );
  nand_x1_sg U63306 ( .A(n31799), .B(n40992), .X(n14618) );
  inv_x1_sg U63307 ( .A(\shifter_0/reg_i_12[6] ), .X(n41014) );
  nand_x1_sg U63308 ( .A(n30088), .B(n41013), .X(n14648) );
  nand_x1_sg U63309 ( .A(n31375), .B(n40991), .X(n14649) );
  inv_x1_sg U63310 ( .A(\shifter_0/reg_i_12[7] ), .X(n41013) );
  nand_x1_sg U63311 ( .A(n30088), .B(n41012), .X(n14741) );
  nand_x1_sg U63312 ( .A(n31375), .B(n40990), .X(n14742) );
  inv_x1_sg U63313 ( .A(\shifter_0/reg_i_12[10] ), .X(n41012) );
  nand_x1_sg U63314 ( .A(n30316), .B(n41011), .X(n14772) );
  nand_x1_sg U63315 ( .A(n31799), .B(n40989), .X(n14773) );
  inv_x1_sg U63316 ( .A(\shifter_0/reg_i_12[11] ), .X(n41011) );
  nand_x1_sg U63317 ( .A(n31378), .B(n41010), .X(n14865) );
  nand_x1_sg U63318 ( .A(n30089), .B(n40988), .X(n14866) );
  inv_x1_sg U63319 ( .A(\shifter_0/reg_i_12[14] ), .X(n41010) );
  nand_x1_sg U63320 ( .A(n34265), .B(n41009), .X(n14896) );
  nand_x1_sg U63321 ( .A(n34269), .B(n40987), .X(n14897) );
  inv_x1_sg U63322 ( .A(\shifter_0/reg_i_12[15] ), .X(n41009) );
  nand_x1_sg U63323 ( .A(n34266), .B(n41008), .X(n15020) );
  nand_x1_sg U63324 ( .A(n31374), .B(n40986), .X(n15021) );
  inv_x1_sg U63325 ( .A(\shifter_0/reg_i_12[19] ), .X(n41008) );
  nor_x1_sg U63326 ( .A(n29725), .B(n35254), .X(\shifter_0/n8938 ) );
  nor_x1_sg U63327 ( .A(n31794), .B(n35253), .X(\shifter_0/n8882 ) );
  nor_x1_sg U63328 ( .A(n42187), .B(n31784), .X(\filter_0/n7589 ) );
  inv_x1_sg U63329 ( .A(\filter_0/reg_i_8[18] ), .X(n42187) );
  nor_x1_sg U63330 ( .A(n42190), .B(n34312), .X(\filter_0/n7577 ) );
  inv_x1_sg U63331 ( .A(\filter_0/reg_i_8[15] ), .X(n42190) );
  nor_x1_sg U63332 ( .A(n42193), .B(n30334), .X(\filter_0/n7565 ) );
  inv_x1_sg U63333 ( .A(\filter_0/reg_i_8[12] ), .X(n42193) );
  nor_x1_sg U63334 ( .A(n42196), .B(n34311), .X(\filter_0/n7553 ) );
  inv_x1_sg U63335 ( .A(\filter_0/reg_i_8[9] ), .X(n42196) );
  nor_x1_sg U63336 ( .A(n42199), .B(n29720), .X(\filter_0/n7541 ) );
  inv_x1_sg U63337 ( .A(\filter_0/reg_i_8[6] ), .X(n42199) );
  nor_x1_sg U63338 ( .A(n42202), .B(n30334), .X(\filter_0/n7529 ) );
  inv_x1_sg U63339 ( .A(\filter_0/reg_i_8[3] ), .X(n42202) );
  nor_x1_sg U63340 ( .A(n42205), .B(n34311), .X(\filter_0/n7517 ) );
  inv_x1_sg U63341 ( .A(\filter_0/reg_i_8[0] ), .X(n42205) );
  nor_x1_sg U63342 ( .A(n42106), .B(n31781), .X(\filter_0/n7193 ) );
  inv_x1_sg U63343 ( .A(\filter_0/reg_i_12[19] ), .X(n42106) );
  nor_x1_sg U63344 ( .A(n42109), .B(n34314), .X(\filter_0/n7181 ) );
  inv_x1_sg U63345 ( .A(\filter_0/reg_i_12[16] ), .X(n42109) );
  nor_x1_sg U63346 ( .A(n42112), .B(n31781), .X(\filter_0/n7169 ) );
  inv_x1_sg U63347 ( .A(\filter_0/reg_i_12[13] ), .X(n42112) );
  nor_x1_sg U63348 ( .A(n42115), .B(n31347), .X(\filter_0/n7157 ) );
  inv_x1_sg U63349 ( .A(\filter_0/reg_i_12[10] ), .X(n42115) );
  nor_x1_sg U63350 ( .A(n42118), .B(n30098), .X(\filter_0/n7145 ) );
  inv_x1_sg U63351 ( .A(\filter_0/reg_i_12[7] ), .X(n42118) );
  nor_x1_sg U63352 ( .A(n42121), .B(n30336), .X(\filter_0/n7133 ) );
  inv_x1_sg U63353 ( .A(\filter_0/reg_i_12[4] ), .X(n42121) );
  nor_x1_sg U63354 ( .A(n42124), .B(n31782), .X(\filter_0/n7121 ) );
  inv_x1_sg U63355 ( .A(\filter_0/reg_i_12[1] ), .X(n42124) );
  nor_x1_sg U63356 ( .A(n41866), .B(n31344), .X(\filter_0/n6277 ) );
  inv_x1_sg U63357 ( .A(\filter_0/reg_w_8[19] ), .X(n41866) );
  nor_x1_sg U63358 ( .A(n41869), .B(n31344), .X(\filter_0/n6265 ) );
  inv_x1_sg U63359 ( .A(\filter_0/reg_w_8[16] ), .X(n41869) );
  nor_x1_sg U63360 ( .A(n41872), .B(n31779), .X(\filter_0/n6253 ) );
  inv_x1_sg U63361 ( .A(\filter_0/reg_w_8[13] ), .X(n41872) );
  nor_x1_sg U63362 ( .A(n41875), .B(n34320), .X(\filter_0/n6241 ) );
  inv_x1_sg U63363 ( .A(\filter_0/reg_w_8[10] ), .X(n41875) );
  nor_x1_sg U63364 ( .A(n41878), .B(n30338), .X(\filter_0/n6229 ) );
  inv_x1_sg U63365 ( .A(\filter_0/reg_w_8[7] ), .X(n41878) );
  nor_x1_sg U63366 ( .A(n41881), .B(n30338), .X(\filter_0/n6217 ) );
  inv_x1_sg U63367 ( .A(\filter_0/reg_w_8[4] ), .X(n41881) );
  nor_x1_sg U63368 ( .A(n41884), .B(n34319), .X(\filter_0/n6205 ) );
  inv_x1_sg U63369 ( .A(\filter_0/reg_w_8[1] ), .X(n41884) );
  nor_x1_sg U63370 ( .A(n41786), .B(n35629), .X(\filter_0/n5877 ) );
  inv_x1_sg U63371 ( .A(\filter_0/reg_w_12[19] ), .X(n41786) );
  nor_x1_sg U63372 ( .A(n41789), .B(n31808), .X(\filter_0/n5865 ) );
  inv_x1_sg U63373 ( .A(\filter_0/reg_w_12[16] ), .X(n41789) );
  nor_x1_sg U63374 ( .A(n41792), .B(n34242), .X(\filter_0/n5853 ) );
  inv_x1_sg U63375 ( .A(\filter_0/reg_w_12[13] ), .X(n41792) );
  nor_x1_sg U63376 ( .A(n41795), .B(n31392), .X(\filter_0/n5841 ) );
  inv_x1_sg U63377 ( .A(\filter_0/reg_w_12[10] ), .X(n41795) );
  nor_x1_sg U63378 ( .A(n41798), .B(n34240), .X(\filter_0/n5829 ) );
  inv_x1_sg U63379 ( .A(\filter_0/reg_w_12[7] ), .X(n41798) );
  nor_x1_sg U63380 ( .A(n41801), .B(n30302), .X(\filter_0/n5817 ) );
  inv_x1_sg U63381 ( .A(\filter_0/reg_w_12[4] ), .X(n41801) );
  nor_x1_sg U63382 ( .A(n41804), .B(n34241), .X(\filter_0/n5805 ) );
  inv_x1_sg U63383 ( .A(\filter_0/reg_w_12[1] ), .X(n41804) );
  nor_x1_sg U63384 ( .A(n42186), .B(n34310), .X(\filter_0/n4981 ) );
  inv_x1_sg U63385 ( .A(\filter_0/reg_i_8[19] ), .X(n42186) );
  nor_x1_sg U63386 ( .A(n42188), .B(n30097), .X(\filter_0/n7585 ) );
  inv_x1_sg U63387 ( .A(\filter_0/reg_i_8[17] ), .X(n42188) );
  nor_x1_sg U63388 ( .A(n42189), .B(n31784), .X(\filter_0/n7581 ) );
  inv_x1_sg U63389 ( .A(\filter_0/reg_i_8[16] ), .X(n42189) );
  nor_x1_sg U63390 ( .A(n42191), .B(n31351), .X(\filter_0/n7573 ) );
  inv_x1_sg U63391 ( .A(\filter_0/reg_i_8[14] ), .X(n42191) );
  nor_x1_sg U63392 ( .A(n42192), .B(n31351), .X(\filter_0/n7569 ) );
  inv_x1_sg U63393 ( .A(\filter_0/reg_i_8[13] ), .X(n42192) );
  nor_x1_sg U63394 ( .A(n42194), .B(n31784), .X(\filter_0/n7561 ) );
  inv_x1_sg U63395 ( .A(\filter_0/reg_i_8[11] ), .X(n42194) );
  nor_x1_sg U63396 ( .A(n42195), .B(n31350), .X(\filter_0/n7557 ) );
  inv_x1_sg U63397 ( .A(\filter_0/reg_i_8[10] ), .X(n42195) );
  nor_x1_sg U63398 ( .A(n42197), .B(n31351), .X(\filter_0/n7549 ) );
  inv_x1_sg U63399 ( .A(\filter_0/reg_i_8[8] ), .X(n42197) );
  nor_x1_sg U63400 ( .A(n42198), .B(n34309), .X(\filter_0/n7545 ) );
  inv_x1_sg U63401 ( .A(\filter_0/reg_i_8[7] ), .X(n42198) );
  nor_x1_sg U63402 ( .A(n42200), .B(n34310), .X(\filter_0/n7537 ) );
  inv_x1_sg U63403 ( .A(\filter_0/reg_i_8[5] ), .X(n42200) );
  nor_x1_sg U63404 ( .A(n42201), .B(n34312), .X(\filter_0/n7533 ) );
  inv_x1_sg U63405 ( .A(\filter_0/reg_i_8[4] ), .X(n42201) );
  nor_x1_sg U63406 ( .A(n42203), .B(n34312), .X(\filter_0/n7525 ) );
  inv_x1_sg U63407 ( .A(\filter_0/reg_i_8[2] ), .X(n42203) );
  nor_x1_sg U63408 ( .A(n42204), .B(n34311), .X(\filter_0/n7521 ) );
  inv_x1_sg U63409 ( .A(\filter_0/reg_i_8[1] ), .X(n42204) );
  nor_x1_sg U63410 ( .A(n42107), .B(n34317), .X(\filter_0/n7189 ) );
  inv_x1_sg U63411 ( .A(\filter_0/reg_i_12[18] ), .X(n42107) );
  nor_x1_sg U63412 ( .A(n42108), .B(n34316), .X(\filter_0/n7185 ) );
  inv_x1_sg U63413 ( .A(\filter_0/reg_i_12[17] ), .X(n42108) );
  nor_x1_sg U63414 ( .A(n42110), .B(n30098), .X(\filter_0/n7177 ) );
  inv_x1_sg U63415 ( .A(\filter_0/reg_i_12[15] ), .X(n42110) );
  nor_x1_sg U63416 ( .A(n42111), .B(n34315), .X(\filter_0/n7173 ) );
  inv_x1_sg U63417 ( .A(\filter_0/reg_i_12[14] ), .X(n42111) );
  nor_x1_sg U63418 ( .A(n42113), .B(n31348), .X(\filter_0/n7165 ) );
  inv_x1_sg U63419 ( .A(\filter_0/reg_i_12[12] ), .X(n42113) );
  nor_x1_sg U63420 ( .A(n42114), .B(n31781), .X(\filter_0/n7161 ) );
  inv_x1_sg U63421 ( .A(\filter_0/reg_i_12[11] ), .X(n42114) );
  nor_x1_sg U63422 ( .A(n42116), .B(n34314), .X(\filter_0/n7153 ) );
  inv_x1_sg U63423 ( .A(\filter_0/reg_i_12[9] ), .X(n42116) );
  nor_x1_sg U63424 ( .A(n42117), .B(n30336), .X(\filter_0/n7149 ) );
  inv_x1_sg U63425 ( .A(\filter_0/reg_i_12[8] ), .X(n42117) );
  nor_x1_sg U63426 ( .A(n42119), .B(n31347), .X(\filter_0/n7141 ) );
  inv_x1_sg U63427 ( .A(\filter_0/reg_i_12[6] ), .X(n42119) );
  nor_x1_sg U63428 ( .A(n42120), .B(n29719), .X(\filter_0/n7137 ) );
  inv_x1_sg U63429 ( .A(\filter_0/reg_i_12[5] ), .X(n42120) );
  nor_x1_sg U63430 ( .A(n42122), .B(n34314), .X(\filter_0/n7129 ) );
  inv_x1_sg U63431 ( .A(\filter_0/reg_i_12[3] ), .X(n42122) );
  nor_x1_sg U63432 ( .A(n42123), .B(n34317), .X(\filter_0/n7125 ) );
  inv_x1_sg U63433 ( .A(\filter_0/reg_i_12[2] ), .X(n42123) );
  nor_x1_sg U63434 ( .A(n42125), .B(n29719), .X(\filter_0/n7117 ) );
  inv_x1_sg U63435 ( .A(\filter_0/reg_i_12[0] ), .X(n42125) );
  nor_x1_sg U63436 ( .A(n15071), .B(n30018), .X(\filter_0/n6304 ) );
  nor_x1_sg U63437 ( .A(n15072), .B(n15073), .X(n15071) );
  nor_x1_sg U63438 ( .A(n35097), .B(n15070), .X(n15072) );
  nor_x1_sg U63439 ( .A(n31593), .B(n30542), .X(n15073) );
  nor_x1_sg U63440 ( .A(n41867), .B(n30099), .X(\filter_0/n6273 ) );
  inv_x1_sg U63441 ( .A(\filter_0/reg_w_8[18] ), .X(n41867) );
  nor_x1_sg U63442 ( .A(n41868), .B(n34322), .X(\filter_0/n6269 ) );
  inv_x1_sg U63443 ( .A(\filter_0/reg_w_8[17] ), .X(n41868) );
  nor_x1_sg U63444 ( .A(n41870), .B(n31345), .X(\filter_0/n6261 ) );
  inv_x1_sg U63445 ( .A(\filter_0/reg_w_8[15] ), .X(n41870) );
  nor_x1_sg U63446 ( .A(n41871), .B(n31779), .X(\filter_0/n6257 ) );
  inv_x1_sg U63447 ( .A(\filter_0/reg_w_8[14] ), .X(n41871) );
  nor_x1_sg U63448 ( .A(n41873), .B(n35597), .X(\filter_0/n6249 ) );
  inv_x1_sg U63449 ( .A(\filter_0/reg_w_8[12] ), .X(n41873) );
  nor_x1_sg U63450 ( .A(n41874), .B(n34321), .X(\filter_0/n6245 ) );
  inv_x1_sg U63451 ( .A(\filter_0/reg_w_8[11] ), .X(n41874) );
  nor_x1_sg U63452 ( .A(n41876), .B(n31345), .X(\filter_0/n6237 ) );
  inv_x1_sg U63453 ( .A(\filter_0/reg_w_8[9] ), .X(n41876) );
  nor_x1_sg U63454 ( .A(n41877), .B(n34322), .X(\filter_0/n6233 ) );
  inv_x1_sg U63455 ( .A(\filter_0/reg_w_8[8] ), .X(n41877) );
  nor_x1_sg U63456 ( .A(n41879), .B(n31780), .X(\filter_0/n6225 ) );
  inv_x1_sg U63457 ( .A(\filter_0/reg_w_8[6] ), .X(n41879) );
  nor_x1_sg U63458 ( .A(n41880), .B(n30338), .X(\filter_0/n6221 ) );
  inv_x1_sg U63459 ( .A(\filter_0/reg_w_8[5] ), .X(n41880) );
  nor_x1_sg U63460 ( .A(n41882), .B(n31345), .X(\filter_0/n6213 ) );
  inv_x1_sg U63461 ( .A(\filter_0/reg_w_8[3] ), .X(n41882) );
  nor_x1_sg U63462 ( .A(n41883), .B(n30099), .X(\filter_0/n6209 ) );
  inv_x1_sg U63463 ( .A(\filter_0/reg_w_8[2] ), .X(n41883) );
  nor_x1_sg U63464 ( .A(n41885), .B(n34319), .X(\filter_0/n6201 ) );
  inv_x1_sg U63465 ( .A(\filter_0/reg_w_8[0] ), .X(n41885) );
  nor_x1_sg U63466 ( .A(n41787), .B(n29730), .X(\filter_0/n5873 ) );
  inv_x1_sg U63467 ( .A(\filter_0/reg_w_12[18] ), .X(n41787) );
  nor_x1_sg U63468 ( .A(n41788), .B(n31807), .X(\filter_0/n5869 ) );
  inv_x1_sg U63469 ( .A(\filter_0/reg_w_12[17] ), .X(n41788) );
  nor_x1_sg U63470 ( .A(n41790), .B(n31808), .X(\filter_0/n5861 ) );
  inv_x1_sg U63471 ( .A(\filter_0/reg_w_12[15] ), .X(n41790) );
  nor_x1_sg U63472 ( .A(n41791), .B(n34241), .X(\filter_0/n5857 ) );
  inv_x1_sg U63473 ( .A(\filter_0/reg_w_12[14] ), .X(n41791) );
  nor_x1_sg U63474 ( .A(n41793), .B(n31393), .X(\filter_0/n5849 ) );
  inv_x1_sg U63475 ( .A(\filter_0/reg_w_12[12] ), .X(n41793) );
  nor_x1_sg U63476 ( .A(n41794), .B(n34240), .X(\filter_0/n5845 ) );
  inv_x1_sg U63477 ( .A(\filter_0/reg_w_12[11] ), .X(n41794) );
  nor_x1_sg U63478 ( .A(n41796), .B(n34241), .X(\filter_0/n5837 ) );
  inv_x1_sg U63479 ( .A(\filter_0/reg_w_12[9] ), .X(n41796) );
  nor_x1_sg U63480 ( .A(n41797), .B(n30302), .X(\filter_0/n5833 ) );
  inv_x1_sg U63481 ( .A(\filter_0/reg_w_12[8] ), .X(n41797) );
  nor_x1_sg U63482 ( .A(n41799), .B(n30083), .X(\filter_0/n5825 ) );
  inv_x1_sg U63483 ( .A(\filter_0/reg_w_12[6] ), .X(n41799) );
  nor_x1_sg U63484 ( .A(n41800), .B(n31392), .X(\filter_0/n5821 ) );
  inv_x1_sg U63485 ( .A(\filter_0/reg_w_12[5] ), .X(n41800) );
  nor_x1_sg U63486 ( .A(n41802), .B(n34242), .X(\filter_0/n5813 ) );
  inv_x1_sg U63487 ( .A(\filter_0/reg_w_12[3] ), .X(n41802) );
  nor_x1_sg U63488 ( .A(n41803), .B(n34239), .X(\filter_0/n5809 ) );
  inv_x1_sg U63489 ( .A(\filter_0/reg_w_12[2] ), .X(n41803) );
  nor_x1_sg U63490 ( .A(n41805), .B(n31808), .X(\filter_0/n5801 ) );
  inv_x1_sg U63491 ( .A(\filter_0/reg_w_12[0] ), .X(n41805) );
  nor_x1_sg U63492 ( .A(n11897), .B(n11800), .X(\shifter_0/n7913 ) );
  nor_x1_sg U63493 ( .A(n11905), .B(n29965), .X(n11897) );
  nor_x1_sg U63494 ( .A(\shifter_0/reg_w_8[0] ), .B(n33814), .X(n11905) );
  nor_x1_sg U63495 ( .A(n11909), .B(n11803), .X(\shifter_0/n7909 ) );
  nor_x1_sg U63496 ( .A(n11917), .B(n33416), .X(n11909) );
  nor_x1_sg U63497 ( .A(\shifter_0/reg_w_8[1] ), .B(n33815), .X(n11917) );
  nor_x1_sg U63498 ( .A(n11920), .B(n11805), .X(\shifter_0/n7905 ) );
  nor_x1_sg U63499 ( .A(n11928), .B(n33416), .X(n11920) );
  nor_x1_sg U63500 ( .A(\shifter_0/reg_w_8[2] ), .B(n33817), .X(n11928) );
  nor_x1_sg U63501 ( .A(n11931), .B(n11807), .X(\shifter_0/n7901 ) );
  nor_x1_sg U63502 ( .A(n11939), .B(n33415), .X(n11931) );
  nor_x1_sg U63503 ( .A(\shifter_0/reg_w_8[3] ), .B(n33816), .X(n11939) );
  nor_x1_sg U63504 ( .A(n11942), .B(n11809), .X(\shifter_0/n7897 ) );
  nor_x1_sg U63505 ( .A(n11950), .B(n29965), .X(n11942) );
  nor_x1_sg U63506 ( .A(\shifter_0/reg_w_8[4] ), .B(n33817), .X(n11950) );
  nor_x1_sg U63507 ( .A(n11953), .B(n11811), .X(\shifter_0/n7893 ) );
  nor_x1_sg U63508 ( .A(n11961), .B(n33417), .X(n11953) );
  nor_x1_sg U63509 ( .A(\shifter_0/reg_w_8[5] ), .B(n33816), .X(n11961) );
  nor_x1_sg U63510 ( .A(n11964), .B(n11813), .X(\shifter_0/n7889 ) );
  nor_x1_sg U63511 ( .A(n11972), .B(n33415), .X(n11964) );
  nor_x1_sg U63512 ( .A(\shifter_0/reg_w_8[6] ), .B(n33814), .X(n11972) );
  nor_x1_sg U63513 ( .A(n11975), .B(n11815), .X(\shifter_0/n7885 ) );
  nor_x1_sg U63514 ( .A(n11983), .B(n29965), .X(n11975) );
  nor_x1_sg U63515 ( .A(\shifter_0/reg_w_8[7] ), .B(n33816), .X(n11983) );
  nor_x1_sg U63516 ( .A(n11986), .B(n11817), .X(\shifter_0/n7881 ) );
  nor_x1_sg U63517 ( .A(n11994), .B(n33417), .X(n11986) );
  nor_x1_sg U63518 ( .A(\shifter_0/reg_w_8[8] ), .B(n33816), .X(n11994) );
  nor_x1_sg U63519 ( .A(n11997), .B(n11819), .X(\shifter_0/n7877 ) );
  nor_x1_sg U63520 ( .A(n12005), .B(n33418), .X(n11997) );
  nor_x1_sg U63521 ( .A(\shifter_0/reg_w_8[9] ), .B(n33817), .X(n12005) );
  nor_x1_sg U63522 ( .A(n12008), .B(n11821), .X(\shifter_0/n7873 ) );
  nor_x1_sg U63523 ( .A(n12016), .B(n33417), .X(n12008) );
  nor_x1_sg U63524 ( .A(\shifter_0/reg_w_8[10] ), .B(n33814), .X(n12016) );
  nor_x1_sg U63525 ( .A(n12019), .B(n11823), .X(\shifter_0/n7869 ) );
  nor_x1_sg U63526 ( .A(n12027), .B(n33418), .X(n12019) );
  nor_x1_sg U63527 ( .A(\shifter_0/reg_w_8[11] ), .B(n33815), .X(n12027) );
  nor_x1_sg U63528 ( .A(n12030), .B(n11825), .X(\shifter_0/n7865 ) );
  nor_x1_sg U63529 ( .A(n12038), .B(n33418), .X(n12030) );
  nor_x1_sg U63530 ( .A(\shifter_0/reg_w_8[12] ), .B(n33815), .X(n12038) );
  nor_x1_sg U63531 ( .A(n12041), .B(n11827), .X(\shifter_0/n7861 ) );
  nor_x1_sg U63532 ( .A(n12049), .B(n33418), .X(n12041) );
  nor_x1_sg U63533 ( .A(n30494), .B(n33815), .X(n12049) );
  nor_x1_sg U63534 ( .A(n12052), .B(n11829), .X(\shifter_0/n7857 ) );
  nor_x1_sg U63535 ( .A(n12060), .B(n33415), .X(n12052) );
  nor_x1_sg U63536 ( .A(n30496), .B(n30976), .X(n12060) );
  nor_x1_sg U63537 ( .A(n12063), .B(n11831), .X(\shifter_0/n7853 ) );
  nor_x1_sg U63538 ( .A(n12071), .B(n33416), .X(n12063) );
  nor_x1_sg U63539 ( .A(\shifter_0/reg_w_8[15] ), .B(n33817), .X(n12071) );
  nor_x1_sg U63540 ( .A(n12074), .B(n11833), .X(\shifter_0/n7849 ) );
  nor_x1_sg U63541 ( .A(n12082), .B(n33417), .X(n12074) );
  nor_x1_sg U63542 ( .A(\shifter_0/reg_w_8[16] ), .B(n30977), .X(n12082) );
  nor_x1_sg U63543 ( .A(n12085), .B(n11835), .X(\shifter_0/n7845 ) );
  nor_x1_sg U63544 ( .A(n12093), .B(n33416), .X(n12085) );
  nor_x1_sg U63545 ( .A(\shifter_0/reg_w_8[17] ), .B(n30976), .X(n12093) );
  nor_x1_sg U63546 ( .A(n12096), .B(n11837), .X(\shifter_0/n7841 ) );
  nor_x1_sg U63547 ( .A(n12104), .B(n33415), .X(n12096) );
  nor_x1_sg U63548 ( .A(\shifter_0/reg_w_8[18] ), .B(n30977), .X(n12104) );
  nor_x1_sg U63549 ( .A(n12107), .B(n11839), .X(\shifter_0/n7837 ) );
  nor_x1_sg U63550 ( .A(n12115), .B(n29965), .X(n12107) );
  nor_x1_sg U63551 ( .A(\shifter_0/reg_w_8[19] ), .B(n30976), .X(n12115) );
  nor_x1_sg U63552 ( .A(n12125), .B(n11848), .X(\shifter_0/n7833 ) );
  nor_x1_sg U63553 ( .A(n12133), .B(n29963), .X(n12125) );
  nor_x1_sg U63554 ( .A(\shifter_0/reg_i_8[0] ), .B(n30983), .X(n12133) );
  nor_x1_sg U63555 ( .A(n12137), .B(n11851), .X(\shifter_0/n7829 ) );
  nor_x1_sg U63556 ( .A(n12145), .B(n33413), .X(n12137) );
  nor_x1_sg U63557 ( .A(\shifter_0/reg_i_8[1] ), .B(n33807), .X(n12145) );
  nor_x1_sg U63558 ( .A(n12159), .B(n11855), .X(\shifter_0/n7821 ) );
  nor_x1_sg U63559 ( .A(n12167), .B(n33411), .X(n12159) );
  nor_x1_sg U63560 ( .A(\shifter_0/reg_i_8[3] ), .B(n33805), .X(n12167) );
  nor_x1_sg U63561 ( .A(n12181), .B(n11859), .X(\shifter_0/n7813 ) );
  nor_x1_sg U63562 ( .A(n12189), .B(n33413), .X(n12181) );
  nor_x1_sg U63563 ( .A(\shifter_0/reg_i_8[5] ), .B(n33804), .X(n12189) );
  nor_x1_sg U63564 ( .A(n12192), .B(n11861), .X(\shifter_0/n7809 ) );
  nor_x1_sg U63565 ( .A(n12200), .B(n33410), .X(n12192) );
  nor_x1_sg U63566 ( .A(n30418), .B(n33804), .X(n12200) );
  nor_x1_sg U63567 ( .A(n12203), .B(n11863), .X(\shifter_0/n7805 ) );
  nor_x1_sg U63568 ( .A(n12211), .B(n33411), .X(n12203) );
  nor_x1_sg U63569 ( .A(\shifter_0/reg_i_8[7] ), .B(n33807), .X(n12211) );
  nor_x1_sg U63570 ( .A(n12214), .B(n11865), .X(\shifter_0/n7801 ) );
  nor_x1_sg U63571 ( .A(n12222), .B(n33410), .X(n12214) );
  nor_x1_sg U63572 ( .A(\shifter_0/reg_i_8[8] ), .B(n30982), .X(n12222) );
  nor_x1_sg U63573 ( .A(n12225), .B(n11867), .X(\shifter_0/n7797 ) );
  nor_x1_sg U63574 ( .A(n12233), .B(n33410), .X(n12225) );
  nor_x1_sg U63575 ( .A(\shifter_0/reg_i_8[9] ), .B(n30982), .X(n12233) );
  nor_x1_sg U63576 ( .A(n12236), .B(n11869), .X(\shifter_0/n7793 ) );
  nor_x1_sg U63577 ( .A(n12244), .B(n33413), .X(n12236) );
  nor_x1_sg U63578 ( .A(n30426), .B(n33807), .X(n12244) );
  nor_x1_sg U63579 ( .A(n12247), .B(n11871), .X(\shifter_0/n7789 ) );
  nor_x1_sg U63580 ( .A(n12255), .B(n33411), .X(n12247) );
  nor_x1_sg U63581 ( .A(\shifter_0/reg_i_8[11] ), .B(n33807), .X(n12255) );
  nor_x1_sg U63582 ( .A(n12258), .B(n11873), .X(\shifter_0/n7785 ) );
  nor_x1_sg U63583 ( .A(n12266), .B(n29963), .X(n12258) );
  nor_x1_sg U63584 ( .A(\shifter_0/reg_i_8[12] ), .B(n33804), .X(n12266) );
  nor_x1_sg U63585 ( .A(n12269), .B(n11875), .X(\shifter_0/n7781 ) );
  nor_x1_sg U63586 ( .A(n12277), .B(n33411), .X(n12269) );
  nor_x1_sg U63587 ( .A(\shifter_0/reg_i_8[13] ), .B(n33806), .X(n12277) );
  nor_x1_sg U63588 ( .A(n12280), .B(n11877), .X(\shifter_0/n7777 ) );
  nor_x1_sg U63589 ( .A(n12288), .B(n33410), .X(n12280) );
  nor_x1_sg U63590 ( .A(n30434), .B(n33806), .X(n12288) );
  nor_x1_sg U63591 ( .A(n12291), .B(n11879), .X(\shifter_0/n7773 ) );
  nor_x1_sg U63592 ( .A(n12299), .B(n33412), .X(n12291) );
  nor_x1_sg U63593 ( .A(n30436), .B(n30983), .X(n12299) );
  nor_x1_sg U63594 ( .A(n12302), .B(n11881), .X(\shifter_0/n7769 ) );
  nor_x1_sg U63595 ( .A(n12310), .B(n33412), .X(n12302) );
  nor_x1_sg U63596 ( .A(n30438), .B(n33806), .X(n12310) );
  nor_x1_sg U63597 ( .A(n12335), .B(n11887), .X(\shifter_0/n7757 ) );
  nor_x1_sg U63598 ( .A(n12343), .B(n33412), .X(n12335) );
  nor_x1_sg U63599 ( .A(\shifter_0/reg_i_8[19] ), .B(n30983), .X(n12343) );
  nor_x1_sg U63600 ( .A(n12148), .B(n11853), .X(\shifter_0/n7825 ) );
  nor_x1_sg U63601 ( .A(n12156), .B(n33412), .X(n12148) );
  nor_x1_sg U63602 ( .A(\shifter_0/reg_i_8[2] ), .B(n33805), .X(n12156) );
  nor_x1_sg U63603 ( .A(n12170), .B(n11857), .X(\shifter_0/n7817 ) );
  nor_x1_sg U63604 ( .A(n12178), .B(n29963), .X(n12170) );
  nor_x1_sg U63605 ( .A(\shifter_0/reg_i_8[4] ), .B(n33805), .X(n12178) );
  nor_x1_sg U63606 ( .A(n12313), .B(n11883), .X(\shifter_0/n7765 ) );
  nor_x1_sg U63607 ( .A(n12321), .B(n29963), .X(n12313) );
  nor_x1_sg U63608 ( .A(\shifter_0/reg_i_8[17] ), .B(n30982), .X(n12321) );
  nor_x1_sg U63609 ( .A(n12324), .B(n11885), .X(\shifter_0/n7761 ) );
  nor_x1_sg U63610 ( .A(n12332), .B(n33413), .X(n12324) );
  nor_x1_sg U63611 ( .A(\shifter_0/reg_i_8[18] ), .B(n33806), .X(n12332) );
  nor_x1_sg U63612 ( .A(n42046), .B(n34229), .X(\filter_0/n7273 ) );
  inv_x1_sg U63613 ( .A(\filter_0/reg_i_15[19] ), .X(n42046) );
  nor_x1_sg U63614 ( .A(n42049), .B(n31398), .X(\filter_0/n7261 ) );
  inv_x1_sg U63615 ( .A(\filter_0/reg_i_15[16] ), .X(n42049) );
  nor_x1_sg U63616 ( .A(n42052), .B(n31812), .X(\filter_0/n7249 ) );
  inv_x1_sg U63617 ( .A(\filter_0/reg_i_15[13] ), .X(n42052) );
  nor_x1_sg U63618 ( .A(n42055), .B(n34232), .X(\filter_0/n7237 ) );
  inv_x1_sg U63619 ( .A(\filter_0/reg_i_15[10] ), .X(n42055) );
  nor_x1_sg U63620 ( .A(n42058), .B(n34230), .X(\filter_0/n7225 ) );
  inv_x1_sg U63621 ( .A(\filter_0/reg_i_15[7] ), .X(n42058) );
  nor_x1_sg U63622 ( .A(n42061), .B(n34231), .X(\filter_0/n7213 ) );
  inv_x1_sg U63623 ( .A(\filter_0/reg_i_15[4] ), .X(n42061) );
  nor_x1_sg U63624 ( .A(n42064), .B(n29732), .X(\filter_0/n7201 ) );
  inv_x1_sg U63625 ( .A(\filter_0/reg_i_15[1] ), .X(n42064) );
  nor_x1_sg U63626 ( .A(n42086), .B(n31803), .X(\filter_0/n7113 ) );
  inv_x1_sg U63627 ( .A(\filter_0/reg_i_13[19] ), .X(n42086) );
  nor_x1_sg U63628 ( .A(n42089), .B(n34250), .X(\filter_0/n7101 ) );
  inv_x1_sg U63629 ( .A(\filter_0/reg_i_13[16] ), .X(n42089) );
  nor_x1_sg U63630 ( .A(n42092), .B(n30085), .X(\filter_0/n7089 ) );
  inv_x1_sg U63631 ( .A(\filter_0/reg_i_13[13] ), .X(n42092) );
  nor_x1_sg U63632 ( .A(n42095), .B(n31804), .X(\filter_0/n7077 ) );
  inv_x1_sg U63633 ( .A(\filter_0/reg_i_13[10] ), .X(n42095) );
  nor_x1_sg U63634 ( .A(n42098), .B(n31803), .X(\filter_0/n7065 ) );
  inv_x1_sg U63635 ( .A(\filter_0/reg_i_13[7] ), .X(n42098) );
  nor_x1_sg U63636 ( .A(n42101), .B(n30085), .X(\filter_0/n7053 ) );
  inv_x1_sg U63637 ( .A(\filter_0/reg_i_13[4] ), .X(n42101) );
  nor_x1_sg U63638 ( .A(n42104), .B(n34251), .X(\filter_0/n7041 ) );
  inv_x1_sg U63639 ( .A(\filter_0/reg_i_13[1] ), .X(n42104) );
  nor_x1_sg U63640 ( .A(n42066), .B(n30350), .X(\filter_0/n7033 ) );
  inv_x1_sg U63641 ( .A(\filter_0/reg_i_14[19] ), .X(n42066) );
  nor_x1_sg U63642 ( .A(n42069), .B(n31327), .X(\filter_0/n7021 ) );
  inv_x1_sg U63643 ( .A(\filter_0/reg_i_14[16] ), .X(n42069) );
  nor_x1_sg U63644 ( .A(n42072), .B(n29712), .X(\filter_0/n7009 ) );
  inv_x1_sg U63645 ( .A(\filter_0/reg_i_14[13] ), .X(n42072) );
  nor_x1_sg U63646 ( .A(n42075), .B(n31327), .X(\filter_0/n6997 ) );
  inv_x1_sg U63647 ( .A(\filter_0/reg_i_14[10] ), .X(n42075) );
  nor_x1_sg U63648 ( .A(n42078), .B(n34350), .X(\filter_0/n6985 ) );
  inv_x1_sg U63649 ( .A(\filter_0/reg_i_14[7] ), .X(n42078) );
  nor_x1_sg U63650 ( .A(n42081), .B(n31767), .X(\filter_0/n6973 ) );
  inv_x1_sg U63651 ( .A(\filter_0/reg_i_14[4] ), .X(n42081) );
  nor_x1_sg U63652 ( .A(n42084), .B(n34349), .X(\filter_0/n6961 ) );
  inv_x1_sg U63653 ( .A(\filter_0/reg_i_14[1] ), .X(n42084) );
  nor_x1_sg U63654 ( .A(n41726), .B(n31806), .X(\filter_0/n5957 ) );
  inv_x1_sg U63655 ( .A(\filter_0/reg_w_15[19] ), .X(n41726) );
  nor_x1_sg U63656 ( .A(n41729), .B(n31390), .X(\filter_0/n5945 ) );
  inv_x1_sg U63657 ( .A(\filter_0/reg_w_15[16] ), .X(n41729) );
  nor_x1_sg U63658 ( .A(n41732), .B(n31390), .X(\filter_0/n5933 ) );
  inv_x1_sg U63659 ( .A(\filter_0/reg_w_15[13] ), .X(n41732) );
  nor_x1_sg U63660 ( .A(n41735), .B(n31389), .X(\filter_0/n5921 ) );
  inv_x1_sg U63661 ( .A(\filter_0/reg_w_15[10] ), .X(n41735) );
  nor_x1_sg U63662 ( .A(n41738), .B(n31389), .X(\filter_0/n5909 ) );
  inv_x1_sg U63663 ( .A(\filter_0/reg_w_15[7] ), .X(n41738) );
  nor_x1_sg U63664 ( .A(n41741), .B(n31390), .X(\filter_0/n5897 ) );
  inv_x1_sg U63665 ( .A(\filter_0/reg_w_15[4] ), .X(n41741) );
  nor_x1_sg U63666 ( .A(n41744), .B(n29729), .X(\filter_0/n5885 ) );
  inv_x1_sg U63667 ( .A(\filter_0/reg_w_15[1] ), .X(n41744) );
  nor_x1_sg U63668 ( .A(n41766), .B(n31341), .X(\filter_0/n5797 ) );
  inv_x1_sg U63669 ( .A(\filter_0/reg_w_13[19] ), .X(n41766) );
  nor_x1_sg U63670 ( .A(n41769), .B(n31341), .X(\filter_0/n5785 ) );
  inv_x1_sg U63671 ( .A(\filter_0/reg_w_13[16] ), .X(n41769) );
  nor_x1_sg U63672 ( .A(n41772), .B(n34327), .X(\filter_0/n5773 ) );
  inv_x1_sg U63673 ( .A(\filter_0/reg_w_13[13] ), .X(n41772) );
  nor_x1_sg U63674 ( .A(n41775), .B(n30340), .X(\filter_0/n5761 ) );
  inv_x1_sg U63675 ( .A(\filter_0/reg_w_13[10] ), .X(n41775) );
  nor_x1_sg U63676 ( .A(n41778), .B(n31342), .X(\filter_0/n5749 ) );
  inv_x1_sg U63677 ( .A(\filter_0/reg_w_13[7] ), .X(n41778) );
  nor_x1_sg U63678 ( .A(n41781), .B(n31342), .X(\filter_0/n5737 ) );
  inv_x1_sg U63679 ( .A(\filter_0/reg_w_13[4] ), .X(n41781) );
  nor_x1_sg U63680 ( .A(n41784), .B(n31777), .X(\filter_0/n5725 ) );
  inv_x1_sg U63681 ( .A(\filter_0/reg_w_13[1] ), .X(n41784) );
  nor_x1_sg U63682 ( .A(n41746), .B(n34330), .X(\filter_0/n5717 ) );
  inv_x1_sg U63683 ( .A(\filter_0/reg_w_14[19] ), .X(n41746) );
  nor_x1_sg U63684 ( .A(n41749), .B(n29716), .X(\filter_0/n5705 ) );
  inv_x1_sg U63685 ( .A(\filter_0/reg_w_14[16] ), .X(n41749) );
  nor_x1_sg U63686 ( .A(n41752), .B(n31339), .X(\filter_0/n5693 ) );
  inv_x1_sg U63687 ( .A(\filter_0/reg_w_14[13] ), .X(n41752) );
  nor_x1_sg U63688 ( .A(n41755), .B(n29716), .X(\filter_0/n5681 ) );
  inv_x1_sg U63689 ( .A(\filter_0/reg_w_14[10] ), .X(n41755) );
  nor_x1_sg U63690 ( .A(n41758), .B(n34332), .X(\filter_0/n5669 ) );
  inv_x1_sg U63691 ( .A(\filter_0/reg_w_14[7] ), .X(n41758) );
  nor_x1_sg U63692 ( .A(n41761), .B(n30101), .X(\filter_0/n5657 ) );
  inv_x1_sg U63693 ( .A(\filter_0/reg_w_14[4] ), .X(n41761) );
  nor_x1_sg U63694 ( .A(n41764), .B(n31339), .X(\filter_0/n5645 ) );
  inv_x1_sg U63695 ( .A(\filter_0/reg_w_14[1] ), .X(n41764) );
  nor_x1_sg U63696 ( .A(n42047), .B(n31811), .X(\filter_0/n7269 ) );
  inv_x1_sg U63697 ( .A(\filter_0/reg_i_15[18] ), .X(n42047) );
  nor_x1_sg U63698 ( .A(n42048), .B(n31811), .X(\filter_0/n7265 ) );
  inv_x1_sg U63699 ( .A(\filter_0/reg_i_15[17] ), .X(n42048) );
  nor_x1_sg U63700 ( .A(n42050), .B(n30298), .X(\filter_0/n7257 ) );
  inv_x1_sg U63701 ( .A(\filter_0/reg_i_15[15] ), .X(n42050) );
  nor_x1_sg U63702 ( .A(n42051), .B(n34232), .X(\filter_0/n7253 ) );
  inv_x1_sg U63703 ( .A(\filter_0/reg_i_15[14] ), .X(n42051) );
  nor_x1_sg U63704 ( .A(n42053), .B(n31399), .X(\filter_0/n7245 ) );
  inv_x1_sg U63705 ( .A(\filter_0/reg_i_15[12] ), .X(n42053) );
  nor_x1_sg U63706 ( .A(n42054), .B(n31398), .X(\filter_0/n7241 ) );
  inv_x1_sg U63707 ( .A(\filter_0/reg_i_15[11] ), .X(n42054) );
  nor_x1_sg U63708 ( .A(n42056), .B(n30298), .X(\filter_0/n7233 ) );
  inv_x1_sg U63709 ( .A(\filter_0/reg_i_15[9] ), .X(n42056) );
  nor_x1_sg U63710 ( .A(n42057), .B(n31398), .X(\filter_0/n7229 ) );
  inv_x1_sg U63711 ( .A(\filter_0/reg_i_15[8] ), .X(n42057) );
  nor_x1_sg U63712 ( .A(n42059), .B(n31399), .X(\filter_0/n7221 ) );
  inv_x1_sg U63713 ( .A(\filter_0/reg_i_15[6] ), .X(n42059) );
  nor_x1_sg U63714 ( .A(n42060), .B(n30081), .X(\filter_0/n7217 ) );
  inv_x1_sg U63715 ( .A(\filter_0/reg_i_15[5] ), .X(n42060) );
  nor_x1_sg U63716 ( .A(n42062), .B(n34232), .X(\filter_0/n7209 ) );
  inv_x1_sg U63717 ( .A(\filter_0/reg_i_15[3] ), .X(n42062) );
  nor_x1_sg U63718 ( .A(n42063), .B(n31398), .X(\filter_0/n7205 ) );
  inv_x1_sg U63719 ( .A(\filter_0/reg_i_15[2] ), .X(n42063) );
  nor_x1_sg U63720 ( .A(n42065), .B(n31811), .X(\filter_0/n7197 ) );
  inv_x1_sg U63721 ( .A(\filter_0/reg_i_15[0] ), .X(n42065) );
  nor_x1_sg U63722 ( .A(n42087), .B(n34251), .X(\filter_0/n7109 ) );
  inv_x1_sg U63723 ( .A(\filter_0/reg_i_13[18] ), .X(n42087) );
  nor_x1_sg U63724 ( .A(n42088), .B(n34251), .X(\filter_0/n7105 ) );
  inv_x1_sg U63725 ( .A(\filter_0/reg_i_13[17] ), .X(n42088) );
  nor_x1_sg U63726 ( .A(n42090), .B(n34252), .X(\filter_0/n7097 ) );
  inv_x1_sg U63727 ( .A(\filter_0/reg_i_13[15] ), .X(n42090) );
  nor_x1_sg U63728 ( .A(n42091), .B(n31803), .X(\filter_0/n7093 ) );
  inv_x1_sg U63729 ( .A(\filter_0/reg_i_13[14] ), .X(n42091) );
  nor_x1_sg U63730 ( .A(n42093), .B(n29728), .X(\filter_0/n7085 ) );
  inv_x1_sg U63731 ( .A(\filter_0/reg_i_13[12] ), .X(n42093) );
  nor_x1_sg U63732 ( .A(n42094), .B(n31804), .X(\filter_0/n7081 ) );
  inv_x1_sg U63733 ( .A(\filter_0/reg_i_13[11] ), .X(n42094) );
  nor_x1_sg U63734 ( .A(n42096), .B(n31387), .X(\filter_0/n7073 ) );
  inv_x1_sg U63735 ( .A(\filter_0/reg_i_13[9] ), .X(n42096) );
  nor_x1_sg U63736 ( .A(n42097), .B(n30306), .X(\filter_0/n7069 ) );
  inv_x1_sg U63737 ( .A(\filter_0/reg_i_13[8] ), .X(n42097) );
  nor_x1_sg U63738 ( .A(n42099), .B(n31804), .X(\filter_0/n7061 ) );
  inv_x1_sg U63739 ( .A(\filter_0/reg_i_13[6] ), .X(n42099) );
  nor_x1_sg U63740 ( .A(n42100), .B(n34249), .X(\filter_0/n7057 ) );
  inv_x1_sg U63741 ( .A(\filter_0/reg_i_13[5] ), .X(n42100) );
  nor_x1_sg U63742 ( .A(n42102), .B(n31386), .X(\filter_0/n7049 ) );
  inv_x1_sg U63743 ( .A(\filter_0/reg_i_13[3] ), .X(n42102) );
  nor_x1_sg U63744 ( .A(n42103), .B(n34250), .X(\filter_0/n7045 ) );
  inv_x1_sg U63745 ( .A(\filter_0/reg_i_13[2] ), .X(n42103) );
  nor_x1_sg U63746 ( .A(n42105), .B(n31387), .X(\filter_0/n7037 ) );
  inv_x1_sg U63747 ( .A(\filter_0/reg_i_13[0] ), .X(n42105) );
  nor_x1_sg U63748 ( .A(n42067), .B(n31768), .X(\filter_0/n7029 ) );
  inv_x1_sg U63749 ( .A(\filter_0/reg_i_14[18] ), .X(n42067) );
  nor_x1_sg U63750 ( .A(n42068), .B(n35631), .X(\filter_0/n7025 ) );
  inv_x1_sg U63751 ( .A(\filter_0/reg_i_14[17] ), .X(n42068) );
  nor_x1_sg U63752 ( .A(n42070), .B(n34349), .X(\filter_0/n7017 ) );
  inv_x1_sg U63753 ( .A(\filter_0/reg_i_14[15] ), .X(n42070) );
  nor_x1_sg U63754 ( .A(n42071), .B(n34351), .X(\filter_0/n7013 ) );
  inv_x1_sg U63755 ( .A(\filter_0/reg_i_14[14] ), .X(n42071) );
  nor_x1_sg U63756 ( .A(n42073), .B(n31326), .X(\filter_0/n7005 ) );
  inv_x1_sg U63757 ( .A(\filter_0/reg_i_14[12] ), .X(n42073) );
  nor_x1_sg U63758 ( .A(n42074), .B(n31768), .X(\filter_0/n7001 ) );
  inv_x1_sg U63759 ( .A(\filter_0/reg_i_14[11] ), .X(n42074) );
  nor_x1_sg U63760 ( .A(n42076), .B(n30350), .X(\filter_0/n6993 ) );
  inv_x1_sg U63761 ( .A(\filter_0/reg_i_14[9] ), .X(n42076) );
  nor_x1_sg U63762 ( .A(n42077), .B(n31326), .X(\filter_0/n6989 ) );
  inv_x1_sg U63763 ( .A(\filter_0/reg_i_14[8] ), .X(n42077) );
  nor_x1_sg U63764 ( .A(n42079), .B(n34349), .X(\filter_0/n6981 ) );
  inv_x1_sg U63765 ( .A(\filter_0/reg_i_14[6] ), .X(n42079) );
  nor_x1_sg U63766 ( .A(n42080), .B(n31326), .X(\filter_0/n6977 ) );
  inv_x1_sg U63767 ( .A(\filter_0/reg_i_14[5] ), .X(n42080) );
  nor_x1_sg U63768 ( .A(n42082), .B(n31767), .X(\filter_0/n6969 ) );
  inv_x1_sg U63769 ( .A(\filter_0/reg_i_14[3] ), .X(n42082) );
  nor_x1_sg U63770 ( .A(n42083), .B(n34349), .X(\filter_0/n6965 ) );
  inv_x1_sg U63771 ( .A(\filter_0/reg_i_14[2] ), .X(n42083) );
  nor_x1_sg U63772 ( .A(n42085), .B(n34351), .X(\filter_0/n6957 ) );
  inv_x1_sg U63773 ( .A(\filter_0/reg_i_14[0] ), .X(n42085) );
  nor_x1_sg U63774 ( .A(n41727), .B(n31389), .X(\filter_0/n5953 ) );
  inv_x1_sg U63775 ( .A(\filter_0/reg_w_15[18] ), .X(n41727) );
  nor_x1_sg U63776 ( .A(n41728), .B(n34244), .X(\filter_0/n5949 ) );
  inv_x1_sg U63777 ( .A(\filter_0/reg_w_15[17] ), .X(n41728) );
  nor_x1_sg U63778 ( .A(n41730), .B(n31390), .X(\filter_0/n5941 ) );
  inv_x1_sg U63779 ( .A(\filter_0/reg_w_15[15] ), .X(n41730) );
  nor_x1_sg U63780 ( .A(n41731), .B(n31805), .X(\filter_0/n5937 ) );
  inv_x1_sg U63781 ( .A(\filter_0/reg_w_15[14] ), .X(n41731) );
  nor_x1_sg U63782 ( .A(n41733), .B(n31806), .X(\filter_0/n5929 ) );
  inv_x1_sg U63783 ( .A(\filter_0/reg_w_15[12] ), .X(n41733) );
  nor_x1_sg U63784 ( .A(n41734), .B(n30084), .X(\filter_0/n5925 ) );
  inv_x1_sg U63785 ( .A(\filter_0/reg_w_15[11] ), .X(n41734) );
  nor_x1_sg U63786 ( .A(n41736), .B(n31805), .X(\filter_0/n5917 ) );
  inv_x1_sg U63787 ( .A(\filter_0/reg_w_15[9] ), .X(n41736) );
  nor_x1_sg U63788 ( .A(n41737), .B(n30304), .X(\filter_0/n5913 ) );
  inv_x1_sg U63789 ( .A(\filter_0/reg_w_15[8] ), .X(n41737) );
  nor_x1_sg U63790 ( .A(n41739), .B(n29729), .X(\filter_0/n5905 ) );
  inv_x1_sg U63791 ( .A(\filter_0/reg_w_15[6] ), .X(n41739) );
  nor_x1_sg U63792 ( .A(n41740), .B(n34244), .X(\filter_0/n5901 ) );
  inv_x1_sg U63793 ( .A(\filter_0/reg_w_15[5] ), .X(n41740) );
  nor_x1_sg U63794 ( .A(n41742), .B(n34247), .X(\filter_0/n5893 ) );
  inv_x1_sg U63795 ( .A(\filter_0/reg_w_15[3] ), .X(n41742) );
  nor_x1_sg U63796 ( .A(n41743), .B(n31805), .X(\filter_0/n5889 ) );
  inv_x1_sg U63797 ( .A(\filter_0/reg_w_15[2] ), .X(n41743) );
  nor_x1_sg U63798 ( .A(n41745), .B(n30084), .X(\filter_0/n5881 ) );
  inv_x1_sg U63799 ( .A(\filter_0/reg_w_15[0] ), .X(n41745) );
  nor_x1_sg U63800 ( .A(n41767), .B(n29717), .X(\filter_0/n5793 ) );
  inv_x1_sg U63801 ( .A(\filter_0/reg_w_13[18] ), .X(n41767) );
  nor_x1_sg U63802 ( .A(n41768), .B(n30100), .X(\filter_0/n5789 ) );
  inv_x1_sg U63803 ( .A(\filter_0/reg_w_13[17] ), .X(n41768) );
  nor_x1_sg U63804 ( .A(n41770), .B(n30100), .X(\filter_0/n5781 ) );
  inv_x1_sg U63805 ( .A(\filter_0/reg_w_13[15] ), .X(n41770) );
  nor_x1_sg U63806 ( .A(n41771), .B(n34324), .X(\filter_0/n5777 ) );
  inv_x1_sg U63807 ( .A(\filter_0/reg_w_13[14] ), .X(n41771) );
  nor_x1_sg U63808 ( .A(n41773), .B(n30340), .X(\filter_0/n5769 ) );
  inv_x1_sg U63809 ( .A(\filter_0/reg_w_13[12] ), .X(n41773) );
  nor_x1_sg U63810 ( .A(n41774), .B(n34326), .X(\filter_0/n5765 ) );
  inv_x1_sg U63811 ( .A(\filter_0/reg_w_13[11] ), .X(n41774) );
  nor_x1_sg U63812 ( .A(n41776), .B(n31778), .X(\filter_0/n5757 ) );
  inv_x1_sg U63813 ( .A(\filter_0/reg_w_13[9] ), .X(n41776) );
  nor_x1_sg U63814 ( .A(n41777), .B(n34324), .X(\filter_0/n5753 ) );
  inv_x1_sg U63815 ( .A(\filter_0/reg_w_13[8] ), .X(n41777) );
  nor_x1_sg U63816 ( .A(n41779), .B(n31778), .X(\filter_0/n5745 ) );
  inv_x1_sg U63817 ( .A(\filter_0/reg_w_13[6] ), .X(n41779) );
  nor_x1_sg U63818 ( .A(n41780), .B(n34325), .X(\filter_0/n5741 ) );
  inv_x1_sg U63819 ( .A(\filter_0/reg_w_13[5] ), .X(n41780) );
  nor_x1_sg U63820 ( .A(n41782), .B(n34326), .X(\filter_0/n5733 ) );
  inv_x1_sg U63821 ( .A(\filter_0/reg_w_13[3] ), .X(n41782) );
  nor_x1_sg U63822 ( .A(n41783), .B(n31777), .X(\filter_0/n5729 ) );
  inv_x1_sg U63823 ( .A(\filter_0/reg_w_13[2] ), .X(n41783) );
  nor_x1_sg U63824 ( .A(n41785), .B(n34327), .X(\filter_0/n5721 ) );
  inv_x1_sg U63825 ( .A(\filter_0/reg_w_13[0] ), .X(n41785) );
  nor_x1_sg U63826 ( .A(n41747), .B(n34331), .X(\filter_0/n5713 ) );
  inv_x1_sg U63827 ( .A(\filter_0/reg_w_14[18] ), .X(n41747) );
  nor_x1_sg U63828 ( .A(n41748), .B(n34332), .X(\filter_0/n5709 ) );
  inv_x1_sg U63829 ( .A(\filter_0/reg_w_14[17] ), .X(n41748) );
  nor_x1_sg U63830 ( .A(n41750), .B(n34329), .X(\filter_0/n5701 ) );
  inv_x1_sg U63831 ( .A(\filter_0/reg_w_14[15] ), .X(n41750) );
  nor_x1_sg U63832 ( .A(n41751), .B(n30342), .X(\filter_0/n5697 ) );
  inv_x1_sg U63833 ( .A(\filter_0/reg_w_14[14] ), .X(n41751) );
  nor_x1_sg U63834 ( .A(n41753), .B(n34332), .X(\filter_0/n5689 ) );
  inv_x1_sg U63835 ( .A(\filter_0/reg_w_14[12] ), .X(n41753) );
  nor_x1_sg U63836 ( .A(n41754), .B(n31776), .X(\filter_0/n5685 ) );
  inv_x1_sg U63837 ( .A(\filter_0/reg_w_14[11] ), .X(n41754) );
  nor_x1_sg U63838 ( .A(n41756), .B(n34329), .X(\filter_0/n5677 ) );
  inv_x1_sg U63839 ( .A(\filter_0/reg_w_14[9] ), .X(n41756) );
  nor_x1_sg U63840 ( .A(n41757), .B(n30342), .X(\filter_0/n5673 ) );
  inv_x1_sg U63841 ( .A(\filter_0/reg_w_14[8] ), .X(n41757) );
  nor_x1_sg U63842 ( .A(n41759), .B(n34331), .X(\filter_0/n5665 ) );
  inv_x1_sg U63843 ( .A(\filter_0/reg_w_14[6] ), .X(n41759) );
  nor_x1_sg U63844 ( .A(n41760), .B(n31339), .X(\filter_0/n5661 ) );
  inv_x1_sg U63845 ( .A(\filter_0/reg_w_14[5] ), .X(n41760) );
  nor_x1_sg U63846 ( .A(n41762), .B(n31775), .X(\filter_0/n5653 ) );
  inv_x1_sg U63847 ( .A(\filter_0/reg_w_14[3] ), .X(n41762) );
  nor_x1_sg U63848 ( .A(n41763), .B(n34330), .X(\filter_0/n5649 ) );
  inv_x1_sg U63849 ( .A(\filter_0/reg_w_14[2] ), .X(n41763) );
  nor_x1_sg U63850 ( .A(n41765), .B(n31776), .X(\filter_0/n5641 ) );
  inv_x1_sg U63851 ( .A(\filter_0/reg_w_14[0] ), .X(n41765) );
  nor_x1_sg U63852 ( .A(n15137), .B(n32002), .X(n15136) );
  nor_x1_sg U63853 ( .A(n32126), .B(\filter_0/reg_xor_i_mask[16] ), .X(n15137)
         );
  nor_x1_sg U63854 ( .A(n15266), .B(n32000), .X(n15265) );
  nor_x1_sg U63855 ( .A(n32126), .B(\filter_0/reg_xor_w_mask[16] ), .X(n15266)
         );
  nor_x1_sg U63856 ( .A(n15087), .B(n15088), .X(n15086) );
  nor_x1_sg U63857 ( .A(n32120), .B(\filter_0/reg_xor_i_mask[1] ), .X(n15087)
         );
  nor_x1_sg U63858 ( .A(n32132), .B(\filter_0/reg_xor_i_mask[4] ), .X(n15088)
         );
  nor_x1_sg U63859 ( .A(n15223), .B(n15224), .X(n15222) );
  nor_x1_sg U63860 ( .A(n32120), .B(\filter_0/reg_xor_w_mask[1] ), .X(n15223)
         );
  nor_x1_sg U63861 ( .A(n32132), .B(\filter_0/reg_xor_w_mask[4] ), .X(n15224)
         );
  nor_x1_sg U63862 ( .A(n42355), .B(n34174), .X(\filter_0/n6597 ) );
  inv_x1_sg U63863 ( .A(\filter_0/reg_i_0[10] ), .X(n42355) );
  nor_x1_sg U63864 ( .A(n42335), .B(n30095), .X(\filter_0/n6517 ) );
  inv_x1_sg U63865 ( .A(\filter_0/reg_i_1[10] ), .X(n42335) );
  nor_x1_sg U63866 ( .A(n42315), .B(n30364), .X(\filter_0/n6437 ) );
  inv_x1_sg U63867 ( .A(\filter_0/reg_i_2[10] ), .X(n42315) );
  nor_x1_sg U63868 ( .A(n42295), .B(n29741), .X(\filter_0/n6357 ) );
  inv_x1_sg U63869 ( .A(\filter_0/reg_i_3[10] ), .X(n42295) );
  nor_x1_sg U63870 ( .A(n42035), .B(n31437), .X(\filter_0/n5281 ) );
  inv_x1_sg U63871 ( .A(\filter_0/reg_w_0[10] ), .X(n42035) );
  nor_x1_sg U63872 ( .A(n42015), .B(n34289), .X(\filter_0/n5201 ) );
  inv_x1_sg U63873 ( .A(\filter_0/reg_w_1[10] ), .X(n42015) );
  nor_x1_sg U63874 ( .A(n41995), .B(n29714), .X(\filter_0/n5121 ) );
  inv_x1_sg U63875 ( .A(\filter_0/reg_w_2[10] ), .X(n41995) );
  nor_x1_sg U63876 ( .A(n41975), .B(n31441), .X(\filter_0/n5041 ) );
  inv_x1_sg U63877 ( .A(\filter_0/reg_w_3[10] ), .X(n41975) );
  nor_x1_sg U63878 ( .A(n42275), .B(n34154), .X(\filter_0/n6917 ) );
  inv_x1_sg U63879 ( .A(\filter_0/reg_i_4[10] ), .X(n42275) );
  nor_x1_sg U63880 ( .A(n42255), .B(n31354), .X(\filter_0/n6837 ) );
  inv_x1_sg U63881 ( .A(\filter_0/reg_i_5[10] ), .X(n42255) );
  nor_x1_sg U63882 ( .A(n42235), .B(n30102), .X(\filter_0/n6757 ) );
  inv_x1_sg U63883 ( .A(\filter_0/reg_i_6[10] ), .X(n42235) );
  nor_x1_sg U63884 ( .A(n42215), .B(n34150), .X(\filter_0/n6677 ) );
  inv_x1_sg U63885 ( .A(\filter_0/reg_i_7[10] ), .X(n42215) );
  nor_x1_sg U63886 ( .A(n41955), .B(n30261), .X(\filter_0/n5601 ) );
  inv_x1_sg U63887 ( .A(\filter_0/reg_w_4[10] ), .X(n41955) );
  nor_x1_sg U63888 ( .A(n41935), .B(n31790), .X(\filter_0/n5521 ) );
  inv_x1_sg U63889 ( .A(\filter_0/reg_w_5[10] ), .X(n41935) );
  nor_x1_sg U63890 ( .A(n41915), .B(n31453), .X(\filter_0/n5441 ) );
  inv_x1_sg U63891 ( .A(\filter_0/reg_w_6[10] ), .X(n41915) );
  nor_x1_sg U63892 ( .A(n41895), .B(n34135), .X(\filter_0/n5361 ) );
  inv_x1_sg U63893 ( .A(\filter_0/reg_w_7[10] ), .X(n41895) );
  nor_x1_sg U63894 ( .A(n42166), .B(n31821), .X(\filter_0/n7513 ) );
  inv_x1_sg U63895 ( .A(\filter_0/reg_i_9[19] ), .X(n42166) );
  nor_x1_sg U63896 ( .A(n42167), .B(n34199), .X(\filter_0/n7509 ) );
  inv_x1_sg U63897 ( .A(\filter_0/reg_i_9[18] ), .X(n42167) );
  nor_x1_sg U63898 ( .A(n42168), .B(n34199), .X(\filter_0/n7505 ) );
  inv_x1_sg U63899 ( .A(\filter_0/reg_i_9[17] ), .X(n42168) );
  nor_x1_sg U63900 ( .A(n42169), .B(n34199), .X(\filter_0/n7501 ) );
  inv_x1_sg U63901 ( .A(\filter_0/reg_i_9[16] ), .X(n42169) );
  nor_x1_sg U63902 ( .A(n42170), .B(n31820), .X(\filter_0/n7497 ) );
  inv_x1_sg U63903 ( .A(\filter_0/reg_i_9[15] ), .X(n42170) );
  nor_x1_sg U63904 ( .A(n42171), .B(n34199), .X(\filter_0/n7493 ) );
  inv_x1_sg U63905 ( .A(\filter_0/reg_i_9[14] ), .X(n42171) );
  nor_x1_sg U63906 ( .A(n42172), .B(n31416), .X(\filter_0/n7489 ) );
  inv_x1_sg U63907 ( .A(\filter_0/reg_i_9[13] ), .X(n42172) );
  nor_x1_sg U63908 ( .A(n42173), .B(n34201), .X(\filter_0/n7485 ) );
  inv_x1_sg U63909 ( .A(\filter_0/reg_i_9[12] ), .X(n42173) );
  nor_x1_sg U63910 ( .A(n42174), .B(n31820), .X(\filter_0/n7481 ) );
  inv_x1_sg U63911 ( .A(\filter_0/reg_i_9[11] ), .X(n42174) );
  nor_x1_sg U63912 ( .A(n42176), .B(n29735), .X(\filter_0/n7473 ) );
  inv_x1_sg U63913 ( .A(\filter_0/reg_i_9[9] ), .X(n42176) );
  nor_x1_sg U63914 ( .A(n42177), .B(n31416), .X(\filter_0/n7469 ) );
  inv_x1_sg U63915 ( .A(\filter_0/reg_i_9[8] ), .X(n42177) );
  nor_x1_sg U63916 ( .A(n42178), .B(n34201), .X(\filter_0/n7465 ) );
  inv_x1_sg U63917 ( .A(\filter_0/reg_i_9[7] ), .X(n42178) );
  nor_x1_sg U63918 ( .A(n42179), .B(n31821), .X(\filter_0/n7461 ) );
  inv_x1_sg U63919 ( .A(\filter_0/reg_i_9[6] ), .X(n42179) );
  nor_x1_sg U63920 ( .A(n42180), .B(n31417), .X(\filter_0/n7457 ) );
  inv_x1_sg U63921 ( .A(\filter_0/reg_i_9[5] ), .X(n42180) );
  nor_x1_sg U63922 ( .A(n42181), .B(n31821), .X(\filter_0/n7453 ) );
  inv_x1_sg U63923 ( .A(\filter_0/reg_i_9[4] ), .X(n42181) );
  nor_x1_sg U63924 ( .A(n42182), .B(n30075), .X(\filter_0/n7449 ) );
  inv_x1_sg U63925 ( .A(\filter_0/reg_i_9[3] ), .X(n42182) );
  nor_x1_sg U63926 ( .A(n42183), .B(n29735), .X(\filter_0/n7445 ) );
  inv_x1_sg U63927 ( .A(\filter_0/reg_i_9[2] ), .X(n42183) );
  nor_x1_sg U63928 ( .A(n42184), .B(n34200), .X(\filter_0/n7441 ) );
  inv_x1_sg U63929 ( .A(\filter_0/reg_i_9[1] ), .X(n42184) );
  nor_x1_sg U63930 ( .A(n42185), .B(n34202), .X(\filter_0/n7437 ) );
  inv_x1_sg U63931 ( .A(\filter_0/reg_i_9[0] ), .X(n42185) );
  nor_x1_sg U63932 ( .A(n42146), .B(n31419), .X(\filter_0/n7433 ) );
  inv_x1_sg U63933 ( .A(\filter_0/reg_i_10[19] ), .X(n42146) );
  nor_x1_sg U63934 ( .A(n42147), .B(n31419), .X(\filter_0/n7429 ) );
  inv_x1_sg U63935 ( .A(\filter_0/reg_i_10[18] ), .X(n42147) );
  nor_x1_sg U63936 ( .A(n42148), .B(n30074), .X(\filter_0/n7425 ) );
  inv_x1_sg U63937 ( .A(\filter_0/reg_i_10[17] ), .X(n42148) );
  nor_x1_sg U63938 ( .A(n42149), .B(n31823), .X(\filter_0/n7421 ) );
  inv_x1_sg U63939 ( .A(\filter_0/reg_i_10[16] ), .X(n42149) );
  nor_x1_sg U63940 ( .A(n42150), .B(n34194), .X(\filter_0/n7417 ) );
  inv_x1_sg U63941 ( .A(\filter_0/reg_i_10[15] ), .X(n42150) );
  nor_x1_sg U63942 ( .A(n42151), .B(n34197), .X(\filter_0/n7413 ) );
  inv_x1_sg U63943 ( .A(\filter_0/reg_i_10[14] ), .X(n42151) );
  nor_x1_sg U63944 ( .A(n42152), .B(n30074), .X(\filter_0/n7409 ) );
  inv_x1_sg U63945 ( .A(\filter_0/reg_i_10[13] ), .X(n42152) );
  nor_x1_sg U63946 ( .A(n42153), .B(n34195), .X(\filter_0/n7405 ) );
  inv_x1_sg U63947 ( .A(\filter_0/reg_i_10[12] ), .X(n42153) );
  nor_x1_sg U63948 ( .A(n42154), .B(n34196), .X(\filter_0/n7401 ) );
  inv_x1_sg U63949 ( .A(\filter_0/reg_i_10[11] ), .X(n42154) );
  nor_x1_sg U63950 ( .A(n42156), .B(n34196), .X(\filter_0/n7393 ) );
  inv_x1_sg U63951 ( .A(\filter_0/reg_i_10[9] ), .X(n42156) );
  nor_x1_sg U63952 ( .A(n42157), .B(n34194), .X(\filter_0/n7389 ) );
  inv_x1_sg U63953 ( .A(\filter_0/reg_i_10[8] ), .X(n42157) );
  nor_x1_sg U63954 ( .A(n42158), .B(n34197), .X(\filter_0/n7385 ) );
  inv_x1_sg U63955 ( .A(\filter_0/reg_i_10[7] ), .X(n42158) );
  nor_x1_sg U63956 ( .A(n42159), .B(n31823), .X(\filter_0/n7381 ) );
  inv_x1_sg U63957 ( .A(\filter_0/reg_i_10[6] ), .X(n42159) );
  nor_x1_sg U63958 ( .A(n42160), .B(n31822), .X(\filter_0/n7377 ) );
  inv_x1_sg U63959 ( .A(\filter_0/reg_i_10[5] ), .X(n42160) );
  nor_x1_sg U63960 ( .A(n42161), .B(n31419), .X(\filter_0/n7373 ) );
  inv_x1_sg U63961 ( .A(\filter_0/reg_i_10[4] ), .X(n42161) );
  nor_x1_sg U63962 ( .A(n42162), .B(n29736), .X(\filter_0/n7369 ) );
  inv_x1_sg U63963 ( .A(\filter_0/reg_i_10[3] ), .X(n42162) );
  nor_x1_sg U63964 ( .A(n42163), .B(n31420), .X(\filter_0/n7365 ) );
  inv_x1_sg U63965 ( .A(\filter_0/reg_i_10[2] ), .X(n42163) );
  nor_x1_sg U63966 ( .A(n42164), .B(n31420), .X(\filter_0/n7361 ) );
  inv_x1_sg U63967 ( .A(\filter_0/reg_i_10[1] ), .X(n42164) );
  nor_x1_sg U63968 ( .A(n42165), .B(n31822), .X(\filter_0/n7357 ) );
  inv_x1_sg U63969 ( .A(\filter_0/reg_i_10[0] ), .X(n42165) );
  nor_x1_sg U63970 ( .A(n42126), .B(n31422), .X(\filter_0/n7353 ) );
  inv_x1_sg U63971 ( .A(\filter_0/reg_i_11[19] ), .X(n42126) );
  nor_x1_sg U63972 ( .A(n42127), .B(n30279), .X(\filter_0/n7349 ) );
  inv_x1_sg U63973 ( .A(\filter_0/reg_i_11[18] ), .X(n42127) );
  nor_x1_sg U63974 ( .A(n42128), .B(n34192), .X(\filter_0/n7345 ) );
  inv_x1_sg U63975 ( .A(\filter_0/reg_i_11[17] ), .X(n42128) );
  nor_x1_sg U63976 ( .A(n42129), .B(n34189), .X(\filter_0/n7341 ) );
  inv_x1_sg U63977 ( .A(\filter_0/reg_i_11[16] ), .X(n42129) );
  nor_x1_sg U63978 ( .A(n42130), .B(n34191), .X(\filter_0/n7337 ) );
  inv_x1_sg U63979 ( .A(\filter_0/reg_i_11[15] ), .X(n42130) );
  nor_x1_sg U63980 ( .A(n42131), .B(n34189), .X(\filter_0/n7333 ) );
  inv_x1_sg U63981 ( .A(\filter_0/reg_i_11[14] ), .X(n42131) );
  nor_x1_sg U63982 ( .A(n42132), .B(n31825), .X(\filter_0/n7329 ) );
  inv_x1_sg U63983 ( .A(\filter_0/reg_i_11[13] ), .X(n42132) );
  nor_x1_sg U63984 ( .A(n42133), .B(n31423), .X(\filter_0/n7325 ) );
  inv_x1_sg U63985 ( .A(\filter_0/reg_i_11[12] ), .X(n42133) );
  nor_x1_sg U63986 ( .A(n42134), .B(n31423), .X(\filter_0/n7321 ) );
  inv_x1_sg U63987 ( .A(\filter_0/reg_i_11[11] ), .X(n42134) );
  nor_x1_sg U63988 ( .A(n42136), .B(n30279), .X(\filter_0/n7313 ) );
  inv_x1_sg U63989 ( .A(\filter_0/reg_i_11[9] ), .X(n42136) );
  nor_x1_sg U63990 ( .A(n42137), .B(n31825), .X(\filter_0/n7309 ) );
  inv_x1_sg U63991 ( .A(\filter_0/reg_i_11[8] ), .X(n42137) );
  nor_x1_sg U63992 ( .A(n42138), .B(n31423), .X(\filter_0/n7305 ) );
  inv_x1_sg U63993 ( .A(\filter_0/reg_i_11[7] ), .X(n42138) );
  nor_x1_sg U63994 ( .A(n42139), .B(n30073), .X(\filter_0/n7301 ) );
  inv_x1_sg U63995 ( .A(\filter_0/reg_i_11[6] ), .X(n42139) );
  nor_x1_sg U63996 ( .A(n42140), .B(n31824), .X(\filter_0/n7297 ) );
  inv_x1_sg U63997 ( .A(\filter_0/reg_i_11[5] ), .X(n42140) );
  nor_x1_sg U63998 ( .A(n42141), .B(n15039), .X(\filter_0/n7293 ) );
  inv_x1_sg U63999 ( .A(\filter_0/reg_i_11[4] ), .X(n42141) );
  nor_x1_sg U64000 ( .A(n42142), .B(n31422), .X(\filter_0/n7289 ) );
  inv_x1_sg U64001 ( .A(\filter_0/reg_i_11[3] ), .X(n42142) );
  nor_x1_sg U64002 ( .A(n42143), .B(n31423), .X(\filter_0/n7285 ) );
  inv_x1_sg U64003 ( .A(\filter_0/reg_i_11[2] ), .X(n42143) );
  nor_x1_sg U64004 ( .A(n42144), .B(n34189), .X(\filter_0/n7281 ) );
  inv_x1_sg U64005 ( .A(\filter_0/reg_i_11[1] ), .X(n42144) );
  nor_x1_sg U64006 ( .A(n42145), .B(n30073), .X(\filter_0/n7277 ) );
  inv_x1_sg U64007 ( .A(\filter_0/reg_i_11[0] ), .X(n42145) );
  nor_x1_sg U64008 ( .A(n41846), .B(n30072), .X(\filter_0/n6197 ) );
  inv_x1_sg U64009 ( .A(\filter_0/reg_w_9[19] ), .X(n41846) );
  nor_x1_sg U64010 ( .A(n41847), .B(n29738), .X(\filter_0/n6193 ) );
  inv_x1_sg U64011 ( .A(\filter_0/reg_w_9[18] ), .X(n41847) );
  nor_x1_sg U64012 ( .A(n41848), .B(n31426), .X(\filter_0/n6189 ) );
  inv_x1_sg U64013 ( .A(\filter_0/reg_w_9[17] ), .X(n41848) );
  nor_x1_sg U64014 ( .A(n41849), .B(n34184), .X(\filter_0/n6185 ) );
  inv_x1_sg U64015 ( .A(\filter_0/reg_w_9[16] ), .X(n41849) );
  nor_x1_sg U64016 ( .A(n41850), .B(n31426), .X(\filter_0/n6181 ) );
  inv_x1_sg U64017 ( .A(\filter_0/reg_w_9[15] ), .X(n41850) );
  nor_x1_sg U64018 ( .A(n41851), .B(n30072), .X(\filter_0/n6177 ) );
  inv_x1_sg U64019 ( .A(\filter_0/reg_w_9[14] ), .X(n41851) );
  nor_x1_sg U64020 ( .A(n41852), .B(n31827), .X(\filter_0/n6173 ) );
  inv_x1_sg U64021 ( .A(\filter_0/reg_w_9[13] ), .X(n41852) );
  nor_x1_sg U64022 ( .A(n41853), .B(n30277), .X(\filter_0/n6169 ) );
  inv_x1_sg U64023 ( .A(\filter_0/reg_w_9[12] ), .X(n41853) );
  nor_x1_sg U64024 ( .A(n41854), .B(n31826), .X(\filter_0/n6165 ) );
  inv_x1_sg U64025 ( .A(\filter_0/reg_w_9[11] ), .X(n41854) );
  nor_x1_sg U64026 ( .A(n41856), .B(n34184), .X(\filter_0/n6157 ) );
  inv_x1_sg U64027 ( .A(\filter_0/reg_w_9[9] ), .X(n41856) );
  nor_x1_sg U64028 ( .A(n41857), .B(n31827), .X(\filter_0/n6153 ) );
  inv_x1_sg U64029 ( .A(\filter_0/reg_w_9[8] ), .X(n41857) );
  nor_x1_sg U64030 ( .A(n41858), .B(n34186), .X(\filter_0/n6149 ) );
  inv_x1_sg U64031 ( .A(\filter_0/reg_w_9[7] ), .X(n41858) );
  nor_x1_sg U64032 ( .A(n41859), .B(n30072), .X(\filter_0/n6145 ) );
  inv_x1_sg U64033 ( .A(\filter_0/reg_w_9[6] ), .X(n41859) );
  nor_x1_sg U64034 ( .A(n41860), .B(n34186), .X(\filter_0/n6141 ) );
  inv_x1_sg U64035 ( .A(\filter_0/reg_w_9[5] ), .X(n41860) );
  nor_x1_sg U64036 ( .A(n41861), .B(n31826), .X(\filter_0/n6137 ) );
  inv_x1_sg U64037 ( .A(\filter_0/reg_w_9[4] ), .X(n41861) );
  nor_x1_sg U64038 ( .A(n41862), .B(n31826), .X(\filter_0/n6133 ) );
  inv_x1_sg U64039 ( .A(\filter_0/reg_w_9[3] ), .X(n41862) );
  nor_x1_sg U64040 ( .A(n41863), .B(n34185), .X(\filter_0/n6129 ) );
  inv_x1_sg U64041 ( .A(\filter_0/reg_w_9[2] ), .X(n41863) );
  nor_x1_sg U64042 ( .A(n41864), .B(n31425), .X(\filter_0/n6125 ) );
  inv_x1_sg U64043 ( .A(\filter_0/reg_w_9[1] ), .X(n41864) );
  nor_x1_sg U64044 ( .A(n41865), .B(n31426), .X(\filter_0/n6121 ) );
  inv_x1_sg U64045 ( .A(\filter_0/reg_w_9[0] ), .X(n41865) );
  nor_x1_sg U64046 ( .A(n41826), .B(n31459), .X(\filter_0/n6117 ) );
  inv_x1_sg U64047 ( .A(\filter_0/reg_w_10[19] ), .X(n41826) );
  nor_x1_sg U64048 ( .A(n41827), .B(n31849), .X(\filter_0/n6113 ) );
  inv_x1_sg U64049 ( .A(\filter_0/reg_w_10[18] ), .X(n41827) );
  nor_x1_sg U64050 ( .A(n41828), .B(n30061), .X(\filter_0/n6109 ) );
  inv_x1_sg U64051 ( .A(\filter_0/reg_w_10[17] ), .X(n41828) );
  nor_x1_sg U64052 ( .A(n41829), .B(n34129), .X(\filter_0/n6105 ) );
  inv_x1_sg U64053 ( .A(\filter_0/reg_w_10[16] ), .X(n41829) );
  nor_x1_sg U64054 ( .A(n41830), .B(n30061), .X(\filter_0/n6101 ) );
  inv_x1_sg U64055 ( .A(\filter_0/reg_w_10[15] ), .X(n41830) );
  nor_x1_sg U64056 ( .A(n41831), .B(n31458), .X(\filter_0/n6097 ) );
  inv_x1_sg U64057 ( .A(\filter_0/reg_w_10[14] ), .X(n41831) );
  nor_x1_sg U64058 ( .A(n41832), .B(n34131), .X(\filter_0/n6093 ) );
  inv_x1_sg U64059 ( .A(\filter_0/reg_w_10[13] ), .X(n41832) );
  nor_x1_sg U64060 ( .A(n41833), .B(n30060), .X(\filter_0/n6089 ) );
  inv_x1_sg U64061 ( .A(\filter_0/reg_w_10[12] ), .X(n41833) );
  nor_x1_sg U64062 ( .A(n41834), .B(n31848), .X(\filter_0/n6085 ) );
  inv_x1_sg U64063 ( .A(\filter_0/reg_w_10[11] ), .X(n41834) );
  nor_x1_sg U64064 ( .A(n41836), .B(n31849), .X(\filter_0/n6077 ) );
  inv_x1_sg U64065 ( .A(\filter_0/reg_w_10[9] ), .X(n41836) );
  nor_x1_sg U64066 ( .A(n41837), .B(n34131), .X(\filter_0/n6073 ) );
  inv_x1_sg U64067 ( .A(\filter_0/reg_w_10[8] ), .X(n41837) );
  nor_x1_sg U64068 ( .A(n41838), .B(n34132), .X(\filter_0/n6069 ) );
  inv_x1_sg U64069 ( .A(\filter_0/reg_w_10[7] ), .X(n41838) );
  nor_x1_sg U64070 ( .A(n41839), .B(n31458), .X(\filter_0/n6065 ) );
  inv_x1_sg U64071 ( .A(\filter_0/reg_w_10[6] ), .X(n41839) );
  nor_x1_sg U64072 ( .A(n41840), .B(n34130), .X(\filter_0/n6061 ) );
  inv_x1_sg U64073 ( .A(\filter_0/reg_w_10[5] ), .X(n41840) );
  nor_x1_sg U64074 ( .A(n41841), .B(n34130), .X(\filter_0/n6057 ) );
  inv_x1_sg U64075 ( .A(\filter_0/reg_w_10[4] ), .X(n41841) );
  nor_x1_sg U64076 ( .A(n41842), .B(n34130), .X(\filter_0/n6053 ) );
  inv_x1_sg U64077 ( .A(\filter_0/reg_w_10[3] ), .X(n41842) );
  nor_x1_sg U64078 ( .A(n41843), .B(n31458), .X(\filter_0/n6049 ) );
  inv_x1_sg U64079 ( .A(\filter_0/reg_w_10[2] ), .X(n41843) );
  nor_x1_sg U64080 ( .A(n41844), .B(n30061), .X(\filter_0/n6045 ) );
  inv_x1_sg U64081 ( .A(\filter_0/reg_w_10[1] ), .X(n41844) );
  nor_x1_sg U64082 ( .A(n41845), .B(n30061), .X(\filter_0/n6041 ) );
  inv_x1_sg U64083 ( .A(\filter_0/reg_w_10[0] ), .X(n41845) );
  nor_x1_sg U64084 ( .A(n41806), .B(n31429), .X(\filter_0/n6037 ) );
  inv_x1_sg U64085 ( .A(\filter_0/reg_w_11[19] ), .X(n41806) );
  nor_x1_sg U64086 ( .A(n41807), .B(n34180), .X(\filter_0/n6033 ) );
  inv_x1_sg U64087 ( .A(\filter_0/reg_w_11[18] ), .X(n41807) );
  nor_x1_sg U64088 ( .A(n41808), .B(n34182), .X(\filter_0/n6029 ) );
  inv_x1_sg U64089 ( .A(\filter_0/reg_w_11[17] ), .X(n41808) );
  nor_x1_sg U64090 ( .A(n41809), .B(n30275), .X(\filter_0/n6025 ) );
  inv_x1_sg U64091 ( .A(\filter_0/reg_w_11[16] ), .X(n41809) );
  nor_x1_sg U64092 ( .A(n41810), .B(n29739), .X(\filter_0/n6021 ) );
  inv_x1_sg U64093 ( .A(\filter_0/reg_w_11[15] ), .X(n41810) );
  nor_x1_sg U64094 ( .A(n41811), .B(n31828), .X(\filter_0/n6017 ) );
  inv_x1_sg U64095 ( .A(\filter_0/reg_w_11[14] ), .X(n41811) );
  nor_x1_sg U64096 ( .A(n41812), .B(n34182), .X(\filter_0/n6013 ) );
  inv_x1_sg U64097 ( .A(\filter_0/reg_w_11[13] ), .X(n41812) );
  nor_x1_sg U64098 ( .A(n41813), .B(n31829), .X(\filter_0/n6009 ) );
  inv_x1_sg U64099 ( .A(\filter_0/reg_w_11[12] ), .X(n41813) );
  nor_x1_sg U64100 ( .A(n41814), .B(n31429), .X(\filter_0/n6005 ) );
  inv_x1_sg U64101 ( .A(\filter_0/reg_w_11[11] ), .X(n41814) );
  nor_x1_sg U64102 ( .A(n41816), .B(n15172), .X(\filter_0/n5997 ) );
  inv_x1_sg U64103 ( .A(\filter_0/reg_w_11[9] ), .X(n41816) );
  nor_x1_sg U64104 ( .A(n41817), .B(n34182), .X(\filter_0/n5993 ) );
  inv_x1_sg U64105 ( .A(\filter_0/reg_w_11[8] ), .X(n41817) );
  nor_x1_sg U64106 ( .A(n41818), .B(n31829), .X(\filter_0/n5989 ) );
  inv_x1_sg U64107 ( .A(\filter_0/reg_w_11[7] ), .X(n41818) );
  nor_x1_sg U64108 ( .A(n41819), .B(n30071), .X(\filter_0/n5985 ) );
  inv_x1_sg U64109 ( .A(\filter_0/reg_w_11[6] ), .X(n41819) );
  nor_x1_sg U64110 ( .A(n41820), .B(n34179), .X(\filter_0/n5981 ) );
  inv_x1_sg U64111 ( .A(\filter_0/reg_w_11[5] ), .X(n41820) );
  nor_x1_sg U64112 ( .A(n41821), .B(n34181), .X(\filter_0/n5977 ) );
  inv_x1_sg U64113 ( .A(\filter_0/reg_w_11[4] ), .X(n41821) );
  nor_x1_sg U64114 ( .A(n41822), .B(n30275), .X(\filter_0/n5973 ) );
  inv_x1_sg U64115 ( .A(\filter_0/reg_w_11[3] ), .X(n41822) );
  nor_x1_sg U64116 ( .A(n41823), .B(n34180), .X(\filter_0/n5969 ) );
  inv_x1_sg U64117 ( .A(\filter_0/reg_w_11[2] ), .X(n41823) );
  nor_x1_sg U64118 ( .A(n41824), .B(n30071), .X(\filter_0/n5965 ) );
  inv_x1_sg U64119 ( .A(\filter_0/reg_w_11[1] ), .X(n41824) );
  nor_x1_sg U64120 ( .A(n41825), .B(n34179), .X(\filter_0/n5961 ) );
  inv_x1_sg U64121 ( .A(\filter_0/reg_w_11[0] ), .X(n41825) );
  nor_x1_sg U64122 ( .A(n42266), .B(n34155), .X(\filter_0/n6953 ) );
  inv_x1_sg U64123 ( .A(\filter_0/reg_i_4[19] ), .X(n42266) );
  nor_x1_sg U64124 ( .A(n42267), .B(n34154), .X(\filter_0/n6949 ) );
  inv_x1_sg U64125 ( .A(\filter_0/reg_i_4[18] ), .X(n42267) );
  nor_x1_sg U64126 ( .A(n42268), .B(n34155), .X(\filter_0/n6945 ) );
  inv_x1_sg U64127 ( .A(\filter_0/reg_i_4[17] ), .X(n42268) );
  nor_x1_sg U64128 ( .A(n42269), .B(n31838), .X(\filter_0/n6941 ) );
  inv_x1_sg U64129 ( .A(\filter_0/reg_i_4[16] ), .X(n42269) );
  nor_x1_sg U64130 ( .A(n42270), .B(n30066), .X(\filter_0/n6937 ) );
  inv_x1_sg U64131 ( .A(\filter_0/reg_i_4[15] ), .X(n42270) );
  nor_x1_sg U64132 ( .A(n42271), .B(n30265), .X(\filter_0/n6933 ) );
  inv_x1_sg U64133 ( .A(\filter_0/reg_i_4[14] ), .X(n42271) );
  nor_x1_sg U64134 ( .A(n42272), .B(n31444), .X(\filter_0/n6929 ) );
  inv_x1_sg U64135 ( .A(\filter_0/reg_i_4[13] ), .X(n42272) );
  nor_x1_sg U64136 ( .A(n42273), .B(n34157), .X(\filter_0/n6925 ) );
  inv_x1_sg U64137 ( .A(\filter_0/reg_i_4[12] ), .X(n42273) );
  nor_x1_sg U64138 ( .A(n42274), .B(n31839), .X(\filter_0/n6921 ) );
  inv_x1_sg U64139 ( .A(\filter_0/reg_i_4[11] ), .X(n42274) );
  nor_x1_sg U64140 ( .A(n42276), .B(n29744), .X(\filter_0/n6913 ) );
  inv_x1_sg U64141 ( .A(\filter_0/reg_i_4[9] ), .X(n42276) );
  nor_x1_sg U64142 ( .A(n42277), .B(n34157), .X(\filter_0/n6909 ) );
  inv_x1_sg U64143 ( .A(\filter_0/reg_i_4[8] ), .X(n42277) );
  nor_x1_sg U64144 ( .A(n42278), .B(n31838), .X(\filter_0/n6905 ) );
  inv_x1_sg U64145 ( .A(\filter_0/reg_i_4[7] ), .X(n42278) );
  nor_x1_sg U64146 ( .A(n42279), .B(n34156), .X(\filter_0/n6901 ) );
  inv_x1_sg U64147 ( .A(\filter_0/reg_i_4[6] ), .X(n42279) );
  nor_x1_sg U64148 ( .A(n42280), .B(n30066), .X(\filter_0/n6897 ) );
  inv_x1_sg U64149 ( .A(\filter_0/reg_i_4[5] ), .X(n42280) );
  nor_x1_sg U64150 ( .A(n42281), .B(n31443), .X(\filter_0/n6893 ) );
  inv_x1_sg U64151 ( .A(\filter_0/reg_i_4[4] ), .X(n42281) );
  nor_x1_sg U64152 ( .A(n42282), .B(n31444), .X(\filter_0/n6889 ) );
  inv_x1_sg U64153 ( .A(\filter_0/reg_i_4[3] ), .X(n42282) );
  nor_x1_sg U64154 ( .A(n42283), .B(n34157), .X(\filter_0/n6885 ) );
  inv_x1_sg U64155 ( .A(\filter_0/reg_i_4[2] ), .X(n42283) );
  nor_x1_sg U64156 ( .A(n42284), .B(n15044), .X(\filter_0/n6881 ) );
  inv_x1_sg U64157 ( .A(\filter_0/reg_i_4[1] ), .X(n42284) );
  nor_x1_sg U64158 ( .A(n42285), .B(n31444), .X(\filter_0/n6877 ) );
  inv_x1_sg U64159 ( .A(\filter_0/reg_i_4[0] ), .X(n42285) );
  nor_x1_sg U64160 ( .A(n42246), .B(n30332), .X(\filter_0/n6873 ) );
  inv_x1_sg U64161 ( .A(\filter_0/reg_i_5[19] ), .X(n42246) );
  nor_x1_sg U64162 ( .A(n42247), .B(n31785), .X(\filter_0/n6869 ) );
  inv_x1_sg U64163 ( .A(\filter_0/reg_i_5[18] ), .X(n42247) );
  nor_x1_sg U64164 ( .A(n42248), .B(n34304), .X(\filter_0/n6865 ) );
  inv_x1_sg U64165 ( .A(\filter_0/reg_i_5[17] ), .X(n42248) );
  nor_x1_sg U64166 ( .A(n42249), .B(n30096), .X(\filter_0/n6861 ) );
  inv_x1_sg U64167 ( .A(\filter_0/reg_i_5[16] ), .X(n42249) );
  nor_x1_sg U64168 ( .A(n42250), .B(n30332), .X(\filter_0/n6857 ) );
  inv_x1_sg U64169 ( .A(\filter_0/reg_i_5[15] ), .X(n42250) );
  nor_x1_sg U64170 ( .A(n42251), .B(n34305), .X(\filter_0/n6853 ) );
  inv_x1_sg U64171 ( .A(\filter_0/reg_i_5[14] ), .X(n42251) );
  nor_x1_sg U64172 ( .A(n42252), .B(n34304), .X(\filter_0/n6849 ) );
  inv_x1_sg U64173 ( .A(\filter_0/reg_i_5[13] ), .X(n42252) );
  nor_x1_sg U64174 ( .A(n42253), .B(n34304), .X(\filter_0/n6845 ) );
  inv_x1_sg U64175 ( .A(\filter_0/reg_i_5[12] ), .X(n42253) );
  nor_x1_sg U64176 ( .A(n42254), .B(n29721), .X(\filter_0/n6841 ) );
  inv_x1_sg U64177 ( .A(\filter_0/reg_i_5[11] ), .X(n42254) );
  nor_x1_sg U64178 ( .A(n42256), .B(n31786), .X(\filter_0/n6833 ) );
  inv_x1_sg U64179 ( .A(\filter_0/reg_i_5[9] ), .X(n42256) );
  nor_x1_sg U64180 ( .A(n42257), .B(n34307), .X(\filter_0/n6829 ) );
  inv_x1_sg U64181 ( .A(\filter_0/reg_i_5[8] ), .X(n42257) );
  nor_x1_sg U64182 ( .A(n42258), .B(n34305), .X(\filter_0/n6825 ) );
  inv_x1_sg U64183 ( .A(\filter_0/reg_i_5[7] ), .X(n42258) );
  nor_x1_sg U64184 ( .A(n42259), .B(n29721), .X(\filter_0/n6821 ) );
  inv_x1_sg U64185 ( .A(\filter_0/reg_i_5[6] ), .X(n42259) );
  nor_x1_sg U64186 ( .A(n42260), .B(n31786), .X(\filter_0/n6817 ) );
  inv_x1_sg U64187 ( .A(\filter_0/reg_i_5[5] ), .X(n42260) );
  nor_x1_sg U64188 ( .A(n42261), .B(n31354), .X(\filter_0/n6813 ) );
  inv_x1_sg U64189 ( .A(\filter_0/reg_i_5[4] ), .X(n42261) );
  nor_x1_sg U64190 ( .A(n42262), .B(n30096), .X(\filter_0/n6809 ) );
  inv_x1_sg U64191 ( .A(\filter_0/reg_i_5[3] ), .X(n42262) );
  nor_x1_sg U64192 ( .A(n42263), .B(n34306), .X(\filter_0/n6805 ) );
  inv_x1_sg U64193 ( .A(\filter_0/reg_i_5[2] ), .X(n42263) );
  nor_x1_sg U64194 ( .A(n42264), .B(n34306), .X(\filter_0/n6801 ) );
  inv_x1_sg U64195 ( .A(\filter_0/reg_i_5[1] ), .X(n42264) );
  nor_x1_sg U64196 ( .A(n42265), .B(n31785), .X(\filter_0/n6797 ) );
  inv_x1_sg U64197 ( .A(\filter_0/reg_i_5[0] ), .X(n42265) );
  nor_x1_sg U64198 ( .A(n42226), .B(n31335), .X(\filter_0/n6793 ) );
  inv_x1_sg U64199 ( .A(\filter_0/reg_i_6[19] ), .X(n42226) );
  nor_x1_sg U64200 ( .A(n42227), .B(n30344), .X(\filter_0/n6789 ) );
  inv_x1_sg U64201 ( .A(\filter_0/reg_i_6[18] ), .X(n42227) );
  nor_x1_sg U64202 ( .A(n42228), .B(n31335), .X(\filter_0/n6785 ) );
  inv_x1_sg U64203 ( .A(\filter_0/reg_i_6[17] ), .X(n42228) );
  nor_x1_sg U64204 ( .A(n42229), .B(n15047), .X(\filter_0/n6781 ) );
  inv_x1_sg U64205 ( .A(\filter_0/reg_i_6[16] ), .X(n42229) );
  nor_x1_sg U64206 ( .A(n42230), .B(n31774), .X(\filter_0/n6777 ) );
  inv_x1_sg U64207 ( .A(\filter_0/reg_i_6[15] ), .X(n42230) );
  nor_x1_sg U64208 ( .A(n42231), .B(n31773), .X(\filter_0/n6773 ) );
  inv_x1_sg U64209 ( .A(\filter_0/reg_i_6[14] ), .X(n42231) );
  nor_x1_sg U64210 ( .A(n42232), .B(n31336), .X(\filter_0/n6769 ) );
  inv_x1_sg U64211 ( .A(\filter_0/reg_i_6[13] ), .X(n42232) );
  nor_x1_sg U64212 ( .A(n42233), .B(n31335), .X(\filter_0/n6765 ) );
  inv_x1_sg U64213 ( .A(\filter_0/reg_i_6[12] ), .X(n42233) );
  nor_x1_sg U64214 ( .A(n42234), .B(n34335), .X(\filter_0/n6761 ) );
  inv_x1_sg U64215 ( .A(\filter_0/reg_i_6[11] ), .X(n42234) );
  nor_x1_sg U64216 ( .A(n42236), .B(n34334), .X(\filter_0/n6753 ) );
  inv_x1_sg U64217 ( .A(\filter_0/reg_i_6[9] ), .X(n42236) );
  nor_x1_sg U64218 ( .A(n42237), .B(n31336), .X(\filter_0/n6749 ) );
  inv_x1_sg U64219 ( .A(\filter_0/reg_i_6[8] ), .X(n42237) );
  nor_x1_sg U64220 ( .A(n42238), .B(n31773), .X(\filter_0/n6745 ) );
  inv_x1_sg U64221 ( .A(\filter_0/reg_i_6[7] ), .X(n42238) );
  nor_x1_sg U64222 ( .A(n42239), .B(n34335), .X(\filter_0/n6741 ) );
  inv_x1_sg U64223 ( .A(\filter_0/reg_i_6[6] ), .X(n42239) );
  nor_x1_sg U64224 ( .A(n42240), .B(n31336), .X(\filter_0/n6737 ) );
  inv_x1_sg U64225 ( .A(\filter_0/reg_i_6[5] ), .X(n42240) );
  nor_x1_sg U64226 ( .A(n42241), .B(n34334), .X(\filter_0/n6733 ) );
  inv_x1_sg U64227 ( .A(\filter_0/reg_i_6[4] ), .X(n42241) );
  nor_x1_sg U64228 ( .A(n42242), .B(n31773), .X(\filter_0/n6729 ) );
  inv_x1_sg U64229 ( .A(\filter_0/reg_i_6[3] ), .X(n42242) );
  nor_x1_sg U64230 ( .A(n42243), .B(n34335), .X(\filter_0/n6725 ) );
  inv_x1_sg U64231 ( .A(\filter_0/reg_i_6[2] ), .X(n42243) );
  nor_x1_sg U64232 ( .A(n42244), .B(n29715), .X(\filter_0/n6721 ) );
  inv_x1_sg U64233 ( .A(\filter_0/reg_i_6[1] ), .X(n42244) );
  nor_x1_sg U64234 ( .A(n42245), .B(n34334), .X(\filter_0/n6717 ) );
  inv_x1_sg U64235 ( .A(\filter_0/reg_i_6[0] ), .X(n42245) );
  nor_x1_sg U64236 ( .A(n42206), .B(n30263), .X(\filter_0/n6713 ) );
  inv_x1_sg U64237 ( .A(\filter_0/reg_i_7[19] ), .X(n42206) );
  nor_x1_sg U64238 ( .A(n42207), .B(n31446), .X(\filter_0/n6709 ) );
  inv_x1_sg U64239 ( .A(\filter_0/reg_i_7[18] ), .X(n42207) );
  nor_x1_sg U64240 ( .A(n42208), .B(n30263), .X(\filter_0/n6705 ) );
  inv_x1_sg U64241 ( .A(\filter_0/reg_i_7[17] ), .X(n42208) );
  nor_x1_sg U64242 ( .A(n42209), .B(n34150), .X(\filter_0/n6701 ) );
  inv_x1_sg U64243 ( .A(\filter_0/reg_i_7[16] ), .X(n42209) );
  nor_x1_sg U64244 ( .A(n42210), .B(n31840), .X(\filter_0/n6697 ) );
  inv_x1_sg U64245 ( .A(\filter_0/reg_i_7[15] ), .X(n42210) );
  nor_x1_sg U64246 ( .A(n42211), .B(n31446), .X(\filter_0/n6693 ) );
  inv_x1_sg U64247 ( .A(\filter_0/reg_i_7[14] ), .X(n42211) );
  nor_x1_sg U64248 ( .A(n42212), .B(n31447), .X(\filter_0/n6689 ) );
  inv_x1_sg U64249 ( .A(\filter_0/reg_i_7[13] ), .X(n42212) );
  nor_x1_sg U64250 ( .A(n42213), .B(n29745), .X(\filter_0/n6685 ) );
  inv_x1_sg U64251 ( .A(\filter_0/reg_i_7[12] ), .X(n42213) );
  nor_x1_sg U64252 ( .A(n42214), .B(n30065), .X(\filter_0/n6681 ) );
  inv_x1_sg U64253 ( .A(\filter_0/reg_i_7[11] ), .X(n42214) );
  nor_x1_sg U64254 ( .A(n42216), .B(n34149), .X(\filter_0/n6673 ) );
  inv_x1_sg U64255 ( .A(\filter_0/reg_i_7[9] ), .X(n42216) );
  nor_x1_sg U64256 ( .A(n42217), .B(n31841), .X(\filter_0/n6669 ) );
  inv_x1_sg U64257 ( .A(\filter_0/reg_i_7[8] ), .X(n42217) );
  nor_x1_sg U64258 ( .A(n42218), .B(n29745), .X(\filter_0/n6665 ) );
  inv_x1_sg U64259 ( .A(\filter_0/reg_i_7[7] ), .X(n42218) );
  nor_x1_sg U64260 ( .A(n42219), .B(n30065), .X(\filter_0/n6661 ) );
  inv_x1_sg U64261 ( .A(\filter_0/reg_i_7[6] ), .X(n42219) );
  nor_x1_sg U64262 ( .A(n42220), .B(n31841), .X(\filter_0/n6657 ) );
  inv_x1_sg U64263 ( .A(\filter_0/reg_i_7[5] ), .X(n42220) );
  nor_x1_sg U64264 ( .A(n42221), .B(n34149), .X(\filter_0/n6653 ) );
  inv_x1_sg U64265 ( .A(\filter_0/reg_i_7[4] ), .X(n42221) );
  nor_x1_sg U64266 ( .A(n42222), .B(n34152), .X(\filter_0/n6649 ) );
  inv_x1_sg U64267 ( .A(\filter_0/reg_i_7[3] ), .X(n42222) );
  nor_x1_sg U64268 ( .A(n42223), .B(n30065), .X(\filter_0/n6645 ) );
  inv_x1_sg U64269 ( .A(\filter_0/reg_i_7[2] ), .X(n42223) );
  nor_x1_sg U64270 ( .A(n42224), .B(n31447), .X(\filter_0/n6641 ) );
  inv_x1_sg U64271 ( .A(\filter_0/reg_i_7[1] ), .X(n42224) );
  nor_x1_sg U64272 ( .A(n42225), .B(n31447), .X(\filter_0/n6637 ) );
  inv_x1_sg U64273 ( .A(\filter_0/reg_i_7[0] ), .X(n42225) );
  nor_x1_sg U64274 ( .A(n42346), .B(n31432), .X(\filter_0/n6633 ) );
  inv_x1_sg U64275 ( .A(\filter_0/reg_i_0[19] ), .X(n42346) );
  nor_x1_sg U64276 ( .A(n42347), .B(n34177), .X(\filter_0/n6629 ) );
  inv_x1_sg U64277 ( .A(\filter_0/reg_i_0[18] ), .X(n42347) );
  nor_x1_sg U64278 ( .A(n42348), .B(n30273), .X(\filter_0/n6625 ) );
  inv_x1_sg U64279 ( .A(\filter_0/reg_i_0[17] ), .X(n42348) );
  nor_x1_sg U64280 ( .A(n42349), .B(n31830), .X(\filter_0/n6621 ) );
  inv_x1_sg U64281 ( .A(\filter_0/reg_i_0[16] ), .X(n42349) );
  nor_x1_sg U64282 ( .A(n42350), .B(n34177), .X(\filter_0/n6617 ) );
  inv_x1_sg U64283 ( .A(\filter_0/reg_i_0[15] ), .X(n42350) );
  nor_x1_sg U64284 ( .A(n42351), .B(n31432), .X(\filter_0/n6613 ) );
  inv_x1_sg U64285 ( .A(\filter_0/reg_i_0[14] ), .X(n42351) );
  nor_x1_sg U64286 ( .A(n42352), .B(n31432), .X(\filter_0/n6609 ) );
  inv_x1_sg U64287 ( .A(\filter_0/reg_i_0[13] ), .X(n42352) );
  nor_x1_sg U64288 ( .A(n42353), .B(n34174), .X(\filter_0/n6605 ) );
  inv_x1_sg U64289 ( .A(\filter_0/reg_i_0[12] ), .X(n42353) );
  nor_x1_sg U64290 ( .A(n42354), .B(n31830), .X(\filter_0/n6601 ) );
  inv_x1_sg U64291 ( .A(\filter_0/reg_i_0[11] ), .X(n42354) );
  nor_x1_sg U64292 ( .A(n42356), .B(n31830), .X(\filter_0/n6593 ) );
  inv_x1_sg U64293 ( .A(\filter_0/reg_i_0[9] ), .X(n42356) );
  nor_x1_sg U64294 ( .A(n42357), .B(n31831), .X(\filter_0/n6589 ) );
  inv_x1_sg U64295 ( .A(\filter_0/reg_i_0[8] ), .X(n42357) );
  nor_x1_sg U64296 ( .A(n42358), .B(n34175), .X(\filter_0/n6585 ) );
  inv_x1_sg U64297 ( .A(\filter_0/reg_i_0[7] ), .X(n42358) );
  nor_x1_sg U64298 ( .A(n42359), .B(n34177), .X(\filter_0/n6581 ) );
  inv_x1_sg U64299 ( .A(\filter_0/reg_i_0[6] ), .X(n42359) );
  nor_x1_sg U64300 ( .A(n42360), .B(n29740), .X(\filter_0/n6577 ) );
  inv_x1_sg U64301 ( .A(\filter_0/reg_i_0[5] ), .X(n42360) );
  nor_x1_sg U64302 ( .A(n42361), .B(n30070), .X(\filter_0/n6573 ) );
  inv_x1_sg U64303 ( .A(\filter_0/reg_i_0[4] ), .X(n42361) );
  nor_x1_sg U64304 ( .A(n42362), .B(n30070), .X(\filter_0/n6569 ) );
  inv_x1_sg U64305 ( .A(\filter_0/reg_i_0[3] ), .X(n42362) );
  nor_x1_sg U64306 ( .A(n42363), .B(n30070), .X(\filter_0/n6565 ) );
  inv_x1_sg U64307 ( .A(\filter_0/reg_i_0[2] ), .X(n42363) );
  nor_x1_sg U64308 ( .A(n42364), .B(n29740), .X(\filter_0/n6561 ) );
  inv_x1_sg U64309 ( .A(\filter_0/reg_i_0[1] ), .X(n42364) );
  nor_x1_sg U64310 ( .A(n42365), .B(n31831), .X(\filter_0/n6557 ) );
  inv_x1_sg U64311 ( .A(\filter_0/reg_i_0[0] ), .X(n42365) );
  nor_x1_sg U64312 ( .A(n42326), .B(n30330), .X(\filter_0/n6553 ) );
  inv_x1_sg U64313 ( .A(\filter_0/reg_i_1[19] ), .X(n42326) );
  nor_x1_sg U64314 ( .A(n42327), .B(n34301), .X(\filter_0/n6549 ) );
  inv_x1_sg U64315 ( .A(\filter_0/reg_i_1[18] ), .X(n42327) );
  nor_x1_sg U64316 ( .A(n42328), .B(n34299), .X(\filter_0/n6545 ) );
  inv_x1_sg U64317 ( .A(\filter_0/reg_i_1[17] ), .X(n42328) );
  nor_x1_sg U64318 ( .A(n42329), .B(n30330), .X(\filter_0/n6541 ) );
  inv_x1_sg U64319 ( .A(\filter_0/reg_i_1[16] ), .X(n42329) );
  nor_x1_sg U64320 ( .A(n42330), .B(n31357), .X(\filter_0/n6537 ) );
  inv_x1_sg U64321 ( .A(\filter_0/reg_i_1[15] ), .X(n42330) );
  nor_x1_sg U64322 ( .A(n42331), .B(n31357), .X(\filter_0/n6533 ) );
  inv_x1_sg U64323 ( .A(\filter_0/reg_i_1[14] ), .X(n42331) );
  nor_x1_sg U64324 ( .A(n42332), .B(n31788), .X(\filter_0/n6529 ) );
  inv_x1_sg U64325 ( .A(\filter_0/reg_i_1[13] ), .X(n42332) );
  nor_x1_sg U64326 ( .A(n42333), .B(n34299), .X(\filter_0/n6525 ) );
  inv_x1_sg U64327 ( .A(\filter_0/reg_i_1[12] ), .X(n42333) );
  nor_x1_sg U64328 ( .A(n42334), .B(n34300), .X(\filter_0/n6521 ) );
  inv_x1_sg U64329 ( .A(\filter_0/reg_i_1[11] ), .X(n42334) );
  nor_x1_sg U64330 ( .A(n42336), .B(n31788), .X(\filter_0/n6513 ) );
  inv_x1_sg U64331 ( .A(\filter_0/reg_i_1[9] ), .X(n42336) );
  nor_x1_sg U64332 ( .A(n42337), .B(n34302), .X(\filter_0/n6509 ) );
  inv_x1_sg U64333 ( .A(\filter_0/reg_i_1[8] ), .X(n42337) );
  nor_x1_sg U64334 ( .A(n42338), .B(n30330), .X(\filter_0/n6505 ) );
  inv_x1_sg U64335 ( .A(\filter_0/reg_i_1[7] ), .X(n42338) );
  nor_x1_sg U64336 ( .A(n42339), .B(n31356), .X(\filter_0/n6501 ) );
  inv_x1_sg U64337 ( .A(\filter_0/reg_i_1[6] ), .X(n42339) );
  nor_x1_sg U64338 ( .A(n42340), .B(n34302), .X(\filter_0/n6497 ) );
  inv_x1_sg U64339 ( .A(\filter_0/reg_i_1[5] ), .X(n42340) );
  nor_x1_sg U64340 ( .A(n42341), .B(n34300), .X(\filter_0/n6493 ) );
  inv_x1_sg U64341 ( .A(\filter_0/reg_i_1[4] ), .X(n42341) );
  nor_x1_sg U64342 ( .A(n42342), .B(n34302), .X(\filter_0/n6489 ) );
  inv_x1_sg U64343 ( .A(\filter_0/reg_i_1[3] ), .X(n42342) );
  nor_x1_sg U64344 ( .A(n42343), .B(n34299), .X(\filter_0/n6485 ) );
  inv_x1_sg U64345 ( .A(\filter_0/reg_i_1[2] ), .X(n42343) );
  nor_x1_sg U64346 ( .A(n42344), .B(n29722), .X(\filter_0/n6481 ) );
  inv_x1_sg U64347 ( .A(\filter_0/reg_i_1[1] ), .X(n42344) );
  nor_x1_sg U64348 ( .A(n42345), .B(n34301), .X(\filter_0/n6477 ) );
  inv_x1_sg U64349 ( .A(\filter_0/reg_i_1[0] ), .X(n42345) );
  nor_x1_sg U64350 ( .A(n42306), .B(n31306), .X(\filter_0/n6473 ) );
  inv_x1_sg U64351 ( .A(\filter_0/reg_i_2[19] ), .X(n42306) );
  nor_x1_sg U64352 ( .A(n42307), .B(n34385), .X(\filter_0/n6469 ) );
  inv_x1_sg U64353 ( .A(\filter_0/reg_i_2[18] ), .X(n42307) );
  nor_x1_sg U64354 ( .A(n42308), .B(n31306), .X(\filter_0/n6465 ) );
  inv_x1_sg U64355 ( .A(\filter_0/reg_i_2[17] ), .X(n42308) );
  nor_x1_sg U64356 ( .A(n42309), .B(n31754), .X(\filter_0/n6461 ) );
  inv_x1_sg U64357 ( .A(\filter_0/reg_i_2[16] ), .X(n42309) );
  nor_x1_sg U64358 ( .A(n42310), .B(n31305), .X(\filter_0/n6457 ) );
  inv_x1_sg U64359 ( .A(\filter_0/reg_i_2[15] ), .X(n42310) );
  nor_x1_sg U64360 ( .A(n42311), .B(n34385), .X(\filter_0/n6453 ) );
  inv_x1_sg U64361 ( .A(\filter_0/reg_i_2[14] ), .X(n42311) );
  nor_x1_sg U64362 ( .A(n42312), .B(n31754), .X(\filter_0/n6449 ) );
  inv_x1_sg U64363 ( .A(\filter_0/reg_i_2[13] ), .X(n42312) );
  nor_x1_sg U64364 ( .A(n42313), .B(n30364), .X(\filter_0/n6445 ) );
  inv_x1_sg U64365 ( .A(\filter_0/reg_i_2[12] ), .X(n42313) );
  nor_x1_sg U64366 ( .A(n42314), .B(n30112), .X(\filter_0/n6441 ) );
  inv_x1_sg U64367 ( .A(\filter_0/reg_i_2[11] ), .X(n42314) );
  nor_x1_sg U64368 ( .A(n42316), .B(n34384), .X(\filter_0/n6433 ) );
  inv_x1_sg U64369 ( .A(\filter_0/reg_i_2[9] ), .X(n42316) );
  nor_x1_sg U64370 ( .A(n42317), .B(n34387), .X(\filter_0/n6429 ) );
  inv_x1_sg U64371 ( .A(\filter_0/reg_i_2[8] ), .X(n42317) );
  nor_x1_sg U64372 ( .A(n42318), .B(n31305), .X(\filter_0/n6425 ) );
  inv_x1_sg U64373 ( .A(\filter_0/reg_i_2[7] ), .X(n42318) );
  nor_x1_sg U64374 ( .A(n42319), .B(n34387), .X(\filter_0/n6421 ) );
  inv_x1_sg U64375 ( .A(\filter_0/reg_i_2[6] ), .X(n42319) );
  nor_x1_sg U64376 ( .A(n42320), .B(n34386), .X(\filter_0/n6417 ) );
  inv_x1_sg U64377 ( .A(\filter_0/reg_i_2[5] ), .X(n42320) );
  nor_x1_sg U64378 ( .A(n42321), .B(n31753), .X(\filter_0/n6413 ) );
  inv_x1_sg U64379 ( .A(\filter_0/reg_i_2[4] ), .X(n42321) );
  nor_x1_sg U64380 ( .A(n42322), .B(n34384), .X(\filter_0/n6409 ) );
  inv_x1_sg U64381 ( .A(\filter_0/reg_i_2[3] ), .X(n42322) );
  nor_x1_sg U64382 ( .A(n42323), .B(n31305), .X(\filter_0/n6405 ) );
  inv_x1_sg U64383 ( .A(\filter_0/reg_i_2[2] ), .X(n42323) );
  nor_x1_sg U64384 ( .A(n42324), .B(n34386), .X(\filter_0/n6401 ) );
  inv_x1_sg U64385 ( .A(\filter_0/reg_i_2[1] ), .X(n42324) );
  nor_x1_sg U64386 ( .A(n42325), .B(n30112), .X(\filter_0/n6397 ) );
  inv_x1_sg U64387 ( .A(\filter_0/reg_i_2[0] ), .X(n42325) );
  nor_x1_sg U64388 ( .A(n42286), .B(n34172), .X(\filter_0/n6393 ) );
  inv_x1_sg U64389 ( .A(\filter_0/reg_i_3[19] ), .X(n42286) );
  nor_x1_sg U64390 ( .A(n42287), .B(n30069), .X(\filter_0/n6389 ) );
  inv_x1_sg U64391 ( .A(\filter_0/reg_i_3[18] ), .X(n42287) );
  nor_x1_sg U64392 ( .A(n42288), .B(n30069), .X(\filter_0/n6385 ) );
  inv_x1_sg U64393 ( .A(\filter_0/reg_i_3[17] ), .X(n42288) );
  nor_x1_sg U64394 ( .A(n42289), .B(n34169), .X(\filter_0/n6381 ) );
  inv_x1_sg U64395 ( .A(\filter_0/reg_i_3[16] ), .X(n42289) );
  nor_x1_sg U64396 ( .A(n42290), .B(n29741), .X(\filter_0/n6377 ) );
  inv_x1_sg U64397 ( .A(\filter_0/reg_i_3[15] ), .X(n42290) );
  nor_x1_sg U64398 ( .A(n42291), .B(n31833), .X(\filter_0/n6373 ) );
  inv_x1_sg U64399 ( .A(\filter_0/reg_i_3[14] ), .X(n42291) );
  nor_x1_sg U64400 ( .A(n42292), .B(n31833), .X(\filter_0/n6369 ) );
  inv_x1_sg U64401 ( .A(\filter_0/reg_i_3[13] ), .X(n42292) );
  nor_x1_sg U64402 ( .A(n42293), .B(n31435), .X(\filter_0/n6365 ) );
  inv_x1_sg U64403 ( .A(\filter_0/reg_i_3[12] ), .X(n42293) );
  nor_x1_sg U64404 ( .A(n42294), .B(n31435), .X(\filter_0/n6361 ) );
  inv_x1_sg U64405 ( .A(\filter_0/reg_i_3[11] ), .X(n42294) );
  nor_x1_sg U64406 ( .A(n42296), .B(n34169), .X(\filter_0/n6353 ) );
  inv_x1_sg U64407 ( .A(\filter_0/reg_i_3[9] ), .X(n42296) );
  nor_x1_sg U64408 ( .A(n42297), .B(n31833), .X(\filter_0/n6349 ) );
  inv_x1_sg U64409 ( .A(\filter_0/reg_i_3[8] ), .X(n42297) );
  nor_x1_sg U64410 ( .A(n42298), .B(n31435), .X(\filter_0/n6345 ) );
  inv_x1_sg U64411 ( .A(\filter_0/reg_i_3[7] ), .X(n42298) );
  nor_x1_sg U64412 ( .A(n42299), .B(n30271), .X(\filter_0/n6341 ) );
  inv_x1_sg U64413 ( .A(\filter_0/reg_i_3[6] ), .X(n42299) );
  nor_x1_sg U64414 ( .A(n42300), .B(n34171), .X(\filter_0/n6337 ) );
  inv_x1_sg U64415 ( .A(\filter_0/reg_i_3[5] ), .X(n42300) );
  nor_x1_sg U64416 ( .A(n42301), .B(n31434), .X(\filter_0/n6333 ) );
  inv_x1_sg U64417 ( .A(\filter_0/reg_i_3[4] ), .X(n42301) );
  nor_x1_sg U64418 ( .A(n42302), .B(n31434), .X(\filter_0/n6329 ) );
  inv_x1_sg U64419 ( .A(\filter_0/reg_i_3[3] ), .X(n42302) );
  nor_x1_sg U64420 ( .A(n42303), .B(n31833), .X(\filter_0/n6325 ) );
  inv_x1_sg U64421 ( .A(\filter_0/reg_i_3[2] ), .X(n42303) );
  nor_x1_sg U64422 ( .A(n42304), .B(n34171), .X(\filter_0/n6321 ) );
  inv_x1_sg U64423 ( .A(\filter_0/reg_i_3[1] ), .X(n42304) );
  nor_x1_sg U64424 ( .A(n42305), .B(n30069), .X(\filter_0/n6317 ) );
  inv_x1_sg U64425 ( .A(\filter_0/reg_i_3[0] ), .X(n42305) );
  nor_x1_sg U64426 ( .A(n41946), .B(n34146), .X(\filter_0/n5637 ) );
  inv_x1_sg U64427 ( .A(\filter_0/reg_w_4[19] ), .X(n41946) );
  nor_x1_sg U64428 ( .A(n41947), .B(n31843), .X(\filter_0/n5633 ) );
  inv_x1_sg U64429 ( .A(\filter_0/reg_w_4[18] ), .X(n41947) );
  nor_x1_sg U64430 ( .A(n41948), .B(n34145), .X(\filter_0/n5629 ) );
  inv_x1_sg U64431 ( .A(\filter_0/reg_w_4[17] ), .X(n41948) );
  nor_x1_sg U64432 ( .A(n41949), .B(n31450), .X(\filter_0/n5625 ) );
  inv_x1_sg U64433 ( .A(\filter_0/reg_w_4[16] ), .X(n41949) );
  nor_x1_sg U64434 ( .A(n41950), .B(n30261), .X(\filter_0/n5621 ) );
  inv_x1_sg U64435 ( .A(\filter_0/reg_w_4[15] ), .X(n41950) );
  nor_x1_sg U64436 ( .A(n41951), .B(n30064), .X(\filter_0/n5617 ) );
  inv_x1_sg U64437 ( .A(\filter_0/reg_w_4[14] ), .X(n41951) );
  nor_x1_sg U64438 ( .A(n41952), .B(n31843), .X(\filter_0/n5613 ) );
  inv_x1_sg U64439 ( .A(\filter_0/reg_w_4[13] ), .X(n41952) );
  nor_x1_sg U64440 ( .A(n41953), .B(n31449), .X(\filter_0/n5609 ) );
  inv_x1_sg U64441 ( .A(\filter_0/reg_w_4[12] ), .X(n41953) );
  nor_x1_sg U64442 ( .A(n41954), .B(n34145), .X(\filter_0/n5605 ) );
  inv_x1_sg U64443 ( .A(\filter_0/reg_w_4[11] ), .X(n41954) );
  nor_x1_sg U64444 ( .A(n41956), .B(n34144), .X(\filter_0/n5597 ) );
  inv_x1_sg U64445 ( .A(\filter_0/reg_w_4[9] ), .X(n41956) );
  nor_x1_sg U64446 ( .A(n41957), .B(n31843), .X(\filter_0/n5593 ) );
  inv_x1_sg U64447 ( .A(\filter_0/reg_w_4[8] ), .X(n41957) );
  nor_x1_sg U64448 ( .A(n41958), .B(n34144), .X(\filter_0/n5589 ) );
  inv_x1_sg U64449 ( .A(\filter_0/reg_w_4[7] ), .X(n41958) );
  nor_x1_sg U64450 ( .A(n41959), .B(n34145), .X(\filter_0/n5585 ) );
  inv_x1_sg U64451 ( .A(\filter_0/reg_w_4[6] ), .X(n41959) );
  nor_x1_sg U64452 ( .A(n41960), .B(n31450), .X(\filter_0/n5581 ) );
  inv_x1_sg U64453 ( .A(\filter_0/reg_w_4[5] ), .X(n41960) );
  nor_x1_sg U64454 ( .A(n41961), .B(n30064), .X(\filter_0/n5577 ) );
  inv_x1_sg U64455 ( .A(\filter_0/reg_w_4[4] ), .X(n41961) );
  nor_x1_sg U64456 ( .A(n41962), .B(n34147), .X(\filter_0/n5573 ) );
  inv_x1_sg U64457 ( .A(\filter_0/reg_w_4[3] ), .X(n41962) );
  nor_x1_sg U64458 ( .A(n41963), .B(n30261), .X(\filter_0/n5569 ) );
  inv_x1_sg U64459 ( .A(\filter_0/reg_w_4[2] ), .X(n41963) );
  nor_x1_sg U64460 ( .A(n41964), .B(n31449), .X(\filter_0/n5565 ) );
  inv_x1_sg U64461 ( .A(\filter_0/reg_w_4[1] ), .X(n41964) );
  nor_x1_sg U64462 ( .A(n41965), .B(n31449), .X(\filter_0/n5561 ) );
  inv_x1_sg U64463 ( .A(\filter_0/reg_w_4[0] ), .X(n41965) );
  nor_x1_sg U64464 ( .A(n41926), .B(n34294), .X(\filter_0/n5557 ) );
  inv_x1_sg U64465 ( .A(\filter_0/reg_w_5[19] ), .X(n41926) );
  nor_x1_sg U64466 ( .A(n41927), .B(n31790), .X(\filter_0/n5553 ) );
  inv_x1_sg U64467 ( .A(\filter_0/reg_w_5[18] ), .X(n41927) );
  nor_x1_sg U64468 ( .A(n41928), .B(n31789), .X(\filter_0/n5549 ) );
  inv_x1_sg U64469 ( .A(\filter_0/reg_w_5[17] ), .X(n41928) );
  nor_x1_sg U64470 ( .A(n41929), .B(n31359), .X(\filter_0/n5545 ) );
  inv_x1_sg U64471 ( .A(\filter_0/reg_w_5[16] ), .X(n41929) );
  nor_x1_sg U64472 ( .A(n41930), .B(n31360), .X(\filter_0/n5541 ) );
  inv_x1_sg U64473 ( .A(\filter_0/reg_w_5[15] ), .X(n41930) );
  nor_x1_sg U64474 ( .A(n41931), .B(n34297), .X(\filter_0/n5537 ) );
  inv_x1_sg U64475 ( .A(\filter_0/reg_w_5[14] ), .X(n41931) );
  nor_x1_sg U64476 ( .A(n41932), .B(n31360), .X(\filter_0/n5533 ) );
  inv_x1_sg U64477 ( .A(\filter_0/reg_w_5[13] ), .X(n41932) );
  nor_x1_sg U64478 ( .A(n41933), .B(n34296), .X(\filter_0/n5529 ) );
  inv_x1_sg U64479 ( .A(\filter_0/reg_w_5[12] ), .X(n41933) );
  nor_x1_sg U64480 ( .A(n41934), .B(n31360), .X(\filter_0/n5525 ) );
  inv_x1_sg U64481 ( .A(\filter_0/reg_w_5[11] ), .X(n41934) );
  nor_x1_sg U64482 ( .A(n41936), .B(n31790), .X(\filter_0/n5517 ) );
  inv_x1_sg U64483 ( .A(\filter_0/reg_w_5[9] ), .X(n41936) );
  nor_x1_sg U64484 ( .A(n41937), .B(n34295), .X(\filter_0/n5513 ) );
  inv_x1_sg U64485 ( .A(\filter_0/reg_w_5[8] ), .X(n41937) );
  nor_x1_sg U64486 ( .A(n41938), .B(n29723), .X(\filter_0/n5509 ) );
  inv_x1_sg U64487 ( .A(\filter_0/reg_w_5[7] ), .X(n41938) );
  nor_x1_sg U64488 ( .A(n41939), .B(n30328), .X(\filter_0/n5505 ) );
  inv_x1_sg U64489 ( .A(\filter_0/reg_w_5[6] ), .X(n41939) );
  nor_x1_sg U64490 ( .A(n41940), .B(n34294), .X(\filter_0/n5501 ) );
  inv_x1_sg U64491 ( .A(\filter_0/reg_w_5[5] ), .X(n41940) );
  nor_x1_sg U64492 ( .A(n41941), .B(n34296), .X(\filter_0/n5497 ) );
  inv_x1_sg U64493 ( .A(\filter_0/reg_w_5[4] ), .X(n41941) );
  nor_x1_sg U64494 ( .A(n41942), .B(n30094), .X(\filter_0/n5493 ) );
  inv_x1_sg U64495 ( .A(\filter_0/reg_w_5[3] ), .X(n41942) );
  nor_x1_sg U64496 ( .A(n41943), .B(n29723), .X(\filter_0/n5489 ) );
  inv_x1_sg U64497 ( .A(\filter_0/reg_w_5[2] ), .X(n41943) );
  nor_x1_sg U64498 ( .A(n41944), .B(n30094), .X(\filter_0/n5485 ) );
  inv_x1_sg U64499 ( .A(\filter_0/reg_w_5[1] ), .X(n41944) );
  nor_x1_sg U64500 ( .A(n41945), .B(n30094), .X(\filter_0/n5481 ) );
  inv_x1_sg U64501 ( .A(\filter_0/reg_w_5[0] ), .X(n41945) );
  nor_x1_sg U64502 ( .A(n41906), .B(n31453), .X(\filter_0/n5477 ) );
  inv_x1_sg U64503 ( .A(\filter_0/reg_w_6[19] ), .X(n41906) );
  nor_x1_sg U64504 ( .A(n41907), .B(n34140), .X(\filter_0/n5473 ) );
  inv_x1_sg U64505 ( .A(\filter_0/reg_w_6[18] ), .X(n41907) );
  nor_x1_sg U64506 ( .A(n41908), .B(n30063), .X(\filter_0/n5469 ) );
  inv_x1_sg U64507 ( .A(\filter_0/reg_w_6[17] ), .X(n41908) );
  nor_x1_sg U64508 ( .A(n41909), .B(n30063), .X(\filter_0/n5465 ) );
  inv_x1_sg U64509 ( .A(\filter_0/reg_w_6[16] ), .X(n41909) );
  nor_x1_sg U64510 ( .A(n41910), .B(n31845), .X(\filter_0/n5461 ) );
  inv_x1_sg U64511 ( .A(\filter_0/reg_w_6[15] ), .X(n41910) );
  nor_x1_sg U64512 ( .A(n41911), .B(n34141), .X(\filter_0/n5457 ) );
  inv_x1_sg U64513 ( .A(\filter_0/reg_w_6[14] ), .X(n41911) );
  nor_x1_sg U64514 ( .A(n41912), .B(n31845), .X(\filter_0/n5453 ) );
  inv_x1_sg U64515 ( .A(\filter_0/reg_w_6[13] ), .X(n41912) );
  nor_x1_sg U64516 ( .A(n41913), .B(n31452), .X(\filter_0/n5449 ) );
  inv_x1_sg U64517 ( .A(\filter_0/reg_w_6[12] ), .X(n41913) );
  nor_x1_sg U64518 ( .A(n41914), .B(n34140), .X(\filter_0/n5445 ) );
  inv_x1_sg U64519 ( .A(\filter_0/reg_w_6[11] ), .X(n41914) );
  nor_x1_sg U64520 ( .A(n41916), .B(n34139), .X(\filter_0/n5437 ) );
  inv_x1_sg U64521 ( .A(\filter_0/reg_w_6[9] ), .X(n41916) );
  nor_x1_sg U64522 ( .A(n41917), .B(n30063), .X(\filter_0/n5433 ) );
  inv_x1_sg U64523 ( .A(\filter_0/reg_w_6[8] ), .X(n41917) );
  nor_x1_sg U64524 ( .A(n41918), .B(n31452), .X(\filter_0/n5429 ) );
  inv_x1_sg U64525 ( .A(\filter_0/reg_w_6[7] ), .X(n41918) );
  nor_x1_sg U64526 ( .A(n41919), .B(n31452), .X(\filter_0/n5425 ) );
  inv_x1_sg U64527 ( .A(\filter_0/reg_w_6[6] ), .X(n41919) );
  nor_x1_sg U64528 ( .A(n41920), .B(n34140), .X(\filter_0/n5421 ) );
  inv_x1_sg U64529 ( .A(\filter_0/reg_w_6[5] ), .X(n41920) );
  nor_x1_sg U64530 ( .A(n41921), .B(n29747), .X(\filter_0/n5417 ) );
  inv_x1_sg U64531 ( .A(\filter_0/reg_w_6[4] ), .X(n41921) );
  nor_x1_sg U64532 ( .A(n41922), .B(n31844), .X(\filter_0/n5413 ) );
  inv_x1_sg U64533 ( .A(\filter_0/reg_w_6[3] ), .X(n41922) );
  nor_x1_sg U64534 ( .A(n41923), .B(n31452), .X(\filter_0/n5409 ) );
  inv_x1_sg U64535 ( .A(\filter_0/reg_w_6[2] ), .X(n41923) );
  nor_x1_sg U64536 ( .A(n41924), .B(n34141), .X(\filter_0/n5405 ) );
  inv_x1_sg U64537 ( .A(\filter_0/reg_w_6[1] ), .X(n41924) );
  nor_x1_sg U64538 ( .A(n41925), .B(n34139), .X(\filter_0/n5401 ) );
  inv_x1_sg U64539 ( .A(\filter_0/reg_w_6[0] ), .X(n41925) );
  nor_x1_sg U64540 ( .A(n41886), .B(n34137), .X(\filter_0/n5397 ) );
  inv_x1_sg U64541 ( .A(\filter_0/reg_w_7[19] ), .X(n41886) );
  nor_x1_sg U64542 ( .A(n41887), .B(n30062), .X(\filter_0/n5393 ) );
  inv_x1_sg U64543 ( .A(\filter_0/reg_w_7[18] ), .X(n41887) );
  nor_x1_sg U64544 ( .A(n41888), .B(n30257), .X(\filter_0/n5389 ) );
  inv_x1_sg U64545 ( .A(\filter_0/reg_w_7[17] ), .X(n41888) );
  nor_x1_sg U64546 ( .A(n41889), .B(n34137), .X(\filter_0/n5385 ) );
  inv_x1_sg U64547 ( .A(\filter_0/reg_w_7[16] ), .X(n41889) );
  nor_x1_sg U64548 ( .A(n41890), .B(n31847), .X(\filter_0/n5381 ) );
  inv_x1_sg U64549 ( .A(\filter_0/reg_w_7[15] ), .X(n41890) );
  nor_x1_sg U64550 ( .A(n41891), .B(n34136), .X(\filter_0/n5377 ) );
  inv_x1_sg U64551 ( .A(\filter_0/reg_w_7[14] ), .X(n41891) );
  nor_x1_sg U64552 ( .A(n41892), .B(n31847), .X(\filter_0/n5373 ) );
  inv_x1_sg U64553 ( .A(\filter_0/reg_w_7[13] ), .X(n41892) );
  nor_x1_sg U64554 ( .A(n41893), .B(n31455), .X(\filter_0/n5369 ) );
  inv_x1_sg U64555 ( .A(\filter_0/reg_w_7[12] ), .X(n41893) );
  nor_x1_sg U64556 ( .A(n41894), .B(n34135), .X(\filter_0/n5365 ) );
  inv_x1_sg U64557 ( .A(\filter_0/reg_w_7[11] ), .X(n41894) );
  nor_x1_sg U64558 ( .A(n41896), .B(n34134), .X(\filter_0/n5357 ) );
  inv_x1_sg U64559 ( .A(\filter_0/reg_w_7[9] ), .X(n41896) );
  nor_x1_sg U64560 ( .A(n41897), .B(n34135), .X(\filter_0/n5353 ) );
  inv_x1_sg U64561 ( .A(\filter_0/reg_w_7[8] ), .X(n41897) );
  nor_x1_sg U64562 ( .A(n41898), .B(n29748), .X(\filter_0/n5349 ) );
  inv_x1_sg U64563 ( .A(\filter_0/reg_w_7[7] ), .X(n41898) );
  nor_x1_sg U64564 ( .A(n41899), .B(n30062), .X(\filter_0/n5345 ) );
  inv_x1_sg U64565 ( .A(\filter_0/reg_w_7[6] ), .X(n41899) );
  nor_x1_sg U64566 ( .A(n41900), .B(n29748), .X(\filter_0/n5341 ) );
  inv_x1_sg U64567 ( .A(\filter_0/reg_w_7[5] ), .X(n41900) );
  nor_x1_sg U64568 ( .A(n41901), .B(n34136), .X(\filter_0/n5337 ) );
  inv_x1_sg U64569 ( .A(\filter_0/reg_w_7[4] ), .X(n41901) );
  nor_x1_sg U64570 ( .A(n41902), .B(n31846), .X(\filter_0/n5333 ) );
  inv_x1_sg U64571 ( .A(\filter_0/reg_w_7[3] ), .X(n41902) );
  nor_x1_sg U64572 ( .A(n41903), .B(n31846), .X(\filter_0/n5329 ) );
  inv_x1_sg U64573 ( .A(\filter_0/reg_w_7[2] ), .X(n41903) );
  nor_x1_sg U64574 ( .A(n41904), .B(n34136), .X(\filter_0/n5325 ) );
  inv_x1_sg U64575 ( .A(\filter_0/reg_w_7[1] ), .X(n41904) );
  nor_x1_sg U64576 ( .A(n41905), .B(n34134), .X(\filter_0/n5321 ) );
  inv_x1_sg U64577 ( .A(\filter_0/reg_w_7[0] ), .X(n41905) );
  nor_x1_sg U64578 ( .A(n42026), .B(n34165), .X(\filter_0/n5317 ) );
  inv_x1_sg U64579 ( .A(\filter_0/reg_w_0[19] ), .X(n42026) );
  nor_x1_sg U64580 ( .A(n42027), .B(n30269), .X(\filter_0/n5313 ) );
  inv_x1_sg U64581 ( .A(\filter_0/reg_w_0[18] ), .X(n42027) );
  nor_x1_sg U64582 ( .A(n42028), .B(n34166), .X(\filter_0/n5309 ) );
  inv_x1_sg U64583 ( .A(\filter_0/reg_w_0[17] ), .X(n42028) );
  nor_x1_sg U64584 ( .A(n42029), .B(n31834), .X(\filter_0/n5305 ) );
  inv_x1_sg U64585 ( .A(\filter_0/reg_w_0[16] ), .X(n42029) );
  nor_x1_sg U64586 ( .A(n42030), .B(n34167), .X(\filter_0/n5301 ) );
  inv_x1_sg U64587 ( .A(\filter_0/reg_w_0[15] ), .X(n42030) );
  nor_x1_sg U64588 ( .A(n42031), .B(n31438), .X(\filter_0/n5297 ) );
  inv_x1_sg U64589 ( .A(\filter_0/reg_w_0[14] ), .X(n42031) );
  nor_x1_sg U64590 ( .A(n42032), .B(n34167), .X(\filter_0/n5293 ) );
  inv_x1_sg U64591 ( .A(\filter_0/reg_w_0[13] ), .X(n42032) );
  nor_x1_sg U64592 ( .A(n42033), .B(n30269), .X(\filter_0/n5289 ) );
  inv_x1_sg U64593 ( .A(\filter_0/reg_w_0[12] ), .X(n42033) );
  nor_x1_sg U64594 ( .A(n42034), .B(n30068), .X(\filter_0/n5285 ) );
  inv_x1_sg U64595 ( .A(\filter_0/reg_w_0[11] ), .X(n42034) );
  nor_x1_sg U64596 ( .A(n42036), .B(n34167), .X(\filter_0/n5277 ) );
  inv_x1_sg U64597 ( .A(\filter_0/reg_w_0[9] ), .X(n42036) );
  nor_x1_sg U64598 ( .A(n42037), .B(n31835), .X(\filter_0/n5273 ) );
  inv_x1_sg U64599 ( .A(\filter_0/reg_w_0[8] ), .X(n42037) );
  nor_x1_sg U64600 ( .A(n42038), .B(n31437), .X(\filter_0/n5269 ) );
  inv_x1_sg U64601 ( .A(\filter_0/reg_w_0[7] ), .X(n42038) );
  nor_x1_sg U64602 ( .A(n42039), .B(n31834), .X(\filter_0/n5265 ) );
  inv_x1_sg U64603 ( .A(\filter_0/reg_w_0[6] ), .X(n42039) );
  nor_x1_sg U64604 ( .A(n42040), .B(n31835), .X(\filter_0/n5261 ) );
  inv_x1_sg U64605 ( .A(\filter_0/reg_w_0[5] ), .X(n42040) );
  nor_x1_sg U64606 ( .A(n42041), .B(n34164), .X(\filter_0/n5257 ) );
  inv_x1_sg U64607 ( .A(\filter_0/reg_w_0[4] ), .X(n42041) );
  nor_x1_sg U64608 ( .A(n42042), .B(n31437), .X(\filter_0/n5253 ) );
  inv_x1_sg U64609 ( .A(\filter_0/reg_w_0[3] ), .X(n42042) );
  nor_x1_sg U64610 ( .A(n42043), .B(n31835), .X(\filter_0/n5249 ) );
  inv_x1_sg U64611 ( .A(\filter_0/reg_w_0[2] ), .X(n42043) );
  nor_x1_sg U64612 ( .A(n42044), .B(n30068), .X(\filter_0/n5245 ) );
  inv_x1_sg U64613 ( .A(\filter_0/reg_w_0[1] ), .X(n42044) );
  nor_x1_sg U64614 ( .A(n42045), .B(n34165), .X(\filter_0/n5241 ) );
  inv_x1_sg U64615 ( .A(\filter_0/reg_w_0[0] ), .X(n42045) );
  nor_x1_sg U64616 ( .A(n42006), .B(n29724), .X(\filter_0/n5237 ) );
  inv_x1_sg U64617 ( .A(\filter_0/reg_w_1[19] ), .X(n42006) );
  nor_x1_sg U64618 ( .A(n42007), .B(n31791), .X(\filter_0/n5233 ) );
  inv_x1_sg U64619 ( .A(\filter_0/reg_w_1[18] ), .X(n42007) );
  nor_x1_sg U64620 ( .A(n42008), .B(n34292), .X(\filter_0/n5229 ) );
  inv_x1_sg U64621 ( .A(\filter_0/reg_w_1[17] ), .X(n42008) );
  nor_x1_sg U64622 ( .A(n42009), .B(n30093), .X(\filter_0/n5225 ) );
  inv_x1_sg U64623 ( .A(\filter_0/reg_w_1[16] ), .X(n42009) );
  nor_x1_sg U64624 ( .A(n42010), .B(n30093), .X(\filter_0/n5221 ) );
  inv_x1_sg U64625 ( .A(\filter_0/reg_w_1[15] ), .X(n42010) );
  nor_x1_sg U64626 ( .A(n42011), .B(n29724), .X(\filter_0/n5217 ) );
  inv_x1_sg U64627 ( .A(\filter_0/reg_w_1[14] ), .X(n42011) );
  nor_x1_sg U64628 ( .A(n42012), .B(n31792), .X(\filter_0/n5213 ) );
  inv_x1_sg U64629 ( .A(\filter_0/reg_w_1[13] ), .X(n42012) );
  nor_x1_sg U64630 ( .A(n42013), .B(n31791), .X(\filter_0/n5209 ) );
  inv_x1_sg U64631 ( .A(\filter_0/reg_w_1[12] ), .X(n42013) );
  nor_x1_sg U64632 ( .A(n42014), .B(n30326), .X(\filter_0/n5205 ) );
  inv_x1_sg U64633 ( .A(\filter_0/reg_w_1[11] ), .X(n42014) );
  nor_x1_sg U64634 ( .A(n42016), .B(n31791), .X(\filter_0/n5197 ) );
  inv_x1_sg U64635 ( .A(\filter_0/reg_w_1[9] ), .X(n42016) );
  nor_x1_sg U64636 ( .A(n42017), .B(n34292), .X(\filter_0/n5193 ) );
  inv_x1_sg U64637 ( .A(\filter_0/reg_w_1[8] ), .X(n42017) );
  nor_x1_sg U64638 ( .A(n42018), .B(n34290), .X(\filter_0/n5189 ) );
  inv_x1_sg U64639 ( .A(\filter_0/reg_w_1[7] ), .X(n42018) );
  nor_x1_sg U64640 ( .A(n42019), .B(n34291), .X(\filter_0/n5185 ) );
  inv_x1_sg U64641 ( .A(\filter_0/reg_w_1[6] ), .X(n42019) );
  nor_x1_sg U64642 ( .A(n42020), .B(n34292), .X(\filter_0/n5181 ) );
  inv_x1_sg U64643 ( .A(\filter_0/reg_w_1[5] ), .X(n42020) );
  nor_x1_sg U64644 ( .A(n42021), .B(n31363), .X(\filter_0/n5177 ) );
  inv_x1_sg U64645 ( .A(\filter_0/reg_w_1[4] ), .X(n42021) );
  nor_x1_sg U64646 ( .A(n42022), .B(n31363), .X(\filter_0/n5173 ) );
  inv_x1_sg U64647 ( .A(\filter_0/reg_w_1[3] ), .X(n42022) );
  nor_x1_sg U64648 ( .A(n42023), .B(n34289), .X(\filter_0/n5169 ) );
  inv_x1_sg U64649 ( .A(\filter_0/reg_w_1[2] ), .X(n42023) );
  nor_x1_sg U64650 ( .A(n42024), .B(n31791), .X(\filter_0/n5165 ) );
  inv_x1_sg U64651 ( .A(\filter_0/reg_w_1[1] ), .X(n42024) );
  nor_x1_sg U64652 ( .A(n42025), .B(n30093), .X(\filter_0/n5161 ) );
  inv_x1_sg U64653 ( .A(\filter_0/reg_w_1[0] ), .X(n42025) );
  nor_x1_sg U64654 ( .A(n41986), .B(n34342), .X(\filter_0/n5157 ) );
  inv_x1_sg U64655 ( .A(\filter_0/reg_w_2[19] ), .X(n41986) );
  nor_x1_sg U64656 ( .A(n41987), .B(n30103), .X(\filter_0/n5153 ) );
  inv_x1_sg U64657 ( .A(\filter_0/reg_w_2[18] ), .X(n41987) );
  nor_x1_sg U64658 ( .A(n41988), .B(n30103), .X(\filter_0/n5149 ) );
  inv_x1_sg U64659 ( .A(\filter_0/reg_w_2[17] ), .X(n41988) );
  nor_x1_sg U64660 ( .A(n41989), .B(n34339), .X(\filter_0/n5145 ) );
  inv_x1_sg U64661 ( .A(\filter_0/reg_w_2[16] ), .X(n41989) );
  nor_x1_sg U64662 ( .A(n41990), .B(n29714), .X(\filter_0/n5141 ) );
  inv_x1_sg U64663 ( .A(\filter_0/reg_w_2[15] ), .X(n41990) );
  nor_x1_sg U64664 ( .A(n41991), .B(n31772), .X(\filter_0/n5137 ) );
  inv_x1_sg U64665 ( .A(\filter_0/reg_w_2[14] ), .X(n41991) );
  nor_x1_sg U64666 ( .A(n41992), .B(n31772), .X(\filter_0/n5133 ) );
  inv_x1_sg U64667 ( .A(\filter_0/reg_w_2[13] ), .X(n41992) );
  nor_x1_sg U64668 ( .A(n41993), .B(n31333), .X(\filter_0/n5129 ) );
  inv_x1_sg U64669 ( .A(\filter_0/reg_w_2[12] ), .X(n41993) );
  nor_x1_sg U64670 ( .A(n41994), .B(n31333), .X(\filter_0/n5125 ) );
  inv_x1_sg U64671 ( .A(\filter_0/reg_w_2[11] ), .X(n41994) );
  nor_x1_sg U64672 ( .A(n41996), .B(n34339), .X(\filter_0/n5117 ) );
  inv_x1_sg U64673 ( .A(\filter_0/reg_w_2[9] ), .X(n41996) );
  nor_x1_sg U64674 ( .A(n41997), .B(n31772), .X(\filter_0/n5113 ) );
  inv_x1_sg U64675 ( .A(\filter_0/reg_w_2[8] ), .X(n41997) );
  nor_x1_sg U64676 ( .A(n41998), .B(n31333), .X(\filter_0/n5109 ) );
  inv_x1_sg U64677 ( .A(\filter_0/reg_w_2[7] ), .X(n41998) );
  nor_x1_sg U64678 ( .A(n41999), .B(n30346), .X(\filter_0/n5105 ) );
  inv_x1_sg U64679 ( .A(\filter_0/reg_w_2[6] ), .X(n41999) );
  nor_x1_sg U64680 ( .A(n42000), .B(n34341), .X(\filter_0/n5101 ) );
  inv_x1_sg U64681 ( .A(\filter_0/reg_w_2[5] ), .X(n42000) );
  nor_x1_sg U64682 ( .A(n42001), .B(n31332), .X(\filter_0/n5097 ) );
  inv_x1_sg U64683 ( .A(\filter_0/reg_w_2[4] ), .X(n42001) );
  nor_x1_sg U64684 ( .A(n42002), .B(n31332), .X(\filter_0/n5093 ) );
  inv_x1_sg U64685 ( .A(\filter_0/reg_w_2[3] ), .X(n42002) );
  nor_x1_sg U64686 ( .A(n42003), .B(n31772), .X(\filter_0/n5089 ) );
  inv_x1_sg U64687 ( .A(\filter_0/reg_w_2[2] ), .X(n42003) );
  nor_x1_sg U64688 ( .A(n42004), .B(n34341), .X(\filter_0/n5085 ) );
  inv_x1_sg U64689 ( .A(\filter_0/reg_w_2[1] ), .X(n42004) );
  nor_x1_sg U64690 ( .A(n42005), .B(n30103), .X(\filter_0/n5081 ) );
  inv_x1_sg U64691 ( .A(\filter_0/reg_w_2[0] ), .X(n42005) );
  nor_x1_sg U64692 ( .A(n41966), .B(n31837), .X(\filter_0/n5077 ) );
  inv_x1_sg U64693 ( .A(\filter_0/reg_w_3[19] ), .X(n41966) );
  nor_x1_sg U64694 ( .A(n41967), .B(n34162), .X(\filter_0/n5073 ) );
  inv_x1_sg U64695 ( .A(\filter_0/reg_w_3[18] ), .X(n41967) );
  nor_x1_sg U64696 ( .A(n41968), .B(n34160), .X(\filter_0/n5069 ) );
  inv_x1_sg U64697 ( .A(\filter_0/reg_w_3[17] ), .X(n41968) );
  nor_x1_sg U64698 ( .A(n41969), .B(n31836), .X(\filter_0/n5065 ) );
  inv_x1_sg U64699 ( .A(\filter_0/reg_w_3[16] ), .X(n41969) );
  nor_x1_sg U64700 ( .A(n41970), .B(n30067), .X(\filter_0/n5061 ) );
  inv_x1_sg U64701 ( .A(\filter_0/reg_w_3[15] ), .X(n41970) );
  nor_x1_sg U64702 ( .A(n41971), .B(n31441), .X(\filter_0/n5057 ) );
  inv_x1_sg U64703 ( .A(\filter_0/reg_w_3[14] ), .X(n41971) );
  nor_x1_sg U64704 ( .A(n41972), .B(n31440), .X(\filter_0/n5053 ) );
  inv_x1_sg U64705 ( .A(\filter_0/reg_w_3[13] ), .X(n41972) );
  nor_x1_sg U64706 ( .A(n41973), .B(n31441), .X(\filter_0/n5049 ) );
  inv_x1_sg U64707 ( .A(\filter_0/reg_w_3[12] ), .X(n41973) );
  nor_x1_sg U64708 ( .A(n41974), .B(n29743), .X(\filter_0/n5045 ) );
  inv_x1_sg U64709 ( .A(\filter_0/reg_w_3[11] ), .X(n41974) );
  nor_x1_sg U64710 ( .A(n41976), .B(n30067), .X(\filter_0/n5037 ) );
  inv_x1_sg U64711 ( .A(\filter_0/reg_w_3[9] ), .X(n41976) );
  nor_x1_sg U64712 ( .A(n41977), .B(n30267), .X(\filter_0/n5033 ) );
  inv_x1_sg U64713 ( .A(\filter_0/reg_w_3[8] ), .X(n41977) );
  nor_x1_sg U64714 ( .A(n41978), .B(n31837), .X(\filter_0/n5029 ) );
  inv_x1_sg U64715 ( .A(\filter_0/reg_w_3[7] ), .X(n41978) );
  nor_x1_sg U64716 ( .A(n41979), .B(n31836), .X(\filter_0/n5025 ) );
  inv_x1_sg U64717 ( .A(\filter_0/reg_w_3[6] ), .X(n41979) );
  nor_x1_sg U64718 ( .A(n41980), .B(n31836), .X(\filter_0/n5021 ) );
  inv_x1_sg U64719 ( .A(\filter_0/reg_w_3[5] ), .X(n41980) );
  nor_x1_sg U64720 ( .A(n41981), .B(n34160), .X(\filter_0/n5017 ) );
  inv_x1_sg U64721 ( .A(\filter_0/reg_w_3[4] ), .X(n41981) );
  nor_x1_sg U64722 ( .A(n41982), .B(n34160), .X(\filter_0/n5013 ) );
  inv_x1_sg U64723 ( .A(\filter_0/reg_w_3[3] ), .X(n41982) );
  nor_x1_sg U64724 ( .A(n41983), .B(n34159), .X(\filter_0/n5009 ) );
  inv_x1_sg U64725 ( .A(\filter_0/reg_w_3[2] ), .X(n41983) );
  nor_x1_sg U64726 ( .A(n41984), .B(n34160), .X(\filter_0/n5005 ) );
  inv_x1_sg U64727 ( .A(\filter_0/reg_w_3[1] ), .X(n41984) );
  nor_x1_sg U64728 ( .A(n41985), .B(n30267), .X(\filter_0/n5001 ) );
  inv_x1_sg U64729 ( .A(\filter_0/reg_w_3[0] ), .X(n41985) );
  nor_x1_sg U64730 ( .A(n42175), .B(n34202), .X(\filter_0/n7477 ) );
  inv_x1_sg U64731 ( .A(\filter_0/reg_i_9[10] ), .X(n42175) );
  nor_x1_sg U64732 ( .A(n42155), .B(n30281), .X(\filter_0/n7397 ) );
  inv_x1_sg U64733 ( .A(\filter_0/reg_i_10[10] ), .X(n42155) );
  nor_x1_sg U64734 ( .A(n42135), .B(n34190), .X(\filter_0/n7317 ) );
  inv_x1_sg U64735 ( .A(\filter_0/reg_i_11[10] ), .X(n42135) );
  nor_x1_sg U64736 ( .A(n41855), .B(n31827), .X(\filter_0/n6161 ) );
  inv_x1_sg U64737 ( .A(\filter_0/reg_w_9[10] ), .X(n41855) );
  nor_x1_sg U64738 ( .A(n41835), .B(n30060), .X(\filter_0/n6081 ) );
  inv_x1_sg U64739 ( .A(\filter_0/reg_w_10[10] ), .X(n41835) );
  nor_x1_sg U64740 ( .A(n41815), .B(n31429), .X(\filter_0/n6001 ) );
  inv_x1_sg U64741 ( .A(\filter_0/reg_w_11[10] ), .X(n41815) );
  nand_x1_sg U64742 ( .A(n41140), .B(n33878), .X(n12458) );
  nand_x1_sg U64743 ( .A(n30949), .B(n35255), .X(n12459) );
  nand_x1_sg U64744 ( .A(n33728), .B(n11853), .X(n12146) );
  nand_x1_sg U64745 ( .A(n30410), .B(n33428), .X(n12147) );
  nand_x1_sg U64746 ( .A(n33729), .B(n11857), .X(n12168) );
  nand_x1_sg U64747 ( .A(n30414), .B(n33425), .X(n12169) );
  nand_x1_sg U64748 ( .A(n33728), .B(n11883), .X(n12311) );
  nand_x1_sg U64749 ( .A(n30440), .B(n29969), .X(n12312) );
  nand_x1_sg U64750 ( .A(n33731), .B(n11885), .X(n12322) );
  nand_x1_sg U64751 ( .A(n30442), .B(n33426), .X(n12323) );
  nand_x1_sg U64752 ( .A(n30940), .B(n12448), .X(n12446) );
  nand_x1_sg U64753 ( .A(\shifter_0/reg_i_7[2] ), .B(n30950), .X(n12447) );
  nand_x1_sg U64754 ( .A(n33875), .B(n12510), .X(n12508) );
  nand_x1_sg U64755 ( .A(\shifter_0/reg_i_7[17] ), .B(n33862), .X(n12509) );
  nand_x1_sg U64756 ( .A(n30941), .B(n12515), .X(n12513) );
  nand_x1_sg U64757 ( .A(\shifter_0/reg_i_7[18] ), .B(n33863), .X(n12514) );
  nand_x1_sg U64758 ( .A(n33712), .B(n11800), .X(n11893) );
  nand_x1_sg U64759 ( .A(n30468), .B(n33421), .X(n11894) );
  nand_x1_sg U64760 ( .A(n33711), .B(n11803), .X(n11907) );
  nand_x1_sg U64761 ( .A(n30470), .B(n33421), .X(n11908) );
  nand_x1_sg U64762 ( .A(n30999), .B(n11805), .X(n11918) );
  nand_x1_sg U64763 ( .A(n30472), .B(n33420), .X(n11919) );
  nand_x1_sg U64764 ( .A(n33713), .B(n11807), .X(n11929) );
  nand_x1_sg U64765 ( .A(n30474), .B(n33421), .X(n11930) );
  nand_x1_sg U64766 ( .A(n33712), .B(n11809), .X(n11940) );
  nand_x1_sg U64767 ( .A(n30476), .B(n33423), .X(n11941) );
  nand_x1_sg U64768 ( .A(n33714), .B(n11811), .X(n11951) );
  nand_x1_sg U64769 ( .A(n30478), .B(n33422), .X(n11952) );
  nand_x1_sg U64770 ( .A(n33711), .B(n11813), .X(n11962) );
  nand_x1_sg U64771 ( .A(n30480), .B(n33420), .X(n11963) );
  nand_x1_sg U64772 ( .A(n33713), .B(n11815), .X(n11973) );
  nand_x1_sg U64773 ( .A(n30482), .B(n29967), .X(n11974) );
  nand_x1_sg U64774 ( .A(n33712), .B(n11817), .X(n11984) );
  nand_x1_sg U64775 ( .A(n30484), .B(n33423), .X(n11985) );
  nand_x1_sg U64776 ( .A(n33711), .B(n11819), .X(n11995) );
  nand_x1_sg U64777 ( .A(n30486), .B(n33420), .X(n11996) );
  nand_x1_sg U64778 ( .A(n33712), .B(n11821), .X(n12006) );
  nand_x1_sg U64779 ( .A(n30488), .B(n33422), .X(n12007) );
  nand_x1_sg U64780 ( .A(n30999), .B(n11823), .X(n12017) );
  nand_x1_sg U64781 ( .A(n30490), .B(n33420), .X(n12018) );
  nand_x1_sg U64782 ( .A(n33713), .B(n11825), .X(n12028) );
  nand_x1_sg U64783 ( .A(n30492), .B(n29967), .X(n12029) );
  nand_x1_sg U64784 ( .A(n33714), .B(n11827), .X(n12039) );
  nand_x1_sg U64785 ( .A(n30494), .B(n33421), .X(n12040) );
  nand_x1_sg U64786 ( .A(n33813), .B(n11829), .X(n12050) );
  nand_x1_sg U64787 ( .A(n30496), .B(n29967), .X(n12051) );
  nand_x1_sg U64788 ( .A(n30999), .B(n11831), .X(n12061) );
  nand_x1_sg U64789 ( .A(n30498), .B(n29967), .X(n12062) );
  nand_x1_sg U64790 ( .A(n30999), .B(n11833), .X(n12072) );
  nand_x1_sg U64791 ( .A(n30500), .B(n33423), .X(n12073) );
  nand_x1_sg U64792 ( .A(n33714), .B(n11835), .X(n12083) );
  nand_x1_sg U64793 ( .A(n30502), .B(n33422), .X(n12084) );
  nand_x1_sg U64794 ( .A(n33714), .B(n11837), .X(n12094) );
  nand_x1_sg U64795 ( .A(n30504), .B(n33423), .X(n12095) );
  nand_x1_sg U64796 ( .A(n33713), .B(n11839), .X(n12105) );
  nand_x1_sg U64797 ( .A(n30506), .B(n33422), .X(n12106) );
  nand_x1_sg U64798 ( .A(n33731), .B(n11848), .X(n12121) );
  nand_x1_sg U64799 ( .A(n30406), .B(n33425), .X(n12122) );
  nand_x1_sg U64800 ( .A(n33730), .B(n11851), .X(n12135) );
  nand_x1_sg U64801 ( .A(n30408), .B(n33425), .X(n12136) );
  nand_x1_sg U64802 ( .A(n30995), .B(n11855), .X(n12157) );
  nand_x1_sg U64803 ( .A(n30412), .B(n33426), .X(n12158) );
  nand_x1_sg U64804 ( .A(n30995), .B(n11859), .X(n12179) );
  nand_x1_sg U64805 ( .A(n30416), .B(n33427), .X(n12180) );
  nand_x1_sg U64806 ( .A(n33730), .B(n11861), .X(n12190) );
  nand_x1_sg U64807 ( .A(n30418), .B(n33426), .X(n12191) );
  nand_x1_sg U64808 ( .A(n33731), .B(n11863), .X(n12201) );
  nand_x1_sg U64809 ( .A(n30420), .B(n33427), .X(n12202) );
  nand_x1_sg U64810 ( .A(n33730), .B(n11865), .X(n12212) );
  nand_x1_sg U64811 ( .A(n30422), .B(n33425), .X(n12213) );
  nand_x1_sg U64812 ( .A(n33729), .B(n11867), .X(n12223) );
  nand_x1_sg U64813 ( .A(n30424), .B(n29969), .X(n12224) );
  nand_x1_sg U64814 ( .A(n33731), .B(n11869), .X(n12234) );
  nand_x1_sg U64815 ( .A(n30426), .B(n33428), .X(n12235) );
  nand_x1_sg U64816 ( .A(n33730), .B(n11871), .X(n12245) );
  nand_x1_sg U64817 ( .A(n30428), .B(n29969), .X(n12246) );
  nand_x1_sg U64818 ( .A(n33803), .B(n11873), .X(n12256) );
  nand_x1_sg U64819 ( .A(n30430), .B(n29969), .X(n12257) );
  nand_x1_sg U64820 ( .A(n33728), .B(n11875), .X(n12267) );
  nand_x1_sg U64821 ( .A(n30432), .B(n33426), .X(n12268) );
  nand_x1_sg U64822 ( .A(n33729), .B(n11877), .X(n12278) );
  nand_x1_sg U64823 ( .A(n30434), .B(n33427), .X(n12279) );
  nand_x1_sg U64824 ( .A(n33729), .B(n11879), .X(n12289) );
  nand_x1_sg U64825 ( .A(n30436), .B(n33428), .X(n12290) );
  nand_x1_sg U64826 ( .A(n30995), .B(n11881), .X(n12300) );
  nand_x1_sg U64827 ( .A(n30438), .B(n33428), .X(n12301) );
  nand_x1_sg U64828 ( .A(n30995), .B(n11887), .X(n12333) );
  nand_x1_sg U64829 ( .A(n30444), .B(n33427), .X(n12334) );
  nand_x1_sg U64830 ( .A(n30551), .B(n33748), .X(n12347) );
  nand_x1_sg U64831 ( .A(n31161), .B(n33281), .X(n12348) );
  nand_x1_sg U64832 ( .A(n30566), .B(n30991), .X(n12354) );
  nand_x1_sg U64833 ( .A(n31163), .B(n33282), .X(n12355) );
  nand_x1_sg U64834 ( .A(n30552), .B(n33746), .X(n12358) );
  nand_x1_sg U64835 ( .A(n31165), .B(n29911), .X(n12359) );
  nand_x1_sg U64836 ( .A(n30571), .B(n33745), .X(n12362) );
  nand_x1_sg U64837 ( .A(n31167), .B(n33280), .X(n12363) );
  nand_x1_sg U64838 ( .A(n30559), .B(n33747), .X(n12366) );
  nand_x1_sg U64839 ( .A(n31169), .B(n33283), .X(n12367) );
  nand_x1_sg U64840 ( .A(n30546), .B(n33747), .X(n12370) );
  nand_x1_sg U64841 ( .A(n31171), .B(n33280), .X(n12371) );
  nand_x1_sg U64842 ( .A(n30572), .B(n33748), .X(n12374) );
  nand_x1_sg U64843 ( .A(n31173), .B(n33283), .X(n12375) );
  nand_x1_sg U64844 ( .A(n30547), .B(n30991), .X(n12378) );
  nand_x1_sg U64845 ( .A(n31175), .B(n33282), .X(n12379) );
  nand_x1_sg U64846 ( .A(n30553), .B(n30991), .X(n12382) );
  nand_x1_sg U64847 ( .A(n31177), .B(n29911), .X(n12383) );
  nand_x1_sg U64848 ( .A(n30548), .B(n33746), .X(n12386) );
  nand_x1_sg U64849 ( .A(n31179), .B(n29911), .X(n12387) );
  nand_x1_sg U64850 ( .A(n30561), .B(n33747), .X(n12390) );
  nand_x1_sg U64851 ( .A(n31181), .B(n33281), .X(n12391) );
  nand_x1_sg U64852 ( .A(n30549), .B(n33747), .X(n12394) );
  nand_x1_sg U64853 ( .A(n31183), .B(n33280), .X(n12395) );
  nand_x1_sg U64854 ( .A(n30554), .B(n33748), .X(n12398) );
  nand_x1_sg U64855 ( .A(n31185), .B(n33282), .X(n12399) );
  nand_x1_sg U64856 ( .A(n30550), .B(n33808), .X(n12402) );
  nand_x1_sg U64857 ( .A(n31187), .B(n33280), .X(n12403) );
  nand_x1_sg U64858 ( .A(n30555), .B(n33745), .X(n12406) );
  nand_x1_sg U64859 ( .A(n31189), .B(n33283), .X(n12407) );
  nand_x1_sg U64860 ( .A(n30556), .B(n33746), .X(n12410) );
  nand_x1_sg U64861 ( .A(n31191), .B(n33283), .X(n12411) );
  nand_x1_sg U64862 ( .A(n30562), .B(n30991), .X(n12414) );
  nand_x1_sg U64863 ( .A(n31193), .B(n33281), .X(n12415) );
  nand_x1_sg U64864 ( .A(n30557), .B(n33746), .X(n12418) );
  nand_x1_sg U64865 ( .A(n31195), .B(n33282), .X(n12419) );
  nand_x1_sg U64866 ( .A(n30558), .B(n33745), .X(n12422) );
  nand_x1_sg U64867 ( .A(n31197), .B(n33281), .X(n12423) );
  nand_x1_sg U64868 ( .A(n30560), .B(n33748), .X(n12426) );
  nand_x1_sg U64869 ( .A(n31199), .B(n29911), .X(n12427) );
  nand_x1_sg U64870 ( .A(n30569), .B(n32909), .X(n12435) );
  nand_x1_sg U64871 ( .A(n31126), .B(n30949), .X(n12436) );
  nand_x1_sg U64872 ( .A(n30565), .B(n29775), .X(n12442) );
  nand_x1_sg U64873 ( .A(n31128), .B(n33860), .X(n12443) );
  nand_x1_sg U64874 ( .A(n30583), .B(n32907), .X(n12451) );
  nand_x1_sg U64875 ( .A(n31130), .B(n33862), .X(n12452) );
  nand_x1_sg U64876 ( .A(n30582), .B(n32909), .X(n12460) );
  nand_x1_sg U64877 ( .A(n31133), .B(n33862), .X(n12461) );
  nand_x1_sg U64878 ( .A(n30581), .B(n32908), .X(n12464) );
  nand_x1_sg U64879 ( .A(n31135), .B(n33861), .X(n12465) );
  nand_x1_sg U64880 ( .A(n30567), .B(n32907), .X(n12468) );
  nand_x1_sg U64881 ( .A(n31137), .B(n33861), .X(n12469) );
  nand_x1_sg U64882 ( .A(n30580), .B(n32906), .X(n12472) );
  nand_x1_sg U64883 ( .A(n31139), .B(n33860), .X(n12473) );
  nand_x1_sg U64884 ( .A(n30579), .B(n32908), .X(n12476) );
  nand_x1_sg U64885 ( .A(n31141), .B(n33860), .X(n12477) );
  nand_x1_sg U64886 ( .A(n30573), .B(n32906), .X(n12480) );
  nand_x1_sg U64887 ( .A(n31143), .B(n30950), .X(n12481) );
  nand_x1_sg U64888 ( .A(n30578), .B(n32909), .X(n12484) );
  nand_x1_sg U64889 ( .A(n31145), .B(n30949), .X(n12485) );
  nand_x1_sg U64890 ( .A(n30577), .B(n32906), .X(n12488) );
  nand_x1_sg U64891 ( .A(n31147), .B(n33863), .X(n12489) );
  nand_x1_sg U64892 ( .A(n30574), .B(n32907), .X(n12492) );
  nand_x1_sg U64893 ( .A(n31149), .B(n30950), .X(n12493) );
  nand_x1_sg U64894 ( .A(n30576), .B(n32909), .X(n12496) );
  nand_x1_sg U64895 ( .A(n31151), .B(n30949), .X(n12497) );
  nand_x1_sg U64896 ( .A(n30575), .B(n32907), .X(n12500) );
  nand_x1_sg U64897 ( .A(n31153), .B(n33860), .X(n12501) );
  nand_x1_sg U64898 ( .A(n30570), .B(n32908), .X(n12504) );
  nand_x1_sg U64899 ( .A(n31155), .B(n33863), .X(n12505) );
  nand_x1_sg U64900 ( .A(n30568), .B(n32908), .X(n12518) );
  nand_x1_sg U64901 ( .A(n31157), .B(n33862), .X(n12519) );
  nand_x1_sg U64902 ( .A(n30941), .B(n12457), .X(n12455) );
  nand_x1_sg U64903 ( .A(n31131), .B(n33863), .X(n12456) );
endmodule

